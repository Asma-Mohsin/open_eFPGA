magic
tech sky130A
magscale 1 2
timestamp 1733268179
<< obsli1 >>
rect 1104 1071 24840 8721
<< obsm1 >>
rect 198 552 25654 9988
<< metal2 >>
rect 202 9840 258 10000
rect 478 9840 534 10000
rect 754 9840 810 10000
rect 1030 9840 1086 10000
rect 1306 9840 1362 10000
rect 1582 9840 1638 10000
rect 1858 9840 1914 10000
rect 2134 9840 2190 10000
rect 2410 9840 2466 10000
rect 2686 9840 2742 10000
rect 2962 9840 3018 10000
rect 3238 9840 3294 10000
rect 3514 9840 3570 10000
rect 3790 9840 3846 10000
rect 4066 9840 4122 10000
rect 4342 9840 4398 10000
rect 4618 9840 4674 10000
rect 4894 9840 4950 10000
rect 5170 9840 5226 10000
rect 5446 9840 5502 10000
rect 5722 9840 5778 10000
rect 5998 9840 6054 10000
rect 6274 9840 6330 10000
rect 6550 9840 6606 10000
rect 6826 9840 6882 10000
rect 7102 9840 7158 10000
rect 7378 9840 7434 10000
rect 7654 9840 7710 10000
rect 7930 9840 7986 10000
rect 8206 9840 8262 10000
rect 8482 9840 8538 10000
rect 8758 9840 8814 10000
rect 9034 9840 9090 10000
rect 9310 9840 9366 10000
rect 9586 9840 9642 10000
rect 9862 9840 9918 10000
rect 10138 9840 10194 10000
rect 10414 9840 10470 10000
rect 10690 9840 10746 10000
rect 10966 9840 11022 10000
rect 11242 9840 11298 10000
rect 11518 9840 11574 10000
rect 11794 9840 11850 10000
rect 12070 9840 12126 10000
rect 12346 9840 12402 10000
rect 12622 9840 12678 10000
rect 12898 9840 12954 10000
rect 13174 9840 13230 10000
rect 13450 9840 13506 10000
rect 13726 9840 13782 10000
rect 14002 9840 14058 10000
rect 14278 9840 14334 10000
rect 14554 9840 14610 10000
rect 14830 9840 14886 10000
rect 15106 9840 15162 10000
rect 15382 9840 15438 10000
rect 15658 9840 15714 10000
rect 15934 9840 15990 10000
rect 16210 9840 16266 10000
rect 16486 9840 16542 10000
rect 16762 9840 16818 10000
rect 17038 9840 17094 10000
rect 17314 9840 17370 10000
rect 17590 9840 17646 10000
rect 17866 9840 17922 10000
rect 18142 9840 18198 10000
rect 18418 9840 18474 10000
rect 18694 9840 18750 10000
rect 18970 9840 19026 10000
rect 19246 9840 19302 10000
rect 19522 9840 19578 10000
rect 19798 9840 19854 10000
rect 20074 9840 20130 10000
rect 20350 9840 20406 10000
rect 20626 9840 20682 10000
rect 20902 9840 20958 10000
rect 21178 9840 21234 10000
rect 21454 9840 21510 10000
rect 21730 9840 21786 10000
rect 22006 9840 22062 10000
rect 22282 9840 22338 10000
rect 22558 9840 22614 10000
rect 22834 9840 22890 10000
rect 23110 9840 23166 10000
rect 23386 9840 23442 10000
rect 23662 9840 23718 10000
rect 23938 9840 23994 10000
rect 24214 9840 24270 10000
rect 24490 9840 24546 10000
rect 24766 9840 24822 10000
rect 25042 9840 25098 10000
rect 25318 9840 25374 10000
rect 25594 9840 25650 10000
rect 938 0 994 160
rect 2134 0 2190 160
rect 3330 0 3386 160
rect 4526 0 4582 160
rect 5722 0 5778 160
rect 6918 0 6974 160
rect 8114 0 8170 160
rect 9310 0 9366 160
rect 10506 0 10562 160
rect 11702 0 11758 160
rect 12898 0 12954 160
rect 14094 0 14150 160
rect 15290 0 15346 160
rect 16486 0 16542 160
rect 17682 0 17738 160
rect 18878 0 18934 160
rect 20074 0 20130 160
rect 21270 0 21326 160
rect 22466 0 22522 160
rect 23662 0 23718 160
rect 24858 0 24914 160
<< obsm2 >>
rect 314 9784 422 9994
rect 590 9784 698 9994
rect 866 9784 974 9994
rect 1142 9784 1250 9994
rect 1418 9784 1526 9994
rect 1694 9784 1802 9994
rect 1970 9784 2078 9994
rect 2246 9784 2354 9994
rect 2522 9784 2630 9994
rect 2798 9784 2906 9994
rect 3074 9784 3182 9994
rect 3350 9784 3458 9994
rect 3626 9784 3734 9994
rect 3902 9784 4010 9994
rect 4178 9784 4286 9994
rect 4454 9784 4562 9994
rect 4730 9784 4838 9994
rect 5006 9784 5114 9994
rect 5282 9784 5390 9994
rect 5558 9784 5666 9994
rect 5834 9784 5942 9994
rect 6110 9784 6218 9994
rect 6386 9784 6494 9994
rect 6662 9784 6770 9994
rect 6938 9784 7046 9994
rect 7214 9784 7322 9994
rect 7490 9784 7598 9994
rect 7766 9784 7874 9994
rect 8042 9784 8150 9994
rect 8318 9784 8426 9994
rect 8594 9784 8702 9994
rect 8870 9784 8978 9994
rect 9146 9784 9254 9994
rect 9422 9784 9530 9994
rect 9698 9784 9806 9994
rect 9974 9784 10082 9994
rect 10250 9784 10358 9994
rect 10526 9784 10634 9994
rect 10802 9784 10910 9994
rect 11078 9784 11186 9994
rect 11354 9784 11462 9994
rect 11630 9784 11738 9994
rect 11906 9784 12014 9994
rect 12182 9784 12290 9994
rect 12458 9784 12566 9994
rect 12734 9784 12842 9994
rect 13010 9784 13118 9994
rect 13286 9784 13394 9994
rect 13562 9784 13670 9994
rect 13838 9784 13946 9994
rect 14114 9784 14222 9994
rect 14390 9784 14498 9994
rect 14666 9784 14774 9994
rect 14942 9784 15050 9994
rect 15218 9784 15326 9994
rect 15494 9784 15602 9994
rect 15770 9784 15878 9994
rect 16046 9784 16154 9994
rect 16322 9784 16430 9994
rect 16598 9784 16706 9994
rect 16874 9784 16982 9994
rect 17150 9784 17258 9994
rect 17426 9784 17534 9994
rect 17702 9784 17810 9994
rect 17978 9784 18086 9994
rect 18254 9784 18362 9994
rect 18530 9784 18638 9994
rect 18806 9784 18914 9994
rect 19082 9784 19190 9994
rect 19358 9784 19466 9994
rect 19634 9784 19742 9994
rect 19910 9784 20018 9994
rect 20186 9784 20294 9994
rect 20462 9784 20570 9994
rect 20738 9784 20846 9994
rect 21014 9784 21122 9994
rect 21290 9784 21398 9994
rect 21566 9784 21674 9994
rect 21842 9784 21950 9994
rect 22118 9784 22226 9994
rect 22394 9784 22502 9994
rect 22670 9784 22778 9994
rect 22946 9784 23054 9994
rect 23222 9784 23330 9994
rect 23498 9784 23606 9994
rect 23774 9784 23882 9994
rect 24050 9784 24158 9994
rect 24326 9784 24434 9994
rect 24602 9784 24710 9994
rect 24878 9784 24986 9994
rect 25154 9784 25262 9994
rect 25430 9784 25538 9994
rect 204 216 25648 9784
rect 204 54 882 216
rect 1050 54 2078 216
rect 2246 54 3274 216
rect 3442 54 4470 216
rect 4638 54 5666 216
rect 5834 54 6862 216
rect 7030 54 8058 216
rect 8226 54 9254 216
rect 9422 54 10450 216
rect 10618 54 11646 216
rect 11814 54 12842 216
rect 13010 54 14038 216
rect 14206 54 15234 216
rect 15402 54 16430 216
rect 16598 54 17626 216
rect 17794 54 18822 216
rect 18990 54 20018 216
rect 20186 54 21214 216
rect 21382 54 22410 216
rect 22578 54 23606 216
rect 23774 54 24802 216
rect 24970 54 25648 216
<< obsm3 >>
rect 1945 1055 24998 9485
<< metal4 >>
rect 3911 1040 4231 8752
rect 6878 1040 7198 8752
rect 9845 1040 10165 8752
rect 12812 1040 13132 8752
rect 15779 1040 16099 8752
rect 18746 1040 19066 8752
rect 21713 1040 22033 8752
rect 24680 1040 25000 8752
<< labels >>
rlabel metal2 s 2134 0 2190 160 6 FrameStrobe[0]
port 1 nsew signal input
rlabel metal2 s 14094 0 14150 160 6 FrameStrobe[10]
port 2 nsew signal input
rlabel metal2 s 15290 0 15346 160 6 FrameStrobe[11]
port 3 nsew signal input
rlabel metal2 s 16486 0 16542 160 6 FrameStrobe[12]
port 4 nsew signal input
rlabel metal2 s 17682 0 17738 160 6 FrameStrobe[13]
port 5 nsew signal input
rlabel metal2 s 18878 0 18934 160 6 FrameStrobe[14]
port 6 nsew signal input
rlabel metal2 s 20074 0 20130 160 6 FrameStrobe[15]
port 7 nsew signal input
rlabel metal2 s 21270 0 21326 160 6 FrameStrobe[16]
port 8 nsew signal input
rlabel metal2 s 22466 0 22522 160 6 FrameStrobe[17]
port 9 nsew signal input
rlabel metal2 s 23662 0 23718 160 6 FrameStrobe[18]
port 10 nsew signal input
rlabel metal2 s 24858 0 24914 160 6 FrameStrobe[19]
port 11 nsew signal input
rlabel metal2 s 3330 0 3386 160 6 FrameStrobe[1]
port 12 nsew signal input
rlabel metal2 s 4526 0 4582 160 6 FrameStrobe[2]
port 13 nsew signal input
rlabel metal2 s 5722 0 5778 160 6 FrameStrobe[3]
port 14 nsew signal input
rlabel metal2 s 6918 0 6974 160 6 FrameStrobe[4]
port 15 nsew signal input
rlabel metal2 s 8114 0 8170 160 6 FrameStrobe[5]
port 16 nsew signal input
rlabel metal2 s 9310 0 9366 160 6 FrameStrobe[6]
port 17 nsew signal input
rlabel metal2 s 10506 0 10562 160 6 FrameStrobe[7]
port 18 nsew signal input
rlabel metal2 s 11702 0 11758 160 6 FrameStrobe[8]
port 19 nsew signal input
rlabel metal2 s 12898 0 12954 160 6 FrameStrobe[9]
port 20 nsew signal input
rlabel metal2 s 20350 9840 20406 10000 6 FrameStrobe_O[0]
port 21 nsew signal output
rlabel metal2 s 23110 9840 23166 10000 6 FrameStrobe_O[10]
port 22 nsew signal output
rlabel metal2 s 23386 9840 23442 10000 6 FrameStrobe_O[11]
port 23 nsew signal output
rlabel metal2 s 23662 9840 23718 10000 6 FrameStrobe_O[12]
port 24 nsew signal output
rlabel metal2 s 23938 9840 23994 10000 6 FrameStrobe_O[13]
port 25 nsew signal output
rlabel metal2 s 24214 9840 24270 10000 6 FrameStrobe_O[14]
port 26 nsew signal output
rlabel metal2 s 24490 9840 24546 10000 6 FrameStrobe_O[15]
port 27 nsew signal output
rlabel metal2 s 24766 9840 24822 10000 6 FrameStrobe_O[16]
port 28 nsew signal output
rlabel metal2 s 25042 9840 25098 10000 6 FrameStrobe_O[17]
port 29 nsew signal output
rlabel metal2 s 25318 9840 25374 10000 6 FrameStrobe_O[18]
port 30 nsew signal output
rlabel metal2 s 25594 9840 25650 10000 6 FrameStrobe_O[19]
port 31 nsew signal output
rlabel metal2 s 20626 9840 20682 10000 6 FrameStrobe_O[1]
port 32 nsew signal output
rlabel metal2 s 20902 9840 20958 10000 6 FrameStrobe_O[2]
port 33 nsew signal output
rlabel metal2 s 21178 9840 21234 10000 6 FrameStrobe_O[3]
port 34 nsew signal output
rlabel metal2 s 21454 9840 21510 10000 6 FrameStrobe_O[4]
port 35 nsew signal output
rlabel metal2 s 21730 9840 21786 10000 6 FrameStrobe_O[5]
port 36 nsew signal output
rlabel metal2 s 22006 9840 22062 10000 6 FrameStrobe_O[6]
port 37 nsew signal output
rlabel metal2 s 22282 9840 22338 10000 6 FrameStrobe_O[7]
port 38 nsew signal output
rlabel metal2 s 22558 9840 22614 10000 6 FrameStrobe_O[8]
port 39 nsew signal output
rlabel metal2 s 22834 9840 22890 10000 6 FrameStrobe_O[9]
port 40 nsew signal output
rlabel metal2 s 202 9840 258 10000 6 N1BEG[0]
port 41 nsew signal output
rlabel metal2 s 478 9840 534 10000 6 N1BEG[1]
port 42 nsew signal output
rlabel metal2 s 754 9840 810 10000 6 N1BEG[2]
port 43 nsew signal output
rlabel metal2 s 1030 9840 1086 10000 6 N1BEG[3]
port 44 nsew signal output
rlabel metal2 s 1306 9840 1362 10000 6 N2BEG[0]
port 45 nsew signal output
rlabel metal2 s 1582 9840 1638 10000 6 N2BEG[1]
port 46 nsew signal output
rlabel metal2 s 1858 9840 1914 10000 6 N2BEG[2]
port 47 nsew signal output
rlabel metal2 s 2134 9840 2190 10000 6 N2BEG[3]
port 48 nsew signal output
rlabel metal2 s 2410 9840 2466 10000 6 N2BEG[4]
port 49 nsew signal output
rlabel metal2 s 2686 9840 2742 10000 6 N2BEG[5]
port 50 nsew signal output
rlabel metal2 s 2962 9840 3018 10000 6 N2BEG[6]
port 51 nsew signal output
rlabel metal2 s 3238 9840 3294 10000 6 N2BEG[7]
port 52 nsew signal output
rlabel metal2 s 3514 9840 3570 10000 6 N2BEGb[0]
port 53 nsew signal output
rlabel metal2 s 3790 9840 3846 10000 6 N2BEGb[1]
port 54 nsew signal output
rlabel metal2 s 4066 9840 4122 10000 6 N2BEGb[2]
port 55 nsew signal output
rlabel metal2 s 4342 9840 4398 10000 6 N2BEGb[3]
port 56 nsew signal output
rlabel metal2 s 4618 9840 4674 10000 6 N2BEGb[4]
port 57 nsew signal output
rlabel metal2 s 4894 9840 4950 10000 6 N2BEGb[5]
port 58 nsew signal output
rlabel metal2 s 5170 9840 5226 10000 6 N2BEGb[6]
port 59 nsew signal output
rlabel metal2 s 5446 9840 5502 10000 6 N2BEGb[7]
port 60 nsew signal output
rlabel metal2 s 5722 9840 5778 10000 6 N4BEG[0]
port 61 nsew signal output
rlabel metal2 s 8482 9840 8538 10000 6 N4BEG[10]
port 62 nsew signal output
rlabel metal2 s 8758 9840 8814 10000 6 N4BEG[11]
port 63 nsew signal output
rlabel metal2 s 9034 9840 9090 10000 6 N4BEG[12]
port 64 nsew signal output
rlabel metal2 s 9310 9840 9366 10000 6 N4BEG[13]
port 65 nsew signal output
rlabel metal2 s 9586 9840 9642 10000 6 N4BEG[14]
port 66 nsew signal output
rlabel metal2 s 9862 9840 9918 10000 6 N4BEG[15]
port 67 nsew signal output
rlabel metal2 s 5998 9840 6054 10000 6 N4BEG[1]
port 68 nsew signal output
rlabel metal2 s 6274 9840 6330 10000 6 N4BEG[2]
port 69 nsew signal output
rlabel metal2 s 6550 9840 6606 10000 6 N4BEG[3]
port 70 nsew signal output
rlabel metal2 s 6826 9840 6882 10000 6 N4BEG[4]
port 71 nsew signal output
rlabel metal2 s 7102 9840 7158 10000 6 N4BEG[5]
port 72 nsew signal output
rlabel metal2 s 7378 9840 7434 10000 6 N4BEG[6]
port 73 nsew signal output
rlabel metal2 s 7654 9840 7710 10000 6 N4BEG[7]
port 74 nsew signal output
rlabel metal2 s 7930 9840 7986 10000 6 N4BEG[8]
port 75 nsew signal output
rlabel metal2 s 8206 9840 8262 10000 6 N4BEG[9]
port 76 nsew signal output
rlabel metal2 s 10138 9840 10194 10000 6 S1END[0]
port 77 nsew signal input
rlabel metal2 s 10414 9840 10470 10000 6 S1END[1]
port 78 nsew signal input
rlabel metal2 s 10690 9840 10746 10000 6 S1END[2]
port 79 nsew signal input
rlabel metal2 s 10966 9840 11022 10000 6 S1END[3]
port 80 nsew signal input
rlabel metal2 s 11242 9840 11298 10000 6 S2END[0]
port 81 nsew signal input
rlabel metal2 s 11518 9840 11574 10000 6 S2END[1]
port 82 nsew signal input
rlabel metal2 s 11794 9840 11850 10000 6 S2END[2]
port 83 nsew signal input
rlabel metal2 s 12070 9840 12126 10000 6 S2END[3]
port 84 nsew signal input
rlabel metal2 s 12346 9840 12402 10000 6 S2END[4]
port 85 nsew signal input
rlabel metal2 s 12622 9840 12678 10000 6 S2END[5]
port 86 nsew signal input
rlabel metal2 s 12898 9840 12954 10000 6 S2END[6]
port 87 nsew signal input
rlabel metal2 s 13174 9840 13230 10000 6 S2END[7]
port 88 nsew signal input
rlabel metal2 s 13450 9840 13506 10000 6 S2MID[0]
port 89 nsew signal input
rlabel metal2 s 13726 9840 13782 10000 6 S2MID[1]
port 90 nsew signal input
rlabel metal2 s 14002 9840 14058 10000 6 S2MID[2]
port 91 nsew signal input
rlabel metal2 s 14278 9840 14334 10000 6 S2MID[3]
port 92 nsew signal input
rlabel metal2 s 14554 9840 14610 10000 6 S2MID[4]
port 93 nsew signal input
rlabel metal2 s 14830 9840 14886 10000 6 S2MID[5]
port 94 nsew signal input
rlabel metal2 s 15106 9840 15162 10000 6 S2MID[6]
port 95 nsew signal input
rlabel metal2 s 15382 9840 15438 10000 6 S2MID[7]
port 96 nsew signal input
rlabel metal2 s 15658 9840 15714 10000 6 S4END[0]
port 97 nsew signal input
rlabel metal2 s 18418 9840 18474 10000 6 S4END[10]
port 98 nsew signal input
rlabel metal2 s 18694 9840 18750 10000 6 S4END[11]
port 99 nsew signal input
rlabel metal2 s 18970 9840 19026 10000 6 S4END[12]
port 100 nsew signal input
rlabel metal2 s 19246 9840 19302 10000 6 S4END[13]
port 101 nsew signal input
rlabel metal2 s 19522 9840 19578 10000 6 S4END[14]
port 102 nsew signal input
rlabel metal2 s 19798 9840 19854 10000 6 S4END[15]
port 103 nsew signal input
rlabel metal2 s 15934 9840 15990 10000 6 S4END[1]
port 104 nsew signal input
rlabel metal2 s 16210 9840 16266 10000 6 S4END[2]
port 105 nsew signal input
rlabel metal2 s 16486 9840 16542 10000 6 S4END[3]
port 106 nsew signal input
rlabel metal2 s 16762 9840 16818 10000 6 S4END[4]
port 107 nsew signal input
rlabel metal2 s 17038 9840 17094 10000 6 S4END[5]
port 108 nsew signal input
rlabel metal2 s 17314 9840 17370 10000 6 S4END[6]
port 109 nsew signal input
rlabel metal2 s 17590 9840 17646 10000 6 S4END[7]
port 110 nsew signal input
rlabel metal2 s 17866 9840 17922 10000 6 S4END[8]
port 111 nsew signal input
rlabel metal2 s 18142 9840 18198 10000 6 S4END[9]
port 112 nsew signal input
rlabel metal2 s 938 0 994 160 6 UserCLK
port 113 nsew signal input
rlabel metal2 s 20074 9840 20130 10000 6 UserCLKo
port 114 nsew signal output
rlabel metal4 s 6878 1040 7198 8752 6 VGND
port 115 nsew ground bidirectional
rlabel metal4 s 12812 1040 13132 8752 6 VGND
port 115 nsew ground bidirectional
rlabel metal4 s 18746 1040 19066 8752 6 VGND
port 115 nsew ground bidirectional
rlabel metal4 s 24680 1040 25000 8752 6 VGND
port 115 nsew ground bidirectional
rlabel metal4 s 3911 1040 4231 8752 6 VPWR
port 116 nsew power bidirectional
rlabel metal4 s 9845 1040 10165 8752 6 VPWR
port 116 nsew power bidirectional
rlabel metal4 s 15779 1040 16099 8752 6 VPWR
port 116 nsew power bidirectional
rlabel metal4 s 21713 1040 22033 8752 6 VPWR
port 116 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 26000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 432184
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/S_term_RAM_IO/runs/24_12_03_23_21/results/signoff/S_term_RAM_IO.magic.gds
string GDS_START 41360
<< end >>

