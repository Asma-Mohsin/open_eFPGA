VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO S_term_DSP
  CLASS BLOCK ;
  FOREIGN S_term_DSP ;
  ORIGIN 0.000 0.000 ;
  SIZE 225.000 BY 50.000 ;
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 0.800 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 0.800 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 0.800 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 0.800 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 0.800 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 0.800 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 0.800 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 0.800 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 0.800 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 0.800 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 0.800 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 0.800 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 0.800 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 0.800 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 0.800 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 0.800 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 0.800 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 0.800 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 0.800 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 0.800 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 171.670 49.200 171.950 50.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 185.470 49.200 185.750 50.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 186.850 49.200 187.130 50.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 188.230 49.200 188.510 50.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 189.610 49.200 189.890 50.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 190.990 49.200 191.270 50.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 192.370 49.200 192.650 50.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 193.750 49.200 194.030 50.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 195.130 49.200 195.410 50.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 196.510 49.200 196.790 50.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 197.890 49.200 198.170 50.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 173.050 49.200 173.330 50.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 174.430 49.200 174.710 50.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 175.810 49.200 176.090 50.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 177.190 49.200 177.470 50.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 178.570 49.200 178.850 50.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 179.950 49.200 180.230 50.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 181.330 49.200 181.610 50.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 182.710 49.200 182.990 50.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 184.090 49.200 184.370 50.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 26.770 49.200 27.050 50.000 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 28.150 49.200 28.430 50.000 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.530 49.200 29.810 50.000 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 30.910 49.200 31.190 50.000 ;
    END
  END N1BEG[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 49.200 32.570 50.000 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 33.670 49.200 33.950 50.000 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.050 49.200 35.330 50.000 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 36.430 49.200 36.710 50.000 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 37.810 49.200 38.090 50.000 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 39.190 49.200 39.470 50.000 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 40.570 49.200 40.850 50.000 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.950 49.200 42.230 50.000 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 43.330 49.200 43.610 50.000 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 44.710 49.200 44.990 50.000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 46.090 49.200 46.370 50.000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 47.470 49.200 47.750 50.000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.850 49.200 49.130 50.000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 50.230 49.200 50.510 50.000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 49.200 51.890 50.000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 52.990 49.200 53.270 50.000 ;
    END
  END N2BEGb[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.370 49.200 54.650 50.000 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 68.170 49.200 68.450 50.000 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 69.550 49.200 69.830 50.000 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.930 49.200 71.210 50.000 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 72.310 49.200 72.590 50.000 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 73.690 49.200 73.970 50.000 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 75.070 49.200 75.350 50.000 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 55.750 49.200 56.030 50.000 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 57.130 49.200 57.410 50.000 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 58.510 49.200 58.790 50.000 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 59.890 49.200 60.170 50.000 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.270 49.200 61.550 50.000 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 62.650 49.200 62.930 50.000 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.030 49.200 64.310 50.000 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.410 49.200 65.690 50.000 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 66.790 49.200 67.070 50.000 ;
    END
  END N4BEG[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 76.450 49.200 76.730 50.000 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.250 49.200 90.530 50.000 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 91.630 49.200 91.910 50.000 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.010 49.200 93.290 50.000 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 94.390 49.200 94.670 50.000 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 95.770 49.200 96.050 50.000 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 97.150 49.200 97.430 50.000 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.830 49.200 78.110 50.000 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 79.210 49.200 79.490 50.000 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 49.200 80.870 50.000 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 81.970 49.200 82.250 50.000 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.350 49.200 83.630 50.000 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 84.730 49.200 85.010 50.000 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 86.110 49.200 86.390 50.000 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.490 49.200 87.770 50.000 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 88.870 49.200 89.150 50.000 ;
    END
  END NN4BEG[9]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 98.530 49.200 98.810 50.000 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 49.200 100.190 50.000 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 101.290 49.200 101.570 50.000 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 102.670 49.200 102.950 50.000 ;
    END
  END S1END[3]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 104.050 49.200 104.330 50.000 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 105.430 49.200 105.710 50.000 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 106.810 49.200 107.090 50.000 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 108.190 49.200 108.470 50.000 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 49.200 109.850 50.000 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 110.950 49.200 111.230 50.000 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 112.330 49.200 112.610 50.000 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 113.710 49.200 113.990 50.000 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 115.090 49.200 115.370 50.000 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.470 49.200 116.750 50.000 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 117.850 49.200 118.130 50.000 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 49.200 119.510 50.000 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 120.610 49.200 120.890 50.000 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 121.990 49.200 122.270 50.000 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 123.370 49.200 123.650 50.000 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 124.750 49.200 125.030 50.000 ;
    END
  END S2MID[7]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 126.130 49.200 126.410 50.000 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 139.930 49.200 140.210 50.000 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 141.310 49.200 141.590 50.000 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 142.690 49.200 142.970 50.000 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.070 49.200 144.350 50.000 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 145.450 49.200 145.730 50.000 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 146.830 49.200 147.110 50.000 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 127.510 49.200 127.790 50.000 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 49.200 129.170 50.000 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 130.270 49.200 130.550 50.000 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 131.650 49.200 131.930 50.000 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 133.030 49.200 133.310 50.000 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 134.410 49.200 134.690 50.000 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 135.790 49.200 136.070 50.000 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 137.170 49.200 137.450 50.000 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 49.200 138.830 50.000 ;
    END
  END S4END[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 148.210 49.200 148.490 50.000 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 162.010 49.200 162.290 50.000 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 163.390 49.200 163.670 50.000 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 164.770 49.200 165.050 50.000 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 166.150 49.200 166.430 50.000 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 49.200 167.810 50.000 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 168.910 49.200 169.190 50.000 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 149.590 49.200 149.870 50.000 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 150.970 49.200 151.250 50.000 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 152.350 49.200 152.630 50.000 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 153.730 49.200 154.010 50.000 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 155.110 49.200 155.390 50.000 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 156.490 49.200 156.770 50.000 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 157.870 49.200 158.150 50.000 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 159.250 49.200 159.530 50.000 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 160.630 49.200 160.910 50.000 ;
    END
  END SS4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 0.800 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 170.290 49.200 170.570 50.000 ;
    END
  END UserCLKo
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 31.455 5.200 33.055 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.925 5.200 86.525 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.395 5.200 139.995 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 191.865 5.200 193.465 43.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 58.190 5.200 59.790 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.660 5.200 113.260 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 165.130 5.200 166.730 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 218.600 5.200 220.200 43.760 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 39.385 219.610 42.215 ;
        RECT 5.330 33.945 219.610 36.775 ;
        RECT 5.330 28.505 219.610 31.335 ;
        RECT 5.330 23.065 219.610 25.895 ;
        RECT 5.330 17.625 219.610 20.455 ;
        RECT 5.330 12.185 219.610 15.015 ;
        RECT 5.330 6.745 219.610 9.575 ;
      LAYER li1 ;
        RECT 5.520 5.355 219.420 43.605 ;
      LAYER met1 ;
        RECT 5.520 4.460 220.200 49.940 ;
      LAYER met2 ;
        RECT 6.540 48.920 26.490 49.970 ;
        RECT 27.330 48.920 27.870 49.970 ;
        RECT 28.710 48.920 29.250 49.970 ;
        RECT 30.090 48.920 30.630 49.970 ;
        RECT 31.470 48.920 32.010 49.970 ;
        RECT 32.850 48.920 33.390 49.970 ;
        RECT 34.230 48.920 34.770 49.970 ;
        RECT 35.610 48.920 36.150 49.970 ;
        RECT 36.990 48.920 37.530 49.970 ;
        RECT 38.370 48.920 38.910 49.970 ;
        RECT 39.750 48.920 40.290 49.970 ;
        RECT 41.130 48.920 41.670 49.970 ;
        RECT 42.510 48.920 43.050 49.970 ;
        RECT 43.890 48.920 44.430 49.970 ;
        RECT 45.270 48.920 45.810 49.970 ;
        RECT 46.650 48.920 47.190 49.970 ;
        RECT 48.030 48.920 48.570 49.970 ;
        RECT 49.410 48.920 49.950 49.970 ;
        RECT 50.790 48.920 51.330 49.970 ;
        RECT 52.170 48.920 52.710 49.970 ;
        RECT 53.550 48.920 54.090 49.970 ;
        RECT 54.930 48.920 55.470 49.970 ;
        RECT 56.310 48.920 56.850 49.970 ;
        RECT 57.690 48.920 58.230 49.970 ;
        RECT 59.070 48.920 59.610 49.970 ;
        RECT 60.450 48.920 60.990 49.970 ;
        RECT 61.830 48.920 62.370 49.970 ;
        RECT 63.210 48.920 63.750 49.970 ;
        RECT 64.590 48.920 65.130 49.970 ;
        RECT 65.970 48.920 66.510 49.970 ;
        RECT 67.350 48.920 67.890 49.970 ;
        RECT 68.730 48.920 69.270 49.970 ;
        RECT 70.110 48.920 70.650 49.970 ;
        RECT 71.490 48.920 72.030 49.970 ;
        RECT 72.870 48.920 73.410 49.970 ;
        RECT 74.250 48.920 74.790 49.970 ;
        RECT 75.630 48.920 76.170 49.970 ;
        RECT 77.010 48.920 77.550 49.970 ;
        RECT 78.390 48.920 78.930 49.970 ;
        RECT 79.770 48.920 80.310 49.970 ;
        RECT 81.150 48.920 81.690 49.970 ;
        RECT 82.530 48.920 83.070 49.970 ;
        RECT 83.910 48.920 84.450 49.970 ;
        RECT 85.290 48.920 85.830 49.970 ;
        RECT 86.670 48.920 87.210 49.970 ;
        RECT 88.050 48.920 88.590 49.970 ;
        RECT 89.430 48.920 89.970 49.970 ;
        RECT 90.810 48.920 91.350 49.970 ;
        RECT 92.190 48.920 92.730 49.970 ;
        RECT 93.570 48.920 94.110 49.970 ;
        RECT 94.950 48.920 95.490 49.970 ;
        RECT 96.330 48.920 96.870 49.970 ;
        RECT 97.710 48.920 98.250 49.970 ;
        RECT 99.090 48.920 99.630 49.970 ;
        RECT 100.470 48.920 101.010 49.970 ;
        RECT 101.850 48.920 102.390 49.970 ;
        RECT 103.230 48.920 103.770 49.970 ;
        RECT 104.610 48.920 105.150 49.970 ;
        RECT 105.990 48.920 106.530 49.970 ;
        RECT 107.370 48.920 107.910 49.970 ;
        RECT 108.750 48.920 109.290 49.970 ;
        RECT 110.130 48.920 110.670 49.970 ;
        RECT 111.510 48.920 112.050 49.970 ;
        RECT 112.890 48.920 113.430 49.970 ;
        RECT 114.270 48.920 114.810 49.970 ;
        RECT 115.650 48.920 116.190 49.970 ;
        RECT 117.030 48.920 117.570 49.970 ;
        RECT 118.410 48.920 118.950 49.970 ;
        RECT 119.790 48.920 120.330 49.970 ;
        RECT 121.170 48.920 121.710 49.970 ;
        RECT 122.550 48.920 123.090 49.970 ;
        RECT 123.930 48.920 124.470 49.970 ;
        RECT 125.310 48.920 125.850 49.970 ;
        RECT 126.690 48.920 127.230 49.970 ;
        RECT 128.070 48.920 128.610 49.970 ;
        RECT 129.450 48.920 129.990 49.970 ;
        RECT 130.830 48.920 131.370 49.970 ;
        RECT 132.210 48.920 132.750 49.970 ;
        RECT 133.590 48.920 134.130 49.970 ;
        RECT 134.970 48.920 135.510 49.970 ;
        RECT 136.350 48.920 136.890 49.970 ;
        RECT 137.730 48.920 138.270 49.970 ;
        RECT 139.110 48.920 139.650 49.970 ;
        RECT 140.490 48.920 141.030 49.970 ;
        RECT 141.870 48.920 142.410 49.970 ;
        RECT 143.250 48.920 143.790 49.970 ;
        RECT 144.630 48.920 145.170 49.970 ;
        RECT 146.010 48.920 146.550 49.970 ;
        RECT 147.390 48.920 147.930 49.970 ;
        RECT 148.770 48.920 149.310 49.970 ;
        RECT 150.150 48.920 150.690 49.970 ;
        RECT 151.530 48.920 152.070 49.970 ;
        RECT 152.910 48.920 153.450 49.970 ;
        RECT 154.290 48.920 154.830 49.970 ;
        RECT 155.670 48.920 156.210 49.970 ;
        RECT 157.050 48.920 157.590 49.970 ;
        RECT 158.430 48.920 158.970 49.970 ;
        RECT 159.810 48.920 160.350 49.970 ;
        RECT 161.190 48.920 161.730 49.970 ;
        RECT 162.570 48.920 163.110 49.970 ;
        RECT 163.950 48.920 164.490 49.970 ;
        RECT 165.330 48.920 165.870 49.970 ;
        RECT 166.710 48.920 167.250 49.970 ;
        RECT 168.090 48.920 168.630 49.970 ;
        RECT 169.470 48.920 170.010 49.970 ;
        RECT 170.850 48.920 171.390 49.970 ;
        RECT 172.230 48.920 172.770 49.970 ;
        RECT 173.610 48.920 174.150 49.970 ;
        RECT 174.990 48.920 175.530 49.970 ;
        RECT 176.370 48.920 176.910 49.970 ;
        RECT 177.750 48.920 178.290 49.970 ;
        RECT 179.130 48.920 179.670 49.970 ;
        RECT 180.510 48.920 181.050 49.970 ;
        RECT 181.890 48.920 182.430 49.970 ;
        RECT 183.270 48.920 183.810 49.970 ;
        RECT 184.650 48.920 185.190 49.970 ;
        RECT 186.030 48.920 186.570 49.970 ;
        RECT 187.410 48.920 187.950 49.970 ;
        RECT 188.790 48.920 189.330 49.970 ;
        RECT 190.170 48.920 190.710 49.970 ;
        RECT 191.550 48.920 192.090 49.970 ;
        RECT 192.930 48.920 193.470 49.970 ;
        RECT 194.310 48.920 194.850 49.970 ;
        RECT 195.690 48.920 196.230 49.970 ;
        RECT 197.070 48.920 197.610 49.970 ;
        RECT 198.450 48.920 220.170 49.970 ;
        RECT 6.540 1.080 220.170 48.920 ;
        RECT 7.090 0.270 16.830 1.080 ;
        RECT 17.670 0.270 27.410 1.080 ;
        RECT 28.250 0.270 37.990 1.080 ;
        RECT 38.830 0.270 48.570 1.080 ;
        RECT 49.410 0.270 59.150 1.080 ;
        RECT 59.990 0.270 69.730 1.080 ;
        RECT 70.570 0.270 80.310 1.080 ;
        RECT 81.150 0.270 90.890 1.080 ;
        RECT 91.730 0.270 101.470 1.080 ;
        RECT 102.310 0.270 112.050 1.080 ;
        RECT 112.890 0.270 122.630 1.080 ;
        RECT 123.470 0.270 133.210 1.080 ;
        RECT 134.050 0.270 143.790 1.080 ;
        RECT 144.630 0.270 154.370 1.080 ;
        RECT 155.210 0.270 164.950 1.080 ;
        RECT 165.790 0.270 175.530 1.080 ;
        RECT 176.370 0.270 186.110 1.080 ;
        RECT 186.950 0.270 196.690 1.080 ;
        RECT 197.530 0.270 207.270 1.080 ;
        RECT 208.110 0.270 217.850 1.080 ;
        RECT 218.690 0.270 220.170 1.080 ;
      LAYER met3 ;
        RECT 24.445 5.275 220.190 49.465 ;
      LAYER met4 ;
        RECT 96.895 34.855 100.905 49.465 ;
  END
END S_term_DSP
END LIBRARY

