magic
tech sky130A
magscale 1 2
timestamp 1733308228
<< viali >>
rect 5181 8585 5215 8619
rect 5733 8585 5767 8619
rect 7297 8585 7331 8619
rect 8309 8585 8343 8619
rect 9781 8585 9815 8619
rect 10149 8585 10183 8619
rect 10701 8585 10735 8619
rect 11253 8585 11287 8619
rect 12357 8585 12391 8619
rect 13277 8585 13311 8619
rect 13829 8585 13863 8619
rect 14381 8585 14415 8619
rect 15301 8585 15335 8619
rect 15853 8585 15887 8619
rect 16405 8585 16439 8619
rect 16957 8585 16991 8619
rect 17325 8585 17359 8619
rect 17877 8585 17911 8619
rect 18245 8585 18279 8619
rect 18613 8585 18647 8619
rect 18981 8585 19015 8619
rect 19533 8585 19567 8619
rect 20085 8585 20119 8619
rect 21189 8585 21223 8619
rect 22293 8585 22327 8619
rect 22845 8585 22879 8619
rect 30297 8585 30331 8619
rect 31125 8585 31159 8619
rect 31401 8585 31435 8619
rect 31677 8585 31711 8619
rect 33701 8585 33735 8619
rect 34345 8585 34379 8619
rect 34897 8585 34931 8619
rect 36001 8585 36035 8619
rect 36553 8585 36587 8619
rect 39129 8585 39163 8619
rect 41153 8585 41187 8619
rect 4537 8517 4571 8551
rect 4905 8517 4939 8551
rect 6837 8517 6871 8551
rect 7205 8517 7239 8551
rect 10425 8517 10459 8551
rect 12081 8517 12115 8551
rect 13553 8517 13587 8551
rect 17601 8517 17635 8551
rect 37381 8517 37415 8551
rect 37933 8517 37967 8551
rect 38485 8517 38519 8551
rect 38853 8517 38887 8551
rect 40877 8517 40911 8551
rect 5457 8449 5491 8483
rect 5917 8449 5951 8483
rect 8033 8449 8067 8483
rect 8493 8449 8527 8483
rect 9045 8449 9079 8483
rect 9505 8449 9539 8483
rect 9965 8449 9999 8483
rect 10977 8449 11011 8483
rect 11621 8449 11655 8483
rect 12817 8449 12851 8483
rect 13093 8449 13127 8483
rect 14197 8449 14231 8483
rect 14565 8449 14599 8483
rect 15025 8449 15059 8483
rect 15669 8449 15703 8483
rect 16129 8449 16163 8483
rect 16773 8449 16807 8483
rect 17141 8449 17175 8483
rect 18061 8449 18095 8483
rect 18429 8449 18463 8483
rect 18797 8449 18831 8483
rect 19441 8449 19475 8483
rect 19993 8449 20027 8483
rect 20821 8449 20855 8483
rect 21097 8449 21131 8483
rect 21373 8449 21407 8483
rect 21649 8449 21683 8483
rect 22201 8449 22235 8483
rect 22477 8449 22511 8483
rect 22753 8449 22787 8483
rect 23029 8449 23063 8483
rect 23305 8449 23339 8483
rect 23581 8449 23615 8483
rect 23857 8449 23891 8483
rect 24133 8449 24167 8483
rect 24593 8449 24627 8483
rect 24869 8449 24903 8483
rect 25145 8449 25179 8483
rect 25421 8449 25455 8483
rect 25697 8449 25731 8483
rect 25973 8449 26007 8483
rect 26249 8449 26283 8483
rect 26525 8449 26559 8483
rect 26801 8449 26835 8483
rect 27169 8449 27203 8483
rect 27445 8449 27479 8483
rect 27721 8449 27755 8483
rect 27997 8449 28031 8483
rect 28273 8449 28307 8483
rect 28549 8449 28583 8483
rect 28825 8449 28859 8483
rect 29101 8449 29135 8483
rect 29377 8449 29411 8483
rect 29745 8449 29779 8483
rect 30021 8449 30055 8483
rect 30113 8449 30147 8483
rect 30389 8449 30423 8483
rect 30665 8449 30699 8483
rect 30941 8449 30975 8483
rect 31217 8449 31251 8483
rect 31493 8449 31527 8483
rect 31769 8449 31803 8483
rect 32137 8449 32171 8483
rect 32413 8449 32447 8483
rect 32689 8449 32723 8483
rect 32965 8449 32999 8483
rect 33241 8449 33275 8483
rect 33517 8449 33551 8483
rect 33793 8449 33827 8483
rect 34161 8449 34195 8483
rect 34805 8449 34839 8483
rect 35265 8449 35299 8483
rect 35909 8449 35943 8483
rect 36461 8449 36495 8483
rect 39037 8449 39071 8483
rect 39957 8449 39991 8483
rect 40509 8449 40543 8483
rect 41061 8449 41095 8483
rect 6101 8313 6135 8347
rect 8677 8313 8711 8347
rect 9229 8313 9263 8347
rect 11805 8313 11839 8347
rect 14749 8313 14783 8347
rect 22569 8313 22603 8347
rect 28917 8313 28951 8347
rect 29193 8313 29227 8347
rect 30573 8313 30607 8347
rect 30849 8313 30883 8347
rect 31953 8313 31987 8347
rect 32597 8313 32631 8347
rect 32873 8313 32907 8347
rect 33977 8313 34011 8347
rect 35449 8313 35483 8347
rect 37565 8313 37599 8347
rect 38117 8313 38151 8347
rect 40141 8313 40175 8347
rect 20637 8245 20671 8279
rect 20913 8245 20947 8279
rect 21465 8245 21499 8279
rect 22017 8245 22051 8279
rect 23121 8245 23155 8279
rect 23397 8245 23431 8279
rect 23673 8245 23707 8279
rect 23949 8245 23983 8279
rect 24409 8245 24443 8279
rect 24685 8245 24719 8279
rect 24961 8245 24995 8279
rect 25237 8245 25271 8279
rect 25513 8245 25547 8279
rect 25789 8245 25823 8279
rect 26065 8245 26099 8279
rect 26341 8245 26375 8279
rect 26617 8245 26651 8279
rect 26985 8245 27019 8279
rect 27261 8245 27295 8279
rect 27537 8245 27571 8279
rect 27813 8245 27847 8279
rect 28089 8245 28123 8279
rect 28365 8245 28399 8279
rect 28641 8245 28675 8279
rect 29561 8245 29595 8279
rect 29837 8245 29871 8279
rect 32321 8245 32355 8279
rect 33149 8245 33183 8279
rect 33425 8245 33459 8279
rect 5733 8041 5767 8075
rect 6285 8041 6319 8075
rect 7573 8041 7607 8075
rect 7941 8041 7975 8075
rect 8493 8041 8527 8075
rect 9321 8041 9355 8075
rect 10149 8041 10183 8075
rect 11253 8041 11287 8075
rect 11805 8041 11839 8075
rect 13277 8041 13311 8075
rect 13829 8041 13863 8075
rect 14565 8041 14599 8075
rect 15117 8041 15151 8075
rect 15669 8041 15703 8075
rect 17049 8041 17083 8075
rect 17417 8041 17451 8075
rect 18889 8041 18923 8075
rect 20177 8041 20211 8075
rect 20453 8041 20487 8075
rect 21373 8041 21407 8075
rect 22937 8041 22971 8075
rect 23213 8041 23247 8075
rect 24593 8041 24627 8075
rect 25421 8041 25455 8075
rect 25697 8041 25731 8075
rect 26525 8041 26559 8075
rect 27629 8041 27663 8075
rect 27905 8041 27939 8075
rect 28181 8041 28215 8075
rect 35633 8041 35667 8075
rect 36277 8041 36311 8075
rect 36829 8041 36863 8075
rect 37657 8041 37691 8075
rect 38209 8041 38243 8075
rect 38761 8041 38795 8075
rect 39313 8041 39347 8075
rect 40601 8041 40635 8075
rect 6929 7973 6963 8007
rect 12449 7973 12483 8007
rect 16589 7973 16623 8007
rect 17969 7973 18003 8007
rect 18337 7973 18371 8007
rect 19441 7973 19475 8007
rect 20821 7973 20855 8007
rect 22661 7973 22695 8007
rect 24041 7973 24075 8007
rect 6193 7837 6227 7871
rect 7389 7837 7423 7871
rect 11161 7837 11195 7871
rect 13001 7837 13035 7871
rect 14933 7837 14967 7871
rect 16957 7837 16991 7871
rect 17601 7837 17635 7871
rect 18521 7837 18555 7871
rect 18797 7837 18831 7871
rect 19073 7837 19107 7871
rect 19625 7837 19659 7871
rect 19901 7837 19935 7871
rect 19993 7837 20027 7871
rect 20269 7813 20303 7847
rect 20545 7837 20579 7871
rect 21005 7837 21039 7871
rect 21097 7837 21131 7871
rect 21557 7837 21591 7871
rect 21649 7837 21683 7871
rect 21925 7837 21959 7871
rect 22201 7837 22235 7871
rect 22477 7837 22511 7871
rect 22753 7837 22787 7871
rect 23029 7837 23063 7871
rect 23297 7837 23331 7871
rect 23581 7837 23615 7871
rect 23857 7837 23891 7871
rect 24409 7837 24443 7871
rect 24685 7837 24719 7871
rect 24961 7837 24995 7871
rect 25237 7837 25271 7871
rect 25513 7837 25547 7871
rect 25789 7837 25823 7871
rect 26065 7837 26099 7871
rect 26341 7837 26375 7871
rect 26617 7837 26651 7871
rect 26893 7837 26927 7871
rect 27169 7837 27203 7871
rect 27445 7837 27479 7871
rect 27721 7837 27755 7871
rect 27997 7837 28031 7871
rect 33609 7837 33643 7871
rect 33885 7837 33919 7871
rect 35449 7837 35483 7871
rect 5641 7769 5675 7803
rect 6745 7769 6779 7803
rect 7849 7769 7883 7803
rect 8401 7769 8435 7803
rect 9229 7769 9263 7803
rect 10057 7769 10091 7803
rect 11713 7769 11747 7803
rect 12265 7769 12299 7803
rect 13553 7769 13587 7803
rect 14473 7769 14507 7803
rect 15577 7769 15611 7803
rect 16405 7769 16439 7803
rect 17785 7769 17819 7803
rect 36185 7769 36219 7803
rect 36737 7769 36771 7803
rect 37565 7769 37599 7803
rect 38117 7769 38151 7803
rect 38669 7769 38703 7803
rect 39221 7769 39255 7803
rect 39957 7769 39991 7803
rect 40509 7769 40543 7803
rect 18613 7701 18647 7735
rect 19717 7701 19751 7735
rect 20729 7701 20763 7735
rect 21281 7701 21315 7735
rect 21833 7701 21867 7735
rect 22109 7701 22143 7735
rect 22385 7701 22419 7735
rect 23489 7701 23523 7735
rect 23765 7701 23799 7735
rect 24869 7701 24903 7735
rect 25145 7701 25179 7735
rect 25973 7701 26007 7735
rect 26249 7701 26283 7735
rect 26801 7701 26835 7735
rect 27077 7701 27111 7735
rect 27353 7701 27387 7735
rect 33793 7701 33827 7735
rect 34069 7701 34103 7735
rect 40049 7701 40083 7735
rect 6101 7497 6135 7531
rect 7205 7497 7239 7531
rect 8033 7497 8067 7531
rect 11989 7497 12023 7531
rect 12909 7497 12943 7531
rect 17509 7497 17543 7531
rect 18153 7497 18187 7531
rect 18705 7497 18739 7531
rect 19901 7497 19935 7531
rect 22937 7497 22971 7531
rect 23489 7497 23523 7531
rect 6561 7429 6595 7463
rect 5917 7361 5951 7395
rect 7021 7361 7055 7395
rect 7389 7361 7423 7395
rect 11805 7361 11839 7395
rect 12725 7361 12759 7395
rect 17693 7361 17727 7395
rect 17969 7361 18003 7395
rect 18337 7361 18371 7395
rect 18613 7361 18647 7395
rect 18889 7361 18923 7395
rect 19165 7361 19199 7395
rect 19441 7361 19475 7395
rect 19717 7361 19751 7395
rect 19993 7361 20027 7395
rect 20545 7361 20579 7395
rect 20821 7361 20855 7395
rect 21281 7361 21315 7395
rect 21373 7361 21407 7395
rect 22017 7361 22051 7395
rect 22293 7361 22327 7395
rect 22753 7361 22787 7395
rect 23305 7361 23339 7395
rect 26433 7361 26467 7395
rect 7573 7225 7607 7259
rect 19349 7225 19383 7259
rect 19625 7225 19659 7259
rect 20361 7225 20395 7259
rect 21097 7225 21131 7259
rect 21833 7225 21867 7259
rect 22109 7225 22143 7259
rect 17785 7157 17819 7191
rect 18429 7157 18463 7191
rect 20177 7157 20211 7191
rect 21005 7157 21039 7191
rect 21557 7157 21591 7191
rect 26617 7157 26651 7191
rect 20085 6953 20119 6987
rect 7021 6749 7055 6783
rect 18797 6749 18831 6783
rect 19993 6749 20027 6783
rect 20269 6749 20303 6783
rect 18613 6613 18647 6647
rect 19809 6613 19843 6647
rect 37473 5321 37507 5355
rect 37657 5185 37691 5219
rect 22753 4777 22787 4811
rect 26065 4777 26099 4811
rect 28181 4777 28215 4811
rect 36645 4777 36679 4811
rect 38209 4777 38243 4811
rect 21833 4709 21867 4743
rect 23029 4709 23063 4743
rect 32413 4709 32447 4743
rect 21649 4573 21683 4607
rect 22569 4573 22603 4607
rect 22845 4573 22879 4607
rect 23121 4573 23155 4607
rect 23397 4573 23431 4607
rect 25881 4573 25915 4607
rect 27997 4573 28031 4607
rect 32229 4573 32263 4607
rect 36829 4573 36863 4607
rect 38393 4573 38427 4607
rect 23305 4437 23339 4471
rect 23581 4437 23615 4471
rect 20913 4233 20947 4267
rect 22109 4233 22143 4267
rect 22661 4233 22695 4267
rect 25145 4233 25179 4267
rect 37657 4233 37691 4267
rect 21097 4097 21131 4131
rect 22017 4097 22051 4131
rect 22293 4097 22327 4131
rect 22569 4097 22603 4131
rect 22845 4097 22879 4131
rect 23765 4097 23799 4131
rect 25329 4097 25363 4131
rect 27445 4097 27479 4131
rect 31677 4097 31711 4131
rect 37841 4097 37875 4131
rect 21833 3961 21867 3995
rect 27261 3961 27295 3995
rect 31493 3961 31527 3995
rect 22385 3893 22419 3927
rect 23949 3893 23983 3927
rect 23029 3689 23063 3723
rect 30297 3689 30331 3723
rect 37289 3689 37323 3723
rect 39957 3689 39991 3723
rect 19717 3621 19751 3655
rect 19533 3485 19567 3519
rect 23213 3485 23247 3519
rect 30113 3485 30147 3519
rect 37473 3485 37507 3519
rect 40141 3485 40175 3519
rect 18797 3145 18831 3179
rect 22569 3145 22603 3179
rect 29377 3145 29411 3179
rect 36185 3145 36219 3179
rect 40693 3145 40727 3179
rect 18981 3009 19015 3043
rect 22017 3009 22051 3043
rect 22385 3009 22419 3043
rect 29561 3009 29595 3043
rect 36369 3009 36403 3043
rect 40877 3009 40911 3043
rect 22201 2873 22235 2907
rect 21281 2601 21315 2635
rect 39865 2601 39899 2635
rect 21557 2533 21591 2567
rect 38945 2533 38979 2567
rect 21465 2397 21499 2431
rect 21741 2397 21775 2431
rect 22845 2397 22879 2431
rect 39129 2397 39163 2431
rect 40049 2397 40083 2431
rect 23029 2261 23063 2295
rect 22109 2057 22143 2091
rect 39221 2057 39255 2091
rect 40049 2057 40083 2091
rect 21833 1921 21867 1955
rect 22293 1921 22327 1955
rect 39405 1921 39439 1955
rect 40233 1921 40267 1955
rect 22017 1785 22051 1819
rect 1593 1513 1627 1547
rect 3985 1513 4019 1547
rect 39497 1513 39531 1547
rect 43361 1513 43395 1547
rect 12173 1445 12207 1479
rect 16221 1445 16255 1479
rect 1409 1309 1443 1343
rect 3801 1309 3835 1343
rect 5641 1309 5675 1343
rect 7757 1309 7791 1343
rect 9873 1309 9907 1343
rect 11989 1309 12023 1343
rect 14289 1309 14323 1343
rect 16405 1309 16439 1343
rect 18521 1309 18555 1343
rect 20637 1309 20671 1343
rect 22753 1309 22787 1343
rect 24869 1309 24903 1343
rect 27169 1309 27203 1343
rect 29101 1309 29135 1343
rect 31217 1309 31251 1343
rect 33333 1309 33367 1343
rect 35449 1309 35483 1343
rect 37565 1309 37599 1343
rect 39681 1309 39715 1343
rect 41797 1309 41831 1343
rect 43545 1309 43579 1343
rect 5825 1173 5859 1207
rect 7941 1173 7975 1207
rect 10057 1173 10091 1207
rect 14105 1173 14139 1207
rect 18337 1173 18371 1207
rect 20453 1173 20487 1207
rect 22569 1173 22603 1207
rect 24685 1173 24719 1207
rect 26985 1173 27019 1207
rect 28917 1173 28951 1207
rect 31033 1173 31067 1207
rect 33149 1173 33183 1207
rect 35265 1173 35299 1207
rect 37381 1173 37415 1207
rect 41613 1173 41647 1207
<< metal1 >>
rect 17586 9976 17592 9988
rect 9048 9948 17592 9976
rect 9048 9784 9076 9948
rect 17586 9936 17592 9948
rect 17644 9936 17650 9988
rect 19058 9936 19064 9988
rect 19116 9976 19122 9988
rect 31662 9976 31668 9988
rect 19116 9948 31668 9976
rect 19116 9936 19122 9948
rect 31662 9936 31668 9948
rect 31720 9936 31726 9988
rect 17678 9868 17684 9920
rect 17736 9908 17742 9920
rect 21450 9908 21456 9920
rect 17736 9880 21456 9908
rect 17736 9868 17742 9880
rect 21450 9868 21456 9880
rect 21508 9868 21514 9920
rect 22922 9840 22928 9852
rect 17236 9812 22928 9840
rect 9030 9732 9036 9784
rect 9088 9732 9094 9784
rect 17034 9704 17040 9716
rect 8312 9676 17040 9704
rect 8312 9376 8340 9676
rect 17034 9664 17040 9676
rect 17092 9664 17098 9716
rect 17236 9636 17264 9812
rect 22922 9800 22928 9812
rect 22980 9800 22986 9852
rect 27338 9772 27344 9784
rect 10428 9608 17264 9636
rect 17328 9744 27344 9772
rect 10428 9444 10456 9608
rect 13170 9528 13176 9580
rect 13228 9568 13234 9580
rect 17328 9568 17356 9744
rect 27338 9732 27344 9744
rect 27396 9732 27402 9784
rect 17586 9664 17592 9716
rect 17644 9704 17650 9716
rect 20530 9704 20536 9716
rect 17644 9676 20536 9704
rect 17644 9664 17650 9676
rect 20530 9664 20536 9676
rect 20588 9664 20594 9716
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 25590 9704 25596 9716
rect 20772 9676 25596 9704
rect 20772 9664 20778 9676
rect 25590 9664 25596 9676
rect 25648 9664 25654 9716
rect 17402 9596 17408 9648
rect 17460 9636 17466 9648
rect 23198 9636 23204 9648
rect 17460 9608 23204 9636
rect 17460 9596 17466 9608
rect 23198 9596 23204 9608
rect 23256 9596 23262 9648
rect 29270 9596 29276 9648
rect 29328 9636 29334 9648
rect 37550 9636 37556 9648
rect 29328 9608 37556 9636
rect 29328 9596 29334 9608
rect 37550 9596 37556 9608
rect 37608 9596 37614 9648
rect 13228 9540 17356 9568
rect 13228 9528 13234 9540
rect 19610 9528 19616 9580
rect 19668 9568 19674 9580
rect 32858 9568 32864 9580
rect 19668 9540 32864 9568
rect 19668 9528 19674 9540
rect 32858 9528 32864 9540
rect 32916 9528 32922 9580
rect 25406 9500 25412 9512
rect 14384 9472 25412 9500
rect 14384 9444 14412 9472
rect 25406 9460 25412 9472
rect 25464 9460 25470 9512
rect 10410 9392 10416 9444
rect 10468 9392 10474 9444
rect 14366 9392 14372 9444
rect 14424 9392 14430 9444
rect 16022 9392 16028 9444
rect 16080 9432 16086 9444
rect 25682 9432 25688 9444
rect 16080 9404 25688 9432
rect 16080 9392 16086 9404
rect 25682 9392 25688 9404
rect 25740 9392 25746 9444
rect 26786 9392 26792 9444
rect 26844 9432 26850 9444
rect 32030 9432 32036 9444
rect 26844 9404 32036 9432
rect 26844 9392 26850 9404
rect 32030 9392 32036 9404
rect 32088 9392 32094 9444
rect 8294 9324 8300 9376
rect 8352 9324 8358 9376
rect 19978 9364 19984 9376
rect 9968 9336 19984 9364
rect 9968 9240 9996 9336
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 20162 9324 20168 9376
rect 20220 9364 20226 9376
rect 21266 9364 21272 9376
rect 20220 9336 21272 9364
rect 20220 9324 20226 9336
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 21358 9324 21364 9376
rect 21416 9364 21422 9376
rect 32766 9364 32772 9376
rect 21416 9336 32772 9364
rect 21416 9324 21422 9336
rect 32766 9324 32772 9336
rect 32824 9324 32830 9376
rect 17034 9256 17040 9308
rect 17092 9296 17098 9308
rect 19058 9296 19064 9308
rect 17092 9268 19064 9296
rect 17092 9256 17098 9268
rect 19058 9256 19064 9268
rect 19116 9256 19122 9308
rect 19150 9256 19156 9308
rect 19208 9296 19214 9308
rect 31386 9296 31392 9308
rect 19208 9268 31392 9296
rect 19208 9256 19214 9268
rect 31386 9256 31392 9268
rect 31444 9256 31450 9308
rect 9950 9188 9956 9240
rect 10008 9188 10014 9240
rect 28166 9228 28172 9240
rect 12406 9200 28172 9228
rect 12066 8916 12072 8968
rect 12124 8956 12130 8968
rect 12406 8956 12434 9200
rect 28166 9188 28172 9200
rect 28224 9188 28230 9240
rect 31478 9188 31484 9240
rect 31536 9228 31542 9240
rect 36630 9228 36636 9240
rect 31536 9200 36636 9228
rect 31536 9188 31542 9200
rect 36630 9188 36636 9200
rect 36688 9188 36694 9240
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 17402 9160 17408 9172
rect 15160 9132 17408 9160
rect 15160 9120 15166 9132
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 17586 9120 17592 9172
rect 17644 9160 17650 9172
rect 31110 9160 31116 9172
rect 17644 9132 31116 9160
rect 17644 9120 17650 9132
rect 31110 9120 31116 9132
rect 31168 9120 31174 9172
rect 33594 9160 33600 9172
rect 31220 9132 33600 9160
rect 13446 9052 13452 9104
rect 13504 9092 13510 9104
rect 20714 9092 20720 9104
rect 13504 9064 20720 9092
rect 13504 9052 13510 9064
rect 20714 9052 20720 9064
rect 20772 9052 20778 9104
rect 21450 9052 21456 9104
rect 21508 9092 21514 9104
rect 26786 9092 26792 9104
rect 21508 9064 26792 9092
rect 21508 9052 21514 9064
rect 26786 9052 26792 9064
rect 26844 9052 26850 9104
rect 26878 9052 26884 9104
rect 26936 9092 26942 9104
rect 31220 9092 31248 9132
rect 33594 9120 33600 9132
rect 33652 9120 33658 9172
rect 37458 9092 37464 9104
rect 26936 9064 31248 9092
rect 31312 9064 37464 9092
rect 26936 9052 26942 9064
rect 14642 8984 14648 9036
rect 14700 9024 14706 9036
rect 15838 9024 15844 9036
rect 14700 8996 15844 9024
rect 14700 8984 14706 8996
rect 15838 8984 15844 8996
rect 15896 8984 15902 9036
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 18690 9024 18696 9036
rect 16632 8996 18696 9024
rect 16632 8984 16638 8996
rect 18690 8984 18696 8996
rect 18748 8984 18754 9036
rect 30558 9024 30564 9036
rect 18984 8996 30564 9024
rect 18984 8968 19012 8996
rect 30558 8984 30564 8996
rect 30616 8984 30622 9036
rect 30650 8984 30656 9036
rect 30708 9024 30714 9036
rect 31312 9024 31340 9064
rect 37458 9052 37464 9064
rect 37516 9052 37522 9104
rect 33686 9024 33692 9036
rect 30708 8996 31340 9024
rect 31726 8996 33692 9024
rect 30708 8984 30714 8996
rect 12124 8928 12434 8956
rect 12124 8916 12130 8928
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 18414 8956 18420 8968
rect 14976 8928 18420 8956
rect 14976 8916 14982 8928
rect 18414 8916 18420 8928
rect 18472 8916 18478 8968
rect 18966 8916 18972 8968
rect 19024 8916 19030 8968
rect 19058 8916 19064 8968
rect 19116 8956 19122 8968
rect 19116 8928 23244 8956
rect 19116 8916 19122 8928
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 20714 8888 20720 8900
rect 8260 8860 20720 8888
rect 8260 8848 8266 8860
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 16574 8820 16580 8832
rect 9916 8792 16580 8820
rect 9916 8780 9922 8792
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 16758 8780 16764 8832
rect 16816 8820 16822 8832
rect 20162 8820 20168 8832
rect 16816 8792 20168 8820
rect 16816 8780 16822 8792
rect 20162 8780 20168 8792
rect 20220 8780 20226 8832
rect 20530 8780 20536 8832
rect 20588 8820 20594 8832
rect 20990 8820 20996 8832
rect 20588 8792 20996 8820
rect 20588 8780 20594 8792
rect 20990 8780 20996 8792
rect 21048 8780 21054 8832
rect 23216 8820 23244 8928
rect 24578 8916 24584 8968
rect 24636 8956 24642 8968
rect 31726 8956 31754 8996
rect 33686 8984 33692 8996
rect 33744 8984 33750 9036
rect 24636 8928 31754 8956
rect 24636 8916 24642 8928
rect 28994 8848 29000 8900
rect 29052 8888 29058 8900
rect 35250 8888 35256 8900
rect 29052 8860 35256 8888
rect 29052 8848 29058 8860
rect 35250 8848 35256 8860
rect 35308 8848 35314 8900
rect 36078 8848 36084 8900
rect 36136 8888 36142 8900
rect 39022 8888 39028 8900
rect 36136 8860 39028 8888
rect 36136 8848 36142 8860
rect 39022 8848 39028 8860
rect 39080 8848 39086 8900
rect 30282 8820 30288 8832
rect 23216 8792 30288 8820
rect 30282 8780 30288 8792
rect 30340 8780 30346 8832
rect 30374 8780 30380 8832
rect 30432 8820 30438 8832
rect 34974 8820 34980 8832
rect 30432 8792 34980 8820
rect 30432 8780 30438 8792
rect 34974 8780 34980 8792
rect 35032 8780 35038 8832
rect 36814 8780 36820 8832
rect 36872 8820 36878 8832
rect 38654 8820 38660 8832
rect 36872 8792 38660 8820
rect 36872 8780 36878 8792
rect 38654 8780 38660 8792
rect 38712 8780 38718 8832
rect 1104 8730 44040 8752
rect 1104 8678 11644 8730
rect 11696 8678 11708 8730
rect 11760 8678 11772 8730
rect 11824 8678 11836 8730
rect 11888 8678 11900 8730
rect 11952 8678 22338 8730
rect 22390 8678 22402 8730
rect 22454 8678 22466 8730
rect 22518 8678 22530 8730
rect 22582 8678 22594 8730
rect 22646 8678 33032 8730
rect 33084 8678 33096 8730
rect 33148 8678 33160 8730
rect 33212 8678 33224 8730
rect 33276 8678 33288 8730
rect 33340 8678 43726 8730
rect 43778 8678 43790 8730
rect 43842 8678 43854 8730
rect 43906 8678 43918 8730
rect 43970 8678 43982 8730
rect 44034 8678 44040 8730
rect 1104 8656 44040 8678
rect 5169 8619 5227 8625
rect 5169 8585 5181 8619
rect 5215 8616 5227 8619
rect 5350 8616 5356 8628
rect 5215 8588 5356 8616
rect 5215 8585 5227 8588
rect 5169 8579 5227 8585
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 5902 8616 5908 8628
rect 5767 8588 5908 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 7285 8619 7343 8625
rect 7285 8616 7297 8619
rect 7064 8588 7297 8616
rect 7064 8576 7070 8588
rect 7285 8585 7297 8588
rect 7331 8585 7343 8619
rect 7285 8579 7343 8585
rect 8202 8576 8208 8628
rect 8260 8576 8266 8628
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8616 8355 8619
rect 8662 8616 8668 8628
rect 8343 8588 8668 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 9490 8576 9496 8628
rect 9548 8576 9554 8628
rect 9766 8576 9772 8628
rect 9824 8576 9830 8628
rect 10137 8619 10195 8625
rect 10137 8585 10149 8619
rect 10183 8616 10195 8619
rect 10594 8616 10600 8628
rect 10183 8588 10600 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 10689 8619 10747 8625
rect 10689 8585 10701 8619
rect 10735 8616 10747 8619
rect 10870 8616 10876 8628
rect 10735 8588 10876 8616
rect 10735 8585 10747 8588
rect 10689 8579 10747 8585
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 11241 8619 11299 8625
rect 11241 8585 11253 8619
rect 11287 8616 11299 8619
rect 11422 8616 11428 8628
rect 11287 8588 11428 8616
rect 11287 8585 11299 8588
rect 11241 8579 11299 8585
rect 11422 8576 11428 8588
rect 11480 8576 11486 8628
rect 12345 8619 12403 8625
rect 12345 8585 12357 8619
rect 12391 8616 12403 8619
rect 12434 8616 12440 8628
rect 12391 8588 12440 8616
rect 12391 8585 12403 8588
rect 12345 8579 12403 8585
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 13170 8576 13176 8628
rect 13228 8576 13234 8628
rect 13265 8619 13323 8625
rect 13265 8585 13277 8619
rect 13311 8616 13323 8619
rect 13630 8616 13636 8628
rect 13311 8588 13636 8616
rect 13311 8585 13323 8588
rect 13265 8579 13323 8585
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 13817 8619 13875 8625
rect 13817 8585 13829 8619
rect 13863 8616 13875 8619
rect 14182 8616 14188 8628
rect 13863 8588 14188 8616
rect 13863 8585 13875 8588
rect 13817 8579 13875 8585
rect 14182 8576 14188 8588
rect 14240 8576 14246 8628
rect 14369 8619 14427 8625
rect 14369 8585 14381 8619
rect 14415 8616 14427 8619
rect 15010 8616 15016 8628
rect 14415 8588 15016 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 15286 8576 15292 8628
rect 15344 8576 15350 8628
rect 15841 8619 15899 8625
rect 15841 8585 15853 8619
rect 15887 8616 15899 8619
rect 16114 8616 16120 8628
rect 15887 8588 16120 8616
rect 15887 8585 15899 8588
rect 15841 8579 15899 8585
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16393 8619 16451 8625
rect 16393 8585 16405 8619
rect 16439 8616 16451 8619
rect 16482 8616 16488 8628
rect 16439 8588 16488 8616
rect 16439 8585 16451 8588
rect 16393 8579 16451 8585
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 16758 8576 16764 8628
rect 16816 8576 16822 8628
rect 16945 8619 17003 8625
rect 16945 8585 16957 8619
rect 16991 8616 17003 8619
rect 17218 8616 17224 8628
rect 16991 8588 17224 8616
rect 16991 8585 17003 8588
rect 16945 8579 17003 8585
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 17313 8619 17371 8625
rect 17313 8585 17325 8619
rect 17359 8616 17371 8619
rect 17494 8616 17500 8628
rect 17359 8588 17500 8616
rect 17359 8585 17371 8588
rect 17313 8579 17371 8585
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 17862 8576 17868 8628
rect 17920 8576 17926 8628
rect 18233 8619 18291 8625
rect 18233 8585 18245 8619
rect 18279 8616 18291 8619
rect 18322 8616 18328 8628
rect 18279 8588 18328 8616
rect 18279 8585 18291 8588
rect 18233 8579 18291 8585
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 18414 8576 18420 8628
rect 18472 8576 18478 8628
rect 18598 8576 18604 8628
rect 18656 8576 18662 8628
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 18969 8619 19027 8625
rect 18969 8616 18981 8619
rect 18932 8588 18981 8616
rect 18932 8576 18938 8588
rect 18969 8585 18981 8588
rect 19015 8585 19027 8619
rect 18969 8579 19027 8585
rect 19518 8576 19524 8628
rect 19576 8576 19582 8628
rect 20073 8619 20131 8625
rect 20073 8585 20085 8619
rect 20119 8585 20131 8619
rect 20073 8579 20131 8585
rect 4525 8551 4583 8557
rect 4525 8517 4537 8551
rect 4571 8548 4583 8551
rect 4890 8548 4896 8560
rect 4571 8520 4896 8548
rect 4571 8517 4583 8520
rect 4525 8511 4583 8517
rect 4890 8508 4896 8520
rect 4948 8508 4954 8560
rect 6825 8551 6883 8557
rect 6825 8517 6837 8551
rect 6871 8548 6883 8551
rect 7193 8551 7251 8557
rect 7193 8548 7205 8551
rect 6871 8520 7205 8548
rect 6871 8517 6883 8520
rect 6825 8511 6883 8517
rect 7193 8517 7205 8520
rect 7239 8548 7251 8551
rect 8220 8548 8248 8576
rect 9508 8548 9536 8576
rect 7239 8520 8248 8548
rect 8680 8520 9536 8548
rect 7239 8517 7251 8520
rect 7193 8511 7251 8517
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 5810 8480 5816 8492
rect 5491 8452 5816 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 5951 8452 6914 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 6886 8412 6914 8452
rect 7466 8440 7472 8492
rect 7524 8440 7530 8492
rect 8018 8440 8024 8492
rect 8076 8440 8082 8492
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 8352 8452 8493 8480
rect 8352 8440 8358 8452
rect 8481 8449 8493 8452
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 7484 8412 7512 8440
rect 6886 8384 7512 8412
rect 6089 8347 6147 8353
rect 6089 8313 6101 8347
rect 6135 8344 6147 8347
rect 8478 8344 8484 8356
rect 6135 8316 8484 8344
rect 6135 8313 6147 8316
rect 6089 8307 6147 8313
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 8680 8353 8708 8520
rect 10410 8508 10416 8560
rect 10468 8508 10474 8560
rect 12066 8508 12072 8560
rect 12124 8508 12130 8560
rect 13188 8548 13216 8576
rect 12406 8520 13216 8548
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 9858 8480 9864 8492
rect 9539 8452 9864 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 9858 8440 9864 8452
rect 9916 8440 9922 8492
rect 9950 8440 9956 8492
rect 10008 8440 10014 8492
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8449 11023 8483
rect 10965 8443 11023 8449
rect 11609 8483 11667 8489
rect 11609 8449 11621 8483
rect 11655 8480 11667 8483
rect 12406 8480 12434 8520
rect 13446 8508 13452 8560
rect 13504 8508 13510 8560
rect 13541 8551 13599 8557
rect 13541 8517 13553 8551
rect 13587 8548 13599 8551
rect 16022 8548 16028 8560
rect 13587 8520 16028 8548
rect 13587 8517 13599 8520
rect 13541 8511 13599 8517
rect 16022 8508 16028 8520
rect 16080 8508 16086 8560
rect 16776 8548 16804 8576
rect 16132 8520 16804 8548
rect 17589 8551 17647 8557
rect 11655 8452 12434 8480
rect 12805 8483 12863 8489
rect 11655 8449 11667 8452
rect 11609 8443 11667 8449
rect 12805 8449 12817 8483
rect 12851 8480 12863 8483
rect 13081 8483 13139 8489
rect 13081 8480 13093 8483
rect 12851 8452 13093 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 13081 8449 13093 8452
rect 13127 8480 13139 8483
rect 13464 8480 13492 8508
rect 13127 8452 13492 8480
rect 14185 8483 14243 8489
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 14185 8449 14197 8483
rect 14231 8480 14243 8483
rect 14366 8480 14372 8492
rect 14231 8452 14372 8480
rect 14231 8449 14243 8452
rect 14185 8443 14243 8449
rect 10980 8412 11008 8443
rect 14366 8440 14372 8452
rect 14424 8440 14430 8492
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8480 14611 8483
rect 14918 8480 14924 8492
rect 14599 8452 14924 8480
rect 14599 8449 14611 8452
rect 14553 8443 14611 8449
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 16132 8489 16160 8520
rect 17589 8517 17601 8551
rect 17635 8548 17647 8551
rect 18138 8548 18144 8560
rect 17635 8520 18144 8548
rect 17635 8517 17647 8520
rect 17589 8511 17647 8517
rect 18138 8508 18144 8520
rect 18196 8508 18202 8560
rect 18432 8548 18460 8576
rect 18432 8520 18644 8548
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8480 15071 8483
rect 15657 8483 15715 8489
rect 15059 8452 15608 8480
rect 15059 8449 15071 8452
rect 15013 8443 15071 8449
rect 14826 8412 14832 8424
rect 10980 8384 14832 8412
rect 14826 8372 14832 8384
rect 14884 8372 14890 8424
rect 8665 8347 8723 8353
rect 8665 8313 8677 8347
rect 8711 8313 8723 8347
rect 8665 8307 8723 8313
rect 9217 8347 9275 8353
rect 9217 8313 9229 8347
rect 9263 8344 9275 8347
rect 9398 8344 9404 8356
rect 9263 8316 9404 8344
rect 9263 8313 9275 8316
rect 9217 8307 9275 8313
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 11793 8347 11851 8353
rect 11793 8313 11805 8347
rect 11839 8344 11851 8347
rect 12434 8344 12440 8356
rect 11839 8316 12440 8344
rect 11839 8313 11851 8316
rect 11793 8307 11851 8313
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 14642 8304 14648 8356
rect 14700 8344 14706 8356
rect 14737 8347 14795 8353
rect 14737 8344 14749 8347
rect 14700 8316 14749 8344
rect 14700 8304 14706 8316
rect 14737 8313 14749 8316
rect 14783 8313 14795 8347
rect 15580 8344 15608 8452
rect 15657 8449 15669 8483
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 15672 8412 15700 8443
rect 16758 8440 16764 8492
rect 16816 8440 16822 8492
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8480 17187 8483
rect 17494 8480 17500 8492
rect 17175 8452 17500 8480
rect 17175 8449 17187 8452
rect 17129 8443 17187 8449
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8480 18107 8483
rect 18322 8480 18328 8492
rect 18095 8452 18328 8480
rect 18095 8449 18107 8452
rect 18049 8443 18107 8449
rect 18322 8440 18328 8452
rect 18380 8440 18386 8492
rect 18417 8483 18475 8489
rect 18417 8449 18429 8483
rect 18463 8449 18475 8483
rect 18417 8443 18475 8449
rect 15672 8384 17356 8412
rect 17126 8344 17132 8356
rect 15580 8316 17132 8344
rect 14737 8307 14795 8313
rect 17126 8304 17132 8316
rect 17184 8304 17190 8356
rect 17328 8344 17356 8384
rect 17402 8372 17408 8424
rect 17460 8412 17466 8424
rect 18432 8412 18460 8443
rect 17460 8384 18460 8412
rect 18616 8412 18644 8520
rect 19334 8508 19340 8560
rect 19392 8548 19398 8560
rect 20088 8548 20116 8579
rect 20162 8576 20168 8628
rect 20220 8616 20226 8628
rect 21177 8619 21235 8625
rect 21177 8616 21189 8619
rect 20220 8588 21189 8616
rect 20220 8576 20226 8588
rect 21177 8585 21189 8588
rect 21223 8585 21235 8619
rect 21177 8579 21235 8585
rect 22281 8619 22339 8625
rect 22281 8585 22293 8619
rect 22327 8616 22339 8619
rect 22327 8588 22416 8616
rect 22327 8585 22339 8588
rect 22281 8579 22339 8585
rect 22094 8548 22100 8560
rect 19392 8520 20116 8548
rect 21008 8520 22100 8548
rect 19392 8508 19398 8520
rect 18690 8440 18696 8492
rect 18748 8480 18754 8492
rect 18785 8483 18843 8489
rect 18785 8480 18797 8483
rect 18748 8452 18797 8480
rect 18748 8440 18754 8452
rect 18785 8449 18797 8452
rect 18831 8449 18843 8483
rect 18785 8443 18843 8449
rect 18874 8440 18880 8492
rect 18932 8480 18938 8492
rect 19429 8483 19487 8489
rect 19429 8480 19441 8483
rect 18932 8452 19441 8480
rect 18932 8440 18938 8452
rect 19429 8449 19441 8452
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19576 8452 19993 8480
rect 19576 8440 19582 8452
rect 19981 8449 19993 8452
rect 20027 8449 20039 8483
rect 19981 8443 20039 8449
rect 20070 8440 20076 8492
rect 20128 8480 20134 8492
rect 20530 8480 20536 8492
rect 20128 8452 20536 8480
rect 20128 8440 20134 8452
rect 20530 8440 20536 8452
rect 20588 8440 20594 8492
rect 20806 8440 20812 8492
rect 20864 8440 20870 8492
rect 20622 8412 20628 8424
rect 18616 8384 20628 8412
rect 17460 8372 17466 8384
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 21008 8344 21036 8520
rect 22094 8508 22100 8520
rect 22152 8508 22158 8560
rect 21082 8440 21088 8492
rect 21140 8440 21146 8492
rect 21358 8440 21364 8492
rect 21416 8440 21422 8492
rect 21634 8440 21640 8492
rect 21692 8440 21698 8492
rect 22002 8440 22008 8492
rect 22060 8480 22066 8492
rect 22189 8483 22247 8489
rect 22189 8480 22201 8483
rect 22060 8452 22201 8480
rect 22060 8440 22066 8452
rect 22189 8449 22201 8452
rect 22235 8449 22247 8483
rect 22189 8443 22247 8449
rect 22388 8412 22416 8588
rect 22554 8576 22560 8628
rect 22612 8616 22618 8628
rect 22833 8619 22891 8625
rect 22833 8616 22845 8619
rect 22612 8588 22845 8616
rect 22612 8576 22618 8588
rect 22833 8585 22845 8588
rect 22879 8585 22891 8619
rect 22833 8579 22891 8585
rect 22922 8576 22928 8628
rect 22980 8576 22986 8628
rect 24762 8576 24768 8628
rect 24820 8616 24826 8628
rect 24820 8588 25176 8616
rect 24820 8576 24826 8588
rect 22646 8508 22652 8560
rect 22704 8548 22710 8560
rect 22940 8548 22968 8576
rect 22704 8520 22968 8548
rect 22704 8508 22710 8520
rect 24394 8508 24400 8560
rect 24452 8548 24458 8560
rect 24452 8520 24900 8548
rect 24452 8508 24458 8520
rect 22462 8440 22468 8492
rect 22520 8440 22526 8492
rect 22738 8440 22744 8492
rect 22796 8440 22802 8492
rect 23014 8440 23020 8492
rect 23072 8440 23078 8492
rect 23106 8440 23112 8492
rect 23164 8480 23170 8492
rect 23293 8483 23351 8489
rect 23293 8480 23305 8483
rect 23164 8452 23305 8480
rect 23164 8440 23170 8452
rect 23293 8449 23305 8452
rect 23339 8449 23351 8483
rect 23293 8443 23351 8449
rect 23566 8440 23572 8492
rect 23624 8440 23630 8492
rect 23842 8440 23848 8492
rect 23900 8440 23906 8492
rect 24118 8440 24124 8492
rect 24176 8440 24182 8492
rect 24302 8440 24308 8492
rect 24360 8480 24366 8492
rect 24872 8489 24900 8520
rect 25148 8489 25176 8588
rect 25498 8576 25504 8628
rect 25556 8616 25562 8628
rect 25556 8588 26004 8616
rect 25556 8576 25562 8588
rect 25222 8508 25228 8560
rect 25280 8548 25286 8560
rect 25280 8520 25728 8548
rect 25280 8508 25286 8520
rect 25700 8489 25728 8520
rect 25976 8489 26004 8588
rect 26326 8576 26332 8628
rect 26384 8616 26390 8628
rect 26384 8588 26832 8616
rect 26384 8576 26390 8588
rect 26142 8508 26148 8560
rect 26200 8548 26206 8560
rect 26200 8520 26556 8548
rect 26200 8508 26206 8520
rect 24581 8483 24639 8489
rect 24581 8480 24593 8483
rect 24360 8452 24593 8480
rect 24360 8440 24366 8452
rect 24581 8449 24593 8452
rect 24627 8449 24639 8483
rect 24581 8443 24639 8449
rect 24857 8483 24915 8489
rect 24857 8449 24869 8483
rect 24903 8449 24915 8483
rect 24857 8443 24915 8449
rect 25133 8483 25191 8489
rect 25133 8449 25145 8483
rect 25179 8449 25191 8483
rect 25133 8443 25191 8449
rect 25409 8483 25467 8489
rect 25409 8449 25421 8483
rect 25455 8449 25467 8483
rect 25409 8443 25467 8449
rect 25685 8483 25743 8489
rect 25685 8449 25697 8483
rect 25731 8449 25743 8483
rect 25685 8443 25743 8449
rect 25961 8483 26019 8489
rect 25961 8449 25973 8483
rect 26007 8449 26019 8483
rect 25961 8443 26019 8449
rect 17328 8316 21036 8344
rect 21100 8384 22416 8412
rect 21100 8288 21128 8384
rect 24946 8372 24952 8424
rect 25004 8412 25010 8424
rect 25424 8412 25452 8443
rect 26050 8440 26056 8492
rect 26108 8480 26114 8492
rect 26528 8489 26556 8520
rect 26804 8489 26832 8588
rect 27154 8576 27160 8628
rect 27212 8616 27218 8628
rect 27212 8588 27752 8616
rect 27212 8576 27218 8588
rect 27062 8508 27068 8560
rect 27120 8548 27126 8560
rect 27120 8520 27476 8548
rect 27120 8508 27126 8520
rect 26237 8483 26295 8489
rect 26237 8480 26249 8483
rect 26108 8452 26249 8480
rect 26108 8440 26114 8452
rect 26237 8449 26249 8452
rect 26283 8449 26295 8483
rect 26237 8443 26295 8449
rect 26513 8483 26571 8489
rect 26513 8449 26525 8483
rect 26559 8449 26571 8483
rect 26513 8443 26571 8449
rect 26789 8483 26847 8489
rect 26789 8449 26801 8483
rect 26835 8449 26847 8483
rect 26789 8443 26847 8449
rect 26878 8440 26884 8492
rect 26936 8480 26942 8492
rect 27448 8489 27476 8520
rect 27724 8489 27752 8588
rect 27982 8576 27988 8628
rect 28040 8616 28046 8628
rect 28040 8588 28212 8616
rect 28040 8576 28046 8588
rect 27798 8508 27804 8560
rect 27856 8548 27862 8560
rect 28184 8548 28212 8588
rect 28258 8576 28264 8628
rect 28316 8616 28322 8628
rect 28316 8588 28856 8616
rect 28316 8576 28322 8588
rect 27856 8520 28120 8548
rect 28184 8520 28396 8548
rect 27856 8508 27862 8520
rect 27157 8483 27215 8489
rect 27157 8480 27169 8483
rect 26936 8452 27169 8480
rect 26936 8440 26942 8452
rect 27157 8449 27169 8452
rect 27203 8449 27215 8483
rect 27157 8443 27215 8449
rect 27433 8483 27491 8489
rect 27433 8449 27445 8483
rect 27479 8449 27491 8483
rect 27433 8443 27491 8449
rect 27709 8483 27767 8489
rect 27709 8449 27721 8483
rect 27755 8449 27767 8483
rect 27709 8443 27767 8449
rect 27985 8483 28043 8489
rect 27985 8449 27997 8483
rect 28031 8449 28043 8483
rect 28092 8480 28120 8520
rect 28261 8483 28319 8489
rect 28261 8480 28273 8483
rect 28092 8452 28273 8480
rect 27985 8443 28043 8449
rect 28261 8449 28273 8452
rect 28307 8449 28319 8483
rect 28368 8480 28396 8520
rect 28828 8489 28856 8588
rect 29086 8576 29092 8628
rect 29144 8616 29150 8628
rect 29144 8588 29500 8616
rect 29144 8576 29150 8588
rect 28902 8508 28908 8560
rect 28960 8548 28966 8560
rect 28960 8520 29408 8548
rect 28960 8508 28966 8520
rect 29380 8489 29408 8520
rect 28537 8483 28595 8489
rect 28537 8480 28549 8483
rect 28368 8452 28549 8480
rect 28261 8443 28319 8449
rect 28537 8449 28549 8452
rect 28583 8449 28595 8483
rect 28537 8443 28595 8449
rect 28813 8483 28871 8489
rect 28813 8449 28825 8483
rect 28859 8449 28871 8483
rect 28813 8443 28871 8449
rect 29089 8483 29147 8489
rect 29089 8449 29101 8483
rect 29135 8449 29147 8483
rect 29089 8443 29147 8449
rect 29365 8483 29423 8489
rect 29365 8449 29377 8483
rect 29411 8449 29423 8483
rect 29472 8480 29500 8588
rect 30282 8576 30288 8628
rect 30340 8576 30346 8628
rect 30466 8576 30472 8628
rect 30524 8616 30530 8628
rect 30524 8588 30972 8616
rect 30524 8576 30530 8588
rect 29638 8508 29644 8560
rect 29696 8548 29702 8560
rect 29696 8520 30144 8548
rect 29696 8508 29702 8520
rect 30116 8489 30144 8520
rect 30190 8508 30196 8560
rect 30248 8548 30254 8560
rect 30248 8520 30696 8548
rect 30248 8508 30254 8520
rect 29733 8483 29791 8489
rect 29733 8480 29745 8483
rect 29472 8452 29745 8480
rect 29365 8443 29423 8449
rect 29733 8449 29745 8452
rect 29779 8449 29791 8483
rect 30009 8483 30067 8489
rect 30009 8480 30021 8483
rect 29733 8443 29791 8449
rect 29840 8452 30021 8480
rect 25004 8384 25452 8412
rect 25004 8372 25010 8384
rect 27522 8372 27528 8424
rect 27580 8412 27586 8424
rect 28000 8412 28028 8443
rect 29104 8412 29132 8443
rect 27580 8384 28028 8412
rect 28092 8384 28764 8412
rect 27580 8372 27586 8384
rect 21634 8304 21640 8356
rect 21692 8344 21698 8356
rect 22557 8347 22615 8353
rect 22557 8344 22569 8347
rect 21692 8316 22569 8344
rect 21692 8304 21698 8316
rect 22557 8313 22569 8316
rect 22603 8313 22615 8347
rect 22557 8307 22615 8313
rect 23290 8304 23296 8356
rect 23348 8344 23354 8356
rect 28092 8344 28120 8384
rect 23348 8316 28120 8344
rect 23348 8304 23354 8316
rect 7374 8236 7380 8288
rect 7432 8276 7438 8288
rect 15102 8276 15108 8288
rect 7432 8248 15108 8276
rect 7432 8236 7438 8248
rect 15102 8236 15108 8248
rect 15160 8236 15166 8288
rect 18506 8236 18512 8288
rect 18564 8276 18570 8288
rect 20346 8276 20352 8288
rect 18564 8248 20352 8276
rect 18564 8236 18570 8248
rect 20346 8236 20352 8248
rect 20404 8236 20410 8288
rect 20438 8236 20444 8288
rect 20496 8276 20502 8288
rect 20625 8279 20683 8285
rect 20625 8276 20637 8279
rect 20496 8248 20637 8276
rect 20496 8236 20502 8248
rect 20625 8245 20637 8248
rect 20671 8245 20683 8279
rect 20625 8239 20683 8245
rect 20898 8236 20904 8288
rect 20956 8236 20962 8288
rect 21082 8236 21088 8288
rect 21140 8236 21146 8288
rect 21450 8236 21456 8288
rect 21508 8236 21514 8288
rect 21726 8236 21732 8288
rect 21784 8276 21790 8288
rect 22005 8279 22063 8285
rect 22005 8276 22017 8279
rect 21784 8248 22017 8276
rect 21784 8236 21790 8248
rect 22005 8245 22017 8248
rect 22051 8245 22063 8279
rect 22005 8239 22063 8245
rect 22186 8236 22192 8288
rect 22244 8276 22250 8288
rect 23014 8276 23020 8288
rect 22244 8248 23020 8276
rect 22244 8236 22250 8248
rect 23014 8236 23020 8248
rect 23072 8236 23078 8288
rect 23106 8236 23112 8288
rect 23164 8236 23170 8288
rect 23382 8236 23388 8288
rect 23440 8236 23446 8288
rect 23658 8236 23664 8288
rect 23716 8236 23722 8288
rect 23934 8236 23940 8288
rect 23992 8236 23998 8288
rect 24394 8236 24400 8288
rect 24452 8236 24458 8288
rect 24486 8236 24492 8288
rect 24544 8276 24550 8288
rect 24673 8279 24731 8285
rect 24673 8276 24685 8279
rect 24544 8248 24685 8276
rect 24544 8236 24550 8248
rect 24673 8245 24685 8248
rect 24719 8245 24731 8279
rect 24673 8239 24731 8245
rect 24854 8236 24860 8288
rect 24912 8276 24918 8288
rect 24949 8279 25007 8285
rect 24949 8276 24961 8279
rect 24912 8248 24961 8276
rect 24912 8236 24918 8248
rect 24949 8245 24961 8248
rect 24995 8245 25007 8279
rect 24949 8239 25007 8245
rect 25038 8236 25044 8288
rect 25096 8276 25102 8288
rect 25225 8279 25283 8285
rect 25225 8276 25237 8279
rect 25096 8248 25237 8276
rect 25096 8236 25102 8248
rect 25225 8245 25237 8248
rect 25271 8245 25283 8279
rect 25225 8239 25283 8245
rect 25314 8236 25320 8288
rect 25372 8276 25378 8288
rect 25501 8279 25559 8285
rect 25501 8276 25513 8279
rect 25372 8248 25513 8276
rect 25372 8236 25378 8248
rect 25501 8245 25513 8248
rect 25547 8245 25559 8279
rect 25501 8239 25559 8245
rect 25774 8236 25780 8288
rect 25832 8236 25838 8288
rect 26050 8236 26056 8288
rect 26108 8236 26114 8288
rect 26326 8236 26332 8288
rect 26384 8236 26390 8288
rect 26602 8236 26608 8288
rect 26660 8236 26666 8288
rect 26970 8236 26976 8288
rect 27028 8236 27034 8288
rect 27246 8236 27252 8288
rect 27304 8236 27310 8288
rect 27522 8236 27528 8288
rect 27580 8236 27586 8288
rect 27801 8279 27859 8285
rect 27801 8245 27813 8279
rect 27847 8276 27859 8279
rect 27982 8276 27988 8288
rect 27847 8248 27988 8276
rect 27847 8245 27859 8248
rect 27801 8239 27859 8245
rect 27982 8236 27988 8248
rect 28040 8236 28046 8288
rect 28077 8279 28135 8285
rect 28077 8245 28089 8279
rect 28123 8276 28135 8279
rect 28166 8276 28172 8288
rect 28123 8248 28172 8276
rect 28123 8245 28135 8248
rect 28077 8239 28135 8245
rect 28166 8236 28172 8248
rect 28224 8236 28230 8288
rect 28350 8236 28356 8288
rect 28408 8236 28414 8288
rect 28442 8236 28448 8288
rect 28500 8276 28506 8288
rect 28629 8279 28687 8285
rect 28629 8276 28641 8279
rect 28500 8248 28641 8276
rect 28500 8236 28506 8248
rect 28629 8245 28641 8248
rect 28675 8245 28687 8279
rect 28736 8276 28764 8384
rect 28828 8384 29132 8412
rect 28828 8356 28856 8384
rect 29546 8372 29552 8424
rect 29604 8412 29610 8424
rect 29840 8412 29868 8452
rect 30009 8449 30021 8452
rect 30055 8449 30067 8483
rect 30009 8443 30067 8449
rect 30101 8483 30159 8489
rect 30101 8449 30113 8483
rect 30147 8449 30159 8483
rect 30101 8443 30159 8449
rect 30377 8483 30435 8489
rect 30377 8449 30389 8483
rect 30423 8449 30435 8483
rect 30377 8443 30435 8449
rect 29604 8384 29868 8412
rect 29604 8372 29610 8384
rect 29914 8372 29920 8424
rect 29972 8412 29978 8424
rect 30392 8412 30420 8443
rect 30558 8440 30564 8492
rect 30616 8440 30622 8492
rect 30668 8489 30696 8520
rect 30944 8489 30972 8588
rect 31110 8576 31116 8628
rect 31168 8576 31174 8628
rect 31386 8576 31392 8628
rect 31444 8576 31450 8628
rect 31662 8576 31668 8628
rect 31720 8576 31726 8628
rect 31846 8576 31852 8628
rect 31904 8616 31910 8628
rect 31904 8588 32444 8616
rect 31904 8576 31910 8588
rect 31018 8508 31024 8560
rect 31076 8548 31082 8560
rect 31076 8520 31524 8548
rect 31076 8508 31082 8520
rect 31496 8489 31524 8520
rect 31570 8508 31576 8560
rect 31628 8548 31634 8560
rect 31628 8520 32168 8548
rect 31628 8508 31634 8520
rect 30653 8483 30711 8489
rect 30653 8449 30665 8483
rect 30699 8449 30711 8483
rect 30653 8443 30711 8449
rect 30929 8483 30987 8489
rect 30929 8449 30941 8483
rect 30975 8449 30987 8483
rect 30929 8443 30987 8449
rect 31205 8483 31263 8489
rect 31205 8449 31217 8483
rect 31251 8449 31263 8483
rect 31205 8443 31263 8449
rect 31481 8483 31539 8489
rect 31481 8449 31493 8483
rect 31527 8449 31539 8483
rect 31481 8443 31539 8449
rect 31757 8483 31815 8489
rect 31757 8449 31769 8483
rect 31803 8449 31815 8483
rect 31757 8443 31815 8449
rect 29972 8384 30420 8412
rect 29972 8372 29978 8384
rect 28810 8304 28816 8356
rect 28868 8304 28874 8356
rect 28902 8304 28908 8356
rect 28960 8304 28966 8356
rect 30576 8353 30604 8440
rect 30742 8372 30748 8424
rect 30800 8412 30806 8424
rect 31220 8412 31248 8443
rect 30800 8384 31248 8412
rect 30800 8372 30806 8384
rect 31294 8372 31300 8424
rect 31352 8412 31358 8424
rect 31772 8412 31800 8443
rect 32030 8440 32036 8492
rect 32088 8440 32094 8492
rect 32140 8489 32168 8520
rect 32214 8508 32220 8560
rect 32272 8508 32278 8560
rect 32125 8483 32183 8489
rect 32125 8449 32137 8483
rect 32171 8449 32183 8483
rect 32125 8443 32183 8449
rect 31352 8384 31800 8412
rect 31352 8372 31358 8384
rect 29181 8347 29239 8353
rect 29181 8344 29193 8347
rect 29012 8316 29193 8344
rect 29012 8276 29040 8316
rect 29181 8313 29193 8316
rect 29227 8313 29239 8347
rect 29181 8307 29239 8313
rect 30561 8347 30619 8353
rect 30561 8313 30573 8347
rect 30607 8313 30619 8347
rect 30561 8307 30619 8313
rect 30834 8304 30840 8356
rect 30892 8304 30898 8356
rect 31938 8304 31944 8356
rect 31996 8304 32002 8356
rect 32048 8344 32076 8440
rect 32232 8344 32260 8508
rect 32416 8489 32444 8588
rect 32674 8576 32680 8628
rect 32732 8616 32738 8628
rect 32732 8588 33272 8616
rect 32732 8576 32738 8588
rect 32582 8508 32588 8560
rect 32640 8548 32646 8560
rect 32640 8520 32996 8548
rect 32640 8508 32646 8520
rect 32401 8483 32459 8489
rect 32401 8449 32413 8483
rect 32447 8449 32459 8483
rect 32401 8443 32459 8449
rect 32677 8483 32735 8489
rect 32677 8449 32689 8483
rect 32723 8449 32735 8483
rect 32677 8443 32735 8449
rect 32306 8372 32312 8424
rect 32364 8412 32370 8424
rect 32692 8412 32720 8443
rect 32766 8440 32772 8492
rect 32824 8440 32830 8492
rect 32968 8489 32996 8520
rect 33244 8489 33272 8588
rect 33686 8576 33692 8628
rect 33744 8576 33750 8628
rect 34054 8576 34060 8628
rect 34112 8616 34118 8628
rect 34333 8619 34391 8625
rect 34333 8616 34345 8619
rect 34112 8588 34345 8616
rect 34112 8576 34118 8588
rect 34333 8585 34345 8588
rect 34379 8585 34391 8619
rect 34333 8579 34391 8585
rect 34422 8576 34428 8628
rect 34480 8616 34486 8628
rect 34885 8619 34943 8625
rect 34885 8616 34897 8619
rect 34480 8588 34897 8616
rect 34480 8576 34486 8588
rect 34885 8585 34897 8588
rect 34931 8585 34943 8619
rect 34885 8579 34943 8585
rect 35158 8576 35164 8628
rect 35216 8616 35222 8628
rect 35989 8619 36047 8625
rect 35989 8616 36001 8619
rect 35216 8588 36001 8616
rect 35216 8576 35222 8588
rect 35989 8585 36001 8588
rect 36035 8585 36047 8619
rect 35989 8579 36047 8585
rect 36541 8619 36599 8625
rect 36541 8585 36553 8619
rect 36587 8585 36599 8619
rect 36541 8579 36599 8585
rect 33410 8508 33416 8560
rect 33468 8548 33474 8560
rect 33468 8520 33824 8548
rect 33468 8508 33474 8520
rect 32953 8483 33011 8489
rect 32953 8449 32965 8483
rect 32999 8449 33011 8483
rect 32953 8443 33011 8449
rect 33229 8483 33287 8489
rect 33229 8449 33241 8483
rect 33275 8449 33287 8483
rect 33229 8443 33287 8449
rect 33318 8440 33324 8492
rect 33376 8480 33382 8492
rect 33796 8489 33824 8520
rect 35434 8508 35440 8560
rect 35492 8548 35498 8560
rect 36556 8548 36584 8579
rect 36630 8576 36636 8628
rect 36688 8616 36694 8628
rect 36688 8588 37412 8616
rect 36688 8576 36694 8588
rect 37384 8557 37412 8588
rect 37458 8576 37464 8628
rect 37516 8576 37522 8628
rect 37550 8576 37556 8628
rect 37608 8616 37614 8628
rect 39117 8619 39175 8625
rect 39117 8616 39129 8619
rect 37608 8588 38516 8616
rect 37608 8576 37614 8588
rect 35492 8520 36584 8548
rect 37369 8551 37427 8557
rect 35492 8508 35498 8520
rect 37369 8517 37381 8551
rect 37415 8517 37427 8551
rect 37476 8548 37504 8576
rect 38488 8557 38516 8588
rect 38580 8588 39129 8616
rect 37921 8551 37979 8557
rect 37921 8548 37933 8551
rect 37476 8520 37933 8548
rect 37369 8511 37427 8517
rect 37921 8517 37933 8520
rect 37967 8517 37979 8551
rect 37921 8511 37979 8517
rect 38473 8551 38531 8557
rect 38473 8517 38485 8551
rect 38519 8517 38531 8551
rect 38473 8511 38531 8517
rect 33505 8483 33563 8489
rect 33505 8480 33517 8483
rect 33376 8452 33517 8480
rect 33376 8440 33382 8452
rect 33505 8449 33517 8452
rect 33551 8449 33563 8483
rect 33505 8443 33563 8449
rect 33781 8483 33839 8489
rect 33781 8449 33793 8483
rect 33827 8449 33839 8483
rect 33781 8443 33839 8449
rect 34146 8440 34152 8492
rect 34204 8440 34210 8492
rect 34793 8483 34851 8489
rect 34793 8449 34805 8483
rect 34839 8449 34851 8483
rect 34793 8443 34851 8449
rect 32364 8384 32720 8412
rect 32784 8412 32812 8440
rect 34808 8412 34836 8443
rect 35250 8440 35256 8492
rect 35308 8440 35314 8492
rect 35897 8483 35955 8489
rect 35897 8449 35909 8483
rect 35943 8449 35955 8483
rect 35897 8443 35955 8449
rect 32784 8384 33088 8412
rect 32364 8372 32370 8384
rect 32585 8347 32643 8353
rect 32585 8344 32597 8347
rect 32048 8316 32168 8344
rect 32232 8316 32597 8344
rect 28736 8248 29040 8276
rect 28629 8239 28687 8245
rect 29546 8236 29552 8288
rect 29604 8236 29610 8288
rect 29822 8236 29828 8288
rect 29880 8236 29886 8288
rect 32140 8276 32168 8316
rect 32585 8313 32597 8316
rect 32631 8313 32643 8347
rect 32585 8307 32643 8313
rect 32858 8304 32864 8356
rect 32916 8304 32922 8356
rect 32309 8279 32367 8285
rect 32309 8276 32321 8279
rect 32140 8248 32321 8276
rect 32309 8245 32321 8248
rect 32355 8245 32367 8279
rect 33060 8276 33088 8384
rect 33612 8384 34836 8412
rect 33226 8304 33232 8356
rect 33284 8344 33290 8356
rect 33612 8344 33640 8384
rect 34974 8372 34980 8424
rect 35032 8412 35038 8424
rect 35912 8412 35940 8443
rect 36446 8440 36452 8492
rect 36504 8440 36510 8492
rect 37642 8440 37648 8492
rect 37700 8480 37706 8492
rect 38580 8480 38608 8588
rect 39117 8585 39129 8588
rect 39163 8585 39175 8619
rect 39117 8579 39175 8585
rect 39298 8576 39304 8628
rect 39356 8616 39362 8628
rect 41141 8619 41199 8625
rect 41141 8616 41153 8619
rect 39356 8588 41153 8616
rect 39356 8576 39362 8588
rect 41141 8585 41153 8588
rect 41187 8585 41199 8619
rect 41141 8579 41199 8585
rect 38654 8508 38660 8560
rect 38712 8548 38718 8560
rect 38841 8551 38899 8557
rect 38841 8548 38853 8551
rect 38712 8520 38853 8548
rect 38712 8508 38718 8520
rect 38841 8517 38853 8520
rect 38887 8517 38899 8551
rect 38841 8511 38899 8517
rect 39206 8508 39212 8560
rect 39264 8548 39270 8560
rect 40865 8551 40923 8557
rect 40865 8548 40877 8551
rect 39264 8520 40877 8548
rect 39264 8508 39270 8520
rect 40865 8517 40877 8520
rect 40911 8517 40923 8551
rect 40865 8511 40923 8517
rect 37700 8452 38608 8480
rect 37700 8440 37706 8452
rect 39022 8440 39028 8492
rect 39080 8440 39086 8492
rect 39298 8440 39304 8492
rect 39356 8480 39362 8492
rect 39945 8483 40003 8489
rect 39945 8480 39957 8483
rect 39356 8452 39957 8480
rect 39356 8440 39362 8452
rect 39945 8449 39957 8452
rect 39991 8449 40003 8483
rect 39945 8443 40003 8449
rect 40494 8440 40500 8492
rect 40552 8440 40558 8492
rect 41046 8440 41052 8492
rect 41104 8440 41110 8492
rect 35032 8384 35940 8412
rect 35032 8372 35038 8384
rect 36538 8372 36544 8424
rect 36596 8412 36602 8424
rect 36596 8384 38148 8412
rect 36596 8372 36602 8384
rect 33284 8316 33640 8344
rect 33284 8304 33290 8316
rect 33686 8304 33692 8356
rect 33744 8304 33750 8356
rect 33962 8304 33968 8356
rect 34020 8304 34026 8356
rect 34606 8304 34612 8356
rect 34664 8344 34670 8356
rect 35437 8347 35495 8353
rect 35437 8344 35449 8347
rect 34664 8316 35449 8344
rect 34664 8304 34670 8316
rect 35437 8313 35449 8316
rect 35483 8313 35495 8347
rect 35437 8307 35495 8313
rect 35710 8304 35716 8356
rect 35768 8344 35774 8356
rect 38120 8353 38148 8384
rect 37553 8347 37611 8353
rect 37553 8344 37565 8347
rect 35768 8316 37565 8344
rect 35768 8304 35774 8316
rect 37553 8313 37565 8316
rect 37599 8313 37611 8347
rect 37553 8307 37611 8313
rect 38105 8347 38163 8353
rect 38105 8313 38117 8347
rect 38151 8313 38163 8347
rect 40129 8347 40187 8353
rect 40129 8344 40141 8347
rect 38105 8307 38163 8313
rect 38212 8316 40141 8344
rect 33137 8279 33195 8285
rect 33137 8276 33149 8279
rect 33060 8248 33149 8276
rect 32309 8239 32367 8245
rect 33137 8245 33149 8248
rect 33183 8245 33195 8279
rect 33137 8239 33195 8245
rect 33413 8279 33471 8285
rect 33413 8245 33425 8279
rect 33459 8276 33471 8279
rect 33704 8276 33732 8304
rect 33459 8248 33732 8276
rect 33459 8245 33471 8248
rect 33413 8239 33471 8245
rect 38010 8236 38016 8288
rect 38068 8276 38074 8288
rect 38212 8276 38240 8316
rect 40129 8313 40141 8316
rect 40175 8313 40187 8347
rect 40129 8307 40187 8313
rect 38068 8248 38240 8276
rect 38068 8236 38074 8248
rect 1104 8186 43884 8208
rect 1104 8134 6297 8186
rect 6349 8134 6361 8186
rect 6413 8134 6425 8186
rect 6477 8134 6489 8186
rect 6541 8134 6553 8186
rect 6605 8134 16991 8186
rect 17043 8134 17055 8186
rect 17107 8134 17119 8186
rect 17171 8134 17183 8186
rect 17235 8134 17247 8186
rect 17299 8134 27685 8186
rect 27737 8134 27749 8186
rect 27801 8134 27813 8186
rect 27865 8134 27877 8186
rect 27929 8134 27941 8186
rect 27993 8134 38379 8186
rect 38431 8134 38443 8186
rect 38495 8134 38507 8186
rect 38559 8134 38571 8186
rect 38623 8134 38635 8186
rect 38687 8134 43884 8186
rect 1104 8112 43884 8134
rect 5718 8032 5724 8084
rect 5776 8032 5782 8084
rect 6178 8032 6184 8084
rect 6236 8072 6242 8084
rect 6273 8075 6331 8081
rect 6273 8072 6285 8075
rect 6236 8044 6285 8072
rect 6236 8032 6242 8044
rect 6273 8041 6285 8044
rect 6319 8041 6331 8075
rect 6273 8035 6331 8041
rect 7558 8032 7564 8084
rect 7616 8032 7622 8084
rect 7926 8032 7932 8084
rect 7984 8032 7990 8084
rect 8478 8032 8484 8084
rect 8536 8032 8542 8084
rect 9306 8032 9312 8084
rect 9364 8032 9370 8084
rect 10134 8032 10140 8084
rect 10192 8032 10198 8084
rect 11238 8032 11244 8084
rect 11296 8032 11302 8084
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 11793 8075 11851 8081
rect 11793 8072 11805 8075
rect 11572 8044 11805 8072
rect 11572 8032 11578 8044
rect 11793 8041 11805 8044
rect 11839 8041 11851 8075
rect 13265 8075 13323 8081
rect 11793 8035 11851 8041
rect 12360 8044 13216 8072
rect 6914 7964 6920 8016
rect 6972 7964 6978 8016
rect 12360 8004 12388 8044
rect 11164 7976 12388 8004
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7868 6239 7871
rect 7377 7871 7435 7877
rect 6227 7840 6914 7868
rect 6227 7837 6239 7840
rect 6181 7831 6239 7837
rect 5629 7803 5687 7809
rect 5629 7769 5641 7803
rect 5675 7769 5687 7803
rect 5629 7763 5687 7769
rect 5644 7732 5672 7763
rect 6730 7760 6736 7812
rect 6788 7760 6794 7812
rect 6886 7800 6914 7840
rect 7377 7837 7389 7871
rect 7423 7868 7435 7871
rect 8202 7868 8208 7880
rect 7423 7840 8208 7868
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 11164 7877 11192 7976
rect 12434 7964 12440 8016
rect 12492 7964 12498 8016
rect 13188 8004 13216 8044
rect 13265 8041 13277 8075
rect 13311 8072 13323 8075
rect 13354 8072 13360 8084
rect 13311 8044 13360 8072
rect 13311 8041 13323 8044
rect 13265 8035 13323 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 13817 8075 13875 8081
rect 13817 8041 13829 8075
rect 13863 8072 13875 8075
rect 13906 8072 13912 8084
rect 13863 8044 13912 8072
rect 13863 8041 13875 8044
rect 13817 8035 13875 8041
rect 13906 8032 13912 8044
rect 13964 8032 13970 8084
rect 14550 8032 14556 8084
rect 14608 8032 14614 8084
rect 14734 8032 14740 8084
rect 14792 8072 14798 8084
rect 15105 8075 15163 8081
rect 15105 8072 15117 8075
rect 14792 8044 15117 8072
rect 14792 8032 14798 8044
rect 15105 8041 15117 8044
rect 15151 8041 15163 8075
rect 15105 8035 15163 8041
rect 15654 8032 15660 8084
rect 15712 8032 15718 8084
rect 15764 8044 16804 8072
rect 15764 8004 15792 8044
rect 13188 7976 15792 8004
rect 16574 7964 16580 8016
rect 16632 7964 16638 8016
rect 16776 8004 16804 8044
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 17037 8075 17095 8081
rect 17037 8072 17049 8075
rect 16908 8044 17049 8072
rect 16908 8032 16914 8044
rect 17037 8041 17049 8044
rect 17083 8041 17095 8075
rect 17037 8035 17095 8041
rect 17402 8032 17408 8084
rect 17460 8032 17466 8084
rect 18782 8072 18788 8084
rect 17512 8044 18788 8072
rect 17512 8004 17540 8044
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 18874 8032 18880 8084
rect 18932 8032 18938 8084
rect 19978 8032 19984 8084
rect 20036 8072 20042 8084
rect 20165 8075 20223 8081
rect 20165 8072 20177 8075
rect 20036 8044 20177 8072
rect 20036 8032 20042 8044
rect 20165 8041 20177 8044
rect 20211 8041 20223 8075
rect 20165 8035 20223 8041
rect 20441 8075 20499 8081
rect 20441 8041 20453 8075
rect 20487 8072 20499 8075
rect 20990 8072 20996 8084
rect 20487 8044 20996 8072
rect 20487 8041 20499 8044
rect 20441 8035 20499 8041
rect 20990 8032 20996 8044
rect 21048 8032 21054 8084
rect 21358 8032 21364 8084
rect 21416 8032 21422 8084
rect 21450 8032 21456 8084
rect 21508 8032 21514 8084
rect 22925 8075 22983 8081
rect 22925 8072 22937 8075
rect 22480 8044 22937 8072
rect 16776 7976 17540 8004
rect 17954 7964 17960 8016
rect 18012 7964 18018 8016
rect 18322 7964 18328 8016
rect 18380 7964 18386 8016
rect 19429 8007 19487 8013
rect 19429 7973 19441 8007
rect 19475 8004 19487 8007
rect 19475 7976 19564 8004
rect 19475 7973 19487 7976
rect 19429 7967 19487 7973
rect 11716 7908 16896 7936
rect 11149 7871 11207 7877
rect 8312 7840 11100 7868
rect 7742 7800 7748 7812
rect 6886 7772 7748 7800
rect 7742 7760 7748 7772
rect 7800 7760 7806 7812
rect 7837 7803 7895 7809
rect 7837 7769 7849 7803
rect 7883 7800 7895 7803
rect 8312 7800 8340 7840
rect 7883 7772 8340 7800
rect 7883 7769 7895 7772
rect 7837 7763 7895 7769
rect 8386 7760 8392 7812
rect 8444 7760 8450 7812
rect 9214 7760 9220 7812
rect 9272 7760 9278 7812
rect 10042 7760 10048 7812
rect 10100 7760 10106 7812
rect 9582 7732 9588 7744
rect 5644 7704 9588 7732
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 11072 7732 11100 7840
rect 11149 7837 11161 7871
rect 11195 7837 11207 7871
rect 11149 7831 11207 7837
rect 11716 7809 11744 7908
rect 12986 7828 12992 7880
rect 13044 7828 13050 7880
rect 14918 7828 14924 7880
rect 14976 7828 14982 7880
rect 16666 7868 16672 7880
rect 15488 7840 16672 7868
rect 11701 7803 11759 7809
rect 11701 7769 11713 7803
rect 11747 7769 11759 7803
rect 11701 7763 11759 7769
rect 12250 7760 12256 7812
rect 12308 7760 12314 7812
rect 13541 7803 13599 7809
rect 13541 7769 13553 7803
rect 13587 7800 13599 7803
rect 14461 7803 14519 7809
rect 13587 7772 14412 7800
rect 13587 7769 13599 7772
rect 13541 7763 13599 7769
rect 13722 7732 13728 7744
rect 11072 7704 13728 7732
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 14384 7732 14412 7772
rect 14461 7769 14473 7803
rect 14507 7800 14519 7803
rect 15488 7800 15516 7840
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 14507 7772 15516 7800
rect 15565 7803 15623 7809
rect 14507 7769 14519 7772
rect 14461 7763 14519 7769
rect 15565 7769 15577 7803
rect 15611 7769 15623 7803
rect 15565 7763 15623 7769
rect 15470 7732 15476 7744
rect 14384 7704 15476 7732
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 15580 7732 15608 7763
rect 16390 7760 16396 7812
rect 16448 7760 16454 7812
rect 16868 7800 16896 7908
rect 16960 7908 19334 7936
rect 16960 7877 16988 7908
rect 19306 7884 19334 7908
rect 19536 7884 19564 7976
rect 19610 7964 19616 8016
rect 19668 7964 19674 8016
rect 20809 8007 20867 8013
rect 20809 8004 20821 8007
rect 19720 7976 20821 8004
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7837 17003 7871
rect 16945 7831 17003 7837
rect 17586 7828 17592 7880
rect 17644 7828 17650 7880
rect 17954 7868 17960 7880
rect 17696 7840 17960 7868
rect 17696 7800 17724 7840
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 18506 7828 18512 7880
rect 18564 7828 18570 7880
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7868 18843 7871
rect 18966 7868 18972 7880
rect 18831 7840 18972 7868
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 18966 7828 18972 7840
rect 19024 7828 19030 7880
rect 19058 7828 19064 7880
rect 19116 7828 19122 7880
rect 19306 7856 19564 7884
rect 19628 7877 19656 7964
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 16868 7772 17724 7800
rect 17770 7760 17776 7812
rect 17828 7760 17834 7812
rect 19720 7800 19748 7976
rect 20809 7973 20821 7976
rect 20855 7973 20867 8007
rect 20809 7967 20867 7973
rect 21468 7936 21496 8032
rect 21818 7964 21824 8016
rect 21876 8004 21882 8016
rect 22480 8004 22508 8044
rect 22925 8041 22937 8044
rect 22971 8041 22983 8075
rect 22925 8035 22983 8041
rect 23014 8032 23020 8084
rect 23072 8072 23078 8084
rect 23201 8075 23259 8081
rect 23201 8072 23213 8075
rect 23072 8044 23213 8072
rect 23072 8032 23078 8044
rect 23201 8041 23213 8044
rect 23247 8041 23259 8075
rect 23201 8035 23259 8041
rect 23658 8032 23664 8084
rect 23716 8032 23722 8084
rect 24394 8032 24400 8084
rect 24452 8032 24458 8084
rect 24581 8075 24639 8081
rect 24581 8041 24593 8075
rect 24627 8072 24639 8075
rect 24670 8072 24676 8084
rect 24627 8044 24676 8072
rect 24627 8041 24639 8044
rect 24581 8035 24639 8041
rect 24670 8032 24676 8044
rect 24728 8032 24734 8084
rect 25406 8032 25412 8084
rect 25464 8032 25470 8084
rect 25498 8032 25504 8084
rect 25556 8072 25562 8084
rect 25685 8075 25743 8081
rect 25685 8072 25697 8075
rect 25556 8044 25697 8072
rect 25556 8032 25562 8044
rect 25685 8041 25697 8044
rect 25731 8041 25743 8075
rect 25685 8035 25743 8041
rect 25866 8032 25872 8084
rect 25924 8072 25930 8084
rect 26513 8075 26571 8081
rect 26513 8072 26525 8075
rect 25924 8044 26525 8072
rect 25924 8032 25930 8044
rect 26513 8041 26525 8044
rect 26559 8041 26571 8075
rect 26513 8035 26571 8041
rect 27154 8032 27160 8084
rect 27212 8072 27218 8084
rect 27617 8075 27675 8081
rect 27617 8072 27629 8075
rect 27212 8044 27629 8072
rect 27212 8032 27218 8044
rect 27617 8041 27629 8044
rect 27663 8041 27675 8075
rect 27617 8035 27675 8041
rect 27706 8032 27712 8084
rect 27764 8072 27770 8084
rect 27893 8075 27951 8081
rect 27893 8072 27905 8075
rect 27764 8044 27905 8072
rect 27764 8032 27770 8044
rect 27893 8041 27905 8044
rect 27939 8041 27951 8075
rect 27893 8035 27951 8041
rect 28169 8075 28227 8081
rect 28169 8041 28181 8075
rect 28215 8072 28227 8075
rect 28258 8072 28264 8084
rect 28215 8044 28264 8072
rect 28215 8041 28227 8044
rect 28169 8035 28227 8041
rect 28258 8032 28264 8044
rect 28316 8032 28322 8084
rect 28442 8032 28448 8084
rect 28500 8032 28506 8084
rect 34882 8032 34888 8084
rect 34940 8072 34946 8084
rect 35621 8075 35679 8081
rect 35621 8072 35633 8075
rect 34940 8044 35633 8072
rect 34940 8032 34946 8044
rect 35621 8041 35633 8044
rect 35667 8041 35679 8075
rect 35621 8035 35679 8041
rect 35986 8032 35992 8084
rect 36044 8072 36050 8084
rect 36265 8075 36323 8081
rect 36265 8072 36277 8075
rect 36044 8044 36277 8072
rect 36044 8032 36050 8044
rect 36265 8041 36277 8044
rect 36311 8041 36323 8075
rect 36265 8035 36323 8041
rect 36354 8032 36360 8084
rect 36412 8072 36418 8084
rect 36817 8075 36875 8081
rect 36817 8072 36829 8075
rect 36412 8044 36829 8072
rect 36412 8032 36418 8044
rect 36817 8041 36829 8044
rect 36863 8041 36875 8075
rect 36817 8035 36875 8041
rect 37366 8032 37372 8084
rect 37424 8072 37430 8084
rect 37645 8075 37703 8081
rect 37645 8072 37657 8075
rect 37424 8044 37657 8072
rect 37424 8032 37430 8044
rect 37645 8041 37657 8044
rect 37691 8041 37703 8075
rect 37645 8035 37703 8041
rect 38197 8075 38255 8081
rect 38197 8041 38209 8075
rect 38243 8041 38255 8075
rect 38197 8035 38255 8041
rect 21876 7976 22508 8004
rect 21876 7964 21882 7976
rect 22554 7964 22560 8016
rect 22612 7964 22618 8016
rect 22646 7964 22652 8016
rect 22704 7964 22710 8016
rect 23676 8004 23704 8032
rect 22756 7976 23704 8004
rect 22572 7936 22600 7964
rect 20548 7908 21496 7936
rect 21928 7908 22600 7936
rect 19886 7828 19892 7880
rect 19944 7828 19950 7880
rect 19981 7871 20039 7877
rect 19981 7837 19993 7871
rect 20027 7837 20039 7871
rect 19981 7831 20039 7837
rect 20257 7847 20315 7853
rect 19996 7800 20024 7831
rect 20257 7813 20269 7847
rect 20303 7844 20315 7847
rect 20438 7844 20444 7880
rect 20303 7828 20444 7844
rect 20496 7828 20502 7880
rect 20548 7877 20576 7908
rect 20533 7871 20591 7877
rect 20533 7837 20545 7871
rect 20579 7837 20591 7871
rect 20533 7831 20591 7837
rect 20990 7828 20996 7880
rect 21048 7828 21054 7880
rect 21082 7828 21088 7880
rect 21140 7828 21146 7880
rect 21542 7828 21548 7880
rect 21600 7828 21606 7880
rect 21634 7828 21640 7880
rect 21692 7828 21698 7880
rect 21928 7877 21956 7908
rect 21913 7871 21971 7877
rect 21913 7837 21925 7871
rect 21959 7837 21971 7871
rect 21913 7831 21971 7837
rect 22189 7871 22247 7877
rect 22189 7837 22201 7871
rect 22235 7837 22247 7871
rect 22189 7831 22247 7837
rect 22465 7871 22523 7877
rect 22465 7837 22477 7871
rect 22511 7868 22523 7871
rect 22646 7868 22652 7880
rect 22511 7840 22652 7868
rect 22511 7837 22523 7840
rect 22465 7831 22523 7837
rect 20303 7816 20484 7828
rect 20303 7813 20315 7816
rect 20257 7807 20315 7813
rect 18524 7772 19748 7800
rect 19912 7772 20024 7800
rect 18524 7732 18552 7772
rect 15580 7704 18552 7732
rect 18601 7735 18659 7741
rect 18601 7701 18613 7735
rect 18647 7732 18659 7735
rect 19518 7732 19524 7744
rect 18647 7704 19524 7732
rect 18647 7701 18659 7704
rect 18601 7695 18659 7701
rect 19518 7692 19524 7704
rect 19576 7692 19582 7744
rect 19705 7735 19763 7741
rect 19705 7701 19717 7735
rect 19751 7732 19763 7735
rect 19912 7732 19940 7772
rect 20622 7760 20628 7812
rect 20680 7800 20686 7812
rect 22204 7800 22232 7831
rect 22646 7828 22652 7840
rect 22704 7828 22710 7880
rect 22756 7877 22784 7976
rect 24026 7964 24032 8016
rect 24084 7964 24090 8016
rect 24412 7936 24440 8032
rect 28460 8004 28488 8032
rect 23032 7908 23244 7936
rect 23032 7877 23060 7908
rect 22741 7871 22799 7877
rect 22741 7837 22753 7871
rect 22787 7837 22799 7871
rect 22741 7831 22799 7837
rect 23017 7871 23075 7877
rect 23017 7837 23029 7871
rect 23063 7837 23075 7871
rect 23017 7831 23075 7837
rect 23106 7828 23112 7880
rect 23164 7828 23170 7880
rect 23124 7800 23152 7828
rect 20680 7772 20852 7800
rect 22204 7772 23152 7800
rect 23216 7800 23244 7908
rect 23584 7908 24440 7936
rect 25516 7976 28488 8004
rect 23290 7877 23296 7880
rect 23285 7831 23296 7877
rect 23348 7868 23354 7880
rect 23584 7877 23612 7908
rect 23569 7871 23627 7877
rect 23348 7840 23385 7868
rect 23290 7828 23296 7831
rect 23348 7828 23354 7840
rect 23569 7837 23581 7871
rect 23615 7837 23627 7871
rect 23569 7831 23627 7837
rect 23845 7871 23903 7877
rect 23845 7837 23857 7871
rect 23891 7868 23903 7871
rect 24302 7868 24308 7880
rect 23891 7840 24308 7868
rect 23891 7837 23903 7840
rect 23845 7831 23903 7837
rect 24302 7828 24308 7840
rect 24360 7828 24366 7880
rect 24397 7871 24455 7877
rect 24397 7837 24409 7871
rect 24443 7868 24455 7871
rect 24486 7868 24492 7880
rect 24443 7840 24492 7868
rect 24443 7837 24455 7840
rect 24397 7831 24455 7837
rect 24486 7828 24492 7840
rect 24544 7828 24550 7880
rect 24673 7871 24731 7877
rect 24673 7837 24685 7871
rect 24719 7868 24731 7871
rect 24854 7868 24860 7880
rect 24719 7840 24860 7868
rect 24719 7837 24731 7840
rect 24673 7831 24731 7837
rect 24854 7828 24860 7840
rect 24912 7828 24918 7880
rect 24949 7871 25007 7877
rect 24949 7837 24961 7871
rect 24995 7868 25007 7871
rect 25038 7868 25044 7880
rect 24995 7840 25044 7868
rect 24995 7837 25007 7840
rect 24949 7831 25007 7837
rect 25038 7828 25044 7840
rect 25096 7828 25102 7880
rect 25225 7871 25283 7877
rect 25225 7837 25237 7871
rect 25271 7868 25283 7871
rect 25314 7868 25320 7880
rect 25271 7840 25320 7868
rect 25271 7837 25283 7840
rect 25225 7831 25283 7837
rect 25314 7828 25320 7840
rect 25372 7828 25378 7880
rect 25516 7877 25544 7976
rect 37274 7964 37280 8016
rect 37332 8004 37338 8016
rect 38212 8004 38240 8035
rect 38746 8032 38752 8084
rect 38804 8032 38810 8084
rect 38838 8032 38844 8084
rect 38896 8072 38902 8084
rect 39301 8075 39359 8081
rect 39301 8072 39313 8075
rect 38896 8044 39313 8072
rect 38896 8032 38902 8044
rect 39301 8041 39313 8044
rect 39347 8041 39359 8075
rect 39301 8035 39359 8041
rect 40034 8032 40040 8084
rect 40092 8072 40098 8084
rect 40589 8075 40647 8081
rect 40589 8072 40601 8075
rect 40092 8044 40601 8072
rect 40092 8032 40098 8044
rect 40589 8041 40601 8044
rect 40635 8041 40647 8075
rect 40589 8035 40647 8041
rect 37332 7976 38240 8004
rect 37332 7964 37338 7976
rect 25590 7896 25596 7948
rect 25648 7936 25654 7948
rect 28166 7936 28172 7948
rect 25648 7908 27108 7936
rect 25648 7896 25654 7908
rect 25501 7871 25559 7877
rect 25501 7837 25513 7871
rect 25547 7837 25559 7871
rect 25501 7831 25559 7837
rect 25774 7828 25780 7880
rect 25832 7828 25838 7880
rect 26050 7828 26056 7880
rect 26108 7828 26114 7880
rect 26326 7828 26332 7880
rect 26384 7828 26390 7880
rect 26602 7828 26608 7880
rect 26660 7828 26666 7880
rect 26881 7871 26939 7877
rect 26881 7837 26893 7871
rect 26927 7868 26939 7871
rect 26970 7868 26976 7880
rect 26927 7840 26976 7868
rect 26927 7837 26939 7840
rect 26881 7831 26939 7837
rect 26970 7828 26976 7840
rect 27028 7828 27034 7880
rect 23216 7772 24072 7800
rect 20680 7760 20686 7772
rect 19751 7704 19940 7732
rect 19751 7701 19763 7704
rect 19705 7695 19763 7701
rect 20530 7692 20536 7744
rect 20588 7732 20594 7744
rect 20717 7735 20775 7741
rect 20717 7732 20729 7735
rect 20588 7704 20729 7732
rect 20588 7692 20594 7704
rect 20717 7701 20729 7704
rect 20763 7701 20775 7735
rect 20824 7732 20852 7772
rect 21082 7732 21088 7744
rect 20824 7704 21088 7732
rect 20717 7695 20775 7701
rect 21082 7692 21088 7704
rect 21140 7692 21146 7744
rect 21266 7692 21272 7744
rect 21324 7692 21330 7744
rect 21358 7692 21364 7744
rect 21416 7732 21422 7744
rect 21821 7735 21879 7741
rect 21821 7732 21833 7735
rect 21416 7704 21833 7732
rect 21416 7692 21422 7704
rect 21821 7701 21833 7704
rect 21867 7701 21879 7735
rect 21821 7695 21879 7701
rect 22094 7692 22100 7744
rect 22152 7692 22158 7744
rect 22373 7735 22431 7741
rect 22373 7701 22385 7735
rect 22419 7732 22431 7735
rect 22830 7732 22836 7744
rect 22419 7704 22836 7732
rect 22419 7701 22431 7704
rect 22373 7695 22431 7701
rect 22830 7692 22836 7704
rect 22888 7692 22894 7744
rect 23290 7692 23296 7744
rect 23348 7732 23354 7744
rect 23477 7735 23535 7741
rect 23477 7732 23489 7735
rect 23348 7704 23489 7732
rect 23348 7692 23354 7704
rect 23477 7701 23489 7704
rect 23523 7701 23535 7735
rect 23477 7695 23535 7701
rect 23750 7692 23756 7744
rect 23808 7692 23814 7744
rect 24044 7732 24072 7772
rect 26142 7760 26148 7812
rect 26200 7800 26206 7812
rect 26200 7772 26832 7800
rect 26200 7760 26206 7772
rect 24486 7732 24492 7744
rect 24044 7704 24492 7732
rect 24486 7692 24492 7704
rect 24544 7692 24550 7744
rect 24854 7692 24860 7744
rect 24912 7692 24918 7744
rect 25130 7692 25136 7744
rect 25188 7692 25194 7744
rect 25958 7692 25964 7744
rect 26016 7692 26022 7744
rect 26234 7692 26240 7744
rect 26292 7692 26298 7744
rect 26804 7741 26832 7772
rect 27080 7741 27108 7908
rect 28000 7908 28172 7936
rect 27157 7871 27215 7877
rect 27157 7837 27169 7871
rect 27203 7868 27215 7871
rect 27246 7868 27252 7880
rect 27203 7840 27252 7868
rect 27203 7837 27215 7840
rect 27157 7831 27215 7837
rect 27246 7828 27252 7840
rect 27304 7828 27310 7880
rect 27338 7828 27344 7880
rect 27396 7828 27402 7880
rect 27433 7871 27491 7877
rect 27433 7837 27445 7871
rect 27479 7868 27491 7871
rect 27522 7868 27528 7880
rect 27479 7840 27528 7868
rect 27479 7837 27491 7840
rect 27433 7831 27491 7837
rect 27522 7828 27528 7840
rect 27580 7828 27586 7880
rect 28000 7877 28028 7908
rect 28166 7896 28172 7908
rect 28224 7896 28230 7948
rect 34606 7896 34612 7948
rect 34664 7936 34670 7948
rect 34664 7908 35894 7936
rect 34664 7896 34670 7908
rect 27709 7871 27767 7877
rect 27709 7837 27721 7871
rect 27755 7837 27767 7871
rect 27709 7831 27767 7837
rect 27985 7871 28043 7877
rect 27985 7837 27997 7871
rect 28031 7837 28043 7871
rect 27985 7831 28043 7837
rect 27356 7741 27384 7828
rect 27724 7800 27752 7831
rect 28074 7828 28080 7880
rect 28132 7828 28138 7880
rect 28258 7828 28264 7880
rect 28316 7868 28322 7880
rect 28902 7868 28908 7880
rect 28316 7840 28908 7868
rect 28316 7828 28322 7840
rect 28902 7828 28908 7840
rect 28960 7828 28966 7880
rect 33594 7828 33600 7880
rect 33652 7828 33658 7880
rect 33870 7828 33876 7880
rect 33928 7828 33934 7880
rect 35434 7828 35440 7880
rect 35492 7828 35498 7880
rect 35866 7868 35894 7908
rect 36262 7896 36268 7948
rect 36320 7936 36326 7948
rect 36320 7908 38148 7936
rect 36320 7896 36326 7908
rect 35866 7840 36768 7868
rect 28092 7800 28120 7828
rect 27724 7772 28120 7800
rect 34514 7760 34520 7812
rect 34572 7800 34578 7812
rect 34572 7772 35894 7800
rect 34572 7760 34578 7772
rect 26789 7735 26847 7741
rect 26789 7701 26801 7735
rect 26835 7701 26847 7735
rect 26789 7695 26847 7701
rect 27065 7735 27123 7741
rect 27065 7701 27077 7735
rect 27111 7701 27123 7735
rect 27065 7695 27123 7701
rect 27341 7735 27399 7741
rect 27341 7701 27353 7735
rect 27387 7701 27399 7735
rect 27341 7695 27399 7701
rect 33778 7692 33784 7744
rect 33836 7692 33842 7744
rect 34054 7692 34060 7744
rect 34112 7692 34118 7744
rect 35866 7732 35894 7772
rect 35986 7760 35992 7812
rect 36044 7800 36050 7812
rect 36740 7809 36768 7840
rect 38120 7809 38148 7908
rect 38194 7828 38200 7880
rect 38252 7868 38258 7880
rect 38252 7840 39252 7868
rect 38252 7828 38258 7840
rect 36173 7803 36231 7809
rect 36173 7800 36185 7803
rect 36044 7772 36185 7800
rect 36044 7760 36050 7772
rect 36173 7769 36185 7772
rect 36219 7769 36231 7803
rect 36173 7763 36231 7769
rect 36725 7803 36783 7809
rect 36725 7769 36737 7803
rect 36771 7769 36783 7803
rect 37553 7803 37611 7809
rect 37553 7800 37565 7803
rect 36725 7763 36783 7769
rect 36832 7772 37565 7800
rect 36832 7732 36860 7772
rect 37553 7769 37565 7772
rect 37599 7769 37611 7803
rect 37553 7763 37611 7769
rect 38105 7803 38163 7809
rect 38105 7769 38117 7803
rect 38151 7769 38163 7803
rect 38105 7763 38163 7769
rect 38286 7760 38292 7812
rect 38344 7800 38350 7812
rect 39224 7809 39252 7840
rect 39850 7828 39856 7880
rect 39908 7868 39914 7880
rect 39908 7840 40540 7868
rect 39908 7828 39914 7840
rect 40512 7809 40540 7840
rect 38657 7803 38715 7809
rect 38657 7800 38669 7803
rect 38344 7772 38669 7800
rect 38344 7760 38350 7772
rect 38657 7769 38669 7772
rect 38703 7769 38715 7803
rect 38657 7763 38715 7769
rect 39209 7803 39267 7809
rect 39209 7769 39221 7803
rect 39255 7769 39267 7803
rect 39945 7803 40003 7809
rect 39945 7800 39957 7803
rect 39209 7763 39267 7769
rect 39316 7772 39957 7800
rect 35866 7704 36860 7732
rect 37458 7692 37464 7744
rect 37516 7732 37522 7744
rect 39316 7732 39344 7772
rect 39945 7769 39957 7772
rect 39991 7769 40003 7803
rect 39945 7763 40003 7769
rect 40497 7803 40555 7809
rect 40497 7769 40509 7803
rect 40543 7769 40555 7803
rect 40497 7763 40555 7769
rect 37516 7704 39344 7732
rect 37516 7692 37522 7704
rect 39390 7692 39396 7744
rect 39448 7732 39454 7744
rect 40037 7735 40095 7741
rect 40037 7732 40049 7735
rect 39448 7704 40049 7732
rect 39448 7692 39454 7704
rect 40037 7701 40049 7704
rect 40083 7701 40095 7735
rect 40037 7695 40095 7701
rect 1104 7642 44040 7664
rect 1104 7590 11644 7642
rect 11696 7590 11708 7642
rect 11760 7590 11772 7642
rect 11824 7590 11836 7642
rect 11888 7590 11900 7642
rect 11952 7590 22338 7642
rect 22390 7590 22402 7642
rect 22454 7590 22466 7642
rect 22518 7590 22530 7642
rect 22582 7590 22594 7642
rect 22646 7590 33032 7642
rect 33084 7590 33096 7642
rect 33148 7590 33160 7642
rect 33212 7590 33224 7642
rect 33276 7590 33288 7642
rect 33340 7590 43726 7642
rect 43778 7590 43790 7642
rect 43842 7590 43854 7642
rect 43906 7590 43918 7642
rect 43970 7590 43982 7642
rect 44034 7590 44040 7642
rect 1104 7568 44040 7590
rect 5810 7488 5816 7540
rect 5868 7488 5874 7540
rect 6089 7531 6147 7537
rect 6089 7497 6101 7531
rect 6135 7528 6147 7531
rect 6638 7528 6644 7540
rect 6135 7500 6644 7528
rect 6135 7497 6147 7500
rect 6089 7491 6147 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7193 7531 7251 7537
rect 7193 7497 7205 7531
rect 7239 7528 7251 7531
rect 7282 7528 7288 7540
rect 7239 7500 7288 7528
rect 7239 7497 7251 7500
rect 7193 7491 7251 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 8018 7488 8024 7540
rect 8076 7488 8082 7540
rect 11974 7488 11980 7540
rect 12032 7488 12038 7540
rect 12897 7531 12955 7537
rect 12897 7497 12909 7531
rect 12943 7528 12955 7531
rect 13078 7528 13084 7540
rect 12943 7500 13084 7528
rect 12943 7497 12955 7500
rect 12897 7491 12955 7497
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 14918 7488 14924 7540
rect 14976 7528 14982 7540
rect 14976 7500 16344 7528
rect 14976 7488 14982 7500
rect 5828 7460 5856 7488
rect 6546 7460 6552 7472
rect 5828 7432 6552 7460
rect 6546 7420 6552 7432
rect 6604 7420 6610 7472
rect 15102 7460 15108 7472
rect 11808 7432 15108 7460
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 7006 7352 7012 7404
rect 7064 7352 7070 7404
rect 7374 7352 7380 7404
rect 7432 7352 7438 7404
rect 11808 7401 11836 7432
rect 15102 7420 15108 7432
rect 15160 7420 15166 7472
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7361 11851 7395
rect 11793 7355 11851 7361
rect 12710 7352 12716 7404
rect 12768 7352 12774 7404
rect 16316 7392 16344 7500
rect 16390 7488 16396 7540
rect 16448 7488 16454 7540
rect 17494 7488 17500 7540
rect 17552 7488 17558 7540
rect 17770 7488 17776 7540
rect 17828 7528 17834 7540
rect 18141 7531 18199 7537
rect 18141 7528 18153 7531
rect 17828 7500 18153 7528
rect 17828 7488 17834 7500
rect 18141 7497 18153 7500
rect 18187 7497 18199 7531
rect 18141 7491 18199 7497
rect 18322 7488 18328 7540
rect 18380 7488 18386 7540
rect 18414 7488 18420 7540
rect 18472 7528 18478 7540
rect 18693 7531 18751 7537
rect 18693 7528 18705 7531
rect 18472 7500 18705 7528
rect 18472 7488 18478 7500
rect 18693 7497 18705 7500
rect 18739 7497 18751 7531
rect 18693 7491 18751 7497
rect 19886 7488 19892 7540
rect 19944 7488 19950 7540
rect 20898 7488 20904 7540
rect 20956 7488 20962 7540
rect 20990 7488 20996 7540
rect 21048 7528 21054 7540
rect 22925 7531 22983 7537
rect 21048 7500 22508 7528
rect 21048 7488 21054 7500
rect 16408 7460 16436 7488
rect 18340 7460 18368 7488
rect 16408 7432 18276 7460
rect 18340 7432 20024 7460
rect 17586 7392 17592 7404
rect 16316 7364 17592 7392
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 17862 7392 17868 7404
rect 17727 7364 17868 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 17957 7395 18015 7401
rect 17957 7361 17969 7395
rect 18003 7392 18015 7395
rect 18138 7392 18144 7404
rect 18003 7364 18144 7392
rect 18003 7361 18015 7364
rect 17957 7355 18015 7361
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 8110 7324 8116 7336
rect 7576 7296 8116 7324
rect 7576 7265 7604 7296
rect 8110 7284 8116 7296
rect 8168 7284 8174 7336
rect 9214 7284 9220 7336
rect 9272 7324 9278 7336
rect 16482 7324 16488 7336
rect 9272 7296 16488 7324
rect 9272 7284 9278 7296
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 18248 7324 18276 7432
rect 18325 7395 18383 7401
rect 18325 7361 18337 7395
rect 18371 7392 18383 7395
rect 18506 7392 18512 7404
rect 18371 7364 18512 7392
rect 18371 7361 18383 7364
rect 18325 7355 18383 7361
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 18598 7352 18604 7404
rect 18656 7352 18662 7404
rect 18877 7395 18935 7401
rect 18877 7361 18889 7395
rect 18923 7392 18935 7395
rect 19058 7392 19064 7404
rect 18923 7364 19064 7392
rect 18923 7361 18935 7364
rect 18877 7355 18935 7361
rect 19058 7352 19064 7364
rect 19116 7352 19122 7404
rect 19150 7352 19156 7404
rect 19208 7352 19214 7404
rect 19334 7392 19340 7404
rect 19306 7352 19340 7392
rect 19392 7352 19398 7404
rect 19429 7395 19487 7401
rect 19429 7361 19441 7395
rect 19475 7392 19487 7395
rect 19518 7392 19524 7404
rect 19475 7364 19524 7392
rect 19475 7361 19487 7364
rect 19429 7355 19487 7361
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 19996 7401 20024 7432
rect 19705 7395 19763 7401
rect 19705 7361 19717 7395
rect 19751 7392 19763 7395
rect 19981 7395 20039 7401
rect 19751 7364 19840 7392
rect 19751 7361 19763 7364
rect 19705 7355 19763 7361
rect 19306 7324 19334 7352
rect 18248 7296 19334 7324
rect 7561 7259 7619 7265
rect 7561 7225 7573 7259
rect 7607 7225 7619 7259
rect 7561 7219 7619 7225
rect 8386 7216 8392 7268
rect 8444 7256 8450 7268
rect 15562 7256 15568 7268
rect 8444 7228 15568 7256
rect 8444 7216 8450 7228
rect 15562 7216 15568 7228
rect 15620 7216 15626 7268
rect 19337 7259 19395 7265
rect 19337 7256 19349 7259
rect 15856 7228 19349 7256
rect 7742 7148 7748 7200
rect 7800 7188 7806 7200
rect 15856 7188 15884 7228
rect 19337 7225 19349 7228
rect 19383 7225 19395 7259
rect 19337 7219 19395 7225
rect 19610 7216 19616 7268
rect 19668 7216 19674 7268
rect 7800 7160 15884 7188
rect 7800 7148 7806 7160
rect 16758 7148 16764 7200
rect 16816 7188 16822 7200
rect 17773 7191 17831 7197
rect 17773 7188 17785 7191
rect 16816 7160 17785 7188
rect 16816 7148 16822 7160
rect 17773 7157 17785 7160
rect 17819 7157 17831 7191
rect 17773 7151 17831 7157
rect 18046 7148 18052 7200
rect 18104 7188 18110 7200
rect 18417 7191 18475 7197
rect 18417 7188 18429 7191
rect 18104 7160 18429 7188
rect 18104 7148 18110 7160
rect 18417 7157 18429 7160
rect 18463 7157 18475 7191
rect 18417 7151 18475 7157
rect 18598 7148 18604 7200
rect 18656 7188 18662 7200
rect 19242 7188 19248 7200
rect 18656 7160 19248 7188
rect 18656 7148 18662 7160
rect 19242 7148 19248 7160
rect 19300 7148 19306 7200
rect 19812 7188 19840 7364
rect 19981 7361 19993 7395
rect 20027 7361 20039 7395
rect 19981 7355 20039 7361
rect 20254 7352 20260 7404
rect 20312 7392 20318 7404
rect 20533 7395 20591 7401
rect 20533 7392 20545 7395
rect 20312 7364 20545 7392
rect 20312 7352 20318 7364
rect 20533 7361 20545 7364
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 20809 7395 20867 7401
rect 20809 7361 20821 7395
rect 20855 7392 20867 7395
rect 20916 7392 20944 7488
rect 21082 7420 21088 7472
rect 21140 7420 21146 7472
rect 21910 7460 21916 7472
rect 21284 7432 21916 7460
rect 20855 7364 20944 7392
rect 20855 7361 20867 7364
rect 20809 7355 20867 7361
rect 21100 7324 21128 7420
rect 21284 7401 21312 7432
rect 21910 7420 21916 7432
rect 21968 7420 21974 7472
rect 22480 7460 22508 7500
rect 22925 7497 22937 7531
rect 22971 7528 22983 7531
rect 23198 7528 23204 7540
rect 22971 7500 23204 7528
rect 22971 7497 22983 7500
rect 22925 7491 22983 7497
rect 23198 7488 23204 7500
rect 23256 7488 23262 7540
rect 23382 7488 23388 7540
rect 23440 7488 23446 7540
rect 23474 7488 23480 7540
rect 23532 7488 23538 7540
rect 23934 7488 23940 7540
rect 23992 7488 23998 7540
rect 24302 7488 24308 7540
rect 24360 7528 24366 7540
rect 28258 7528 28264 7540
rect 24360 7500 28264 7528
rect 24360 7488 24366 7500
rect 28258 7488 28264 7500
rect 28316 7488 28322 7540
rect 29546 7528 29552 7540
rect 28460 7500 29552 7528
rect 23400 7460 23428 7488
rect 22480 7432 22692 7460
rect 21269 7395 21327 7401
rect 21269 7361 21281 7395
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 21726 7392 21732 7404
rect 21407 7364 21732 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 21726 7352 21732 7364
rect 21784 7352 21790 7404
rect 22002 7352 22008 7404
rect 22060 7352 22066 7404
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7392 22339 7395
rect 22462 7392 22468 7404
rect 22327 7364 22468 7392
rect 22327 7361 22339 7364
rect 22281 7355 22339 7361
rect 22462 7352 22468 7364
rect 22520 7352 22526 7404
rect 21100 7296 21220 7324
rect 20349 7259 20407 7265
rect 20349 7256 20361 7259
rect 20088 7228 20361 7256
rect 20088 7188 20116 7228
rect 20349 7225 20361 7228
rect 20395 7225 20407 7259
rect 20349 7219 20407 7225
rect 21082 7216 21088 7268
rect 21140 7216 21146 7268
rect 21192 7256 21220 7296
rect 21542 7284 21548 7336
rect 21600 7324 21606 7336
rect 22370 7324 22376 7336
rect 21600 7296 22376 7324
rect 21600 7284 21606 7296
rect 22370 7284 22376 7296
rect 22428 7284 22434 7336
rect 22664 7324 22692 7432
rect 22848 7432 23428 7460
rect 22741 7396 22799 7401
rect 22848 7396 22876 7432
rect 22741 7395 22876 7396
rect 22741 7361 22753 7395
rect 22787 7368 22876 7395
rect 23293 7395 23351 7401
rect 22787 7361 22799 7368
rect 22741 7355 22799 7361
rect 23293 7361 23305 7395
rect 23339 7392 23351 7395
rect 23952 7392 23980 7488
rect 24486 7420 24492 7472
rect 24544 7460 24550 7472
rect 28460 7460 28488 7500
rect 29546 7488 29552 7500
rect 29604 7488 29610 7540
rect 33778 7488 33784 7540
rect 33836 7488 33842 7540
rect 34054 7488 34060 7540
rect 34112 7488 34118 7540
rect 24544 7432 28488 7460
rect 24544 7420 24550 7432
rect 23339 7364 23980 7392
rect 26421 7395 26479 7401
rect 23339 7361 23351 7364
rect 23293 7355 23351 7361
rect 26421 7361 26433 7395
rect 26467 7392 26479 7395
rect 28350 7392 28356 7404
rect 26467 7364 28356 7392
rect 26467 7361 26479 7364
rect 26421 7355 26479 7361
rect 28350 7352 28356 7364
rect 28408 7352 28414 7404
rect 33796 7324 33824 7488
rect 22664 7296 33824 7324
rect 21821 7259 21879 7265
rect 21821 7256 21833 7259
rect 21192 7228 21833 7256
rect 21821 7225 21833 7228
rect 21867 7225 21879 7259
rect 21821 7219 21879 7225
rect 22097 7259 22155 7265
rect 22097 7225 22109 7259
rect 22143 7256 22155 7259
rect 22186 7256 22192 7268
rect 22143 7228 22192 7256
rect 22143 7225 22155 7228
rect 22097 7219 22155 7225
rect 22186 7216 22192 7228
rect 22244 7216 22250 7268
rect 22462 7216 22468 7268
rect 22520 7216 22526 7268
rect 22554 7216 22560 7268
rect 22612 7256 22618 7268
rect 34072 7256 34100 7488
rect 37274 7284 37280 7336
rect 37332 7324 37338 7336
rect 38286 7324 38292 7336
rect 37332 7296 38292 7324
rect 37332 7284 37338 7296
rect 38286 7284 38292 7296
rect 38344 7284 38350 7336
rect 22612 7228 34100 7256
rect 22612 7216 22618 7228
rect 19812 7160 20116 7188
rect 20162 7148 20168 7200
rect 20220 7148 20226 7200
rect 20990 7148 20996 7200
rect 21048 7148 21054 7200
rect 21450 7148 21456 7200
rect 21508 7188 21514 7200
rect 21545 7191 21603 7197
rect 21545 7188 21557 7191
rect 21508 7160 21557 7188
rect 21508 7148 21514 7160
rect 21545 7157 21557 7160
rect 21591 7157 21603 7191
rect 22480 7188 22508 7216
rect 24578 7188 24584 7200
rect 22480 7160 24584 7188
rect 21545 7151 21603 7157
rect 24578 7148 24584 7160
rect 24636 7148 24642 7200
rect 24854 7148 24860 7200
rect 24912 7188 24918 7200
rect 26605 7191 26663 7197
rect 26605 7188 26617 7191
rect 24912 7160 26617 7188
rect 24912 7148 24918 7160
rect 26605 7157 26617 7160
rect 26651 7157 26663 7191
rect 26605 7151 26663 7157
rect 1104 7098 43884 7120
rect 1104 7046 6297 7098
rect 6349 7046 6361 7098
rect 6413 7046 6425 7098
rect 6477 7046 6489 7098
rect 6541 7046 6553 7098
rect 6605 7046 16991 7098
rect 17043 7046 17055 7098
rect 17107 7046 17119 7098
rect 17171 7046 17183 7098
rect 17235 7046 17247 7098
rect 17299 7046 27685 7098
rect 27737 7046 27749 7098
rect 27801 7046 27813 7098
rect 27865 7046 27877 7098
rect 27929 7046 27941 7098
rect 27993 7046 38379 7098
rect 38431 7046 38443 7098
rect 38495 7046 38507 7098
rect 38559 7046 38571 7098
rect 38623 7046 38635 7098
rect 38687 7046 43884 7098
rect 1104 7024 43884 7046
rect 10042 6944 10048 6996
rect 10100 6984 10106 6996
rect 10100 6956 12434 6984
rect 10100 6944 10106 6956
rect 12406 6916 12434 6956
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 20073 6987 20131 6993
rect 20073 6984 20085 6987
rect 19576 6956 20085 6984
rect 19576 6944 19582 6956
rect 20073 6953 20085 6956
rect 20119 6953 20131 6987
rect 20073 6947 20131 6953
rect 20990 6944 20996 6996
rect 21048 6944 21054 6996
rect 21266 6944 21272 6996
rect 21324 6944 21330 6996
rect 23290 6984 23296 6996
rect 22066 6956 23296 6984
rect 21008 6916 21036 6944
rect 12406 6888 21036 6916
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 10318 6848 10324 6860
rect 9456 6820 10324 6848
rect 9456 6808 9462 6820
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 16482 6808 16488 6860
rect 16540 6848 16546 6860
rect 21284 6848 21312 6944
rect 21450 6876 21456 6928
rect 21508 6916 21514 6928
rect 22066 6916 22094 6956
rect 23290 6944 23296 6956
rect 23348 6944 23354 6996
rect 29822 6944 29828 6996
rect 29880 6944 29886 6996
rect 21508 6888 22094 6916
rect 21508 6876 21514 6888
rect 22738 6876 22744 6928
rect 22796 6916 22802 6928
rect 29840 6916 29868 6944
rect 22796 6888 29868 6916
rect 22796 6876 22802 6888
rect 16540 6820 21312 6848
rect 16540 6808 16546 6820
rect 21910 6808 21916 6860
rect 21968 6848 21974 6860
rect 25130 6848 25136 6860
rect 21968 6820 25136 6848
rect 21968 6808 21974 6820
rect 25130 6808 25136 6820
rect 25188 6808 25194 6860
rect 38102 6808 38108 6860
rect 38160 6848 38166 6860
rect 39390 6848 39396 6860
rect 38160 6820 39396 6848
rect 38160 6808 38166 6820
rect 39390 6808 39396 6820
rect 39448 6808 39454 6860
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 7466 6780 7472 6792
rect 7055 6752 7472 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 18782 6740 18788 6792
rect 18840 6740 18846 6792
rect 19150 6740 19156 6792
rect 19208 6740 19214 6792
rect 19978 6740 19984 6792
rect 20036 6740 20042 6792
rect 20254 6740 20260 6792
rect 20312 6740 20318 6792
rect 21082 6740 21088 6792
rect 21140 6740 21146 6792
rect 18690 6672 18696 6724
rect 18748 6672 18754 6724
rect 18601 6647 18659 6653
rect 18601 6613 18613 6647
rect 18647 6644 18659 6647
rect 18708 6644 18736 6672
rect 18647 6616 18736 6644
rect 19168 6644 19196 6740
rect 19334 6672 19340 6724
rect 19392 6712 19398 6724
rect 21100 6712 21128 6740
rect 19392 6684 21128 6712
rect 19392 6672 19398 6684
rect 19797 6647 19855 6653
rect 19797 6644 19809 6647
rect 19168 6616 19809 6644
rect 18647 6613 18659 6616
rect 18601 6607 18659 6613
rect 19797 6613 19809 6616
rect 19843 6613 19855 6647
rect 19797 6607 19855 6613
rect 1104 6554 44040 6576
rect 1104 6502 11644 6554
rect 11696 6502 11708 6554
rect 11760 6502 11772 6554
rect 11824 6502 11836 6554
rect 11888 6502 11900 6554
rect 11952 6502 22338 6554
rect 22390 6502 22402 6554
rect 22454 6502 22466 6554
rect 22518 6502 22530 6554
rect 22582 6502 22594 6554
rect 22646 6502 33032 6554
rect 33084 6502 33096 6554
rect 33148 6502 33160 6554
rect 33212 6502 33224 6554
rect 33276 6502 33288 6554
rect 33340 6502 43726 6554
rect 43778 6502 43790 6554
rect 43842 6502 43854 6554
rect 43906 6502 43918 6554
rect 43970 6502 43982 6554
rect 44034 6502 44040 6554
rect 1104 6480 44040 6502
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 5960 6412 12434 6440
rect 5960 6400 5966 6412
rect 12406 6372 12434 6412
rect 13722 6400 13728 6452
rect 13780 6440 13786 6452
rect 21818 6440 21824 6452
rect 13780 6412 21824 6440
rect 13780 6400 13786 6412
rect 21818 6400 21824 6412
rect 21876 6400 21882 6452
rect 21910 6372 21916 6384
rect 12406 6344 21916 6372
rect 21910 6332 21916 6344
rect 21968 6332 21974 6384
rect 17586 6264 17592 6316
rect 17644 6304 17650 6316
rect 25958 6304 25964 6316
rect 17644 6276 25964 6304
rect 17644 6264 17650 6276
rect 25958 6264 25964 6276
rect 26016 6264 26022 6316
rect 12250 6196 12256 6248
rect 12308 6236 12314 6248
rect 12308 6208 12434 6236
rect 12308 6196 12314 6208
rect 12406 6100 12434 6208
rect 15470 6196 15476 6248
rect 15528 6236 15534 6248
rect 26142 6236 26148 6248
rect 15528 6208 26148 6236
rect 15528 6196 15534 6208
rect 26142 6196 26148 6208
rect 26200 6196 26206 6248
rect 16666 6128 16672 6180
rect 16724 6168 16730 6180
rect 26234 6168 26240 6180
rect 16724 6140 26240 6168
rect 16724 6128 16730 6140
rect 26234 6128 26240 6140
rect 26292 6128 26298 6180
rect 17310 6100 17316 6112
rect 12406 6072 17316 6100
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 1104 6010 43884 6032
rect 1104 5958 6297 6010
rect 6349 5958 6361 6010
rect 6413 5958 6425 6010
rect 6477 5958 6489 6010
rect 6541 5958 6553 6010
rect 6605 5958 16991 6010
rect 17043 5958 17055 6010
rect 17107 5958 17119 6010
rect 17171 5958 17183 6010
rect 17235 5958 17247 6010
rect 17299 5958 27685 6010
rect 27737 5958 27749 6010
rect 27801 5958 27813 6010
rect 27865 5958 27877 6010
rect 27929 5958 27941 6010
rect 27993 5958 38379 6010
rect 38431 5958 38443 6010
rect 38495 5958 38507 6010
rect 38559 5958 38571 6010
rect 38623 5958 38635 6010
rect 38687 5958 43884 6010
rect 1104 5936 43884 5958
rect 18782 5856 18788 5908
rect 18840 5896 18846 5908
rect 30834 5896 30840 5908
rect 18840 5868 30840 5896
rect 18840 5856 18846 5868
rect 30834 5856 30840 5868
rect 30892 5856 30898 5908
rect 17310 5788 17316 5840
rect 17368 5828 17374 5840
rect 24854 5828 24860 5840
rect 17368 5800 24860 5828
rect 17368 5788 17374 5800
rect 24854 5788 24860 5800
rect 24912 5788 24918 5840
rect 22738 5584 22744 5636
rect 22796 5624 22802 5636
rect 28994 5624 29000 5636
rect 22796 5596 29000 5624
rect 22796 5584 22802 5596
rect 28994 5584 29000 5596
rect 29052 5584 29058 5636
rect 1104 5466 44040 5488
rect 1104 5414 11644 5466
rect 11696 5414 11708 5466
rect 11760 5414 11772 5466
rect 11824 5414 11836 5466
rect 11888 5414 11900 5466
rect 11952 5414 22338 5466
rect 22390 5414 22402 5466
rect 22454 5414 22466 5466
rect 22518 5414 22530 5466
rect 22582 5414 22594 5466
rect 22646 5414 33032 5466
rect 33084 5414 33096 5466
rect 33148 5414 33160 5466
rect 33212 5414 33224 5466
rect 33276 5414 33288 5466
rect 33340 5414 43726 5466
rect 43778 5414 43790 5466
rect 43842 5414 43854 5466
rect 43906 5414 43918 5466
rect 43970 5414 43982 5466
rect 44034 5414 44040 5466
rect 1104 5392 44040 5414
rect 37458 5312 37464 5364
rect 37516 5312 37522 5364
rect 37642 5176 37648 5228
rect 37700 5176 37706 5228
rect 25958 5108 25964 5160
rect 26016 5148 26022 5160
rect 30650 5148 30656 5160
rect 26016 5120 30656 5148
rect 26016 5108 26022 5120
rect 30650 5108 30656 5120
rect 30708 5108 30714 5160
rect 26050 4972 26056 5024
rect 26108 5012 26114 5024
rect 36262 5012 36268 5024
rect 26108 4984 36268 5012
rect 26108 4972 26114 4984
rect 36262 4972 36268 4984
rect 36320 4972 36326 5024
rect 1104 4922 43884 4944
rect 1104 4870 6297 4922
rect 6349 4870 6361 4922
rect 6413 4870 6425 4922
rect 6477 4870 6489 4922
rect 6541 4870 6553 4922
rect 6605 4870 16991 4922
rect 17043 4870 17055 4922
rect 17107 4870 17119 4922
rect 17171 4870 17183 4922
rect 17235 4870 17247 4922
rect 17299 4870 27685 4922
rect 27737 4870 27749 4922
rect 27801 4870 27813 4922
rect 27865 4870 27877 4922
rect 27929 4870 27941 4922
rect 27993 4870 38379 4922
rect 38431 4870 38443 4922
rect 38495 4870 38507 4922
rect 38559 4870 38571 4922
rect 38623 4870 38635 4922
rect 38687 4870 43884 4922
rect 1104 4848 43884 4870
rect 22738 4768 22744 4820
rect 22796 4768 22802 4820
rect 25958 4808 25964 4820
rect 22940 4780 25964 4808
rect 21821 4743 21879 4749
rect 21821 4709 21833 4743
rect 21867 4740 21879 4743
rect 22940 4740 22968 4780
rect 25958 4768 25964 4780
rect 26016 4768 26022 4820
rect 26050 4768 26056 4820
rect 26108 4768 26114 4820
rect 28169 4811 28227 4817
rect 28169 4777 28181 4811
rect 28215 4808 28227 4811
rect 34514 4808 34520 4820
rect 28215 4780 34520 4808
rect 28215 4777 28227 4780
rect 28169 4771 28227 4777
rect 34514 4768 34520 4780
rect 34572 4768 34578 4820
rect 36633 4811 36691 4817
rect 36633 4777 36645 4811
rect 36679 4808 36691 4811
rect 37642 4808 37648 4820
rect 36679 4780 37648 4808
rect 36679 4777 36691 4780
rect 36633 4771 36691 4777
rect 37642 4768 37648 4780
rect 37700 4768 37706 4820
rect 38194 4768 38200 4820
rect 38252 4768 38258 4820
rect 21867 4712 22968 4740
rect 23017 4743 23075 4749
rect 21867 4709 21879 4712
rect 21821 4703 21879 4709
rect 23017 4709 23029 4743
rect 23063 4740 23075 4743
rect 32401 4743 32459 4749
rect 23063 4712 31754 4740
rect 23063 4709 23075 4712
rect 23017 4703 23075 4709
rect 30374 4672 30380 4684
rect 23308 4644 30380 4672
rect 21634 4564 21640 4616
rect 21692 4564 21698 4616
rect 22186 4564 22192 4616
rect 22244 4604 22250 4616
rect 22557 4607 22615 4613
rect 22557 4604 22569 4607
rect 22244 4576 22569 4604
rect 22244 4564 22250 4576
rect 22557 4573 22569 4576
rect 22603 4573 22615 4607
rect 22557 4567 22615 4573
rect 22738 4564 22744 4616
rect 22796 4604 22802 4616
rect 22833 4607 22891 4613
rect 22833 4604 22845 4607
rect 22796 4576 22845 4604
rect 22796 4564 22802 4576
rect 22833 4573 22845 4576
rect 22879 4573 22891 4607
rect 22833 4567 22891 4573
rect 23106 4564 23112 4616
rect 23164 4564 23170 4616
rect 23308 4477 23336 4644
rect 30374 4632 30380 4644
rect 30432 4632 30438 4684
rect 31726 4672 31754 4712
rect 32401 4709 32413 4743
rect 32447 4740 32459 4743
rect 39298 4740 39304 4752
rect 32447 4712 39304 4740
rect 32447 4709 32459 4712
rect 32401 4703 32459 4709
rect 39298 4700 39304 4712
rect 39356 4700 39362 4752
rect 35434 4672 35440 4684
rect 31726 4644 35440 4672
rect 35434 4632 35440 4644
rect 35492 4632 35498 4684
rect 23382 4564 23388 4616
rect 23440 4564 23446 4616
rect 25866 4564 25872 4616
rect 25924 4564 25930 4616
rect 27982 4564 27988 4616
rect 28040 4564 28046 4616
rect 32214 4564 32220 4616
rect 32272 4564 32278 4616
rect 34514 4564 34520 4616
rect 34572 4604 34578 4616
rect 36817 4607 36875 4613
rect 36817 4604 36829 4607
rect 34572 4576 36829 4604
rect 34572 4564 34578 4576
rect 36817 4573 36829 4576
rect 36863 4573 36875 4607
rect 36817 4567 36875 4573
rect 38378 4564 38384 4616
rect 38436 4564 38442 4616
rect 36446 4536 36452 4548
rect 23584 4508 31754 4536
rect 23584 4477 23612 4508
rect 23293 4471 23351 4477
rect 23293 4437 23305 4471
rect 23339 4437 23351 4471
rect 23293 4431 23351 4437
rect 23569 4471 23627 4477
rect 23569 4437 23581 4471
rect 23615 4437 23627 4471
rect 31726 4468 31754 4508
rect 35866 4508 36452 4536
rect 35866 4468 35894 4508
rect 36446 4496 36452 4508
rect 36504 4496 36510 4548
rect 31726 4440 35894 4468
rect 23569 4431 23627 4437
rect 1104 4378 44040 4400
rect 1104 4326 11644 4378
rect 11696 4326 11708 4378
rect 11760 4326 11772 4378
rect 11824 4326 11836 4378
rect 11888 4326 11900 4378
rect 11952 4326 22338 4378
rect 22390 4326 22402 4378
rect 22454 4326 22466 4378
rect 22518 4326 22530 4378
rect 22582 4326 22594 4378
rect 22646 4326 33032 4378
rect 33084 4326 33096 4378
rect 33148 4326 33160 4378
rect 33212 4326 33224 4378
rect 33276 4326 33288 4378
rect 33340 4326 43726 4378
rect 43778 4326 43790 4378
rect 43842 4326 43854 4378
rect 43906 4326 43918 4378
rect 43970 4326 43982 4378
rect 44034 4326 44040 4378
rect 1104 4304 44040 4326
rect 20901 4267 20959 4273
rect 20901 4233 20913 4267
rect 20947 4264 20959 4267
rect 21634 4264 21640 4276
rect 20947 4236 21640 4264
rect 20947 4233 20959 4236
rect 20901 4227 20959 4233
rect 21634 4224 21640 4236
rect 21692 4224 21698 4276
rect 22097 4267 22155 4273
rect 22097 4233 22109 4267
rect 22143 4233 22155 4267
rect 22097 4227 22155 4233
rect 22649 4267 22707 4273
rect 22649 4233 22661 4267
rect 22695 4264 22707 4267
rect 23382 4264 23388 4276
rect 22695 4236 23388 4264
rect 22695 4233 22707 4236
rect 22649 4227 22707 4233
rect 22112 4196 22140 4227
rect 23382 4224 23388 4236
rect 23440 4224 23446 4276
rect 25133 4267 25191 4273
rect 25133 4233 25145 4267
rect 25179 4264 25191 4267
rect 25866 4264 25872 4276
rect 25179 4236 25872 4264
rect 25179 4233 25191 4236
rect 25133 4227 25191 4233
rect 25866 4224 25872 4236
rect 25924 4224 25930 4276
rect 37645 4267 37703 4273
rect 37645 4233 37657 4267
rect 37691 4264 37703 4267
rect 38378 4264 38384 4276
rect 37691 4236 38384 4264
rect 37691 4233 37703 4236
rect 37645 4227 37703 4233
rect 38378 4224 38384 4236
rect 38436 4224 38442 4276
rect 22738 4196 22744 4208
rect 22112 4168 22744 4196
rect 22738 4156 22744 4168
rect 22796 4156 22802 4208
rect 20530 4088 20536 4140
rect 20588 4128 20594 4140
rect 21085 4131 21143 4137
rect 21085 4128 21097 4131
rect 20588 4100 21097 4128
rect 20588 4088 20594 4100
rect 21085 4097 21097 4100
rect 21131 4097 21143 4131
rect 21085 4091 21143 4097
rect 22002 4088 22008 4140
rect 22060 4088 22066 4140
rect 22281 4131 22339 4137
rect 22281 4097 22293 4131
rect 22327 4097 22339 4131
rect 22281 4091 22339 4097
rect 22557 4131 22615 4137
rect 22557 4097 22569 4131
rect 22603 4097 22615 4131
rect 22557 4091 22615 4097
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 22296 4060 22324 4091
rect 7984 4032 22324 4060
rect 7984 4020 7990 4032
rect 21821 3995 21879 4001
rect 21821 3961 21833 3995
rect 21867 3992 21879 3995
rect 22186 3992 22192 4004
rect 21867 3964 22192 3992
rect 21867 3961 21879 3964
rect 21821 3955 21879 3961
rect 22186 3952 22192 3964
rect 22244 3952 22250 4004
rect 22572 3992 22600 4091
rect 22830 4088 22836 4140
rect 22888 4088 22894 4140
rect 23750 4088 23756 4140
rect 23808 4088 23814 4140
rect 24762 4088 24768 4140
rect 24820 4128 24826 4140
rect 25317 4131 25375 4137
rect 25317 4128 25329 4131
rect 24820 4100 25329 4128
rect 24820 4088 24826 4100
rect 25317 4097 25329 4100
rect 25363 4097 25375 4131
rect 25317 4091 25375 4097
rect 27430 4088 27436 4140
rect 27488 4088 27494 4140
rect 31662 4088 31668 4140
rect 31720 4088 31726 4140
rect 37366 4088 37372 4140
rect 37424 4128 37430 4140
rect 37829 4131 37887 4137
rect 37829 4128 37841 4131
rect 37424 4100 37841 4128
rect 37424 4088 37430 4100
rect 37829 4097 37841 4100
rect 37875 4097 37887 4131
rect 37829 4091 37887 4097
rect 27982 4020 27988 4072
rect 28040 4020 28046 4072
rect 32214 4020 32220 4072
rect 32272 4020 32278 4072
rect 22296 3964 22600 3992
rect 18230 3884 18236 3936
rect 18288 3924 18294 3936
rect 22296 3924 22324 3964
rect 23106 3952 23112 4004
rect 23164 3952 23170 4004
rect 27249 3995 27307 4001
rect 27249 3961 27261 3995
rect 27295 3992 27307 3995
rect 28000 3992 28028 4020
rect 27295 3964 28028 3992
rect 27295 3961 27307 3964
rect 27249 3955 27307 3961
rect 29270 3952 29276 4004
rect 29328 3952 29334 4004
rect 31481 3995 31539 4001
rect 31481 3961 31493 3995
rect 31527 3992 31539 3995
rect 32232 3992 32260 4020
rect 31527 3964 32260 3992
rect 31527 3961 31539 3964
rect 31481 3955 31539 3961
rect 18288 3896 22324 3924
rect 22373 3927 22431 3933
rect 18288 3884 18294 3896
rect 22373 3893 22385 3927
rect 22419 3924 22431 3927
rect 23124 3924 23152 3952
rect 22419 3896 23152 3924
rect 23937 3927 23995 3933
rect 22419 3893 22431 3896
rect 22373 3887 22431 3893
rect 23937 3893 23949 3927
rect 23983 3924 23995 3927
rect 29288 3924 29316 3952
rect 23983 3896 29316 3924
rect 23983 3893 23995 3896
rect 23937 3887 23995 3893
rect 1104 3834 43884 3856
rect 1104 3782 6297 3834
rect 6349 3782 6361 3834
rect 6413 3782 6425 3834
rect 6477 3782 6489 3834
rect 6541 3782 6553 3834
rect 6605 3782 16991 3834
rect 17043 3782 17055 3834
rect 17107 3782 17119 3834
rect 17171 3782 17183 3834
rect 17235 3782 17247 3834
rect 17299 3782 27685 3834
rect 27737 3782 27749 3834
rect 27801 3782 27813 3834
rect 27865 3782 27877 3834
rect 27929 3782 27941 3834
rect 27993 3782 38379 3834
rect 38431 3782 38443 3834
rect 38495 3782 38507 3834
rect 38559 3782 38571 3834
rect 38623 3782 38635 3834
rect 38687 3782 43884 3834
rect 1104 3760 43884 3782
rect 22002 3720 22008 3732
rect 6886 3692 22008 3720
rect 5810 3612 5816 3664
rect 5868 3652 5874 3664
rect 6886 3652 6914 3692
rect 22002 3680 22008 3692
rect 22060 3680 22066 3732
rect 23017 3723 23075 3729
rect 23017 3689 23029 3723
rect 23063 3720 23075 3723
rect 23750 3720 23756 3732
rect 23063 3692 23756 3720
rect 23063 3689 23075 3692
rect 23017 3683 23075 3689
rect 23750 3680 23756 3692
rect 23808 3680 23814 3732
rect 30285 3723 30343 3729
rect 30285 3689 30297 3723
rect 30331 3720 30343 3723
rect 36078 3720 36084 3732
rect 30331 3692 36084 3720
rect 30331 3689 30343 3692
rect 30285 3683 30343 3689
rect 36078 3680 36084 3692
rect 36136 3680 36142 3732
rect 37274 3680 37280 3732
rect 37332 3680 37338 3732
rect 39945 3723 40003 3729
rect 39945 3689 39957 3723
rect 39991 3720 40003 3723
rect 41046 3720 41052 3732
rect 39991 3692 41052 3720
rect 39991 3689 40003 3692
rect 39945 3683 40003 3689
rect 41046 3680 41052 3692
rect 41104 3680 41110 3732
rect 5868 3624 6914 3652
rect 19705 3655 19763 3661
rect 5868 3612 5874 3624
rect 19705 3621 19717 3655
rect 19751 3652 19763 3655
rect 34606 3652 34612 3664
rect 19751 3624 34612 3652
rect 19751 3621 19763 3624
rect 19705 3615 19763 3621
rect 34606 3612 34612 3624
rect 34664 3612 34670 3664
rect 19610 3544 19616 3596
rect 19668 3584 19674 3596
rect 22830 3584 22836 3596
rect 19668 3556 22836 3584
rect 19668 3544 19674 3556
rect 22830 3544 22836 3556
rect 22888 3544 22894 3596
rect 19518 3476 19524 3528
rect 19576 3476 19582 3528
rect 23198 3476 23204 3528
rect 23256 3476 23262 3528
rect 30098 3476 30104 3528
rect 30156 3476 30162 3528
rect 37458 3476 37464 3528
rect 37516 3476 37522 3528
rect 40126 3476 40132 3528
rect 40184 3476 40190 3528
rect 1104 3290 44040 3312
rect 1104 3238 11644 3290
rect 11696 3238 11708 3290
rect 11760 3238 11772 3290
rect 11824 3238 11836 3290
rect 11888 3238 11900 3290
rect 11952 3238 22338 3290
rect 22390 3238 22402 3290
rect 22454 3238 22466 3290
rect 22518 3238 22530 3290
rect 22582 3238 22594 3290
rect 22646 3238 33032 3290
rect 33084 3238 33096 3290
rect 33148 3238 33160 3290
rect 33212 3238 33224 3290
rect 33276 3238 33288 3290
rect 33340 3238 43726 3290
rect 43778 3238 43790 3290
rect 43842 3238 43854 3290
rect 43906 3238 43918 3290
rect 43970 3238 43982 3290
rect 44034 3238 44040 3290
rect 1104 3216 44040 3238
rect 18785 3179 18843 3185
rect 18785 3145 18797 3179
rect 18831 3176 18843 3179
rect 19518 3176 19524 3188
rect 18831 3148 19524 3176
rect 18831 3145 18843 3148
rect 18785 3139 18843 3145
rect 19518 3136 19524 3148
rect 19576 3136 19582 3188
rect 22557 3179 22615 3185
rect 22557 3145 22569 3179
rect 22603 3145 22615 3179
rect 22557 3139 22615 3145
rect 29365 3179 29423 3185
rect 29365 3145 29377 3179
rect 29411 3176 29423 3179
rect 30098 3176 30104 3188
rect 29411 3148 30104 3176
rect 29411 3145 29423 3148
rect 29365 3139 29423 3145
rect 22572 3108 22600 3139
rect 30098 3136 30104 3148
rect 30156 3136 30162 3188
rect 31478 3136 31484 3188
rect 31536 3136 31542 3188
rect 36173 3179 36231 3185
rect 36173 3145 36185 3179
rect 36219 3176 36231 3179
rect 37458 3176 37464 3188
rect 36219 3148 37464 3176
rect 36219 3145 36231 3148
rect 36173 3139 36231 3145
rect 37458 3136 37464 3148
rect 37516 3136 37522 3188
rect 40126 3136 40132 3188
rect 40184 3176 40190 3188
rect 40681 3179 40739 3185
rect 40681 3176 40693 3179
rect 40184 3148 40693 3176
rect 40184 3136 40190 3148
rect 40681 3145 40693 3148
rect 40727 3145 40739 3179
rect 40681 3139 40739 3145
rect 31496 3108 31524 3136
rect 22572 3080 31524 3108
rect 18966 3000 18972 3052
rect 19024 3000 19030 3052
rect 22002 3000 22008 3052
rect 22060 3000 22066 3052
rect 22370 3000 22376 3052
rect 22428 3000 22434 3052
rect 28902 3000 28908 3052
rect 28960 3040 28966 3052
rect 29549 3043 29607 3049
rect 29549 3040 29561 3043
rect 28960 3012 29561 3040
rect 28960 3000 28966 3012
rect 29549 3009 29561 3012
rect 29595 3009 29607 3043
rect 29549 3003 29607 3009
rect 35250 3000 35256 3052
rect 35308 3040 35314 3052
rect 36357 3043 36415 3049
rect 36357 3040 36369 3043
rect 35308 3012 36369 3040
rect 35308 3000 35314 3012
rect 36357 3009 36369 3012
rect 36403 3009 36415 3043
rect 36357 3003 36415 3009
rect 40862 3000 40868 3052
rect 40920 3000 40926 3052
rect 35986 2972 35992 2984
rect 31726 2944 35992 2972
rect 22189 2907 22247 2913
rect 22189 2873 22201 2907
rect 22235 2904 22247 2907
rect 31726 2904 31754 2944
rect 35986 2932 35992 2944
rect 36044 2932 36050 2984
rect 22235 2876 31754 2904
rect 22235 2873 22247 2876
rect 22189 2867 22247 2873
rect 1104 2746 43884 2768
rect 1104 2694 6297 2746
rect 6349 2694 6361 2746
rect 6413 2694 6425 2746
rect 6477 2694 6489 2746
rect 6541 2694 6553 2746
rect 6605 2694 16991 2746
rect 17043 2694 17055 2746
rect 17107 2694 17119 2746
rect 17171 2694 17183 2746
rect 17235 2694 17247 2746
rect 17299 2694 27685 2746
rect 27737 2694 27749 2746
rect 27801 2694 27813 2746
rect 27865 2694 27877 2746
rect 27929 2694 27941 2746
rect 27993 2694 38379 2746
rect 38431 2694 38443 2746
rect 38495 2694 38507 2746
rect 38559 2694 38571 2746
rect 38623 2694 38635 2746
rect 38687 2694 43884 2746
rect 1104 2672 43884 2694
rect 21269 2635 21327 2641
rect 21269 2601 21281 2635
rect 21315 2632 21327 2635
rect 22002 2632 22008 2644
rect 21315 2604 22008 2632
rect 21315 2601 21327 2604
rect 21269 2595 21327 2601
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 22370 2592 22376 2644
rect 22428 2592 22434 2644
rect 39850 2592 39856 2644
rect 39908 2592 39914 2644
rect 40494 2592 40500 2644
rect 40552 2592 40558 2644
rect 21545 2567 21603 2573
rect 21545 2533 21557 2567
rect 21591 2564 21603 2567
rect 22388 2564 22416 2592
rect 21591 2536 22416 2564
rect 38933 2567 38991 2573
rect 21591 2533 21603 2536
rect 21545 2527 21603 2533
rect 38933 2533 38945 2567
rect 38979 2564 38991 2567
rect 40512 2564 40540 2592
rect 38979 2536 40540 2564
rect 38979 2533 38991 2536
rect 38933 2527 38991 2533
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 21453 2431 21511 2437
rect 21453 2428 21465 2431
rect 19392 2400 21465 2428
rect 19392 2388 19398 2400
rect 21453 2397 21465 2400
rect 21499 2397 21511 2431
rect 21453 2391 21511 2397
rect 21726 2388 21732 2440
rect 21784 2388 21790 2440
rect 22830 2388 22836 2440
rect 22888 2388 22894 2440
rect 39114 2388 39120 2440
rect 39172 2388 39178 2440
rect 40034 2388 40040 2440
rect 40092 2388 40098 2440
rect 23017 2295 23075 2301
rect 23017 2261 23029 2295
rect 23063 2292 23075 2295
rect 32950 2292 32956 2304
rect 23063 2264 32956 2292
rect 23063 2261 23075 2264
rect 23017 2255 23075 2261
rect 32950 2252 32956 2264
rect 33008 2252 33014 2304
rect 1104 2202 44040 2224
rect 1104 2150 11644 2202
rect 11696 2150 11708 2202
rect 11760 2150 11772 2202
rect 11824 2150 11836 2202
rect 11888 2150 11900 2202
rect 11952 2150 22338 2202
rect 22390 2150 22402 2202
rect 22454 2150 22466 2202
rect 22518 2150 22530 2202
rect 22582 2150 22594 2202
rect 22646 2150 33032 2202
rect 33084 2150 33096 2202
rect 33148 2150 33160 2202
rect 33212 2150 33224 2202
rect 33276 2150 33288 2202
rect 33340 2150 43726 2202
rect 43778 2150 43790 2202
rect 43842 2150 43854 2202
rect 43906 2150 43918 2202
rect 43970 2150 43982 2202
rect 44034 2150 44040 2202
rect 1104 2128 44040 2150
rect 22097 2091 22155 2097
rect 22097 2057 22109 2091
rect 22143 2088 22155 2091
rect 22830 2088 22836 2100
rect 22143 2060 22836 2088
rect 22143 2057 22155 2060
rect 22097 2051 22155 2057
rect 22830 2048 22836 2060
rect 22888 2048 22894 2100
rect 39114 2048 39120 2100
rect 39172 2088 39178 2100
rect 39209 2091 39267 2097
rect 39209 2088 39221 2091
rect 39172 2060 39221 2088
rect 39172 2048 39178 2060
rect 39209 2057 39221 2060
rect 39255 2057 39267 2091
rect 39209 2051 39267 2057
rect 40034 2048 40040 2100
rect 40092 2048 40098 2100
rect 1578 1912 1584 1964
rect 1636 1952 1642 1964
rect 21821 1955 21879 1961
rect 21821 1952 21833 1955
rect 1636 1924 21833 1952
rect 1636 1912 1642 1924
rect 21821 1921 21833 1924
rect 21867 1921 21879 1955
rect 21821 1915 21879 1921
rect 22281 1955 22339 1961
rect 22281 1921 22293 1955
rect 22327 1921 22339 1955
rect 22281 1915 22339 1921
rect 3970 1844 3976 1896
rect 4028 1884 4034 1896
rect 22296 1884 22324 1915
rect 39390 1912 39396 1964
rect 39448 1912 39454 1964
rect 40221 1955 40279 1961
rect 40221 1921 40233 1955
rect 40267 1952 40279 1955
rect 43346 1952 43352 1964
rect 40267 1924 43352 1952
rect 40267 1921 40279 1924
rect 40221 1915 40279 1921
rect 43346 1912 43352 1924
rect 43404 1912 43410 1964
rect 4028 1856 22324 1884
rect 4028 1844 4034 1856
rect 22005 1819 22063 1825
rect 22005 1785 22017 1819
rect 22051 1816 22063 1819
rect 34146 1816 34152 1828
rect 22051 1788 34152 1816
rect 22051 1785 22063 1788
rect 22005 1779 22063 1785
rect 34146 1776 34152 1788
rect 34204 1776 34210 1828
rect 1104 1658 43884 1680
rect 1104 1606 6297 1658
rect 6349 1606 6361 1658
rect 6413 1606 6425 1658
rect 6477 1606 6489 1658
rect 6541 1606 6553 1658
rect 6605 1606 16991 1658
rect 17043 1606 17055 1658
rect 17107 1606 17119 1658
rect 17171 1606 17183 1658
rect 17235 1606 17247 1658
rect 17299 1606 27685 1658
rect 27737 1606 27749 1658
rect 27801 1606 27813 1658
rect 27865 1606 27877 1658
rect 27929 1606 27941 1658
rect 27993 1606 38379 1658
rect 38431 1606 38443 1658
rect 38495 1606 38507 1658
rect 38559 1606 38571 1658
rect 38623 1606 38635 1658
rect 38687 1606 43884 1658
rect 1104 1584 43884 1606
rect 1578 1504 1584 1556
rect 1636 1504 1642 1556
rect 3970 1504 3976 1556
rect 4028 1504 4034 1556
rect 39390 1504 39396 1556
rect 39448 1544 39454 1556
rect 39485 1547 39543 1553
rect 39485 1544 39497 1547
rect 39448 1516 39497 1544
rect 39448 1504 39454 1516
rect 39485 1513 39497 1516
rect 39531 1513 39543 1547
rect 39485 1507 39543 1513
rect 43346 1504 43352 1556
rect 43404 1504 43410 1556
rect 12161 1479 12219 1485
rect 12161 1445 12173 1479
rect 12207 1445 12219 1479
rect 12161 1439 12219 1445
rect 16209 1479 16267 1485
rect 16209 1445 16221 1479
rect 16255 1445 16267 1479
rect 16209 1439 16267 1445
rect 1302 1300 1308 1352
rect 1360 1340 1366 1352
rect 1397 1343 1455 1349
rect 1397 1340 1409 1343
rect 1360 1312 1409 1340
rect 1360 1300 1366 1312
rect 1397 1309 1409 1312
rect 1443 1309 1455 1343
rect 1397 1303 1455 1309
rect 3786 1300 3792 1352
rect 3844 1300 3850 1352
rect 5626 1300 5632 1352
rect 5684 1300 5690 1352
rect 5810 1300 5816 1352
rect 5868 1300 5874 1352
rect 7742 1300 7748 1352
rect 7800 1300 7806 1352
rect 9858 1300 9864 1352
rect 9916 1300 9922 1352
rect 11974 1300 11980 1352
rect 12032 1300 12038 1352
rect 12176 1340 12204 1439
rect 16224 1408 16252 1439
rect 14200 1380 14412 1408
rect 16224 1380 16528 1408
rect 14200 1340 14228 1380
rect 12176 1312 14228 1340
rect 14274 1300 14280 1352
rect 14332 1300 14338 1352
rect 14384 1340 14412 1380
rect 14384 1312 16344 1340
rect 5828 1213 5856 1300
rect 16316 1272 16344 1312
rect 16390 1300 16396 1352
rect 16448 1300 16454 1352
rect 16500 1340 16528 1380
rect 18892 1380 19104 1408
rect 16500 1312 18460 1340
rect 18138 1272 18144 1284
rect 10060 1244 14228 1272
rect 16316 1244 18144 1272
rect 5813 1207 5871 1213
rect 5813 1173 5825 1207
rect 5859 1173 5871 1207
rect 5813 1167 5871 1173
rect 7926 1164 7932 1216
rect 7984 1164 7990 1216
rect 10060 1213 10088 1244
rect 10045 1207 10103 1213
rect 10045 1173 10057 1207
rect 10091 1173 10103 1207
rect 10045 1167 10103 1173
rect 14090 1164 14096 1216
rect 14148 1164 14154 1216
rect 14200 1204 14228 1244
rect 18138 1232 18144 1244
rect 18196 1232 18202 1284
rect 18432 1272 18460 1312
rect 18506 1300 18512 1352
rect 18564 1300 18570 1352
rect 18892 1272 18920 1380
rect 18966 1300 18972 1352
rect 19024 1300 19030 1352
rect 19076 1340 19104 1380
rect 19334 1340 19340 1352
rect 19076 1312 19340 1340
rect 19334 1300 19340 1312
rect 19392 1300 19398 1352
rect 20622 1300 20628 1352
rect 20680 1300 20686 1352
rect 22738 1300 22744 1352
rect 22796 1300 22802 1352
rect 23198 1300 23204 1352
rect 23256 1300 23262 1352
rect 24854 1300 24860 1352
rect 24912 1300 24918 1352
rect 26694 1300 26700 1352
rect 26752 1340 26758 1352
rect 27157 1343 27215 1349
rect 27157 1340 27169 1343
rect 26752 1312 27169 1340
rect 26752 1300 26758 1312
rect 27157 1309 27169 1312
rect 27203 1309 27215 1343
rect 27157 1303 27215 1309
rect 27430 1300 27436 1352
rect 27488 1300 27494 1352
rect 28902 1300 28908 1352
rect 28960 1300 28966 1352
rect 29086 1300 29092 1352
rect 29144 1300 29150 1352
rect 31202 1300 31208 1352
rect 31260 1300 31266 1352
rect 31662 1300 31668 1352
rect 31720 1300 31726 1352
rect 33318 1300 33324 1352
rect 33376 1300 33382 1352
rect 34514 1300 34520 1352
rect 34572 1300 34578 1352
rect 35250 1300 35256 1352
rect 35308 1300 35314 1352
rect 35434 1300 35440 1352
rect 35492 1300 35498 1352
rect 37550 1300 37556 1352
rect 37608 1300 37614 1352
rect 39390 1300 39396 1352
rect 39448 1340 39454 1352
rect 39669 1343 39727 1349
rect 39669 1340 39681 1343
rect 39448 1312 39681 1340
rect 39448 1300 39454 1312
rect 39669 1309 39681 1312
rect 39715 1309 39727 1343
rect 39669 1303 39727 1309
rect 40862 1300 40868 1352
rect 40920 1300 40926 1352
rect 41782 1300 41788 1352
rect 41840 1300 41846 1352
rect 43530 1300 43536 1352
rect 43588 1300 43594 1352
rect 18432 1244 18920 1272
rect 18230 1204 18236 1216
rect 14200 1176 18236 1204
rect 18230 1164 18236 1176
rect 18288 1164 18294 1216
rect 18325 1207 18383 1213
rect 18325 1173 18337 1207
rect 18371 1204 18383 1207
rect 18984 1204 19012 1300
rect 20530 1232 20536 1284
rect 20588 1232 20594 1284
rect 18371 1176 19012 1204
rect 20441 1207 20499 1213
rect 18371 1173 18383 1176
rect 18325 1167 18383 1173
rect 20441 1173 20453 1207
rect 20487 1204 20499 1207
rect 20548 1204 20576 1232
rect 20487 1176 20576 1204
rect 22557 1207 22615 1213
rect 20487 1173 20499 1176
rect 20441 1167 20499 1173
rect 22557 1173 22569 1207
rect 22603 1204 22615 1207
rect 23216 1204 23244 1300
rect 24762 1232 24768 1284
rect 24820 1232 24826 1284
rect 22603 1176 23244 1204
rect 24673 1207 24731 1213
rect 22603 1173 22615 1176
rect 22557 1167 22615 1173
rect 24673 1173 24685 1207
rect 24719 1204 24731 1207
rect 24780 1204 24808 1232
rect 24719 1176 24808 1204
rect 26973 1207 27031 1213
rect 24719 1173 24731 1176
rect 24673 1167 24731 1173
rect 26973 1173 26985 1207
rect 27019 1204 27031 1207
rect 27448 1204 27476 1300
rect 28920 1213 28948 1300
rect 27019 1176 27476 1204
rect 28905 1207 28963 1213
rect 27019 1173 27031 1176
rect 26973 1167 27031 1173
rect 28905 1173 28917 1207
rect 28951 1173 28963 1207
rect 28905 1167 28963 1173
rect 31021 1207 31079 1213
rect 31021 1173 31033 1207
rect 31067 1204 31079 1207
rect 31680 1204 31708 1300
rect 31067 1176 31708 1204
rect 33137 1207 33195 1213
rect 31067 1173 31079 1176
rect 31021 1167 31079 1173
rect 33137 1173 33149 1207
rect 33183 1204 33195 1207
rect 34532 1204 34560 1300
rect 35268 1213 35296 1300
rect 33183 1176 34560 1204
rect 35253 1207 35311 1213
rect 33183 1173 33195 1176
rect 33137 1167 33195 1173
rect 35253 1173 35265 1207
rect 35299 1173 35311 1207
rect 35253 1167 35311 1173
rect 37366 1164 37372 1216
rect 37424 1164 37430 1216
rect 40880 1204 40908 1300
rect 41601 1207 41659 1213
rect 41601 1204 41613 1207
rect 40880 1176 41613 1204
rect 41601 1173 41613 1176
rect 41647 1173 41659 1207
rect 41601 1167 41659 1173
rect 1104 1114 44040 1136
rect 1104 1062 11644 1114
rect 11696 1062 11708 1114
rect 11760 1062 11772 1114
rect 11824 1062 11836 1114
rect 11888 1062 11900 1114
rect 11952 1062 22338 1114
rect 22390 1062 22402 1114
rect 22454 1062 22466 1114
rect 22518 1062 22530 1114
rect 22582 1062 22594 1114
rect 22646 1062 33032 1114
rect 33084 1062 33096 1114
rect 33148 1062 33160 1114
rect 33212 1062 33224 1114
rect 33276 1062 33288 1114
rect 33340 1062 43726 1114
rect 43778 1062 43790 1114
rect 43842 1062 43854 1114
rect 43906 1062 43918 1114
rect 43970 1062 43982 1114
rect 44034 1062 44040 1114
rect 1104 1040 44040 1062
rect 14090 960 14096 1012
rect 14148 1000 14154 1012
rect 21726 1000 21732 1012
rect 14148 972 21732 1000
rect 14148 960 14154 972
rect 21726 960 21732 972
rect 21784 960 21790 1012
rect 18138 892 18144 944
rect 18196 932 18202 944
rect 19610 932 19616 944
rect 18196 904 19616 932
rect 18196 892 18202 904
rect 19610 892 19616 904
rect 19668 892 19674 944
<< via1 >>
rect 17592 9936 17644 9988
rect 19064 9936 19116 9988
rect 31668 9936 31720 9988
rect 17684 9868 17736 9920
rect 21456 9868 21508 9920
rect 9036 9732 9088 9784
rect 17040 9664 17092 9716
rect 22928 9800 22980 9852
rect 13176 9528 13228 9580
rect 27344 9732 27396 9784
rect 17592 9664 17644 9716
rect 20536 9664 20588 9716
rect 20720 9664 20772 9716
rect 25596 9664 25648 9716
rect 17408 9596 17460 9648
rect 23204 9596 23256 9648
rect 29276 9596 29328 9648
rect 37556 9596 37608 9648
rect 19616 9528 19668 9580
rect 32864 9528 32916 9580
rect 25412 9460 25464 9512
rect 10416 9392 10468 9444
rect 14372 9392 14424 9444
rect 16028 9392 16080 9444
rect 25688 9392 25740 9444
rect 26792 9392 26844 9444
rect 32036 9392 32088 9444
rect 8300 9324 8352 9376
rect 19984 9324 20036 9376
rect 20168 9324 20220 9376
rect 21272 9324 21324 9376
rect 21364 9324 21416 9376
rect 32772 9324 32824 9376
rect 17040 9256 17092 9308
rect 19064 9256 19116 9308
rect 19156 9256 19208 9308
rect 31392 9256 31444 9308
rect 9956 9188 10008 9240
rect 12072 8916 12124 8968
rect 28172 9188 28224 9240
rect 31484 9188 31536 9240
rect 36636 9188 36688 9240
rect 15108 9120 15160 9172
rect 17408 9120 17460 9172
rect 17592 9120 17644 9172
rect 31116 9120 31168 9172
rect 13452 9052 13504 9104
rect 20720 9052 20772 9104
rect 21456 9052 21508 9104
rect 26792 9052 26844 9104
rect 26884 9052 26936 9104
rect 33600 9120 33652 9172
rect 14648 8984 14700 9036
rect 15844 8984 15896 9036
rect 16580 8984 16632 9036
rect 18696 8984 18748 9036
rect 30564 8984 30616 9036
rect 30656 8984 30708 9036
rect 37464 9052 37516 9104
rect 14924 8916 14976 8968
rect 18420 8916 18472 8968
rect 18972 8916 19024 8968
rect 19064 8916 19116 8968
rect 8208 8848 8260 8900
rect 20720 8848 20772 8900
rect 9864 8780 9916 8832
rect 16580 8780 16632 8832
rect 16764 8780 16816 8832
rect 20168 8780 20220 8832
rect 20536 8780 20588 8832
rect 20996 8780 21048 8832
rect 24584 8916 24636 8968
rect 33692 8984 33744 9036
rect 29000 8848 29052 8900
rect 35256 8848 35308 8900
rect 36084 8848 36136 8900
rect 39028 8848 39080 8900
rect 30288 8780 30340 8832
rect 30380 8780 30432 8832
rect 34980 8780 35032 8832
rect 36820 8780 36872 8832
rect 38660 8780 38712 8832
rect 11644 8678 11696 8730
rect 11708 8678 11760 8730
rect 11772 8678 11824 8730
rect 11836 8678 11888 8730
rect 11900 8678 11952 8730
rect 22338 8678 22390 8730
rect 22402 8678 22454 8730
rect 22466 8678 22518 8730
rect 22530 8678 22582 8730
rect 22594 8678 22646 8730
rect 33032 8678 33084 8730
rect 33096 8678 33148 8730
rect 33160 8678 33212 8730
rect 33224 8678 33276 8730
rect 33288 8678 33340 8730
rect 43726 8678 43778 8730
rect 43790 8678 43842 8730
rect 43854 8678 43906 8730
rect 43918 8678 43970 8730
rect 43982 8678 44034 8730
rect 5356 8576 5408 8628
rect 5908 8576 5960 8628
rect 7012 8576 7064 8628
rect 8208 8576 8260 8628
rect 8668 8576 8720 8628
rect 9496 8576 9548 8628
rect 9772 8619 9824 8628
rect 9772 8585 9781 8619
rect 9781 8585 9815 8619
rect 9815 8585 9824 8619
rect 9772 8576 9824 8585
rect 10600 8576 10652 8628
rect 10876 8576 10928 8628
rect 11428 8576 11480 8628
rect 12440 8576 12492 8628
rect 13176 8576 13228 8628
rect 13636 8576 13688 8628
rect 14188 8576 14240 8628
rect 15016 8576 15068 8628
rect 15292 8619 15344 8628
rect 15292 8585 15301 8619
rect 15301 8585 15335 8619
rect 15335 8585 15344 8619
rect 15292 8576 15344 8585
rect 16120 8576 16172 8628
rect 16488 8576 16540 8628
rect 16764 8576 16816 8628
rect 17224 8576 17276 8628
rect 17500 8576 17552 8628
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 18328 8576 18380 8628
rect 18420 8576 18472 8628
rect 18604 8619 18656 8628
rect 18604 8585 18613 8619
rect 18613 8585 18647 8619
rect 18647 8585 18656 8619
rect 18604 8576 18656 8585
rect 18880 8576 18932 8628
rect 19524 8619 19576 8628
rect 19524 8585 19533 8619
rect 19533 8585 19567 8619
rect 19567 8585 19576 8619
rect 19524 8576 19576 8585
rect 4896 8551 4948 8560
rect 4896 8517 4905 8551
rect 4905 8517 4939 8551
rect 4939 8517 4948 8551
rect 4896 8508 4948 8517
rect 5816 8440 5868 8492
rect 7472 8440 7524 8492
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 8300 8440 8352 8492
rect 8484 8304 8536 8356
rect 10416 8551 10468 8560
rect 10416 8517 10425 8551
rect 10425 8517 10459 8551
rect 10459 8517 10468 8551
rect 10416 8508 10468 8517
rect 12072 8551 12124 8560
rect 12072 8517 12081 8551
rect 12081 8517 12115 8551
rect 12115 8517 12124 8551
rect 12072 8508 12124 8517
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 9864 8440 9916 8492
rect 9956 8483 10008 8492
rect 9956 8449 9965 8483
rect 9965 8449 9999 8483
rect 9999 8449 10008 8483
rect 9956 8440 10008 8449
rect 13452 8508 13504 8560
rect 16028 8508 16080 8560
rect 14372 8440 14424 8492
rect 14924 8440 14976 8492
rect 18144 8508 18196 8560
rect 14832 8372 14884 8424
rect 9404 8304 9456 8356
rect 12440 8304 12492 8356
rect 14648 8304 14700 8356
rect 16764 8483 16816 8492
rect 16764 8449 16773 8483
rect 16773 8449 16807 8483
rect 16807 8449 16816 8483
rect 16764 8440 16816 8449
rect 17500 8440 17552 8492
rect 18328 8440 18380 8492
rect 17132 8304 17184 8356
rect 17408 8372 17460 8424
rect 19340 8508 19392 8560
rect 20168 8576 20220 8628
rect 18696 8440 18748 8492
rect 18880 8440 18932 8492
rect 19524 8440 19576 8492
rect 20076 8440 20128 8492
rect 20536 8440 20588 8492
rect 20812 8483 20864 8492
rect 20812 8449 20821 8483
rect 20821 8449 20855 8483
rect 20855 8449 20864 8483
rect 20812 8440 20864 8449
rect 20628 8372 20680 8424
rect 22100 8508 22152 8560
rect 21088 8483 21140 8492
rect 21088 8449 21097 8483
rect 21097 8449 21131 8483
rect 21131 8449 21140 8483
rect 21088 8440 21140 8449
rect 21364 8483 21416 8492
rect 21364 8449 21373 8483
rect 21373 8449 21407 8483
rect 21407 8449 21416 8483
rect 21364 8440 21416 8449
rect 21640 8483 21692 8492
rect 21640 8449 21649 8483
rect 21649 8449 21683 8483
rect 21683 8449 21692 8483
rect 21640 8440 21692 8449
rect 22008 8440 22060 8492
rect 22560 8576 22612 8628
rect 22928 8576 22980 8628
rect 24768 8576 24820 8628
rect 22652 8508 22704 8560
rect 24400 8508 24452 8560
rect 22468 8483 22520 8492
rect 22468 8449 22477 8483
rect 22477 8449 22511 8483
rect 22511 8449 22520 8483
rect 22468 8440 22520 8449
rect 22744 8483 22796 8492
rect 22744 8449 22753 8483
rect 22753 8449 22787 8483
rect 22787 8449 22796 8483
rect 22744 8440 22796 8449
rect 23020 8483 23072 8492
rect 23020 8449 23029 8483
rect 23029 8449 23063 8483
rect 23063 8449 23072 8483
rect 23020 8440 23072 8449
rect 23112 8440 23164 8492
rect 23572 8483 23624 8492
rect 23572 8449 23581 8483
rect 23581 8449 23615 8483
rect 23615 8449 23624 8483
rect 23572 8440 23624 8449
rect 23848 8483 23900 8492
rect 23848 8449 23857 8483
rect 23857 8449 23891 8483
rect 23891 8449 23900 8483
rect 23848 8440 23900 8449
rect 24124 8483 24176 8492
rect 24124 8449 24133 8483
rect 24133 8449 24167 8483
rect 24167 8449 24176 8483
rect 24124 8440 24176 8449
rect 24308 8440 24360 8492
rect 25504 8576 25556 8628
rect 25228 8508 25280 8560
rect 26332 8576 26384 8628
rect 26148 8508 26200 8560
rect 24952 8372 25004 8424
rect 26056 8440 26108 8492
rect 27160 8576 27212 8628
rect 27068 8508 27120 8560
rect 26884 8440 26936 8492
rect 27988 8576 28040 8628
rect 27804 8508 27856 8560
rect 28264 8576 28316 8628
rect 29092 8576 29144 8628
rect 28908 8508 28960 8560
rect 30288 8619 30340 8628
rect 30288 8585 30297 8619
rect 30297 8585 30331 8619
rect 30331 8585 30340 8619
rect 30288 8576 30340 8585
rect 30472 8576 30524 8628
rect 29644 8508 29696 8560
rect 30196 8508 30248 8560
rect 27528 8372 27580 8424
rect 21640 8304 21692 8356
rect 23296 8304 23348 8356
rect 7380 8236 7432 8288
rect 15108 8236 15160 8288
rect 18512 8236 18564 8288
rect 20352 8236 20404 8288
rect 20444 8236 20496 8288
rect 20904 8279 20956 8288
rect 20904 8245 20913 8279
rect 20913 8245 20947 8279
rect 20947 8245 20956 8279
rect 20904 8236 20956 8245
rect 21088 8236 21140 8288
rect 21456 8279 21508 8288
rect 21456 8245 21465 8279
rect 21465 8245 21499 8279
rect 21499 8245 21508 8279
rect 21456 8236 21508 8245
rect 21732 8236 21784 8288
rect 22192 8236 22244 8288
rect 23020 8236 23072 8288
rect 23112 8279 23164 8288
rect 23112 8245 23121 8279
rect 23121 8245 23155 8279
rect 23155 8245 23164 8279
rect 23112 8236 23164 8245
rect 23388 8279 23440 8288
rect 23388 8245 23397 8279
rect 23397 8245 23431 8279
rect 23431 8245 23440 8279
rect 23388 8236 23440 8245
rect 23664 8279 23716 8288
rect 23664 8245 23673 8279
rect 23673 8245 23707 8279
rect 23707 8245 23716 8279
rect 23664 8236 23716 8245
rect 23940 8279 23992 8288
rect 23940 8245 23949 8279
rect 23949 8245 23983 8279
rect 23983 8245 23992 8279
rect 23940 8236 23992 8245
rect 24400 8279 24452 8288
rect 24400 8245 24409 8279
rect 24409 8245 24443 8279
rect 24443 8245 24452 8279
rect 24400 8236 24452 8245
rect 24492 8236 24544 8288
rect 24860 8236 24912 8288
rect 25044 8236 25096 8288
rect 25320 8236 25372 8288
rect 25780 8279 25832 8288
rect 25780 8245 25789 8279
rect 25789 8245 25823 8279
rect 25823 8245 25832 8279
rect 25780 8236 25832 8245
rect 26056 8279 26108 8288
rect 26056 8245 26065 8279
rect 26065 8245 26099 8279
rect 26099 8245 26108 8279
rect 26056 8236 26108 8245
rect 26332 8279 26384 8288
rect 26332 8245 26341 8279
rect 26341 8245 26375 8279
rect 26375 8245 26384 8279
rect 26332 8236 26384 8245
rect 26608 8279 26660 8288
rect 26608 8245 26617 8279
rect 26617 8245 26651 8279
rect 26651 8245 26660 8279
rect 26608 8236 26660 8245
rect 26976 8279 27028 8288
rect 26976 8245 26985 8279
rect 26985 8245 27019 8279
rect 27019 8245 27028 8279
rect 26976 8236 27028 8245
rect 27252 8279 27304 8288
rect 27252 8245 27261 8279
rect 27261 8245 27295 8279
rect 27295 8245 27304 8279
rect 27252 8236 27304 8245
rect 27528 8279 27580 8288
rect 27528 8245 27537 8279
rect 27537 8245 27571 8279
rect 27571 8245 27580 8279
rect 27528 8236 27580 8245
rect 27988 8236 28040 8288
rect 28172 8236 28224 8288
rect 28356 8279 28408 8288
rect 28356 8245 28365 8279
rect 28365 8245 28399 8279
rect 28399 8245 28408 8279
rect 28356 8236 28408 8245
rect 28448 8236 28500 8288
rect 29552 8372 29604 8424
rect 29920 8372 29972 8424
rect 30564 8440 30616 8492
rect 31116 8619 31168 8628
rect 31116 8585 31125 8619
rect 31125 8585 31159 8619
rect 31159 8585 31168 8619
rect 31116 8576 31168 8585
rect 31392 8619 31444 8628
rect 31392 8585 31401 8619
rect 31401 8585 31435 8619
rect 31435 8585 31444 8619
rect 31392 8576 31444 8585
rect 31668 8619 31720 8628
rect 31668 8585 31677 8619
rect 31677 8585 31711 8619
rect 31711 8585 31720 8619
rect 31668 8576 31720 8585
rect 31852 8576 31904 8628
rect 31024 8508 31076 8560
rect 31576 8508 31628 8560
rect 28816 8304 28868 8356
rect 28908 8347 28960 8356
rect 28908 8313 28917 8347
rect 28917 8313 28951 8347
rect 28951 8313 28960 8347
rect 28908 8304 28960 8313
rect 30748 8372 30800 8424
rect 31300 8372 31352 8424
rect 32036 8440 32088 8492
rect 32220 8508 32272 8560
rect 30840 8347 30892 8356
rect 30840 8313 30849 8347
rect 30849 8313 30883 8347
rect 30883 8313 30892 8347
rect 30840 8304 30892 8313
rect 31944 8347 31996 8356
rect 31944 8313 31953 8347
rect 31953 8313 31987 8347
rect 31987 8313 31996 8347
rect 31944 8304 31996 8313
rect 32680 8576 32732 8628
rect 32588 8508 32640 8560
rect 32312 8372 32364 8424
rect 32772 8440 32824 8492
rect 33692 8619 33744 8628
rect 33692 8585 33701 8619
rect 33701 8585 33735 8619
rect 33735 8585 33744 8619
rect 33692 8576 33744 8585
rect 34060 8576 34112 8628
rect 34428 8576 34480 8628
rect 35164 8576 35216 8628
rect 33416 8508 33468 8560
rect 33324 8440 33376 8492
rect 35440 8508 35492 8560
rect 36636 8576 36688 8628
rect 37464 8576 37516 8628
rect 37556 8576 37608 8628
rect 34152 8483 34204 8492
rect 34152 8449 34161 8483
rect 34161 8449 34195 8483
rect 34195 8449 34204 8483
rect 34152 8440 34204 8449
rect 35256 8483 35308 8492
rect 35256 8449 35265 8483
rect 35265 8449 35299 8483
rect 35299 8449 35308 8483
rect 35256 8440 35308 8449
rect 29552 8279 29604 8288
rect 29552 8245 29561 8279
rect 29561 8245 29595 8279
rect 29595 8245 29604 8279
rect 29552 8236 29604 8245
rect 29828 8279 29880 8288
rect 29828 8245 29837 8279
rect 29837 8245 29871 8279
rect 29871 8245 29880 8279
rect 29828 8236 29880 8245
rect 32864 8347 32916 8356
rect 32864 8313 32873 8347
rect 32873 8313 32907 8347
rect 32907 8313 32916 8347
rect 32864 8304 32916 8313
rect 33232 8304 33284 8356
rect 34980 8372 35032 8424
rect 36452 8483 36504 8492
rect 36452 8449 36461 8483
rect 36461 8449 36495 8483
rect 36495 8449 36504 8483
rect 36452 8440 36504 8449
rect 37648 8440 37700 8492
rect 39304 8576 39356 8628
rect 38660 8508 38712 8560
rect 39212 8508 39264 8560
rect 39028 8483 39080 8492
rect 39028 8449 39037 8483
rect 39037 8449 39071 8483
rect 39071 8449 39080 8483
rect 39028 8440 39080 8449
rect 39304 8440 39356 8492
rect 40500 8483 40552 8492
rect 40500 8449 40509 8483
rect 40509 8449 40543 8483
rect 40543 8449 40552 8483
rect 40500 8440 40552 8449
rect 41052 8483 41104 8492
rect 41052 8449 41061 8483
rect 41061 8449 41095 8483
rect 41095 8449 41104 8483
rect 41052 8440 41104 8449
rect 36544 8372 36596 8424
rect 33692 8304 33744 8356
rect 33968 8347 34020 8356
rect 33968 8313 33977 8347
rect 33977 8313 34011 8347
rect 34011 8313 34020 8347
rect 33968 8304 34020 8313
rect 34612 8304 34664 8356
rect 35716 8304 35768 8356
rect 38016 8236 38068 8288
rect 6297 8134 6349 8186
rect 6361 8134 6413 8186
rect 6425 8134 6477 8186
rect 6489 8134 6541 8186
rect 6553 8134 6605 8186
rect 16991 8134 17043 8186
rect 17055 8134 17107 8186
rect 17119 8134 17171 8186
rect 17183 8134 17235 8186
rect 17247 8134 17299 8186
rect 27685 8134 27737 8186
rect 27749 8134 27801 8186
rect 27813 8134 27865 8186
rect 27877 8134 27929 8186
rect 27941 8134 27993 8186
rect 38379 8134 38431 8186
rect 38443 8134 38495 8186
rect 38507 8134 38559 8186
rect 38571 8134 38623 8186
rect 38635 8134 38687 8186
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 6184 8032 6236 8084
rect 7564 8075 7616 8084
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 7932 8075 7984 8084
rect 7932 8041 7941 8075
rect 7941 8041 7975 8075
rect 7975 8041 7984 8075
rect 7932 8032 7984 8041
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 9312 8075 9364 8084
rect 9312 8041 9321 8075
rect 9321 8041 9355 8075
rect 9355 8041 9364 8075
rect 9312 8032 9364 8041
rect 10140 8075 10192 8084
rect 10140 8041 10149 8075
rect 10149 8041 10183 8075
rect 10183 8041 10192 8075
rect 10140 8032 10192 8041
rect 11244 8075 11296 8084
rect 11244 8041 11253 8075
rect 11253 8041 11287 8075
rect 11287 8041 11296 8075
rect 11244 8032 11296 8041
rect 11520 8032 11572 8084
rect 6920 8007 6972 8016
rect 6920 7973 6929 8007
rect 6929 7973 6963 8007
rect 6963 7973 6972 8007
rect 6920 7964 6972 7973
rect 6736 7803 6788 7812
rect 6736 7769 6745 7803
rect 6745 7769 6779 7803
rect 6779 7769 6788 7803
rect 6736 7760 6788 7769
rect 8208 7828 8260 7880
rect 12440 8007 12492 8016
rect 12440 7973 12449 8007
rect 12449 7973 12483 8007
rect 12483 7973 12492 8007
rect 12440 7964 12492 7973
rect 13360 8032 13412 8084
rect 13912 8032 13964 8084
rect 14556 8075 14608 8084
rect 14556 8041 14565 8075
rect 14565 8041 14599 8075
rect 14599 8041 14608 8075
rect 14556 8032 14608 8041
rect 14740 8032 14792 8084
rect 15660 8075 15712 8084
rect 15660 8041 15669 8075
rect 15669 8041 15703 8075
rect 15703 8041 15712 8075
rect 15660 8032 15712 8041
rect 16580 8007 16632 8016
rect 16580 7973 16589 8007
rect 16589 7973 16623 8007
rect 16623 7973 16632 8007
rect 16580 7964 16632 7973
rect 16856 8032 16908 8084
rect 17408 8075 17460 8084
rect 17408 8041 17417 8075
rect 17417 8041 17451 8075
rect 17451 8041 17460 8075
rect 17408 8032 17460 8041
rect 18788 8032 18840 8084
rect 18880 8075 18932 8084
rect 18880 8041 18889 8075
rect 18889 8041 18923 8075
rect 18923 8041 18932 8075
rect 18880 8032 18932 8041
rect 19984 8032 20036 8084
rect 20996 8032 21048 8084
rect 21364 8075 21416 8084
rect 21364 8041 21373 8075
rect 21373 8041 21407 8075
rect 21407 8041 21416 8075
rect 21364 8032 21416 8041
rect 21456 8032 21508 8084
rect 17960 8007 18012 8016
rect 17960 7973 17969 8007
rect 17969 7973 18003 8007
rect 18003 7973 18012 8007
rect 17960 7964 18012 7973
rect 18328 8007 18380 8016
rect 18328 7973 18337 8007
rect 18337 7973 18371 8007
rect 18371 7973 18380 8007
rect 18328 7964 18380 7973
rect 7748 7760 7800 7812
rect 8392 7803 8444 7812
rect 8392 7769 8401 7803
rect 8401 7769 8435 7803
rect 8435 7769 8444 7803
rect 8392 7760 8444 7769
rect 9220 7803 9272 7812
rect 9220 7769 9229 7803
rect 9229 7769 9263 7803
rect 9263 7769 9272 7803
rect 9220 7760 9272 7769
rect 10048 7803 10100 7812
rect 10048 7769 10057 7803
rect 10057 7769 10091 7803
rect 10091 7769 10100 7803
rect 10048 7760 10100 7769
rect 9588 7692 9640 7744
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 14924 7871 14976 7880
rect 14924 7837 14933 7871
rect 14933 7837 14967 7871
rect 14967 7837 14976 7871
rect 14924 7828 14976 7837
rect 12256 7803 12308 7812
rect 12256 7769 12265 7803
rect 12265 7769 12299 7803
rect 12299 7769 12308 7803
rect 12256 7760 12308 7769
rect 13728 7692 13780 7744
rect 16672 7828 16724 7880
rect 15476 7692 15528 7744
rect 16396 7803 16448 7812
rect 16396 7769 16405 7803
rect 16405 7769 16439 7803
rect 16439 7769 16448 7803
rect 16396 7760 16448 7769
rect 19616 7964 19668 8016
rect 17592 7871 17644 7880
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 17960 7828 18012 7880
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 18972 7828 19024 7880
rect 19064 7871 19116 7880
rect 19064 7837 19073 7871
rect 19073 7837 19107 7871
rect 19107 7837 19116 7871
rect 19064 7828 19116 7837
rect 17776 7803 17828 7812
rect 17776 7769 17785 7803
rect 17785 7769 17819 7803
rect 17819 7769 17828 7803
rect 17776 7760 17828 7769
rect 21824 7964 21876 8016
rect 23020 8032 23072 8084
rect 23664 8032 23716 8084
rect 24400 8032 24452 8084
rect 24676 8032 24728 8084
rect 25412 8075 25464 8084
rect 25412 8041 25421 8075
rect 25421 8041 25455 8075
rect 25455 8041 25464 8075
rect 25412 8032 25464 8041
rect 25504 8032 25556 8084
rect 25872 8032 25924 8084
rect 27160 8032 27212 8084
rect 27712 8032 27764 8084
rect 28264 8032 28316 8084
rect 28448 8032 28500 8084
rect 34888 8032 34940 8084
rect 35992 8032 36044 8084
rect 36360 8032 36412 8084
rect 37372 8032 37424 8084
rect 22560 7964 22612 8016
rect 22652 8007 22704 8016
rect 22652 7973 22661 8007
rect 22661 7973 22695 8007
rect 22695 7973 22704 8007
rect 22652 7964 22704 7973
rect 19892 7871 19944 7880
rect 19892 7837 19901 7871
rect 19901 7837 19935 7871
rect 19935 7837 19944 7871
rect 19892 7828 19944 7837
rect 20444 7828 20496 7880
rect 20996 7871 21048 7880
rect 20996 7837 21005 7871
rect 21005 7837 21039 7871
rect 21039 7837 21048 7871
rect 20996 7828 21048 7837
rect 21088 7871 21140 7880
rect 21088 7837 21097 7871
rect 21097 7837 21131 7871
rect 21131 7837 21140 7871
rect 21088 7828 21140 7837
rect 21548 7871 21600 7880
rect 21548 7837 21557 7871
rect 21557 7837 21591 7871
rect 21591 7837 21600 7871
rect 21548 7828 21600 7837
rect 21640 7871 21692 7880
rect 21640 7837 21649 7871
rect 21649 7837 21683 7871
rect 21683 7837 21692 7871
rect 21640 7828 21692 7837
rect 19524 7692 19576 7744
rect 20628 7760 20680 7812
rect 22652 7828 22704 7880
rect 24032 8007 24084 8016
rect 24032 7973 24041 8007
rect 24041 7973 24075 8007
rect 24075 7973 24084 8007
rect 24032 7964 24084 7973
rect 23112 7828 23164 7880
rect 23296 7871 23348 7880
rect 23296 7837 23297 7871
rect 23297 7837 23331 7871
rect 23331 7837 23348 7871
rect 23296 7828 23348 7837
rect 24308 7828 24360 7880
rect 24492 7828 24544 7880
rect 24860 7828 24912 7880
rect 25044 7828 25096 7880
rect 25320 7828 25372 7880
rect 37280 7964 37332 8016
rect 38752 8075 38804 8084
rect 38752 8041 38761 8075
rect 38761 8041 38795 8075
rect 38795 8041 38804 8075
rect 38752 8032 38804 8041
rect 38844 8032 38896 8084
rect 40040 8032 40092 8084
rect 25596 7896 25648 7948
rect 25780 7871 25832 7880
rect 25780 7837 25789 7871
rect 25789 7837 25823 7871
rect 25823 7837 25832 7871
rect 25780 7828 25832 7837
rect 26056 7871 26108 7880
rect 26056 7837 26065 7871
rect 26065 7837 26099 7871
rect 26099 7837 26108 7871
rect 26056 7828 26108 7837
rect 26332 7871 26384 7880
rect 26332 7837 26341 7871
rect 26341 7837 26375 7871
rect 26375 7837 26384 7871
rect 26332 7828 26384 7837
rect 26608 7871 26660 7880
rect 26608 7837 26617 7871
rect 26617 7837 26651 7871
rect 26651 7837 26660 7871
rect 26608 7828 26660 7837
rect 26976 7828 27028 7880
rect 20536 7692 20588 7744
rect 21088 7692 21140 7744
rect 21272 7735 21324 7744
rect 21272 7701 21281 7735
rect 21281 7701 21315 7735
rect 21315 7701 21324 7735
rect 21272 7692 21324 7701
rect 21364 7692 21416 7744
rect 22100 7735 22152 7744
rect 22100 7701 22109 7735
rect 22109 7701 22143 7735
rect 22143 7701 22152 7735
rect 22100 7692 22152 7701
rect 22836 7692 22888 7744
rect 23296 7692 23348 7744
rect 23756 7735 23808 7744
rect 23756 7701 23765 7735
rect 23765 7701 23799 7735
rect 23799 7701 23808 7735
rect 23756 7692 23808 7701
rect 26148 7760 26200 7812
rect 24492 7692 24544 7744
rect 24860 7735 24912 7744
rect 24860 7701 24869 7735
rect 24869 7701 24903 7735
rect 24903 7701 24912 7735
rect 24860 7692 24912 7701
rect 25136 7735 25188 7744
rect 25136 7701 25145 7735
rect 25145 7701 25179 7735
rect 25179 7701 25188 7735
rect 25136 7692 25188 7701
rect 25964 7735 26016 7744
rect 25964 7701 25973 7735
rect 25973 7701 26007 7735
rect 26007 7701 26016 7735
rect 25964 7692 26016 7701
rect 26240 7735 26292 7744
rect 26240 7701 26249 7735
rect 26249 7701 26283 7735
rect 26283 7701 26292 7735
rect 26240 7692 26292 7701
rect 27252 7828 27304 7880
rect 27344 7828 27396 7880
rect 27528 7828 27580 7880
rect 28172 7896 28224 7948
rect 34612 7896 34664 7948
rect 28080 7828 28132 7880
rect 28264 7828 28316 7880
rect 28908 7828 28960 7880
rect 33600 7871 33652 7880
rect 33600 7837 33609 7871
rect 33609 7837 33643 7871
rect 33643 7837 33652 7871
rect 33600 7828 33652 7837
rect 33876 7871 33928 7880
rect 33876 7837 33885 7871
rect 33885 7837 33919 7871
rect 33919 7837 33928 7871
rect 33876 7828 33928 7837
rect 35440 7871 35492 7880
rect 35440 7837 35449 7871
rect 35449 7837 35483 7871
rect 35483 7837 35492 7871
rect 35440 7828 35492 7837
rect 36268 7896 36320 7948
rect 34520 7760 34572 7812
rect 33784 7735 33836 7744
rect 33784 7701 33793 7735
rect 33793 7701 33827 7735
rect 33827 7701 33836 7735
rect 33784 7692 33836 7701
rect 34060 7735 34112 7744
rect 34060 7701 34069 7735
rect 34069 7701 34103 7735
rect 34103 7701 34112 7735
rect 34060 7692 34112 7701
rect 35992 7760 36044 7812
rect 38200 7828 38252 7880
rect 38292 7760 38344 7812
rect 39856 7828 39908 7880
rect 37464 7692 37516 7744
rect 39396 7692 39448 7744
rect 11644 7590 11696 7642
rect 11708 7590 11760 7642
rect 11772 7590 11824 7642
rect 11836 7590 11888 7642
rect 11900 7590 11952 7642
rect 22338 7590 22390 7642
rect 22402 7590 22454 7642
rect 22466 7590 22518 7642
rect 22530 7590 22582 7642
rect 22594 7590 22646 7642
rect 33032 7590 33084 7642
rect 33096 7590 33148 7642
rect 33160 7590 33212 7642
rect 33224 7590 33276 7642
rect 33288 7590 33340 7642
rect 43726 7590 43778 7642
rect 43790 7590 43842 7642
rect 43854 7590 43906 7642
rect 43918 7590 43970 7642
rect 43982 7590 44034 7642
rect 5816 7488 5868 7540
rect 6644 7488 6696 7540
rect 7288 7488 7340 7540
rect 8024 7531 8076 7540
rect 8024 7497 8033 7531
rect 8033 7497 8067 7531
rect 8067 7497 8076 7531
rect 8024 7488 8076 7497
rect 11980 7531 12032 7540
rect 11980 7497 11989 7531
rect 11989 7497 12023 7531
rect 12023 7497 12032 7531
rect 11980 7488 12032 7497
rect 13084 7488 13136 7540
rect 14924 7488 14976 7540
rect 6552 7463 6604 7472
rect 6552 7429 6561 7463
rect 6561 7429 6595 7463
rect 6595 7429 6604 7463
rect 6552 7420 6604 7429
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 15108 7420 15160 7472
rect 12716 7395 12768 7404
rect 12716 7361 12725 7395
rect 12725 7361 12759 7395
rect 12759 7361 12768 7395
rect 12716 7352 12768 7361
rect 16396 7488 16448 7540
rect 17500 7531 17552 7540
rect 17500 7497 17509 7531
rect 17509 7497 17543 7531
rect 17543 7497 17552 7531
rect 17500 7488 17552 7497
rect 17776 7488 17828 7540
rect 18328 7488 18380 7540
rect 18420 7488 18472 7540
rect 19892 7531 19944 7540
rect 19892 7497 19901 7531
rect 19901 7497 19935 7531
rect 19935 7497 19944 7531
rect 19892 7488 19944 7497
rect 20904 7488 20956 7540
rect 20996 7488 21048 7540
rect 17592 7352 17644 7404
rect 17868 7352 17920 7404
rect 18144 7352 18196 7404
rect 8116 7284 8168 7336
rect 9220 7284 9272 7336
rect 16488 7284 16540 7336
rect 18512 7352 18564 7404
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 19064 7352 19116 7404
rect 19156 7395 19208 7404
rect 19156 7361 19165 7395
rect 19165 7361 19199 7395
rect 19199 7361 19208 7395
rect 19156 7352 19208 7361
rect 19340 7352 19392 7404
rect 19524 7352 19576 7404
rect 8392 7216 8444 7268
rect 15568 7216 15620 7268
rect 7748 7148 7800 7200
rect 19616 7259 19668 7268
rect 19616 7225 19625 7259
rect 19625 7225 19659 7259
rect 19659 7225 19668 7259
rect 19616 7216 19668 7225
rect 16764 7148 16816 7200
rect 18052 7148 18104 7200
rect 18604 7148 18656 7200
rect 19248 7148 19300 7200
rect 20260 7352 20312 7404
rect 21088 7420 21140 7472
rect 21916 7420 21968 7472
rect 23204 7488 23256 7540
rect 23388 7488 23440 7540
rect 23480 7531 23532 7540
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 23480 7488 23532 7497
rect 23940 7488 23992 7540
rect 24308 7488 24360 7540
rect 28264 7488 28316 7540
rect 21732 7352 21784 7404
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 22468 7352 22520 7404
rect 21088 7259 21140 7268
rect 21088 7225 21097 7259
rect 21097 7225 21131 7259
rect 21131 7225 21140 7259
rect 21088 7216 21140 7225
rect 21548 7284 21600 7336
rect 22376 7284 22428 7336
rect 24492 7420 24544 7472
rect 29552 7488 29604 7540
rect 33784 7488 33836 7540
rect 34060 7488 34112 7540
rect 28356 7352 28408 7404
rect 22192 7216 22244 7268
rect 22468 7216 22520 7268
rect 22560 7216 22612 7268
rect 37280 7284 37332 7336
rect 38292 7284 38344 7336
rect 20168 7191 20220 7200
rect 20168 7157 20177 7191
rect 20177 7157 20211 7191
rect 20211 7157 20220 7191
rect 20168 7148 20220 7157
rect 20996 7191 21048 7200
rect 20996 7157 21005 7191
rect 21005 7157 21039 7191
rect 21039 7157 21048 7191
rect 20996 7148 21048 7157
rect 21456 7148 21508 7200
rect 24584 7148 24636 7200
rect 24860 7148 24912 7200
rect 6297 7046 6349 7098
rect 6361 7046 6413 7098
rect 6425 7046 6477 7098
rect 6489 7046 6541 7098
rect 6553 7046 6605 7098
rect 16991 7046 17043 7098
rect 17055 7046 17107 7098
rect 17119 7046 17171 7098
rect 17183 7046 17235 7098
rect 17247 7046 17299 7098
rect 27685 7046 27737 7098
rect 27749 7046 27801 7098
rect 27813 7046 27865 7098
rect 27877 7046 27929 7098
rect 27941 7046 27993 7098
rect 38379 7046 38431 7098
rect 38443 7046 38495 7098
rect 38507 7046 38559 7098
rect 38571 7046 38623 7098
rect 38635 7046 38687 7098
rect 10048 6944 10100 6996
rect 19524 6944 19576 6996
rect 20996 6944 21048 6996
rect 21272 6944 21324 6996
rect 9404 6808 9456 6860
rect 10324 6808 10376 6860
rect 16488 6808 16540 6860
rect 21456 6876 21508 6928
rect 23296 6944 23348 6996
rect 29828 6944 29880 6996
rect 22744 6876 22796 6928
rect 21916 6808 21968 6860
rect 25136 6808 25188 6860
rect 38108 6808 38160 6860
rect 39396 6808 39448 6860
rect 7472 6740 7524 6792
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 19156 6740 19208 6792
rect 19984 6783 20036 6792
rect 19984 6749 19993 6783
rect 19993 6749 20027 6783
rect 20027 6749 20036 6783
rect 19984 6740 20036 6749
rect 20260 6783 20312 6792
rect 20260 6749 20269 6783
rect 20269 6749 20303 6783
rect 20303 6749 20312 6783
rect 20260 6740 20312 6749
rect 21088 6740 21140 6792
rect 18696 6672 18748 6724
rect 19340 6672 19392 6724
rect 11644 6502 11696 6554
rect 11708 6502 11760 6554
rect 11772 6502 11824 6554
rect 11836 6502 11888 6554
rect 11900 6502 11952 6554
rect 22338 6502 22390 6554
rect 22402 6502 22454 6554
rect 22466 6502 22518 6554
rect 22530 6502 22582 6554
rect 22594 6502 22646 6554
rect 33032 6502 33084 6554
rect 33096 6502 33148 6554
rect 33160 6502 33212 6554
rect 33224 6502 33276 6554
rect 33288 6502 33340 6554
rect 43726 6502 43778 6554
rect 43790 6502 43842 6554
rect 43854 6502 43906 6554
rect 43918 6502 43970 6554
rect 43982 6502 44034 6554
rect 5908 6400 5960 6452
rect 13728 6400 13780 6452
rect 21824 6400 21876 6452
rect 21916 6332 21968 6384
rect 17592 6264 17644 6316
rect 25964 6264 26016 6316
rect 12256 6196 12308 6248
rect 15476 6196 15528 6248
rect 26148 6196 26200 6248
rect 16672 6128 16724 6180
rect 26240 6128 26292 6180
rect 17316 6060 17368 6112
rect 6297 5958 6349 6010
rect 6361 5958 6413 6010
rect 6425 5958 6477 6010
rect 6489 5958 6541 6010
rect 6553 5958 6605 6010
rect 16991 5958 17043 6010
rect 17055 5958 17107 6010
rect 17119 5958 17171 6010
rect 17183 5958 17235 6010
rect 17247 5958 17299 6010
rect 27685 5958 27737 6010
rect 27749 5958 27801 6010
rect 27813 5958 27865 6010
rect 27877 5958 27929 6010
rect 27941 5958 27993 6010
rect 38379 5958 38431 6010
rect 38443 5958 38495 6010
rect 38507 5958 38559 6010
rect 38571 5958 38623 6010
rect 38635 5958 38687 6010
rect 18788 5856 18840 5908
rect 30840 5856 30892 5908
rect 17316 5788 17368 5840
rect 24860 5788 24912 5840
rect 22744 5584 22796 5636
rect 29000 5584 29052 5636
rect 11644 5414 11696 5466
rect 11708 5414 11760 5466
rect 11772 5414 11824 5466
rect 11836 5414 11888 5466
rect 11900 5414 11952 5466
rect 22338 5414 22390 5466
rect 22402 5414 22454 5466
rect 22466 5414 22518 5466
rect 22530 5414 22582 5466
rect 22594 5414 22646 5466
rect 33032 5414 33084 5466
rect 33096 5414 33148 5466
rect 33160 5414 33212 5466
rect 33224 5414 33276 5466
rect 33288 5414 33340 5466
rect 43726 5414 43778 5466
rect 43790 5414 43842 5466
rect 43854 5414 43906 5466
rect 43918 5414 43970 5466
rect 43982 5414 44034 5466
rect 37464 5355 37516 5364
rect 37464 5321 37473 5355
rect 37473 5321 37507 5355
rect 37507 5321 37516 5355
rect 37464 5312 37516 5321
rect 37648 5219 37700 5228
rect 37648 5185 37657 5219
rect 37657 5185 37691 5219
rect 37691 5185 37700 5219
rect 37648 5176 37700 5185
rect 25964 5108 26016 5160
rect 30656 5108 30708 5160
rect 26056 4972 26108 5024
rect 36268 4972 36320 5024
rect 6297 4870 6349 4922
rect 6361 4870 6413 4922
rect 6425 4870 6477 4922
rect 6489 4870 6541 4922
rect 6553 4870 6605 4922
rect 16991 4870 17043 4922
rect 17055 4870 17107 4922
rect 17119 4870 17171 4922
rect 17183 4870 17235 4922
rect 17247 4870 17299 4922
rect 27685 4870 27737 4922
rect 27749 4870 27801 4922
rect 27813 4870 27865 4922
rect 27877 4870 27929 4922
rect 27941 4870 27993 4922
rect 38379 4870 38431 4922
rect 38443 4870 38495 4922
rect 38507 4870 38559 4922
rect 38571 4870 38623 4922
rect 38635 4870 38687 4922
rect 22744 4811 22796 4820
rect 22744 4777 22753 4811
rect 22753 4777 22787 4811
rect 22787 4777 22796 4811
rect 22744 4768 22796 4777
rect 25964 4768 26016 4820
rect 26056 4811 26108 4820
rect 26056 4777 26065 4811
rect 26065 4777 26099 4811
rect 26099 4777 26108 4811
rect 26056 4768 26108 4777
rect 34520 4768 34572 4820
rect 37648 4768 37700 4820
rect 38200 4811 38252 4820
rect 38200 4777 38209 4811
rect 38209 4777 38243 4811
rect 38243 4777 38252 4811
rect 38200 4768 38252 4777
rect 21640 4607 21692 4616
rect 21640 4573 21649 4607
rect 21649 4573 21683 4607
rect 21683 4573 21692 4607
rect 21640 4564 21692 4573
rect 22192 4564 22244 4616
rect 22744 4564 22796 4616
rect 23112 4607 23164 4616
rect 23112 4573 23121 4607
rect 23121 4573 23155 4607
rect 23155 4573 23164 4607
rect 23112 4564 23164 4573
rect 30380 4632 30432 4684
rect 39304 4700 39356 4752
rect 35440 4632 35492 4684
rect 23388 4607 23440 4616
rect 23388 4573 23397 4607
rect 23397 4573 23431 4607
rect 23431 4573 23440 4607
rect 23388 4564 23440 4573
rect 25872 4607 25924 4616
rect 25872 4573 25881 4607
rect 25881 4573 25915 4607
rect 25915 4573 25924 4607
rect 25872 4564 25924 4573
rect 27988 4607 28040 4616
rect 27988 4573 27997 4607
rect 27997 4573 28031 4607
rect 28031 4573 28040 4607
rect 27988 4564 28040 4573
rect 32220 4607 32272 4616
rect 32220 4573 32229 4607
rect 32229 4573 32263 4607
rect 32263 4573 32272 4607
rect 32220 4564 32272 4573
rect 34520 4564 34572 4616
rect 38384 4607 38436 4616
rect 38384 4573 38393 4607
rect 38393 4573 38427 4607
rect 38427 4573 38436 4607
rect 38384 4564 38436 4573
rect 36452 4496 36504 4548
rect 11644 4326 11696 4378
rect 11708 4326 11760 4378
rect 11772 4326 11824 4378
rect 11836 4326 11888 4378
rect 11900 4326 11952 4378
rect 22338 4326 22390 4378
rect 22402 4326 22454 4378
rect 22466 4326 22518 4378
rect 22530 4326 22582 4378
rect 22594 4326 22646 4378
rect 33032 4326 33084 4378
rect 33096 4326 33148 4378
rect 33160 4326 33212 4378
rect 33224 4326 33276 4378
rect 33288 4326 33340 4378
rect 43726 4326 43778 4378
rect 43790 4326 43842 4378
rect 43854 4326 43906 4378
rect 43918 4326 43970 4378
rect 43982 4326 44034 4378
rect 21640 4224 21692 4276
rect 23388 4224 23440 4276
rect 25872 4224 25924 4276
rect 38384 4224 38436 4276
rect 22744 4156 22796 4208
rect 20536 4088 20588 4140
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 7932 4020 7984 4072
rect 22192 3952 22244 4004
rect 22836 4131 22888 4140
rect 22836 4097 22845 4131
rect 22845 4097 22879 4131
rect 22879 4097 22888 4131
rect 22836 4088 22888 4097
rect 23756 4131 23808 4140
rect 23756 4097 23765 4131
rect 23765 4097 23799 4131
rect 23799 4097 23808 4131
rect 23756 4088 23808 4097
rect 24768 4088 24820 4140
rect 27436 4131 27488 4140
rect 27436 4097 27445 4131
rect 27445 4097 27479 4131
rect 27479 4097 27488 4131
rect 27436 4088 27488 4097
rect 31668 4131 31720 4140
rect 31668 4097 31677 4131
rect 31677 4097 31711 4131
rect 31711 4097 31720 4131
rect 31668 4088 31720 4097
rect 37372 4088 37424 4140
rect 27988 4020 28040 4072
rect 32220 4020 32272 4072
rect 18236 3884 18288 3936
rect 23112 3952 23164 4004
rect 29276 3952 29328 4004
rect 6297 3782 6349 3834
rect 6361 3782 6413 3834
rect 6425 3782 6477 3834
rect 6489 3782 6541 3834
rect 6553 3782 6605 3834
rect 16991 3782 17043 3834
rect 17055 3782 17107 3834
rect 17119 3782 17171 3834
rect 17183 3782 17235 3834
rect 17247 3782 17299 3834
rect 27685 3782 27737 3834
rect 27749 3782 27801 3834
rect 27813 3782 27865 3834
rect 27877 3782 27929 3834
rect 27941 3782 27993 3834
rect 38379 3782 38431 3834
rect 38443 3782 38495 3834
rect 38507 3782 38559 3834
rect 38571 3782 38623 3834
rect 38635 3782 38687 3834
rect 5816 3612 5868 3664
rect 22008 3680 22060 3732
rect 23756 3680 23808 3732
rect 36084 3680 36136 3732
rect 37280 3723 37332 3732
rect 37280 3689 37289 3723
rect 37289 3689 37323 3723
rect 37323 3689 37332 3723
rect 37280 3680 37332 3689
rect 41052 3680 41104 3732
rect 34612 3612 34664 3664
rect 19616 3544 19668 3596
rect 22836 3544 22888 3596
rect 19524 3519 19576 3528
rect 19524 3485 19533 3519
rect 19533 3485 19567 3519
rect 19567 3485 19576 3519
rect 19524 3476 19576 3485
rect 23204 3519 23256 3528
rect 23204 3485 23213 3519
rect 23213 3485 23247 3519
rect 23247 3485 23256 3519
rect 23204 3476 23256 3485
rect 30104 3519 30156 3528
rect 30104 3485 30113 3519
rect 30113 3485 30147 3519
rect 30147 3485 30156 3519
rect 30104 3476 30156 3485
rect 37464 3519 37516 3528
rect 37464 3485 37473 3519
rect 37473 3485 37507 3519
rect 37507 3485 37516 3519
rect 37464 3476 37516 3485
rect 40132 3519 40184 3528
rect 40132 3485 40141 3519
rect 40141 3485 40175 3519
rect 40175 3485 40184 3519
rect 40132 3476 40184 3485
rect 11644 3238 11696 3290
rect 11708 3238 11760 3290
rect 11772 3238 11824 3290
rect 11836 3238 11888 3290
rect 11900 3238 11952 3290
rect 22338 3238 22390 3290
rect 22402 3238 22454 3290
rect 22466 3238 22518 3290
rect 22530 3238 22582 3290
rect 22594 3238 22646 3290
rect 33032 3238 33084 3290
rect 33096 3238 33148 3290
rect 33160 3238 33212 3290
rect 33224 3238 33276 3290
rect 33288 3238 33340 3290
rect 43726 3238 43778 3290
rect 43790 3238 43842 3290
rect 43854 3238 43906 3290
rect 43918 3238 43970 3290
rect 43982 3238 44034 3290
rect 19524 3136 19576 3188
rect 30104 3136 30156 3188
rect 31484 3136 31536 3188
rect 37464 3136 37516 3188
rect 40132 3136 40184 3188
rect 18972 3043 19024 3052
rect 18972 3009 18981 3043
rect 18981 3009 19015 3043
rect 19015 3009 19024 3043
rect 18972 3000 19024 3009
rect 22008 3043 22060 3052
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 22376 3043 22428 3052
rect 22376 3009 22385 3043
rect 22385 3009 22419 3043
rect 22419 3009 22428 3043
rect 22376 3000 22428 3009
rect 28908 3000 28960 3052
rect 35256 3000 35308 3052
rect 40868 3043 40920 3052
rect 40868 3009 40877 3043
rect 40877 3009 40911 3043
rect 40911 3009 40920 3043
rect 40868 3000 40920 3009
rect 35992 2932 36044 2984
rect 6297 2694 6349 2746
rect 6361 2694 6413 2746
rect 6425 2694 6477 2746
rect 6489 2694 6541 2746
rect 6553 2694 6605 2746
rect 16991 2694 17043 2746
rect 17055 2694 17107 2746
rect 17119 2694 17171 2746
rect 17183 2694 17235 2746
rect 17247 2694 17299 2746
rect 27685 2694 27737 2746
rect 27749 2694 27801 2746
rect 27813 2694 27865 2746
rect 27877 2694 27929 2746
rect 27941 2694 27993 2746
rect 38379 2694 38431 2746
rect 38443 2694 38495 2746
rect 38507 2694 38559 2746
rect 38571 2694 38623 2746
rect 38635 2694 38687 2746
rect 22008 2592 22060 2644
rect 22376 2592 22428 2644
rect 39856 2635 39908 2644
rect 39856 2601 39865 2635
rect 39865 2601 39899 2635
rect 39899 2601 39908 2635
rect 39856 2592 39908 2601
rect 40500 2592 40552 2644
rect 19340 2388 19392 2440
rect 21732 2431 21784 2440
rect 21732 2397 21741 2431
rect 21741 2397 21775 2431
rect 21775 2397 21784 2431
rect 21732 2388 21784 2397
rect 22836 2431 22888 2440
rect 22836 2397 22845 2431
rect 22845 2397 22879 2431
rect 22879 2397 22888 2431
rect 22836 2388 22888 2397
rect 39120 2431 39172 2440
rect 39120 2397 39129 2431
rect 39129 2397 39163 2431
rect 39163 2397 39172 2431
rect 39120 2388 39172 2397
rect 40040 2431 40092 2440
rect 40040 2397 40049 2431
rect 40049 2397 40083 2431
rect 40083 2397 40092 2431
rect 40040 2388 40092 2397
rect 32956 2252 33008 2304
rect 11644 2150 11696 2202
rect 11708 2150 11760 2202
rect 11772 2150 11824 2202
rect 11836 2150 11888 2202
rect 11900 2150 11952 2202
rect 22338 2150 22390 2202
rect 22402 2150 22454 2202
rect 22466 2150 22518 2202
rect 22530 2150 22582 2202
rect 22594 2150 22646 2202
rect 33032 2150 33084 2202
rect 33096 2150 33148 2202
rect 33160 2150 33212 2202
rect 33224 2150 33276 2202
rect 33288 2150 33340 2202
rect 43726 2150 43778 2202
rect 43790 2150 43842 2202
rect 43854 2150 43906 2202
rect 43918 2150 43970 2202
rect 43982 2150 44034 2202
rect 22836 2048 22888 2100
rect 39120 2048 39172 2100
rect 40040 2091 40092 2100
rect 40040 2057 40049 2091
rect 40049 2057 40083 2091
rect 40083 2057 40092 2091
rect 40040 2048 40092 2057
rect 1584 1912 1636 1964
rect 3976 1844 4028 1896
rect 39396 1955 39448 1964
rect 39396 1921 39405 1955
rect 39405 1921 39439 1955
rect 39439 1921 39448 1955
rect 39396 1912 39448 1921
rect 43352 1912 43404 1964
rect 34152 1776 34204 1828
rect 6297 1606 6349 1658
rect 6361 1606 6413 1658
rect 6425 1606 6477 1658
rect 6489 1606 6541 1658
rect 6553 1606 6605 1658
rect 16991 1606 17043 1658
rect 17055 1606 17107 1658
rect 17119 1606 17171 1658
rect 17183 1606 17235 1658
rect 17247 1606 17299 1658
rect 27685 1606 27737 1658
rect 27749 1606 27801 1658
rect 27813 1606 27865 1658
rect 27877 1606 27929 1658
rect 27941 1606 27993 1658
rect 38379 1606 38431 1658
rect 38443 1606 38495 1658
rect 38507 1606 38559 1658
rect 38571 1606 38623 1658
rect 38635 1606 38687 1658
rect 1584 1547 1636 1556
rect 1584 1513 1593 1547
rect 1593 1513 1627 1547
rect 1627 1513 1636 1547
rect 1584 1504 1636 1513
rect 3976 1547 4028 1556
rect 3976 1513 3985 1547
rect 3985 1513 4019 1547
rect 4019 1513 4028 1547
rect 3976 1504 4028 1513
rect 39396 1504 39448 1556
rect 43352 1547 43404 1556
rect 43352 1513 43361 1547
rect 43361 1513 43395 1547
rect 43395 1513 43404 1547
rect 43352 1504 43404 1513
rect 1308 1300 1360 1352
rect 3792 1343 3844 1352
rect 3792 1309 3801 1343
rect 3801 1309 3835 1343
rect 3835 1309 3844 1343
rect 3792 1300 3844 1309
rect 5632 1343 5684 1352
rect 5632 1309 5641 1343
rect 5641 1309 5675 1343
rect 5675 1309 5684 1343
rect 5632 1300 5684 1309
rect 5816 1300 5868 1352
rect 7748 1343 7800 1352
rect 7748 1309 7757 1343
rect 7757 1309 7791 1343
rect 7791 1309 7800 1343
rect 7748 1300 7800 1309
rect 9864 1343 9916 1352
rect 9864 1309 9873 1343
rect 9873 1309 9907 1343
rect 9907 1309 9916 1343
rect 9864 1300 9916 1309
rect 11980 1343 12032 1352
rect 11980 1309 11989 1343
rect 11989 1309 12023 1343
rect 12023 1309 12032 1343
rect 11980 1300 12032 1309
rect 14280 1343 14332 1352
rect 14280 1309 14289 1343
rect 14289 1309 14323 1343
rect 14323 1309 14332 1343
rect 14280 1300 14332 1309
rect 16396 1343 16448 1352
rect 16396 1309 16405 1343
rect 16405 1309 16439 1343
rect 16439 1309 16448 1343
rect 16396 1300 16448 1309
rect 7932 1207 7984 1216
rect 7932 1173 7941 1207
rect 7941 1173 7975 1207
rect 7975 1173 7984 1207
rect 7932 1164 7984 1173
rect 14096 1207 14148 1216
rect 14096 1173 14105 1207
rect 14105 1173 14139 1207
rect 14139 1173 14148 1207
rect 14096 1164 14148 1173
rect 18144 1232 18196 1284
rect 18512 1343 18564 1352
rect 18512 1309 18521 1343
rect 18521 1309 18555 1343
rect 18555 1309 18564 1343
rect 18512 1300 18564 1309
rect 18972 1300 19024 1352
rect 19340 1300 19392 1352
rect 20628 1343 20680 1352
rect 20628 1309 20637 1343
rect 20637 1309 20671 1343
rect 20671 1309 20680 1343
rect 20628 1300 20680 1309
rect 22744 1343 22796 1352
rect 22744 1309 22753 1343
rect 22753 1309 22787 1343
rect 22787 1309 22796 1343
rect 22744 1300 22796 1309
rect 23204 1300 23256 1352
rect 24860 1343 24912 1352
rect 24860 1309 24869 1343
rect 24869 1309 24903 1343
rect 24903 1309 24912 1343
rect 24860 1300 24912 1309
rect 26700 1300 26752 1352
rect 27436 1300 27488 1352
rect 28908 1300 28960 1352
rect 29092 1343 29144 1352
rect 29092 1309 29101 1343
rect 29101 1309 29135 1343
rect 29135 1309 29144 1343
rect 29092 1300 29144 1309
rect 31208 1343 31260 1352
rect 31208 1309 31217 1343
rect 31217 1309 31251 1343
rect 31251 1309 31260 1343
rect 31208 1300 31260 1309
rect 31668 1300 31720 1352
rect 33324 1343 33376 1352
rect 33324 1309 33333 1343
rect 33333 1309 33367 1343
rect 33367 1309 33376 1343
rect 33324 1300 33376 1309
rect 34520 1300 34572 1352
rect 35256 1300 35308 1352
rect 35440 1343 35492 1352
rect 35440 1309 35449 1343
rect 35449 1309 35483 1343
rect 35483 1309 35492 1343
rect 35440 1300 35492 1309
rect 37556 1343 37608 1352
rect 37556 1309 37565 1343
rect 37565 1309 37599 1343
rect 37599 1309 37608 1343
rect 37556 1300 37608 1309
rect 39396 1300 39448 1352
rect 40868 1300 40920 1352
rect 41788 1343 41840 1352
rect 41788 1309 41797 1343
rect 41797 1309 41831 1343
rect 41831 1309 41840 1343
rect 41788 1300 41840 1309
rect 43536 1343 43588 1352
rect 43536 1309 43545 1343
rect 43545 1309 43579 1343
rect 43579 1309 43588 1343
rect 43536 1300 43588 1309
rect 18236 1164 18288 1216
rect 20536 1232 20588 1284
rect 24768 1232 24820 1284
rect 37372 1207 37424 1216
rect 37372 1173 37381 1207
rect 37381 1173 37415 1207
rect 37415 1173 37424 1207
rect 37372 1164 37424 1173
rect 11644 1062 11696 1114
rect 11708 1062 11760 1114
rect 11772 1062 11824 1114
rect 11836 1062 11888 1114
rect 11900 1062 11952 1114
rect 22338 1062 22390 1114
rect 22402 1062 22454 1114
rect 22466 1062 22518 1114
rect 22530 1062 22582 1114
rect 22594 1062 22646 1114
rect 33032 1062 33084 1114
rect 33096 1062 33148 1114
rect 33160 1062 33212 1114
rect 33224 1062 33276 1114
rect 33288 1062 33340 1114
rect 43726 1062 43778 1114
rect 43790 1062 43842 1114
rect 43854 1062 43906 1114
rect 43918 1062 43970 1114
rect 43982 1062 44034 1114
rect 14096 960 14148 1012
rect 21732 960 21784 1012
rect 18144 892 18196 944
rect 19616 892 19668 944
<< metal2 >>
rect 5354 9840 5410 10000
rect 5630 9840 5686 10000
rect 5906 9840 5962 10000
rect 6182 9840 6238 10000
rect 6458 9840 6514 10000
rect 6734 9840 6790 10000
rect 7010 9840 7066 10000
rect 7286 9840 7342 10000
rect 7562 9840 7618 10000
rect 7838 9840 7894 10000
rect 8114 9840 8170 10000
rect 8390 9840 8446 10000
rect 8666 9840 8722 10000
rect 8942 9840 8998 10000
rect 9218 9840 9274 10000
rect 9494 9840 9550 10000
rect 9770 9840 9826 10000
rect 10046 9840 10102 10000
rect 10322 9840 10378 10000
rect 10598 9840 10654 10000
rect 10874 9840 10930 10000
rect 11150 9840 11206 10000
rect 11426 9840 11482 10000
rect 11702 9840 11758 10000
rect 11978 9840 12034 10000
rect 12254 9840 12310 10000
rect 12530 9840 12586 10000
rect 12636 9846 12756 9874
rect 4894 9072 4950 9081
rect 4894 9007 4950 9016
rect 4908 8566 4936 9007
rect 5368 8634 5396 9840
rect 5644 8786 5672 9840
rect 5644 8758 5764 8786
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 5736 8090 5764 8758
rect 5920 8634 5948 9840
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5828 7546 5856 8434
rect 6196 8090 6224 9840
rect 6472 8378 6500 9840
rect 6472 8350 6684 8378
rect 6297 8188 6605 8197
rect 6297 8186 6303 8188
rect 6359 8186 6383 8188
rect 6439 8186 6463 8188
rect 6519 8186 6543 8188
rect 6599 8186 6605 8188
rect 6359 8134 6361 8186
rect 6541 8134 6543 8186
rect 6297 8132 6303 8134
rect 6359 8132 6383 8134
rect 6439 8132 6463 8134
rect 6519 8132 6543 8134
rect 6599 8132 6605 8134
rect 6297 8123 6605 8132
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6656 7546 6684 8350
rect 6748 8242 6776 9840
rect 7024 8634 7052 9840
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6748 8214 6960 8242
rect 6932 8022 6960 8214
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6734 7848 6790 7857
rect 6734 7783 6736 7792
rect 6788 7783 6790 7792
rect 6736 7754 6788 7760
rect 7300 7546 7328 9840
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 6552 7472 6604 7478
rect 6552 7414 6604 7420
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5920 6458 5948 7346
rect 6564 7313 6592 7414
rect 7392 7410 7420 8230
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 6550 7304 6606 7313
rect 6550 7239 6606 7248
rect 6297 7100 6605 7109
rect 6297 7098 6303 7100
rect 6359 7098 6383 7100
rect 6439 7098 6463 7100
rect 6519 7098 6543 7100
rect 6599 7098 6605 7100
rect 6359 7046 6361 7098
rect 6541 7046 6543 7098
rect 6297 7044 6303 7046
rect 6359 7044 6383 7046
rect 6439 7044 6463 7046
rect 6519 7044 6543 7046
rect 6599 7044 6605 7046
rect 6297 7035 6605 7044
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 7024 6361 7052 7346
rect 7484 6798 7512 8434
rect 7576 8090 7604 9840
rect 7564 8084 7616 8090
rect 7852 8072 7880 9840
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 7932 8084 7984 8090
rect 7852 8044 7932 8072
rect 7564 8026 7616 8032
rect 7932 8026 7984 8032
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7760 7206 7788 7754
rect 8036 7546 8064 8434
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7472 6792 7524 6798
rect 7470 6760 7472 6769
rect 7524 6760 7526 6769
rect 7470 6695 7526 6704
rect 7010 6352 7066 6361
rect 7010 6287 7066 6296
rect 8036 6225 8064 7482
rect 8128 7342 8156 9840
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8220 8634 8248 8842
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8312 8498 8340 9318
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8404 8072 8432 9840
rect 8680 8634 8708 9840
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8956 8514 8984 9840
rect 9036 9784 9088 9790
rect 9036 9726 9088 9732
rect 8496 8486 8984 8514
rect 9048 8498 9076 9726
rect 9036 8492 9088 8498
rect 8496 8362 8524 8486
rect 9036 8434 9088 8440
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8484 8084 8536 8090
rect 8404 8044 8484 8072
rect 9232 8072 9260 9840
rect 9508 8634 9536 9840
rect 9784 8634 9812 9840
rect 9956 9240 10008 9246
rect 9956 9182 10008 9188
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9876 8498 9904 8774
rect 9968 8498 9996 9182
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9312 8084 9364 8090
rect 9232 8044 9312 8072
rect 8484 8026 8536 8032
rect 9312 8026 9364 8032
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8022 6216 8078 6225
rect 8022 6151 8078 6160
rect 6297 6012 6605 6021
rect 6297 6010 6303 6012
rect 6359 6010 6383 6012
rect 6439 6010 6463 6012
rect 6519 6010 6543 6012
rect 6599 6010 6605 6012
rect 6359 5958 6361 6010
rect 6541 5958 6543 6010
rect 6297 5956 6303 5958
rect 6359 5956 6383 5958
rect 6439 5956 6463 5958
rect 6519 5956 6543 5958
rect 6599 5956 6605 5958
rect 6297 5947 6605 5956
rect 8220 5817 8248 7822
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 8404 7274 8432 7754
rect 9232 7342 9260 7754
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 9416 6866 9444 8298
rect 10060 8072 10088 9840
rect 10140 8084 10192 8090
rect 10060 8044 10140 8072
rect 10140 8026 10192 8032
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 7449 9628 7686
rect 9586 7440 9642 7449
rect 9586 7375 9642 7384
rect 10060 7002 10088 7754
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10336 6866 10364 9840
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10428 8566 10456 9386
rect 10612 8634 10640 9840
rect 10888 8634 10916 9840
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 11164 8072 11192 9840
rect 11440 8634 11468 9840
rect 11716 8922 11744 9840
rect 11532 8894 11744 8922
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11532 8090 11560 8894
rect 11644 8732 11952 8741
rect 11644 8730 11650 8732
rect 11706 8730 11730 8732
rect 11786 8730 11810 8732
rect 11866 8730 11890 8732
rect 11946 8730 11952 8732
rect 11706 8678 11708 8730
rect 11888 8678 11890 8730
rect 11644 8676 11650 8678
rect 11706 8676 11730 8678
rect 11786 8676 11810 8678
rect 11866 8676 11890 8678
rect 11946 8676 11952 8678
rect 11644 8667 11952 8676
rect 11244 8084 11296 8090
rect 11164 8044 11244 8072
rect 11244 8026 11296 8032
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11644 7644 11952 7653
rect 11644 7642 11650 7644
rect 11706 7642 11730 7644
rect 11786 7642 11810 7644
rect 11866 7642 11890 7644
rect 11946 7642 11952 7644
rect 11706 7590 11708 7642
rect 11888 7590 11890 7642
rect 11644 7588 11650 7590
rect 11706 7588 11730 7590
rect 11786 7588 11810 7590
rect 11866 7588 11890 7590
rect 11946 7588 11952 7590
rect 11644 7579 11952 7588
rect 11992 7546 12020 9840
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12084 8566 12112 8910
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12268 8004 12296 9840
rect 12440 8628 12492 8634
rect 12544 8616 12572 9840
rect 12492 8588 12572 8616
rect 12440 8570 12492 8576
rect 12636 8514 12664 9846
rect 12728 9840 12756 9846
rect 12806 9840 12862 10000
rect 13082 9840 13138 10000
rect 13358 9840 13414 10000
rect 13634 9840 13690 10000
rect 13910 9840 13966 10000
rect 14186 9840 14242 10000
rect 14462 9840 14518 10000
rect 14738 9840 14794 10000
rect 15014 9840 15070 10000
rect 15290 9840 15346 10000
rect 15566 9840 15622 10000
rect 15842 9840 15898 10000
rect 16118 9840 16174 10000
rect 16394 9840 16450 10000
rect 16500 9846 16620 9874
rect 12728 9812 12848 9840
rect 12714 9208 12770 9217
rect 12714 9143 12770 9152
rect 12452 8486 12664 8514
rect 12452 8362 12480 8486
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12440 8016 12492 8022
rect 12268 7976 12440 8004
rect 12440 7958 12492 7964
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 11644 6556 11952 6565
rect 11644 6554 11650 6556
rect 11706 6554 11730 6556
rect 11786 6554 11810 6556
rect 11866 6554 11890 6556
rect 11946 6554 11952 6556
rect 11706 6502 11708 6554
rect 11888 6502 11890 6554
rect 11644 6500 11650 6502
rect 11706 6500 11730 6502
rect 11786 6500 11810 6502
rect 11866 6500 11890 6502
rect 11946 6500 11952 6502
rect 11644 6491 11952 6500
rect 12268 6254 12296 7754
rect 12728 7410 12756 9143
rect 12990 7984 13046 7993
rect 12990 7919 13046 7928
rect 13004 7886 13032 7919
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13096 7546 13124 9840
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13188 8634 13216 9522
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13372 8090 13400 9840
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13464 8566 13492 9046
rect 13648 8634 13676 9840
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13924 8090 13952 9840
rect 14200 8634 14228 9840
rect 14372 9444 14424 9450
rect 14372 9386 14424 9392
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 14384 8498 14412 9386
rect 14476 8786 14504 9840
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14476 8758 14596 8786
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14568 8090 14596 8758
rect 14660 8362 14688 8978
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14752 8090 14780 9840
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14936 8498 14964 8910
rect 15028 8634 15056 9840
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 13740 6458 13768 7686
rect 14844 6633 14872 8366
rect 15120 8294 15148 9114
rect 15304 8634 15332 9840
rect 15580 8786 15608 9840
rect 15856 9042 15884 9840
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15580 8758 15700 8786
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15672 8090 15700 8758
rect 16040 8566 16068 9386
rect 16132 8634 16160 9840
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 16408 8004 16436 9840
rect 16500 8634 16528 9846
rect 16592 9840 16620 9846
rect 16670 9840 16726 10000
rect 16946 9840 17002 10000
rect 17222 9840 17278 10000
rect 17498 9840 17554 10000
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 16592 9812 16712 9840
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16592 8838 16620 8978
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16764 8832 16816 8838
rect 16960 8786 16988 9840
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 17052 9314 17080 9658
rect 17130 9480 17186 9489
rect 17130 9415 17186 9424
rect 17040 9308 17092 9314
rect 17040 9250 17092 9256
rect 16764 8774 16816 8780
rect 16776 8634 16804 8774
rect 16868 8758 16988 8786
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16580 8016 16632 8022
rect 16408 7976 16580 8004
rect 16580 7958 16632 7964
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 14936 7546 14964 7822
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 15476 7744 15528 7750
rect 15106 7712 15162 7721
rect 15476 7686 15528 7692
rect 15106 7647 15162 7656
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 15120 7478 15148 7647
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 14830 6624 14886 6633
rect 14830 6559 14886 6568
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 15488 6254 15516 7686
rect 16408 7546 16436 7754
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15580 6905 15608 7210
rect 15566 6896 15622 6905
rect 16500 6866 16528 7278
rect 15566 6831 15622 6840
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 16684 6186 16712 7822
rect 16776 7206 16804 8434
rect 16868 8090 16896 8758
rect 17144 8362 17172 9415
rect 17236 8634 17264 9840
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17420 9178 17448 9590
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17512 8634 17540 9840
rect 17604 9722 17632 9930
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 16991 8188 17299 8197
rect 16991 8186 16997 8188
rect 17053 8186 17077 8188
rect 17133 8186 17157 8188
rect 17213 8186 17237 8188
rect 17293 8186 17299 8188
rect 17053 8134 17055 8186
rect 17235 8134 17237 8186
rect 16991 8132 16997 8134
rect 17053 8132 17077 8134
rect 17133 8132 17157 8134
rect 17213 8132 17237 8134
rect 17293 8132 17299 8134
rect 16991 8123 17299 8132
rect 17420 8090 17448 8366
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17512 7546 17540 8434
rect 17604 7886 17632 9114
rect 17696 7936 17724 9862
rect 17774 9840 17830 10000
rect 17880 9846 18000 9874
rect 17788 8004 17816 9840
rect 17880 8634 17908 9846
rect 17972 9840 18000 9846
rect 18050 9840 18106 10000
rect 18326 9840 18382 10000
rect 18602 9840 18658 10000
rect 18878 9840 18934 10000
rect 19064 9988 19116 9994
rect 19064 9930 19116 9936
rect 17972 9812 18092 9840
rect 18340 8634 18368 9840
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18432 8634 18460 8910
rect 18616 8634 18644 9840
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18708 8809 18736 8978
rect 18694 8800 18750 8809
rect 18694 8735 18750 8744
rect 18892 8634 18920 9840
rect 19076 9738 19104 9930
rect 19154 9840 19210 10000
rect 19260 9846 19380 9874
rect 19260 9840 19288 9846
rect 19168 9812 19288 9840
rect 19076 9710 19288 9738
rect 19062 9344 19118 9353
rect 19062 9279 19064 9288
rect 19116 9279 19118 9288
rect 19156 9308 19208 9314
rect 19064 9250 19116 9256
rect 19156 9250 19208 9256
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18234 8528 18290 8537
rect 17960 8016 18012 8022
rect 17788 7976 17960 8004
rect 17960 7958 18012 7964
rect 17696 7908 17908 7936
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17788 7546 17816 7754
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17880 7410 17908 7908
rect 17960 7880 18012 7886
rect 17958 7848 17960 7857
rect 18012 7848 18014 7857
rect 18156 7800 18184 8502
rect 18234 8463 18290 8472
rect 18328 8492 18380 8498
rect 17958 7783 18014 7792
rect 18064 7772 18184 7800
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16991 7100 17299 7109
rect 16991 7098 16997 7100
rect 17053 7098 17077 7100
rect 17133 7098 17157 7100
rect 17213 7098 17237 7100
rect 17293 7098 17299 7100
rect 17053 7046 17055 7098
rect 17235 7046 17237 7098
rect 16991 7044 16997 7046
rect 17053 7044 17077 7046
rect 17133 7044 17157 7046
rect 17213 7044 17237 7046
rect 17293 7044 17299 7046
rect 16991 7035 17299 7044
rect 17604 6322 17632 7346
rect 18064 7206 18092 7772
rect 18248 7426 18276 8463
rect 18696 8492 18748 8498
rect 18380 8452 18460 8480
rect 18328 8434 18380 8440
rect 18328 8016 18380 8022
rect 18328 7958 18380 7964
rect 18340 7546 18368 7958
rect 18432 7546 18460 8452
rect 18696 8434 18748 8440
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18602 8256 18658 8265
rect 18524 7886 18552 8230
rect 18602 8191 18658 8200
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18616 7732 18644 8191
rect 18524 7704 18644 7732
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18156 7410 18276 7426
rect 18524 7410 18552 7704
rect 18144 7404 18276 7410
rect 18196 7398 18276 7404
rect 18512 7404 18564 7410
rect 18144 7346 18196 7352
rect 18512 7346 18564 7352
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18616 7206 18644 7346
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18708 6730 18736 8434
rect 18786 8392 18842 8401
rect 18786 8327 18842 8336
rect 18800 8090 18828 8327
rect 18892 8090 18920 8434
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18984 7886 19012 8910
rect 19076 7886 19104 8910
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19168 7732 19196 9250
rect 19076 7704 19196 7732
rect 19076 7410 19104 7704
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19168 6798 19196 7346
rect 19260 7206 19288 9710
rect 19352 8566 19380 9846
rect 19430 9840 19486 10000
rect 19706 9840 19762 10000
rect 19982 9840 20038 10000
rect 20074 9888 20130 9897
rect 19444 8616 19472 9840
rect 19616 9580 19668 9586
rect 19616 9522 19668 9528
rect 19524 8628 19576 8634
rect 19444 8588 19524 8616
rect 19524 8570 19576 8576
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19536 7750 19564 8434
rect 19628 8022 19656 9522
rect 19720 8265 19748 9840
rect 19996 9832 20074 9840
rect 20258 9840 20314 10000
rect 20364 9846 20484 9874
rect 19996 9823 20130 9832
rect 19996 9812 20116 9823
rect 19984 9376 20036 9382
rect 20168 9376 20220 9382
rect 19984 9318 20036 9324
rect 20166 9344 20168 9353
rect 20220 9344 20222 9353
rect 19706 8256 19762 8265
rect 19706 8191 19762 8200
rect 19996 8090 20024 9318
rect 20166 9279 20222 9288
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20180 8634 20208 8774
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19616 8016 19668 8022
rect 19616 7958 19668 7964
rect 19892 7880 19944 7886
rect 20088 7868 20116 8434
rect 20272 7936 20300 9840
rect 20364 8294 20392 9846
rect 20456 9840 20484 9846
rect 20534 9840 20590 10000
rect 20640 9846 20760 9874
rect 20456 9812 20576 9840
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20548 8838 20576 9658
rect 20536 8832 20588 8838
rect 20442 8800 20498 8809
rect 20536 8774 20588 8780
rect 20442 8735 20498 8744
rect 20456 8378 20484 8735
rect 20640 8650 20668 9846
rect 20732 9840 20760 9846
rect 20810 9840 20866 10000
rect 20916 9846 21036 9874
rect 20732 9812 20852 9840
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20732 9110 20760 9658
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20548 8622 20668 8650
rect 20548 8498 20576 8622
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20628 8424 20680 8430
rect 20456 8350 20576 8378
rect 20628 8366 20680 8372
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 19944 7840 20116 7868
rect 20180 7908 20300 7936
rect 19892 7822 19944 7828
rect 20180 7800 20208 7908
rect 20456 7886 20484 8230
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20180 7772 20300 7800
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 20074 7712 20130 7721
rect 20074 7647 20130 7656
rect 20088 7562 20116 7647
rect 19904 7546 20116 7562
rect 19892 7540 20116 7546
rect 19944 7534 20116 7540
rect 20166 7576 20222 7585
rect 20166 7511 20222 7520
rect 19892 7482 19944 7488
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 18696 6724 18748 6730
rect 18696 6666 18748 6672
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 16991 6012 17299 6021
rect 16991 6010 16997 6012
rect 17053 6010 17077 6012
rect 17133 6010 17157 6012
rect 17213 6010 17237 6012
rect 17293 6010 17299 6012
rect 17053 5958 17055 6010
rect 17235 5958 17237 6010
rect 16991 5956 16997 5958
rect 17053 5956 17077 5958
rect 17133 5956 17157 5958
rect 17213 5956 17237 5958
rect 17293 5956 17299 5958
rect 16991 5947 17299 5956
rect 17328 5846 17356 6054
rect 18800 5914 18828 6734
rect 19352 6730 19380 7346
rect 19536 7002 19564 7346
rect 20180 7313 20208 7511
rect 20272 7410 20300 7772
rect 20548 7750 20576 8350
rect 20640 7818 20668 8366
rect 20732 8265 20760 8842
rect 20812 8492 20864 8498
rect 20916 8480 20944 9846
rect 21008 9840 21036 9846
rect 21086 9840 21142 10000
rect 21192 9846 21312 9874
rect 21008 9812 21128 9840
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 20864 8452 20944 8480
rect 20812 8434 20864 8440
rect 20904 8288 20956 8294
rect 20718 8256 20774 8265
rect 20904 8230 20956 8236
rect 20718 8191 20774 8200
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20916 7546 20944 8230
rect 21008 8090 21036 8774
rect 21088 8492 21140 8498
rect 21192 8480 21220 9846
rect 21284 9840 21312 9846
rect 21362 9840 21418 10000
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 21284 9812 21404 9840
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21140 8452 21220 8480
rect 21088 8434 21140 8440
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21100 7886 21128 8230
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 21284 7834 21312 9318
rect 21376 8498 21404 9318
rect 21468 9110 21496 9862
rect 21638 9840 21694 10000
rect 21914 9840 21970 10000
rect 22190 9840 22246 10000
rect 22466 9840 22522 10000
rect 22742 9840 22798 10000
rect 22928 9852 22980 9858
rect 21546 9480 21602 9489
rect 21546 9415 21602 9424
rect 21456 9104 21508 9110
rect 21456 9046 21508 9052
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21560 8378 21588 9415
rect 21652 8498 21680 9840
rect 21928 9194 21956 9840
rect 21928 9166 22048 9194
rect 21914 9072 21970 9081
rect 21914 9007 21970 9016
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21376 8350 21588 8378
rect 21640 8356 21692 8362
rect 21376 8090 21404 8350
rect 21640 8298 21692 8304
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21468 8090 21496 8230
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21652 7886 21680 8298
rect 21732 8288 21784 8294
rect 21732 8230 21784 8236
rect 21548 7880 21600 7886
rect 21008 7546 21036 7822
rect 21284 7806 21496 7834
rect 21548 7822 21600 7828
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 21100 7478 21128 7686
rect 21088 7472 21140 7478
rect 21088 7414 21140 7420
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 19614 7304 19670 7313
rect 19614 7239 19616 7248
rect 19668 7239 19670 7248
rect 20166 7304 20222 7313
rect 20166 7239 20222 7248
rect 21088 7268 21140 7274
rect 19616 7210 19668 7216
rect 21088 7210 21140 7216
rect 20168 7200 20220 7206
rect 20166 7168 20168 7177
rect 20996 7200 21048 7206
rect 20220 7168 20222 7177
rect 20996 7142 21048 7148
rect 20166 7103 20222 7112
rect 19982 7032 20038 7041
rect 19524 6996 19576 7002
rect 19982 6967 20038 6976
rect 20258 7032 20314 7041
rect 21008 7002 21036 7142
rect 20258 6967 20314 6976
rect 20996 6996 21048 7002
rect 19524 6938 19576 6944
rect 19996 6798 20024 6967
rect 20272 6798 20300 6967
rect 20996 6938 21048 6944
rect 21100 6798 21128 7210
rect 21284 7002 21312 7686
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 21088 6792 21140 6798
rect 21376 6769 21404 7686
rect 21468 7206 21496 7806
rect 21560 7342 21588 7822
rect 21744 7410 21772 8230
rect 21824 8016 21876 8022
rect 21824 7958 21876 7964
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21456 6928 21508 6934
rect 21456 6870 21508 6876
rect 21088 6734 21140 6740
rect 21362 6760 21418 6769
rect 19340 6724 19392 6730
rect 21362 6695 21418 6704
rect 19340 6666 19392 6672
rect 21468 6633 21496 6870
rect 21454 6624 21510 6633
rect 21454 6559 21510 6568
rect 21836 6458 21864 7958
rect 21928 7478 21956 9007
rect 22020 8498 22048 9166
rect 22100 8560 22152 8566
rect 22100 8502 22152 8508
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 22112 7834 22140 8502
rect 22204 8480 22232 9840
rect 22480 9194 22508 9840
rect 22756 9330 22784 9840
rect 23018 9840 23074 10000
rect 23294 9840 23350 10000
rect 23570 9840 23626 10000
rect 23846 9840 23902 10000
rect 24122 9840 24178 10000
rect 24398 9840 24454 10000
rect 24674 9840 24730 10000
rect 24950 9840 25006 10000
rect 25226 9840 25282 10000
rect 25502 9840 25558 10000
rect 25778 9840 25834 10000
rect 26054 9840 26110 10000
rect 26330 9840 26386 10000
rect 26606 9840 26662 10000
rect 26882 9840 26938 10000
rect 27158 9840 27214 10000
rect 27434 9840 27490 10000
rect 27710 9840 27766 10000
rect 27986 9840 28042 10000
rect 28262 9840 28318 10000
rect 28538 9840 28594 10000
rect 28814 9840 28870 10000
rect 29090 9840 29146 10000
rect 29366 9840 29422 10000
rect 29642 9840 29698 10000
rect 29918 9840 29974 10000
rect 30194 9840 30250 10000
rect 30470 9840 30526 10000
rect 30746 9840 30802 10000
rect 31022 9840 31078 10000
rect 31298 9840 31354 10000
rect 31574 9840 31630 10000
rect 31668 9988 31720 9994
rect 31668 9930 31720 9936
rect 22928 9794 22980 9800
rect 22756 9302 22876 9330
rect 22480 9166 22784 9194
rect 22338 8732 22646 8741
rect 22338 8730 22344 8732
rect 22400 8730 22424 8732
rect 22480 8730 22504 8732
rect 22560 8730 22584 8732
rect 22640 8730 22646 8732
rect 22400 8678 22402 8730
rect 22582 8678 22584 8730
rect 22338 8676 22344 8678
rect 22400 8676 22424 8678
rect 22480 8676 22504 8678
rect 22560 8676 22584 8678
rect 22640 8676 22646 8678
rect 22338 8667 22646 8676
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22468 8492 22520 8498
rect 22204 8452 22468 8480
rect 22468 8434 22520 8440
rect 22190 8392 22246 8401
rect 22190 8327 22246 8336
rect 22204 8294 22232 8327
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 22572 8022 22600 8570
rect 22652 8560 22704 8566
rect 22652 8502 22704 8508
rect 22664 8022 22692 8502
rect 22756 8498 22784 9166
rect 22744 8492 22796 8498
rect 22848 8480 22876 9302
rect 22940 8634 22968 9794
rect 23032 9194 23060 9840
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 23032 9166 23152 9194
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 23124 8498 23152 9166
rect 23020 8492 23072 8498
rect 22848 8452 23020 8480
rect 22744 8434 22796 8440
rect 23020 8434 23072 8440
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23112 8288 23164 8294
rect 23112 8230 23164 8236
rect 23032 8090 23060 8230
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 22560 8016 22612 8022
rect 22560 7958 22612 7964
rect 22652 8016 22704 8022
rect 22652 7958 22704 7964
rect 23124 7886 23152 8230
rect 22652 7880 22704 7886
rect 22112 7806 22232 7834
rect 23112 7880 23164 7886
rect 22704 7828 22784 7834
rect 22652 7822 22784 7828
rect 23112 7822 23164 7828
rect 22664 7806 22784 7822
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 21916 7472 21968 7478
rect 21916 7414 21968 7420
rect 22006 7440 22062 7449
rect 22006 7375 22008 7384
rect 22060 7375 22062 7384
rect 22008 7346 22060 7352
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 21928 6390 21956 6802
rect 21916 6384 21968 6390
rect 21916 6326 21968 6332
rect 22112 6225 22140 7686
rect 22204 7274 22232 7806
rect 22338 7644 22646 7653
rect 22338 7642 22344 7644
rect 22400 7642 22424 7644
rect 22480 7642 22504 7644
rect 22560 7642 22584 7644
rect 22640 7642 22646 7644
rect 22400 7590 22402 7642
rect 22582 7590 22584 7642
rect 22338 7588 22344 7590
rect 22400 7588 22424 7590
rect 22480 7588 22504 7590
rect 22560 7588 22584 7590
rect 22640 7588 22646 7590
rect 22338 7579 22646 7588
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 22192 7268 22244 7274
rect 22192 7210 22244 7216
rect 22388 7154 22416 7278
rect 22480 7274 22508 7346
rect 22468 7268 22520 7274
rect 22468 7210 22520 7216
rect 22560 7268 22612 7274
rect 22560 7210 22612 7216
rect 22572 7154 22600 7210
rect 22388 7126 22600 7154
rect 22756 6934 22784 7806
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 22744 6928 22796 6934
rect 22848 6905 22876 7686
rect 23216 7546 23244 9590
rect 23308 9194 23336 9840
rect 23584 9194 23612 9840
rect 23860 9194 23888 9840
rect 24136 9194 24164 9840
rect 23308 9166 23428 9194
rect 23584 9166 23704 9194
rect 23860 9166 23980 9194
rect 24136 9166 24256 9194
rect 23400 8480 23428 9166
rect 23572 8492 23624 8498
rect 23400 8452 23572 8480
rect 23676 8480 23704 9166
rect 23848 8492 23900 8498
rect 23676 8452 23848 8480
rect 23572 8434 23624 8440
rect 23952 8480 23980 9166
rect 24124 8492 24176 8498
rect 23952 8452 24124 8480
rect 23848 8434 23900 8440
rect 24228 8480 24256 9166
rect 24412 8566 24440 9840
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24400 8560 24452 8566
rect 24400 8502 24452 8508
rect 24308 8492 24360 8498
rect 24228 8452 24308 8480
rect 24124 8434 24176 8440
rect 24308 8434 24360 8440
rect 23296 8356 23348 8362
rect 23296 8298 23348 8304
rect 23308 7886 23336 8298
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 23940 8288 23992 8294
rect 23940 8230 23992 8236
rect 24400 8288 24452 8294
rect 24400 8230 24452 8236
rect 24492 8288 24544 8294
rect 24492 8230 24544 8236
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 23308 7002 23336 7686
rect 23400 7546 23428 8230
rect 23676 8090 23704 8230
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 22744 6870 22796 6876
rect 22834 6896 22890 6905
rect 22834 6831 22890 6840
rect 22338 6556 22646 6565
rect 22338 6554 22344 6556
rect 22400 6554 22424 6556
rect 22480 6554 22504 6556
rect 22560 6554 22584 6556
rect 22640 6554 22646 6556
rect 22400 6502 22402 6554
rect 22582 6502 22584 6554
rect 22338 6500 22344 6502
rect 22400 6500 22424 6502
rect 22480 6500 22504 6502
rect 22560 6500 22584 6502
rect 22640 6500 22646 6502
rect 22338 6491 22646 6500
rect 22098 6216 22154 6225
rect 22098 6151 22154 6160
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 17316 5840 17368 5846
rect 8206 5808 8262 5817
rect 23492 5817 23520 7482
rect 23768 6361 23796 7686
rect 23952 7546 23980 8230
rect 24412 8090 24440 8230
rect 24400 8084 24452 8090
rect 24400 8026 24452 8032
rect 24032 8016 24084 8022
rect 24032 7958 24084 7964
rect 24044 7857 24072 7958
rect 24504 7886 24532 8230
rect 24308 7880 24360 7886
rect 24030 7848 24086 7857
rect 24308 7822 24360 7828
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 24030 7783 24086 7792
rect 24320 7546 24348 7822
rect 24492 7744 24544 7750
rect 24492 7686 24544 7692
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 24308 7540 24360 7546
rect 24308 7482 24360 7488
rect 24504 7478 24532 7686
rect 24492 7472 24544 7478
rect 24492 7414 24544 7420
rect 24596 7206 24624 8910
rect 24688 8616 24716 9840
rect 24768 8628 24820 8634
rect 24688 8588 24768 8616
rect 24768 8570 24820 8576
rect 24964 8430 24992 9840
rect 25240 8566 25268 9840
rect 25412 9512 25464 9518
rect 25412 9454 25464 9460
rect 25228 8560 25280 8566
rect 25228 8502 25280 8508
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 24860 8288 24912 8294
rect 24674 8256 24730 8265
rect 24860 8230 24912 8236
rect 25044 8288 25096 8294
rect 25044 8230 25096 8236
rect 25320 8288 25372 8294
rect 25320 8230 25372 8236
rect 24674 8191 24730 8200
rect 24688 8090 24716 8191
rect 24676 8084 24728 8090
rect 24676 8026 24728 8032
rect 24872 7886 24900 8230
rect 25056 7886 25084 8230
rect 25332 7886 25360 8230
rect 25424 8090 25452 9454
rect 25516 8634 25544 9840
rect 25596 9716 25648 9722
rect 25596 9658 25648 9664
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 25502 8120 25558 8129
rect 25412 8084 25464 8090
rect 25502 8055 25504 8064
rect 25412 8026 25464 8032
rect 25556 8055 25558 8064
rect 25504 8026 25556 8032
rect 25608 7954 25636 9658
rect 25688 9444 25740 9450
rect 25688 9386 25740 9392
rect 25700 8378 25728 9386
rect 25792 8480 25820 9840
rect 26068 9194 26096 9840
rect 26068 9166 26188 9194
rect 26160 8566 26188 9166
rect 26344 8634 26372 9840
rect 26332 8628 26384 8634
rect 26332 8570 26384 8576
rect 26148 8560 26200 8566
rect 26148 8502 26200 8508
rect 26056 8492 26108 8498
rect 25792 8452 26056 8480
rect 26620 8480 26648 9840
rect 26792 9444 26844 9450
rect 26792 9386 26844 9392
rect 26804 9110 26832 9386
rect 26896 9194 26924 9840
rect 26896 9166 27108 9194
rect 26792 9104 26844 9110
rect 26884 9104 26936 9110
rect 26792 9046 26844 9052
rect 26882 9072 26884 9081
rect 26936 9072 26938 9081
rect 26882 9007 26938 9016
rect 27080 8566 27108 9166
rect 27172 8634 27200 9840
rect 27344 9784 27396 9790
rect 27344 9726 27396 9732
rect 27250 9208 27306 9217
rect 27250 9143 27306 9152
rect 27160 8628 27212 8634
rect 27160 8570 27212 8576
rect 27068 8560 27120 8566
rect 27068 8502 27120 8508
rect 26884 8492 26936 8498
rect 26620 8452 26884 8480
rect 26056 8434 26108 8440
rect 26884 8434 26936 8440
rect 27264 8378 27292 9143
rect 25700 8350 25912 8378
rect 25780 8288 25832 8294
rect 25780 8230 25832 8236
rect 25596 7948 25648 7954
rect 25596 7890 25648 7896
rect 25792 7886 25820 8230
rect 25884 8090 25912 8350
rect 27172 8350 27292 8378
rect 26056 8288 26108 8294
rect 26056 8230 26108 8236
rect 26332 8288 26384 8294
rect 26332 8230 26384 8236
rect 26608 8288 26660 8294
rect 26608 8230 26660 8236
rect 26976 8288 27028 8294
rect 26976 8230 27028 8236
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 26068 7886 26096 8230
rect 26344 7886 26372 8230
rect 26620 7886 26648 8230
rect 26988 7886 27016 8230
rect 27172 8090 27200 8350
rect 27252 8288 27304 8294
rect 27252 8230 27304 8236
rect 27356 8242 27384 9726
rect 27448 8412 27476 9840
rect 27724 9194 27752 9840
rect 27724 9166 27844 9194
rect 27816 8566 27844 9166
rect 28000 8634 28028 9840
rect 28172 9240 28224 9246
rect 28172 9182 28224 9188
rect 27988 8628 28040 8634
rect 27988 8570 28040 8576
rect 27804 8560 27856 8566
rect 27804 8502 27856 8508
rect 27528 8424 27580 8430
rect 27448 8384 27528 8412
rect 27528 8366 27580 8372
rect 28184 8378 28212 9182
rect 28276 8634 28304 9840
rect 28264 8628 28316 8634
rect 28264 8570 28316 8576
rect 28184 8350 28304 8378
rect 27528 8288 27580 8294
rect 27160 8084 27212 8090
rect 27160 8026 27212 8032
rect 27264 7886 27292 8230
rect 27356 8214 27476 8242
rect 27528 8230 27580 8236
rect 27988 8288 28040 8294
rect 28172 8288 28224 8294
rect 28040 8248 28120 8276
rect 27988 8230 28040 8236
rect 27342 7984 27398 7993
rect 27342 7919 27398 7928
rect 27356 7886 27384 7919
rect 24860 7880 24912 7886
rect 24860 7822 24912 7828
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 25320 7880 25372 7886
rect 25320 7822 25372 7828
rect 25780 7880 25832 7886
rect 25780 7822 25832 7828
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 26332 7880 26384 7886
rect 26332 7822 26384 7828
rect 26608 7880 26660 7886
rect 26608 7822 26660 7828
rect 26976 7880 27028 7886
rect 26976 7822 27028 7828
rect 27252 7880 27304 7886
rect 27252 7822 27304 7828
rect 27344 7880 27396 7886
rect 27344 7822 27396 7828
rect 26148 7812 26200 7818
rect 26148 7754 26200 7760
rect 24860 7744 24912 7750
rect 24860 7686 24912 7692
rect 25136 7744 25188 7750
rect 25136 7686 25188 7692
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 24872 7313 24900 7686
rect 24858 7304 24914 7313
rect 24858 7239 24914 7248
rect 24584 7200 24636 7206
rect 24584 7142 24636 7148
rect 24860 7200 24912 7206
rect 24860 7142 24912 7148
rect 23754 6352 23810 6361
rect 23754 6287 23810 6296
rect 24872 5846 24900 7142
rect 25148 6866 25176 7686
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 25976 6322 26004 7686
rect 25964 6316 26016 6322
rect 25964 6258 26016 6264
rect 26160 6254 26188 7754
rect 26240 7744 26292 7750
rect 26240 7686 26292 7692
rect 27448 7698 27476 8214
rect 27540 7886 27568 8230
rect 27685 8188 27993 8197
rect 27685 8186 27691 8188
rect 27747 8186 27771 8188
rect 27827 8186 27851 8188
rect 27907 8186 27931 8188
rect 27987 8186 27993 8188
rect 27747 8134 27749 8186
rect 27929 8134 27931 8186
rect 27685 8132 27691 8134
rect 27747 8132 27771 8134
rect 27827 8132 27851 8134
rect 27907 8132 27931 8134
rect 27987 8132 27993 8134
rect 27685 8123 27993 8132
rect 27712 8084 27764 8090
rect 27712 8026 27764 8032
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 27724 7698 27752 8026
rect 28092 7886 28120 8248
rect 28172 8230 28224 8236
rect 28184 7954 28212 8230
rect 28276 8090 28304 8350
rect 28552 8344 28580 9840
rect 28828 9194 28856 9840
rect 28828 9166 28948 9194
rect 28920 8566 28948 9166
rect 29000 8900 29052 8906
rect 29000 8842 29052 8848
rect 28908 8560 28960 8566
rect 28908 8502 28960 8508
rect 28816 8356 28868 8362
rect 28552 8316 28816 8344
rect 28816 8298 28868 8304
rect 28908 8356 28960 8362
rect 28908 8298 28960 8304
rect 28356 8288 28408 8294
rect 28356 8230 28408 8236
rect 28448 8288 28500 8294
rect 28448 8230 28500 8236
rect 28264 8084 28316 8090
rect 28264 8026 28316 8032
rect 28172 7948 28224 7954
rect 28172 7890 28224 7896
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 28264 7880 28316 7886
rect 28264 7822 28316 7828
rect 26148 6248 26200 6254
rect 26148 6190 26200 6196
rect 26252 6186 26280 7686
rect 27448 7670 27752 7698
rect 28276 7546 28304 7822
rect 28264 7540 28316 7546
rect 28264 7482 28316 7488
rect 28368 7410 28396 8230
rect 28460 8090 28488 8230
rect 28448 8084 28500 8090
rect 28448 8026 28500 8032
rect 28920 7886 28948 8298
rect 28908 7880 28960 7886
rect 28908 7822 28960 7828
rect 28356 7404 28408 7410
rect 28356 7346 28408 7352
rect 27685 7100 27993 7109
rect 27685 7098 27691 7100
rect 27747 7098 27771 7100
rect 27827 7098 27851 7100
rect 27907 7098 27931 7100
rect 27987 7098 27993 7100
rect 27747 7046 27749 7098
rect 27929 7046 27931 7098
rect 27685 7044 27691 7046
rect 27747 7044 27771 7046
rect 27827 7044 27851 7046
rect 27907 7044 27931 7046
rect 27987 7044 27993 7046
rect 27685 7035 27993 7044
rect 26240 6180 26292 6186
rect 26240 6122 26292 6128
rect 27685 6012 27993 6021
rect 27685 6010 27691 6012
rect 27747 6010 27771 6012
rect 27827 6010 27851 6012
rect 27907 6010 27931 6012
rect 27987 6010 27993 6012
rect 27747 5958 27749 6010
rect 27929 5958 27931 6010
rect 27685 5956 27691 5958
rect 27747 5956 27771 5958
rect 27827 5956 27851 5958
rect 27907 5956 27931 5958
rect 27987 5956 27993 5958
rect 27685 5947 27993 5956
rect 24860 5840 24912 5846
rect 17316 5782 17368 5788
rect 23478 5808 23534 5817
rect 8206 5743 8262 5752
rect 24860 5782 24912 5788
rect 23478 5743 23534 5752
rect 29012 5642 29040 8842
rect 29104 8634 29132 9840
rect 29276 9648 29328 9654
rect 29276 9590 29328 9596
rect 29092 8628 29144 8634
rect 29092 8570 29144 8576
rect 22744 5636 22796 5642
rect 22744 5578 22796 5584
rect 29000 5636 29052 5642
rect 29000 5578 29052 5584
rect 11644 5468 11952 5477
rect 11644 5466 11650 5468
rect 11706 5466 11730 5468
rect 11786 5466 11810 5468
rect 11866 5466 11890 5468
rect 11946 5466 11952 5468
rect 11706 5414 11708 5466
rect 11888 5414 11890 5466
rect 11644 5412 11650 5414
rect 11706 5412 11730 5414
rect 11786 5412 11810 5414
rect 11866 5412 11890 5414
rect 11946 5412 11952 5414
rect 11644 5403 11952 5412
rect 22338 5468 22646 5477
rect 22338 5466 22344 5468
rect 22400 5466 22424 5468
rect 22480 5466 22504 5468
rect 22560 5466 22584 5468
rect 22640 5466 22646 5468
rect 22400 5414 22402 5466
rect 22582 5414 22584 5466
rect 22338 5412 22344 5414
rect 22400 5412 22424 5414
rect 22480 5412 22504 5414
rect 22560 5412 22584 5414
rect 22640 5412 22646 5414
rect 22338 5403 22646 5412
rect 6297 4924 6605 4933
rect 6297 4922 6303 4924
rect 6359 4922 6383 4924
rect 6439 4922 6463 4924
rect 6519 4922 6543 4924
rect 6599 4922 6605 4924
rect 6359 4870 6361 4922
rect 6541 4870 6543 4922
rect 6297 4868 6303 4870
rect 6359 4868 6383 4870
rect 6439 4868 6463 4870
rect 6519 4868 6543 4870
rect 6599 4868 6605 4870
rect 6297 4859 6605 4868
rect 16991 4924 17299 4933
rect 16991 4922 16997 4924
rect 17053 4922 17077 4924
rect 17133 4922 17157 4924
rect 17213 4922 17237 4924
rect 17293 4922 17299 4924
rect 17053 4870 17055 4922
rect 17235 4870 17237 4922
rect 16991 4868 16997 4870
rect 17053 4868 17077 4870
rect 17133 4868 17157 4870
rect 17213 4868 17237 4870
rect 17293 4868 17299 4870
rect 16991 4859 17299 4868
rect 22756 4826 22784 5578
rect 25964 5160 26016 5166
rect 25964 5102 26016 5108
rect 25976 4826 26004 5102
rect 26056 5024 26108 5030
rect 26056 4966 26108 4972
rect 26068 4826 26096 4966
rect 27685 4924 27993 4933
rect 27685 4922 27691 4924
rect 27747 4922 27771 4924
rect 27827 4922 27851 4924
rect 27907 4922 27931 4924
rect 27987 4922 27993 4924
rect 27747 4870 27749 4922
rect 27929 4870 27931 4922
rect 27685 4868 27691 4870
rect 27747 4868 27771 4870
rect 27827 4868 27851 4870
rect 27907 4868 27931 4870
rect 27987 4868 27993 4870
rect 27685 4859 27993 4868
rect 22744 4820 22796 4826
rect 22744 4762 22796 4768
rect 25964 4820 26016 4826
rect 25964 4762 26016 4768
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 25872 4616 25924 4622
rect 25872 4558 25924 4564
rect 27988 4616 28040 4622
rect 27988 4558 28040 4564
rect 11644 4380 11952 4389
rect 11644 4378 11650 4380
rect 11706 4378 11730 4380
rect 11786 4378 11810 4380
rect 11866 4378 11890 4380
rect 11946 4378 11952 4380
rect 11706 4326 11708 4378
rect 11888 4326 11890 4378
rect 11644 4324 11650 4326
rect 11706 4324 11730 4326
rect 11786 4324 11810 4326
rect 11866 4324 11890 4326
rect 11946 4324 11952 4326
rect 11644 4315 11952 4324
rect 21652 4282 21680 4558
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 6297 3836 6605 3845
rect 6297 3834 6303 3836
rect 6359 3834 6383 3836
rect 6439 3834 6463 3836
rect 6519 3834 6543 3836
rect 6599 3834 6605 3836
rect 6359 3782 6361 3834
rect 6541 3782 6543 3834
rect 6297 3780 6303 3782
rect 6359 3780 6383 3782
rect 6439 3780 6463 3782
rect 6519 3780 6543 3782
rect 6599 3780 6605 3782
rect 6297 3771 6605 3780
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 1584 1964 1636 1970
rect 1584 1906 1636 1912
rect 1596 1562 1624 1906
rect 3976 1896 4028 1902
rect 3976 1838 4028 1844
rect 3988 1562 4016 1838
rect 1584 1556 1636 1562
rect 1584 1498 1636 1504
rect 3976 1556 4028 1562
rect 3976 1498 4028 1504
rect 5828 1358 5856 3606
rect 6297 2748 6605 2757
rect 6297 2746 6303 2748
rect 6359 2746 6383 2748
rect 6439 2746 6463 2748
rect 6519 2746 6543 2748
rect 6599 2746 6605 2748
rect 6359 2694 6361 2746
rect 6541 2694 6543 2746
rect 6297 2692 6303 2694
rect 6359 2692 6383 2694
rect 6439 2692 6463 2694
rect 6519 2692 6543 2694
rect 6599 2692 6605 2694
rect 6297 2683 6605 2692
rect 6297 1660 6605 1669
rect 6297 1658 6303 1660
rect 6359 1658 6383 1660
rect 6439 1658 6463 1660
rect 6519 1658 6543 1660
rect 6599 1658 6605 1660
rect 6359 1606 6361 1658
rect 6541 1606 6543 1658
rect 6297 1604 6303 1606
rect 6359 1604 6383 1606
rect 6439 1604 6463 1606
rect 6519 1604 6543 1606
rect 6599 1604 6605 1606
rect 6297 1595 6605 1604
rect 1308 1352 1360 1358
rect 1308 1294 1360 1300
rect 3792 1352 3844 1358
rect 3792 1294 3844 1300
rect 5632 1352 5684 1358
rect 5632 1294 5684 1300
rect 5816 1352 5868 1358
rect 5816 1294 5868 1300
rect 7748 1352 7800 1358
rect 7748 1294 7800 1300
rect 1320 160 1348 1294
rect 1306 0 1362 160
rect 3422 82 3478 160
rect 3804 82 3832 1294
rect 3422 54 3832 82
rect 5538 82 5594 160
rect 5644 82 5672 1294
rect 5538 54 5672 82
rect 7654 82 7710 160
rect 7760 82 7788 1294
rect 7944 1222 7972 4014
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 16991 3836 17299 3845
rect 16991 3834 16997 3836
rect 17053 3834 17077 3836
rect 17133 3834 17157 3836
rect 17213 3834 17237 3836
rect 17293 3834 17299 3836
rect 17053 3782 17055 3834
rect 17235 3782 17237 3834
rect 16991 3780 16997 3782
rect 17053 3780 17077 3782
rect 17133 3780 17157 3782
rect 17213 3780 17237 3782
rect 17293 3780 17299 3782
rect 16991 3771 17299 3780
rect 11644 3292 11952 3301
rect 11644 3290 11650 3292
rect 11706 3290 11730 3292
rect 11786 3290 11810 3292
rect 11866 3290 11890 3292
rect 11946 3290 11952 3292
rect 11706 3238 11708 3290
rect 11888 3238 11890 3290
rect 11644 3236 11650 3238
rect 11706 3236 11730 3238
rect 11786 3236 11810 3238
rect 11866 3236 11890 3238
rect 11946 3236 11952 3238
rect 11644 3227 11952 3236
rect 16991 2748 17299 2757
rect 16991 2746 16997 2748
rect 17053 2746 17077 2748
rect 17133 2746 17157 2748
rect 17213 2746 17237 2748
rect 17293 2746 17299 2748
rect 17053 2694 17055 2746
rect 17235 2694 17237 2746
rect 16991 2692 16997 2694
rect 17053 2692 17077 2694
rect 17133 2692 17157 2694
rect 17213 2692 17237 2694
rect 17293 2692 17299 2694
rect 16991 2683 17299 2692
rect 11644 2204 11952 2213
rect 11644 2202 11650 2204
rect 11706 2202 11730 2204
rect 11786 2202 11810 2204
rect 11866 2202 11890 2204
rect 11946 2202 11952 2204
rect 11706 2150 11708 2202
rect 11888 2150 11890 2202
rect 11644 2148 11650 2150
rect 11706 2148 11730 2150
rect 11786 2148 11810 2150
rect 11866 2148 11890 2150
rect 11946 2148 11952 2150
rect 11644 2139 11952 2148
rect 16991 1660 17299 1669
rect 16991 1658 16997 1660
rect 17053 1658 17077 1660
rect 17133 1658 17157 1660
rect 17213 1658 17237 1660
rect 17293 1658 17299 1660
rect 17053 1606 17055 1658
rect 17235 1606 17237 1658
rect 16991 1604 16997 1606
rect 17053 1604 17077 1606
rect 17133 1604 17157 1606
rect 17213 1604 17237 1606
rect 17293 1604 17299 1606
rect 16991 1595 17299 1604
rect 9864 1352 9916 1358
rect 9864 1294 9916 1300
rect 11980 1352 12032 1358
rect 11980 1294 12032 1300
rect 14280 1352 14332 1358
rect 14280 1294 14332 1300
rect 16396 1352 16448 1358
rect 16396 1294 16448 1300
rect 7932 1216 7984 1222
rect 7932 1158 7984 1164
rect 7654 54 7788 82
rect 9770 82 9826 160
rect 9876 82 9904 1294
rect 11644 1116 11952 1125
rect 11644 1114 11650 1116
rect 11706 1114 11730 1116
rect 11786 1114 11810 1116
rect 11866 1114 11890 1116
rect 11946 1114 11952 1116
rect 11706 1062 11708 1114
rect 11888 1062 11890 1114
rect 11644 1060 11650 1062
rect 11706 1060 11730 1062
rect 11786 1060 11810 1062
rect 11866 1060 11890 1062
rect 11946 1060 11952 1062
rect 11644 1051 11952 1060
rect 9770 54 9904 82
rect 11886 82 11942 160
rect 11992 82 12020 1294
rect 14096 1216 14148 1222
rect 14096 1158 14148 1164
rect 14108 1018 14136 1158
rect 14096 1012 14148 1018
rect 14096 954 14148 960
rect 11886 54 12020 82
rect 14002 82 14058 160
rect 14292 82 14320 1294
rect 14002 54 14320 82
rect 16118 82 16174 160
rect 16408 82 16436 1294
rect 18144 1284 18196 1290
rect 18144 1226 18196 1232
rect 18156 950 18184 1226
rect 18248 1222 18276 3878
rect 19616 3596 19668 3602
rect 19616 3538 19668 3544
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19536 3194 19564 3470
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18984 1358 19012 2994
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19352 1358 19380 2382
rect 18512 1352 18564 1358
rect 18512 1294 18564 1300
rect 18972 1352 19024 1358
rect 18972 1294 19024 1300
rect 19340 1352 19392 1358
rect 19340 1294 19392 1300
rect 18236 1216 18288 1222
rect 18236 1158 18288 1164
rect 18144 944 18196 950
rect 18144 886 18196 892
rect 16118 54 16436 82
rect 18234 82 18290 160
rect 18524 82 18552 1294
rect 19628 950 19656 3538
rect 20548 1290 20576 4082
rect 22020 3738 22048 4082
rect 22204 4010 22232 4558
rect 22338 4380 22646 4389
rect 22338 4378 22344 4380
rect 22400 4378 22424 4380
rect 22480 4378 22504 4380
rect 22560 4378 22584 4380
rect 22640 4378 22646 4380
rect 22400 4326 22402 4378
rect 22582 4326 22584 4378
rect 22338 4324 22344 4326
rect 22400 4324 22424 4326
rect 22480 4324 22504 4326
rect 22560 4324 22584 4326
rect 22640 4324 22646 4326
rect 22338 4315 22646 4324
rect 22756 4214 22784 4558
rect 22744 4208 22796 4214
rect 22744 4150 22796 4156
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 22008 3732 22060 3738
rect 22008 3674 22060 3680
rect 22848 3602 22876 4082
rect 23124 4010 23152 4558
rect 23400 4282 23428 4558
rect 25884 4282 25912 4558
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 25872 4276 25924 4282
rect 25872 4218 25924 4224
rect 23756 4140 23808 4146
rect 23756 4082 23808 4088
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 27436 4140 27488 4146
rect 27436 4082 27488 4088
rect 23112 4004 23164 4010
rect 23112 3946 23164 3952
rect 23768 3738 23796 4082
rect 23756 3732 23808 3738
rect 23756 3674 23808 3680
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 22338 3292 22646 3301
rect 22338 3290 22344 3292
rect 22400 3290 22424 3292
rect 22480 3290 22504 3292
rect 22560 3290 22584 3292
rect 22640 3290 22646 3292
rect 22400 3238 22402 3290
rect 22582 3238 22584 3290
rect 22338 3236 22344 3238
rect 22400 3236 22424 3238
rect 22480 3236 22504 3238
rect 22560 3236 22584 3238
rect 22640 3236 22646 3238
rect 22338 3227 22646 3236
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 22020 2650 22048 2994
rect 22388 2650 22416 2994
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 21732 2440 21784 2446
rect 21732 2382 21784 2388
rect 22836 2440 22888 2446
rect 22836 2382 22888 2388
rect 20628 1352 20680 1358
rect 20628 1294 20680 1300
rect 20536 1284 20588 1290
rect 20536 1226 20588 1232
rect 19616 944 19668 950
rect 19616 886 19668 892
rect 18234 54 18552 82
rect 20350 82 20406 160
rect 20640 82 20668 1294
rect 21744 1018 21772 2382
rect 22338 2204 22646 2213
rect 22338 2202 22344 2204
rect 22400 2202 22424 2204
rect 22480 2202 22504 2204
rect 22560 2202 22584 2204
rect 22640 2202 22646 2204
rect 22400 2150 22402 2202
rect 22582 2150 22584 2202
rect 22338 2148 22344 2150
rect 22400 2148 22424 2150
rect 22480 2148 22504 2150
rect 22560 2148 22584 2150
rect 22640 2148 22646 2150
rect 22338 2139 22646 2148
rect 22848 2106 22876 2382
rect 22836 2100 22888 2106
rect 22836 2042 22888 2048
rect 23216 1358 23244 3470
rect 22744 1352 22796 1358
rect 22744 1294 22796 1300
rect 23204 1352 23256 1358
rect 23204 1294 23256 1300
rect 22338 1116 22646 1125
rect 22338 1114 22344 1116
rect 22400 1114 22424 1116
rect 22480 1114 22504 1116
rect 22560 1114 22584 1116
rect 22640 1114 22646 1116
rect 22400 1062 22402 1114
rect 22582 1062 22584 1114
rect 22338 1060 22344 1062
rect 22400 1060 22424 1062
rect 22480 1060 22504 1062
rect 22560 1060 22584 1062
rect 22640 1060 22646 1062
rect 22338 1051 22646 1060
rect 21732 1012 21784 1018
rect 21732 954 21784 960
rect 20350 54 20668 82
rect 22466 82 22522 160
rect 22756 82 22784 1294
rect 24780 1290 24808 4082
rect 27448 1358 27476 4082
rect 28000 4078 28028 4558
rect 27988 4072 28040 4078
rect 27988 4014 28040 4020
rect 29288 4010 29316 9590
rect 29380 8412 29408 9840
rect 29656 8566 29684 9840
rect 29644 8560 29696 8566
rect 29644 8502 29696 8508
rect 29932 8430 29960 9840
rect 30208 8566 30236 9840
rect 30288 8832 30340 8838
rect 30288 8774 30340 8780
rect 30380 8832 30432 8838
rect 30380 8774 30432 8780
rect 30300 8634 30328 8774
rect 30288 8628 30340 8634
rect 30288 8570 30340 8576
rect 30196 8560 30248 8566
rect 30196 8502 30248 8508
rect 29552 8424 29604 8430
rect 29380 8384 29552 8412
rect 29552 8366 29604 8372
rect 29920 8424 29972 8430
rect 29920 8366 29972 8372
rect 29552 8288 29604 8294
rect 29552 8230 29604 8236
rect 29828 8288 29880 8294
rect 29828 8230 29880 8236
rect 29564 7546 29592 8230
rect 29552 7540 29604 7546
rect 29552 7482 29604 7488
rect 29840 7002 29868 8230
rect 29828 6996 29880 7002
rect 29828 6938 29880 6944
rect 30392 4690 30420 8774
rect 30484 8634 30512 9840
rect 30564 9036 30616 9042
rect 30564 8978 30616 8984
rect 30656 9036 30708 9042
rect 30656 8978 30708 8984
rect 30472 8628 30524 8634
rect 30472 8570 30524 8576
rect 30576 8498 30604 8978
rect 30564 8492 30616 8498
rect 30564 8434 30616 8440
rect 30668 5166 30696 8978
rect 30760 8430 30788 9840
rect 31036 8566 31064 9840
rect 31116 9172 31168 9178
rect 31116 9114 31168 9120
rect 31128 8634 31156 9114
rect 31116 8628 31168 8634
rect 31116 8570 31168 8576
rect 31024 8560 31076 8566
rect 31024 8502 31076 8508
rect 31312 8430 31340 9840
rect 31392 9308 31444 9314
rect 31392 9250 31444 9256
rect 31404 8634 31432 9250
rect 31484 9240 31536 9246
rect 31484 9182 31536 9188
rect 31392 8628 31444 8634
rect 31392 8570 31444 8576
rect 30748 8424 30800 8430
rect 30748 8366 30800 8372
rect 31300 8424 31352 8430
rect 31300 8366 31352 8372
rect 30840 8356 30892 8362
rect 30840 8298 30892 8304
rect 30852 5914 30880 8298
rect 30840 5908 30892 5914
rect 30840 5850 30892 5856
rect 30656 5160 30708 5166
rect 30656 5102 30708 5108
rect 30380 4684 30432 4690
rect 30380 4626 30432 4632
rect 29276 4004 29328 4010
rect 29276 3946 29328 3952
rect 27685 3836 27993 3845
rect 27685 3834 27691 3836
rect 27747 3834 27771 3836
rect 27827 3834 27851 3836
rect 27907 3834 27931 3836
rect 27987 3834 27993 3836
rect 27747 3782 27749 3834
rect 27929 3782 27931 3834
rect 27685 3780 27691 3782
rect 27747 3780 27771 3782
rect 27827 3780 27851 3782
rect 27907 3780 27931 3782
rect 27987 3780 27993 3782
rect 27685 3771 27993 3780
rect 30104 3528 30156 3534
rect 30104 3470 30156 3476
rect 30116 3194 30144 3470
rect 31496 3194 31524 9182
rect 31588 8566 31616 9840
rect 31680 8634 31708 9930
rect 31850 9840 31906 10000
rect 32126 9840 32182 10000
rect 32402 9840 32458 10000
rect 32678 9840 32734 10000
rect 32954 9840 33010 10000
rect 33230 9840 33286 10000
rect 33506 9840 33562 10000
rect 33782 9840 33838 10000
rect 34058 9840 34114 10000
rect 34334 9840 34390 10000
rect 34610 9840 34666 10000
rect 34886 9840 34942 10000
rect 35162 9840 35218 10000
rect 35438 9840 35494 10000
rect 35714 9840 35770 10000
rect 35990 9840 36046 10000
rect 36266 9840 36322 10000
rect 36542 9840 36598 10000
rect 36818 9840 36874 10000
rect 37094 9840 37150 10000
rect 37370 9840 37426 10000
rect 37646 9840 37702 10000
rect 37922 9840 37978 10000
rect 38198 9840 38254 10000
rect 38474 9840 38530 10000
rect 38750 9840 38806 10000
rect 39026 9840 39082 10000
rect 39132 9846 39252 9874
rect 39132 9840 39160 9846
rect 31864 8634 31892 9840
rect 32036 9444 32088 9450
rect 32036 9386 32088 9392
rect 31668 8628 31720 8634
rect 31668 8570 31720 8576
rect 31852 8628 31904 8634
rect 31852 8570 31904 8576
rect 31576 8560 31628 8566
rect 31576 8502 31628 8508
rect 31942 8528 31998 8537
rect 32048 8498 32076 9386
rect 31942 8463 31998 8472
rect 32036 8492 32088 8498
rect 31956 8362 31984 8463
rect 32036 8434 32088 8440
rect 32140 8412 32168 9840
rect 32218 8936 32274 8945
rect 32218 8871 32274 8880
rect 32232 8566 32260 8871
rect 32220 8560 32272 8566
rect 32416 8548 32444 9840
rect 32692 8634 32720 9840
rect 32864 9580 32916 9586
rect 32864 9522 32916 9528
rect 32772 9376 32824 9382
rect 32772 9318 32824 9324
rect 32680 8628 32732 8634
rect 32680 8570 32732 8576
rect 32588 8560 32640 8566
rect 32416 8520 32588 8548
rect 32220 8502 32272 8508
rect 32588 8502 32640 8508
rect 32784 8498 32812 9318
rect 32772 8492 32824 8498
rect 32772 8434 32824 8440
rect 32312 8424 32364 8430
rect 32140 8384 32312 8412
rect 32312 8366 32364 8372
rect 32876 8362 32904 9522
rect 32968 8480 32996 9840
rect 33244 9194 33272 9840
rect 33244 9166 33456 9194
rect 33032 8732 33340 8741
rect 33032 8730 33038 8732
rect 33094 8730 33118 8732
rect 33174 8730 33198 8732
rect 33254 8730 33278 8732
rect 33334 8730 33340 8732
rect 33094 8678 33096 8730
rect 33276 8678 33278 8730
rect 33032 8676 33038 8678
rect 33094 8676 33118 8678
rect 33174 8676 33198 8678
rect 33254 8676 33278 8678
rect 33334 8676 33340 8678
rect 33032 8667 33340 8676
rect 33428 8566 33456 9166
rect 33416 8560 33468 8566
rect 33416 8502 33468 8508
rect 33324 8492 33376 8498
rect 32968 8452 33324 8480
rect 33324 8434 33376 8440
rect 31944 8356 31996 8362
rect 31944 8298 31996 8304
rect 32864 8356 32916 8362
rect 32864 8298 32916 8304
rect 33232 8356 33284 8362
rect 33232 8298 33284 8304
rect 33244 8242 33272 8298
rect 32968 8214 33272 8242
rect 32220 4616 32272 4622
rect 32220 4558 32272 4564
rect 31668 4140 31720 4146
rect 31668 4082 31720 4088
rect 30104 3188 30156 3194
rect 30104 3130 30156 3136
rect 31484 3188 31536 3194
rect 31484 3130 31536 3136
rect 28908 3052 28960 3058
rect 28908 2994 28960 3000
rect 27685 2748 27993 2757
rect 27685 2746 27691 2748
rect 27747 2746 27771 2748
rect 27827 2746 27851 2748
rect 27907 2746 27931 2748
rect 27987 2746 27993 2748
rect 27747 2694 27749 2746
rect 27929 2694 27931 2746
rect 27685 2692 27691 2694
rect 27747 2692 27771 2694
rect 27827 2692 27851 2694
rect 27907 2692 27931 2694
rect 27987 2692 27993 2694
rect 27685 2683 27993 2692
rect 27685 1660 27993 1669
rect 27685 1658 27691 1660
rect 27747 1658 27771 1660
rect 27827 1658 27851 1660
rect 27907 1658 27931 1660
rect 27987 1658 27993 1660
rect 27747 1606 27749 1658
rect 27929 1606 27931 1658
rect 27685 1604 27691 1606
rect 27747 1604 27771 1606
rect 27827 1604 27851 1606
rect 27907 1604 27931 1606
rect 27987 1604 27993 1606
rect 27685 1595 27993 1604
rect 28920 1358 28948 2994
rect 31680 1358 31708 4082
rect 32232 4078 32260 4558
rect 32220 4072 32272 4078
rect 32220 4014 32272 4020
rect 32968 2310 32996 8214
rect 33520 7868 33548 9840
rect 33600 9172 33652 9178
rect 33600 9114 33652 9120
rect 33612 8378 33640 9114
rect 33692 9036 33744 9042
rect 33692 8978 33744 8984
rect 33704 8634 33732 8978
rect 33692 8628 33744 8634
rect 33692 8570 33744 8576
rect 33612 8362 33732 8378
rect 33612 8356 33744 8362
rect 33612 8350 33692 8356
rect 33692 8298 33744 8304
rect 33600 7880 33652 7886
rect 33520 7840 33600 7868
rect 33796 7868 33824 9840
rect 34072 8634 34100 9840
rect 34348 9092 34376 9840
rect 34348 9064 34468 9092
rect 34440 8634 34468 9064
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 34428 8628 34480 8634
rect 34428 8570 34480 8576
rect 34152 8492 34204 8498
rect 34152 8434 34204 8440
rect 33968 8356 34020 8362
rect 33968 8298 34020 8304
rect 33876 7880 33928 7886
rect 33796 7840 33876 7868
rect 33600 7822 33652 7828
rect 33876 7822 33928 7828
rect 33784 7744 33836 7750
rect 33784 7686 33836 7692
rect 33032 7644 33340 7653
rect 33032 7642 33038 7644
rect 33094 7642 33118 7644
rect 33174 7642 33198 7644
rect 33254 7642 33278 7644
rect 33334 7642 33340 7644
rect 33094 7590 33096 7642
rect 33276 7590 33278 7642
rect 33032 7588 33038 7590
rect 33094 7588 33118 7590
rect 33174 7588 33198 7590
rect 33254 7588 33278 7590
rect 33334 7588 33340 7590
rect 33032 7579 33340 7588
rect 33796 7546 33824 7686
rect 33784 7540 33836 7546
rect 33784 7482 33836 7488
rect 33980 7449 34008 8298
rect 34060 7744 34112 7750
rect 34060 7686 34112 7692
rect 34072 7546 34100 7686
rect 34060 7540 34112 7546
rect 34060 7482 34112 7488
rect 33966 7440 34022 7449
rect 33966 7375 34022 7384
rect 33032 6556 33340 6565
rect 33032 6554 33038 6556
rect 33094 6554 33118 6556
rect 33174 6554 33198 6556
rect 33254 6554 33278 6556
rect 33334 6554 33340 6556
rect 33094 6502 33096 6554
rect 33276 6502 33278 6554
rect 33032 6500 33038 6502
rect 33094 6500 33118 6502
rect 33174 6500 33198 6502
rect 33254 6500 33278 6502
rect 33334 6500 33340 6502
rect 33032 6491 33340 6500
rect 33032 5468 33340 5477
rect 33032 5466 33038 5468
rect 33094 5466 33118 5468
rect 33174 5466 33198 5468
rect 33254 5466 33278 5468
rect 33334 5466 33340 5468
rect 33094 5414 33096 5466
rect 33276 5414 33278 5466
rect 33032 5412 33038 5414
rect 33094 5412 33118 5414
rect 33174 5412 33198 5414
rect 33254 5412 33278 5414
rect 33334 5412 33340 5414
rect 33032 5403 33340 5412
rect 33032 4380 33340 4389
rect 33032 4378 33038 4380
rect 33094 4378 33118 4380
rect 33174 4378 33198 4380
rect 33254 4378 33278 4380
rect 33334 4378 33340 4380
rect 33094 4326 33096 4378
rect 33276 4326 33278 4378
rect 33032 4324 33038 4326
rect 33094 4324 33118 4326
rect 33174 4324 33198 4326
rect 33254 4324 33278 4326
rect 33334 4324 33340 4326
rect 33032 4315 33340 4324
rect 33032 3292 33340 3301
rect 33032 3290 33038 3292
rect 33094 3290 33118 3292
rect 33174 3290 33198 3292
rect 33254 3290 33278 3292
rect 33334 3290 33340 3292
rect 33094 3238 33096 3290
rect 33276 3238 33278 3290
rect 33032 3236 33038 3238
rect 33094 3236 33118 3238
rect 33174 3236 33198 3238
rect 33254 3236 33278 3238
rect 33334 3236 33340 3238
rect 33032 3227 33340 3236
rect 32956 2304 33008 2310
rect 32956 2246 33008 2252
rect 33032 2204 33340 2213
rect 33032 2202 33038 2204
rect 33094 2202 33118 2204
rect 33174 2202 33198 2204
rect 33254 2202 33278 2204
rect 33334 2202 33340 2204
rect 33094 2150 33096 2202
rect 33276 2150 33278 2202
rect 33032 2148 33038 2150
rect 33094 2148 33118 2150
rect 33174 2148 33198 2150
rect 33254 2148 33278 2150
rect 33334 2148 33340 2150
rect 33032 2139 33340 2148
rect 34164 1834 34192 8434
rect 34624 8362 34652 9840
rect 34612 8356 34664 8362
rect 34612 8298 34664 8304
rect 34900 8090 34928 9840
rect 34980 8832 35032 8838
rect 34980 8774 35032 8780
rect 34992 8430 35020 8774
rect 35176 8634 35204 9840
rect 35256 8900 35308 8906
rect 35256 8842 35308 8848
rect 35164 8628 35216 8634
rect 35164 8570 35216 8576
rect 35268 8498 35296 8842
rect 35452 8566 35480 9840
rect 35440 8560 35492 8566
rect 35440 8502 35492 8508
rect 35256 8492 35308 8498
rect 35256 8434 35308 8440
rect 34980 8424 35032 8430
rect 34980 8366 35032 8372
rect 35728 8362 35756 9840
rect 35716 8356 35768 8362
rect 35716 8298 35768 8304
rect 36004 8090 36032 9840
rect 36084 8900 36136 8906
rect 36084 8842 36136 8848
rect 34888 8084 34940 8090
rect 34888 8026 34940 8032
rect 35992 8084 36044 8090
rect 35992 8026 36044 8032
rect 34612 7948 34664 7954
rect 34612 7890 34664 7896
rect 34520 7812 34572 7818
rect 34520 7754 34572 7760
rect 34532 4826 34560 7754
rect 34520 4820 34572 4826
rect 34520 4762 34572 4768
rect 34520 4616 34572 4622
rect 34520 4558 34572 4564
rect 34152 1828 34204 1834
rect 34152 1770 34204 1776
rect 34532 1358 34560 4558
rect 34624 3670 34652 7890
rect 35440 7880 35492 7886
rect 35440 7822 35492 7828
rect 35452 4690 35480 7822
rect 35992 7812 36044 7818
rect 35992 7754 36044 7760
rect 35440 4684 35492 4690
rect 35440 4626 35492 4632
rect 34612 3664 34664 3670
rect 34612 3606 34664 3612
rect 35256 3052 35308 3058
rect 35256 2994 35308 3000
rect 35268 1358 35296 2994
rect 36004 2990 36032 7754
rect 36096 3738 36124 8842
rect 36280 8786 36308 9840
rect 36280 8758 36400 8786
rect 36372 8090 36400 8758
rect 36452 8492 36504 8498
rect 36452 8434 36504 8440
rect 36360 8084 36412 8090
rect 36360 8026 36412 8032
rect 36268 7948 36320 7954
rect 36268 7890 36320 7896
rect 36280 5030 36308 7890
rect 36268 5024 36320 5030
rect 36268 4966 36320 4972
rect 36464 4554 36492 8434
rect 36556 8430 36584 9840
rect 36636 9240 36688 9246
rect 36636 9182 36688 9188
rect 36648 8634 36676 9182
rect 36832 8838 36860 9840
rect 36820 8832 36872 8838
rect 36820 8774 36872 8780
rect 36636 8628 36688 8634
rect 36636 8570 36688 8576
rect 36544 8424 36596 8430
rect 36544 8366 36596 8372
rect 37108 8242 37136 9840
rect 37108 8214 37320 8242
rect 37292 8022 37320 8214
rect 37384 8090 37412 9840
rect 37556 9648 37608 9654
rect 37556 9590 37608 9596
rect 37464 9104 37516 9110
rect 37464 9046 37516 9052
rect 37476 8634 37504 9046
rect 37568 8634 37596 9590
rect 37464 8628 37516 8634
rect 37464 8570 37516 8576
rect 37556 8628 37608 8634
rect 37556 8570 37608 8576
rect 37660 8498 37688 9840
rect 37936 9058 37964 9840
rect 38212 9738 38240 9840
rect 38120 9710 38240 9738
rect 37936 9030 38056 9058
rect 37648 8492 37700 8498
rect 37648 8434 37700 8440
rect 38028 8294 38056 9030
rect 38016 8288 38068 8294
rect 38016 8230 38068 8236
rect 37372 8084 37424 8090
rect 37372 8026 37424 8032
rect 37280 8016 37332 8022
rect 37280 7958 37332 7964
rect 37464 7744 37516 7750
rect 37464 7686 37516 7692
rect 37280 7336 37332 7342
rect 37280 7278 37332 7284
rect 36452 4548 36504 4554
rect 36452 4490 36504 4496
rect 37292 3738 37320 7278
rect 37476 5370 37504 7686
rect 38120 6866 38148 9710
rect 38488 8344 38516 9840
rect 38660 8832 38712 8838
rect 38660 8774 38712 8780
rect 38764 8786 38792 9840
rect 39040 9812 39160 9840
rect 39028 8900 39080 8906
rect 39028 8842 39080 8848
rect 38672 8566 38700 8774
rect 38764 8758 38884 8786
rect 38660 8560 38712 8566
rect 38660 8502 38712 8508
rect 38488 8316 38792 8344
rect 38379 8188 38687 8197
rect 38379 8186 38385 8188
rect 38441 8186 38465 8188
rect 38521 8186 38545 8188
rect 38601 8186 38625 8188
rect 38681 8186 38687 8188
rect 38441 8134 38443 8186
rect 38623 8134 38625 8186
rect 38379 8132 38385 8134
rect 38441 8132 38465 8134
rect 38521 8132 38545 8134
rect 38601 8132 38625 8134
rect 38681 8132 38687 8134
rect 38379 8123 38687 8132
rect 38764 8090 38792 8316
rect 38856 8090 38884 8758
rect 39040 8498 39068 8842
rect 39224 8566 39252 9846
rect 39302 9840 39358 10000
rect 39578 9840 39634 10000
rect 39684 9846 39988 9874
rect 39684 9840 39712 9846
rect 39316 8634 39344 9840
rect 39592 9812 39712 9840
rect 39304 8628 39356 8634
rect 39304 8570 39356 8576
rect 39212 8560 39264 8566
rect 39212 8502 39264 8508
rect 39028 8492 39080 8498
rect 39028 8434 39080 8440
rect 39304 8492 39356 8498
rect 39304 8434 39356 8440
rect 38752 8084 38804 8090
rect 38752 8026 38804 8032
rect 38844 8084 38896 8090
rect 38844 8026 38896 8032
rect 38200 7880 38252 7886
rect 38200 7822 38252 7828
rect 38108 6860 38160 6866
rect 38108 6802 38160 6808
rect 37464 5364 37516 5370
rect 37464 5306 37516 5312
rect 37648 5228 37700 5234
rect 37648 5170 37700 5176
rect 37660 4826 37688 5170
rect 38212 4826 38240 7822
rect 38292 7812 38344 7818
rect 38292 7754 38344 7760
rect 38304 7342 38332 7754
rect 38292 7336 38344 7342
rect 38292 7278 38344 7284
rect 38379 7100 38687 7109
rect 38379 7098 38385 7100
rect 38441 7098 38465 7100
rect 38521 7098 38545 7100
rect 38601 7098 38625 7100
rect 38681 7098 38687 7100
rect 38441 7046 38443 7098
rect 38623 7046 38625 7098
rect 38379 7044 38385 7046
rect 38441 7044 38465 7046
rect 38521 7044 38545 7046
rect 38601 7044 38625 7046
rect 38681 7044 38687 7046
rect 38379 7035 38687 7044
rect 38379 6012 38687 6021
rect 38379 6010 38385 6012
rect 38441 6010 38465 6012
rect 38521 6010 38545 6012
rect 38601 6010 38625 6012
rect 38681 6010 38687 6012
rect 38441 5958 38443 6010
rect 38623 5958 38625 6010
rect 38379 5956 38385 5958
rect 38441 5956 38465 5958
rect 38521 5956 38545 5958
rect 38601 5956 38625 5958
rect 38681 5956 38687 5958
rect 38379 5947 38687 5956
rect 38379 4924 38687 4933
rect 38379 4922 38385 4924
rect 38441 4922 38465 4924
rect 38521 4922 38545 4924
rect 38601 4922 38625 4924
rect 38681 4922 38687 4924
rect 38441 4870 38443 4922
rect 38623 4870 38625 4922
rect 38379 4868 38385 4870
rect 38441 4868 38465 4870
rect 38521 4868 38545 4870
rect 38601 4868 38625 4870
rect 38681 4868 38687 4870
rect 38379 4859 38687 4868
rect 37648 4820 37700 4826
rect 37648 4762 37700 4768
rect 38200 4820 38252 4826
rect 38200 4762 38252 4768
rect 39316 4758 39344 8434
rect 39960 8242 39988 9846
rect 43726 8732 44034 8741
rect 43726 8730 43732 8732
rect 43788 8730 43812 8732
rect 43868 8730 43892 8732
rect 43948 8730 43972 8732
rect 44028 8730 44034 8732
rect 43788 8678 43790 8730
rect 43970 8678 43972 8730
rect 43726 8676 43732 8678
rect 43788 8676 43812 8678
rect 43868 8676 43892 8678
rect 43948 8676 43972 8678
rect 44028 8676 44034 8678
rect 43726 8667 44034 8676
rect 40500 8492 40552 8498
rect 40500 8434 40552 8440
rect 41052 8492 41104 8498
rect 41052 8434 41104 8440
rect 39960 8214 40080 8242
rect 40052 8090 40080 8214
rect 40040 8084 40092 8090
rect 40040 8026 40092 8032
rect 39856 7880 39908 7886
rect 39856 7822 39908 7828
rect 39396 7744 39448 7750
rect 39396 7686 39448 7692
rect 39408 6866 39436 7686
rect 39396 6860 39448 6866
rect 39396 6802 39448 6808
rect 39304 4752 39356 4758
rect 39304 4694 39356 4700
rect 38384 4616 38436 4622
rect 38384 4558 38436 4564
rect 38396 4282 38424 4558
rect 38384 4276 38436 4282
rect 38384 4218 38436 4224
rect 37372 4140 37424 4146
rect 37372 4082 37424 4088
rect 36084 3732 36136 3738
rect 36084 3674 36136 3680
rect 37280 3732 37332 3738
rect 37280 3674 37332 3680
rect 35992 2984 36044 2990
rect 35992 2926 36044 2932
rect 24860 1352 24912 1358
rect 24860 1294 24912 1300
rect 26700 1352 26752 1358
rect 26700 1294 26752 1300
rect 27436 1352 27488 1358
rect 27436 1294 27488 1300
rect 28908 1352 28960 1358
rect 28908 1294 28960 1300
rect 29092 1352 29144 1358
rect 29092 1294 29144 1300
rect 31208 1352 31260 1358
rect 31208 1294 31260 1300
rect 31668 1352 31720 1358
rect 31668 1294 31720 1300
rect 33324 1352 33376 1358
rect 34520 1352 34572 1358
rect 33376 1300 33456 1306
rect 33324 1294 33456 1300
rect 34520 1294 34572 1300
rect 35256 1352 35308 1358
rect 35256 1294 35308 1300
rect 35440 1352 35492 1358
rect 35440 1294 35492 1300
rect 24768 1284 24820 1290
rect 24768 1226 24820 1232
rect 22466 54 22784 82
rect 24582 82 24638 160
rect 24872 82 24900 1294
rect 26712 160 26740 1294
rect 24582 54 24900 82
rect 3422 0 3478 54
rect 5538 0 5594 54
rect 7654 0 7710 54
rect 9770 0 9826 54
rect 11886 0 11942 54
rect 14002 0 14058 54
rect 16118 0 16174 54
rect 18234 0 18290 54
rect 20350 0 20406 54
rect 22466 0 22522 54
rect 24582 0 24638 54
rect 26698 0 26754 160
rect 28814 82 28870 160
rect 29104 82 29132 1294
rect 28814 54 29132 82
rect 30930 82 30986 160
rect 31220 82 31248 1294
rect 33336 1278 33456 1294
rect 33032 1116 33340 1125
rect 33032 1114 33038 1116
rect 33094 1114 33118 1116
rect 33174 1114 33198 1116
rect 33254 1114 33278 1116
rect 33334 1114 33340 1116
rect 33094 1062 33096 1114
rect 33276 1062 33278 1114
rect 33032 1060 33038 1062
rect 33094 1060 33118 1062
rect 33174 1060 33198 1062
rect 33254 1060 33278 1062
rect 33334 1060 33340 1062
rect 33032 1051 33340 1060
rect 30930 54 31248 82
rect 33046 82 33102 160
rect 33428 82 33456 1278
rect 33046 54 33456 82
rect 35162 82 35218 160
rect 35452 82 35480 1294
rect 37384 1222 37412 4082
rect 38379 3836 38687 3845
rect 38379 3834 38385 3836
rect 38441 3834 38465 3836
rect 38521 3834 38545 3836
rect 38601 3834 38625 3836
rect 38681 3834 38687 3836
rect 38441 3782 38443 3834
rect 38623 3782 38625 3834
rect 38379 3780 38385 3782
rect 38441 3780 38465 3782
rect 38521 3780 38545 3782
rect 38601 3780 38625 3782
rect 38681 3780 38687 3782
rect 38379 3771 38687 3780
rect 37464 3528 37516 3534
rect 37464 3470 37516 3476
rect 37476 3194 37504 3470
rect 37464 3188 37516 3194
rect 37464 3130 37516 3136
rect 38379 2748 38687 2757
rect 38379 2746 38385 2748
rect 38441 2746 38465 2748
rect 38521 2746 38545 2748
rect 38601 2746 38625 2748
rect 38681 2746 38687 2748
rect 38441 2694 38443 2746
rect 38623 2694 38625 2746
rect 38379 2692 38385 2694
rect 38441 2692 38465 2694
rect 38521 2692 38545 2694
rect 38601 2692 38625 2694
rect 38681 2692 38687 2694
rect 38379 2683 38687 2692
rect 39868 2650 39896 7822
rect 40132 3528 40184 3534
rect 40132 3470 40184 3476
rect 40144 3194 40172 3470
rect 40132 3188 40184 3194
rect 40132 3130 40184 3136
rect 40512 2650 40540 8434
rect 41064 3738 41092 8434
rect 43726 7644 44034 7653
rect 43726 7642 43732 7644
rect 43788 7642 43812 7644
rect 43868 7642 43892 7644
rect 43948 7642 43972 7644
rect 44028 7642 44034 7644
rect 43788 7590 43790 7642
rect 43970 7590 43972 7642
rect 43726 7588 43732 7590
rect 43788 7588 43812 7590
rect 43868 7588 43892 7590
rect 43948 7588 43972 7590
rect 44028 7588 44034 7590
rect 43726 7579 44034 7588
rect 43726 6556 44034 6565
rect 43726 6554 43732 6556
rect 43788 6554 43812 6556
rect 43868 6554 43892 6556
rect 43948 6554 43972 6556
rect 44028 6554 44034 6556
rect 43788 6502 43790 6554
rect 43970 6502 43972 6554
rect 43726 6500 43732 6502
rect 43788 6500 43812 6502
rect 43868 6500 43892 6502
rect 43948 6500 43972 6502
rect 44028 6500 44034 6502
rect 43726 6491 44034 6500
rect 43726 5468 44034 5477
rect 43726 5466 43732 5468
rect 43788 5466 43812 5468
rect 43868 5466 43892 5468
rect 43948 5466 43972 5468
rect 44028 5466 44034 5468
rect 43788 5414 43790 5466
rect 43970 5414 43972 5466
rect 43726 5412 43732 5414
rect 43788 5412 43812 5414
rect 43868 5412 43892 5414
rect 43948 5412 43972 5414
rect 44028 5412 44034 5414
rect 43726 5403 44034 5412
rect 43726 4380 44034 4389
rect 43726 4378 43732 4380
rect 43788 4378 43812 4380
rect 43868 4378 43892 4380
rect 43948 4378 43972 4380
rect 44028 4378 44034 4380
rect 43788 4326 43790 4378
rect 43970 4326 43972 4378
rect 43726 4324 43732 4326
rect 43788 4324 43812 4326
rect 43868 4324 43892 4326
rect 43948 4324 43972 4326
rect 44028 4324 44034 4326
rect 43726 4315 44034 4324
rect 41052 3732 41104 3738
rect 41052 3674 41104 3680
rect 43726 3292 44034 3301
rect 43726 3290 43732 3292
rect 43788 3290 43812 3292
rect 43868 3290 43892 3292
rect 43948 3290 43972 3292
rect 44028 3290 44034 3292
rect 43788 3238 43790 3290
rect 43970 3238 43972 3290
rect 43726 3236 43732 3238
rect 43788 3236 43812 3238
rect 43868 3236 43892 3238
rect 43948 3236 43972 3238
rect 44028 3236 44034 3238
rect 43726 3227 44034 3236
rect 40868 3052 40920 3058
rect 40868 2994 40920 3000
rect 39856 2644 39908 2650
rect 39856 2586 39908 2592
rect 40500 2644 40552 2650
rect 40500 2586 40552 2592
rect 39120 2440 39172 2446
rect 39120 2382 39172 2388
rect 40040 2440 40092 2446
rect 40040 2382 40092 2388
rect 39132 2106 39160 2382
rect 40052 2106 40080 2382
rect 39120 2100 39172 2106
rect 39120 2042 39172 2048
rect 40040 2100 40092 2106
rect 40040 2042 40092 2048
rect 39396 1964 39448 1970
rect 39396 1906 39448 1912
rect 38379 1660 38687 1669
rect 38379 1658 38385 1660
rect 38441 1658 38465 1660
rect 38521 1658 38545 1660
rect 38601 1658 38625 1660
rect 38681 1658 38687 1660
rect 38441 1606 38443 1658
rect 38623 1606 38625 1658
rect 38379 1604 38385 1606
rect 38441 1604 38465 1606
rect 38521 1604 38545 1606
rect 38601 1604 38625 1606
rect 38681 1604 38687 1606
rect 38379 1595 38687 1604
rect 39408 1562 39436 1906
rect 39396 1556 39448 1562
rect 39396 1498 39448 1504
rect 40880 1358 40908 2994
rect 43726 2204 44034 2213
rect 43726 2202 43732 2204
rect 43788 2202 43812 2204
rect 43868 2202 43892 2204
rect 43948 2202 43972 2204
rect 44028 2202 44034 2204
rect 43788 2150 43790 2202
rect 43970 2150 43972 2202
rect 43726 2148 43732 2150
rect 43788 2148 43812 2150
rect 43868 2148 43892 2150
rect 43948 2148 43972 2150
rect 44028 2148 44034 2150
rect 43726 2139 44034 2148
rect 43352 1964 43404 1970
rect 43352 1906 43404 1912
rect 43364 1562 43392 1906
rect 43352 1556 43404 1562
rect 43352 1498 43404 1504
rect 37556 1352 37608 1358
rect 37556 1294 37608 1300
rect 39396 1352 39448 1358
rect 39396 1294 39448 1300
rect 40868 1352 40920 1358
rect 40868 1294 40920 1300
rect 41788 1352 41840 1358
rect 41788 1294 41840 1300
rect 43536 1352 43588 1358
rect 43536 1294 43588 1300
rect 37372 1216 37424 1222
rect 37372 1158 37424 1164
rect 35162 54 35480 82
rect 37278 82 37334 160
rect 37568 82 37596 1294
rect 39408 160 39436 1294
rect 37278 54 37596 82
rect 28814 0 28870 54
rect 30930 0 30986 54
rect 33046 0 33102 54
rect 35162 0 35218 54
rect 37278 0 37334 54
rect 39394 0 39450 160
rect 41510 82 41566 160
rect 41800 82 41828 1294
rect 41510 54 41828 82
rect 43548 82 43576 1294
rect 43726 1116 44034 1125
rect 43726 1114 43732 1116
rect 43788 1114 43812 1116
rect 43868 1114 43892 1116
rect 43948 1114 43972 1116
rect 44028 1114 44034 1116
rect 43788 1062 43790 1114
rect 43970 1062 43972 1114
rect 43726 1060 43732 1062
rect 43788 1060 43812 1062
rect 43868 1060 43892 1062
rect 43948 1060 43972 1062
rect 44028 1060 44034 1062
rect 43726 1051 44034 1060
rect 43626 82 43682 160
rect 43548 54 43682 82
rect 41510 0 41566 54
rect 43626 0 43682 54
<< via2 >>
rect 4894 9016 4950 9072
rect 6303 8186 6359 8188
rect 6383 8186 6439 8188
rect 6463 8186 6519 8188
rect 6543 8186 6599 8188
rect 6303 8134 6349 8186
rect 6349 8134 6359 8186
rect 6383 8134 6413 8186
rect 6413 8134 6425 8186
rect 6425 8134 6439 8186
rect 6463 8134 6477 8186
rect 6477 8134 6489 8186
rect 6489 8134 6519 8186
rect 6543 8134 6553 8186
rect 6553 8134 6599 8186
rect 6303 8132 6359 8134
rect 6383 8132 6439 8134
rect 6463 8132 6519 8134
rect 6543 8132 6599 8134
rect 6734 7812 6790 7848
rect 6734 7792 6736 7812
rect 6736 7792 6788 7812
rect 6788 7792 6790 7812
rect 6550 7248 6606 7304
rect 6303 7098 6359 7100
rect 6383 7098 6439 7100
rect 6463 7098 6519 7100
rect 6543 7098 6599 7100
rect 6303 7046 6349 7098
rect 6349 7046 6359 7098
rect 6383 7046 6413 7098
rect 6413 7046 6425 7098
rect 6425 7046 6439 7098
rect 6463 7046 6477 7098
rect 6477 7046 6489 7098
rect 6489 7046 6519 7098
rect 6543 7046 6553 7098
rect 6553 7046 6599 7098
rect 6303 7044 6359 7046
rect 6383 7044 6439 7046
rect 6463 7044 6519 7046
rect 6543 7044 6599 7046
rect 7470 6740 7472 6760
rect 7472 6740 7524 6760
rect 7524 6740 7526 6760
rect 7470 6704 7526 6740
rect 7010 6296 7066 6352
rect 8022 6160 8078 6216
rect 6303 6010 6359 6012
rect 6383 6010 6439 6012
rect 6463 6010 6519 6012
rect 6543 6010 6599 6012
rect 6303 5958 6349 6010
rect 6349 5958 6359 6010
rect 6383 5958 6413 6010
rect 6413 5958 6425 6010
rect 6425 5958 6439 6010
rect 6463 5958 6477 6010
rect 6477 5958 6489 6010
rect 6489 5958 6519 6010
rect 6543 5958 6553 6010
rect 6553 5958 6599 6010
rect 6303 5956 6359 5958
rect 6383 5956 6439 5958
rect 6463 5956 6519 5958
rect 6543 5956 6599 5958
rect 9586 7384 9642 7440
rect 11650 8730 11706 8732
rect 11730 8730 11786 8732
rect 11810 8730 11866 8732
rect 11890 8730 11946 8732
rect 11650 8678 11696 8730
rect 11696 8678 11706 8730
rect 11730 8678 11760 8730
rect 11760 8678 11772 8730
rect 11772 8678 11786 8730
rect 11810 8678 11824 8730
rect 11824 8678 11836 8730
rect 11836 8678 11866 8730
rect 11890 8678 11900 8730
rect 11900 8678 11946 8730
rect 11650 8676 11706 8678
rect 11730 8676 11786 8678
rect 11810 8676 11866 8678
rect 11890 8676 11946 8678
rect 11650 7642 11706 7644
rect 11730 7642 11786 7644
rect 11810 7642 11866 7644
rect 11890 7642 11946 7644
rect 11650 7590 11696 7642
rect 11696 7590 11706 7642
rect 11730 7590 11760 7642
rect 11760 7590 11772 7642
rect 11772 7590 11786 7642
rect 11810 7590 11824 7642
rect 11824 7590 11836 7642
rect 11836 7590 11866 7642
rect 11890 7590 11900 7642
rect 11900 7590 11946 7642
rect 11650 7588 11706 7590
rect 11730 7588 11786 7590
rect 11810 7588 11866 7590
rect 11890 7588 11946 7590
rect 12714 9152 12770 9208
rect 11650 6554 11706 6556
rect 11730 6554 11786 6556
rect 11810 6554 11866 6556
rect 11890 6554 11946 6556
rect 11650 6502 11696 6554
rect 11696 6502 11706 6554
rect 11730 6502 11760 6554
rect 11760 6502 11772 6554
rect 11772 6502 11786 6554
rect 11810 6502 11824 6554
rect 11824 6502 11836 6554
rect 11836 6502 11866 6554
rect 11890 6502 11900 6554
rect 11900 6502 11946 6554
rect 11650 6500 11706 6502
rect 11730 6500 11786 6502
rect 11810 6500 11866 6502
rect 11890 6500 11946 6502
rect 12990 7928 13046 7984
rect 17130 9424 17186 9480
rect 15106 7656 15162 7712
rect 14830 6568 14886 6624
rect 15566 6840 15622 6896
rect 16997 8186 17053 8188
rect 17077 8186 17133 8188
rect 17157 8186 17213 8188
rect 17237 8186 17293 8188
rect 16997 8134 17043 8186
rect 17043 8134 17053 8186
rect 17077 8134 17107 8186
rect 17107 8134 17119 8186
rect 17119 8134 17133 8186
rect 17157 8134 17171 8186
rect 17171 8134 17183 8186
rect 17183 8134 17213 8186
rect 17237 8134 17247 8186
rect 17247 8134 17293 8186
rect 16997 8132 17053 8134
rect 17077 8132 17133 8134
rect 17157 8132 17213 8134
rect 17237 8132 17293 8134
rect 18694 8744 18750 8800
rect 19062 9308 19118 9344
rect 19062 9288 19064 9308
rect 19064 9288 19116 9308
rect 19116 9288 19118 9308
rect 17958 7828 17960 7848
rect 17960 7828 18012 7848
rect 18012 7828 18014 7848
rect 17958 7792 18014 7828
rect 18234 8472 18290 8528
rect 16997 7098 17053 7100
rect 17077 7098 17133 7100
rect 17157 7098 17213 7100
rect 17237 7098 17293 7100
rect 16997 7046 17043 7098
rect 17043 7046 17053 7098
rect 17077 7046 17107 7098
rect 17107 7046 17119 7098
rect 17119 7046 17133 7098
rect 17157 7046 17171 7098
rect 17171 7046 17183 7098
rect 17183 7046 17213 7098
rect 17237 7046 17247 7098
rect 17247 7046 17293 7098
rect 16997 7044 17053 7046
rect 17077 7044 17133 7046
rect 17157 7044 17213 7046
rect 17237 7044 17293 7046
rect 18602 8200 18658 8256
rect 18786 8336 18842 8392
rect 20074 9832 20130 9888
rect 20166 9324 20168 9344
rect 20168 9324 20220 9344
rect 20220 9324 20222 9344
rect 19706 8200 19762 8256
rect 20166 9288 20222 9324
rect 20442 8744 20498 8800
rect 20074 7656 20130 7712
rect 20166 7520 20222 7576
rect 16997 6010 17053 6012
rect 17077 6010 17133 6012
rect 17157 6010 17213 6012
rect 17237 6010 17293 6012
rect 16997 5958 17043 6010
rect 17043 5958 17053 6010
rect 17077 5958 17107 6010
rect 17107 5958 17119 6010
rect 17119 5958 17133 6010
rect 17157 5958 17171 6010
rect 17171 5958 17183 6010
rect 17183 5958 17213 6010
rect 17237 5958 17247 6010
rect 17247 5958 17293 6010
rect 16997 5956 17053 5958
rect 17077 5956 17133 5958
rect 17157 5956 17213 5958
rect 17237 5956 17293 5958
rect 20718 8200 20774 8256
rect 21546 9424 21602 9480
rect 21914 9016 21970 9072
rect 19614 7268 19670 7304
rect 19614 7248 19616 7268
rect 19616 7248 19668 7268
rect 19668 7248 19670 7268
rect 20166 7248 20222 7304
rect 20166 7148 20168 7168
rect 20168 7148 20220 7168
rect 20220 7148 20222 7168
rect 20166 7112 20222 7148
rect 19982 6976 20038 7032
rect 20258 6976 20314 7032
rect 21362 6704 21418 6760
rect 21454 6568 21510 6624
rect 22344 8730 22400 8732
rect 22424 8730 22480 8732
rect 22504 8730 22560 8732
rect 22584 8730 22640 8732
rect 22344 8678 22390 8730
rect 22390 8678 22400 8730
rect 22424 8678 22454 8730
rect 22454 8678 22466 8730
rect 22466 8678 22480 8730
rect 22504 8678 22518 8730
rect 22518 8678 22530 8730
rect 22530 8678 22560 8730
rect 22584 8678 22594 8730
rect 22594 8678 22640 8730
rect 22344 8676 22400 8678
rect 22424 8676 22480 8678
rect 22504 8676 22560 8678
rect 22584 8676 22640 8678
rect 22190 8336 22246 8392
rect 22006 7404 22062 7440
rect 22006 7384 22008 7404
rect 22008 7384 22060 7404
rect 22060 7384 22062 7404
rect 22344 7642 22400 7644
rect 22424 7642 22480 7644
rect 22504 7642 22560 7644
rect 22584 7642 22640 7644
rect 22344 7590 22390 7642
rect 22390 7590 22400 7642
rect 22424 7590 22454 7642
rect 22454 7590 22466 7642
rect 22466 7590 22480 7642
rect 22504 7590 22518 7642
rect 22518 7590 22530 7642
rect 22530 7590 22560 7642
rect 22584 7590 22594 7642
rect 22594 7590 22640 7642
rect 22344 7588 22400 7590
rect 22424 7588 22480 7590
rect 22504 7588 22560 7590
rect 22584 7588 22640 7590
rect 22834 6840 22890 6896
rect 22344 6554 22400 6556
rect 22424 6554 22480 6556
rect 22504 6554 22560 6556
rect 22584 6554 22640 6556
rect 22344 6502 22390 6554
rect 22390 6502 22400 6554
rect 22424 6502 22454 6554
rect 22454 6502 22466 6554
rect 22466 6502 22480 6554
rect 22504 6502 22518 6554
rect 22518 6502 22530 6554
rect 22530 6502 22560 6554
rect 22584 6502 22594 6554
rect 22594 6502 22640 6554
rect 22344 6500 22400 6502
rect 22424 6500 22480 6502
rect 22504 6500 22560 6502
rect 22584 6500 22640 6502
rect 22098 6160 22154 6216
rect 8206 5752 8262 5808
rect 24030 7792 24086 7848
rect 24674 8200 24730 8256
rect 25502 8084 25558 8120
rect 25502 8064 25504 8084
rect 25504 8064 25556 8084
rect 25556 8064 25558 8084
rect 26882 9052 26884 9072
rect 26884 9052 26936 9072
rect 26936 9052 26938 9072
rect 26882 9016 26938 9052
rect 27250 9152 27306 9208
rect 27342 7928 27398 7984
rect 24858 7248 24914 7304
rect 23754 6296 23810 6352
rect 27691 8186 27747 8188
rect 27771 8186 27827 8188
rect 27851 8186 27907 8188
rect 27931 8186 27987 8188
rect 27691 8134 27737 8186
rect 27737 8134 27747 8186
rect 27771 8134 27801 8186
rect 27801 8134 27813 8186
rect 27813 8134 27827 8186
rect 27851 8134 27865 8186
rect 27865 8134 27877 8186
rect 27877 8134 27907 8186
rect 27931 8134 27941 8186
rect 27941 8134 27987 8186
rect 27691 8132 27747 8134
rect 27771 8132 27827 8134
rect 27851 8132 27907 8134
rect 27931 8132 27987 8134
rect 27691 7098 27747 7100
rect 27771 7098 27827 7100
rect 27851 7098 27907 7100
rect 27931 7098 27987 7100
rect 27691 7046 27737 7098
rect 27737 7046 27747 7098
rect 27771 7046 27801 7098
rect 27801 7046 27813 7098
rect 27813 7046 27827 7098
rect 27851 7046 27865 7098
rect 27865 7046 27877 7098
rect 27877 7046 27907 7098
rect 27931 7046 27941 7098
rect 27941 7046 27987 7098
rect 27691 7044 27747 7046
rect 27771 7044 27827 7046
rect 27851 7044 27907 7046
rect 27931 7044 27987 7046
rect 27691 6010 27747 6012
rect 27771 6010 27827 6012
rect 27851 6010 27907 6012
rect 27931 6010 27987 6012
rect 27691 5958 27737 6010
rect 27737 5958 27747 6010
rect 27771 5958 27801 6010
rect 27801 5958 27813 6010
rect 27813 5958 27827 6010
rect 27851 5958 27865 6010
rect 27865 5958 27877 6010
rect 27877 5958 27907 6010
rect 27931 5958 27941 6010
rect 27941 5958 27987 6010
rect 27691 5956 27747 5958
rect 27771 5956 27827 5958
rect 27851 5956 27907 5958
rect 27931 5956 27987 5958
rect 23478 5752 23534 5808
rect 11650 5466 11706 5468
rect 11730 5466 11786 5468
rect 11810 5466 11866 5468
rect 11890 5466 11946 5468
rect 11650 5414 11696 5466
rect 11696 5414 11706 5466
rect 11730 5414 11760 5466
rect 11760 5414 11772 5466
rect 11772 5414 11786 5466
rect 11810 5414 11824 5466
rect 11824 5414 11836 5466
rect 11836 5414 11866 5466
rect 11890 5414 11900 5466
rect 11900 5414 11946 5466
rect 11650 5412 11706 5414
rect 11730 5412 11786 5414
rect 11810 5412 11866 5414
rect 11890 5412 11946 5414
rect 22344 5466 22400 5468
rect 22424 5466 22480 5468
rect 22504 5466 22560 5468
rect 22584 5466 22640 5468
rect 22344 5414 22390 5466
rect 22390 5414 22400 5466
rect 22424 5414 22454 5466
rect 22454 5414 22466 5466
rect 22466 5414 22480 5466
rect 22504 5414 22518 5466
rect 22518 5414 22530 5466
rect 22530 5414 22560 5466
rect 22584 5414 22594 5466
rect 22594 5414 22640 5466
rect 22344 5412 22400 5414
rect 22424 5412 22480 5414
rect 22504 5412 22560 5414
rect 22584 5412 22640 5414
rect 6303 4922 6359 4924
rect 6383 4922 6439 4924
rect 6463 4922 6519 4924
rect 6543 4922 6599 4924
rect 6303 4870 6349 4922
rect 6349 4870 6359 4922
rect 6383 4870 6413 4922
rect 6413 4870 6425 4922
rect 6425 4870 6439 4922
rect 6463 4870 6477 4922
rect 6477 4870 6489 4922
rect 6489 4870 6519 4922
rect 6543 4870 6553 4922
rect 6553 4870 6599 4922
rect 6303 4868 6359 4870
rect 6383 4868 6439 4870
rect 6463 4868 6519 4870
rect 6543 4868 6599 4870
rect 16997 4922 17053 4924
rect 17077 4922 17133 4924
rect 17157 4922 17213 4924
rect 17237 4922 17293 4924
rect 16997 4870 17043 4922
rect 17043 4870 17053 4922
rect 17077 4870 17107 4922
rect 17107 4870 17119 4922
rect 17119 4870 17133 4922
rect 17157 4870 17171 4922
rect 17171 4870 17183 4922
rect 17183 4870 17213 4922
rect 17237 4870 17247 4922
rect 17247 4870 17293 4922
rect 16997 4868 17053 4870
rect 17077 4868 17133 4870
rect 17157 4868 17213 4870
rect 17237 4868 17293 4870
rect 27691 4922 27747 4924
rect 27771 4922 27827 4924
rect 27851 4922 27907 4924
rect 27931 4922 27987 4924
rect 27691 4870 27737 4922
rect 27737 4870 27747 4922
rect 27771 4870 27801 4922
rect 27801 4870 27813 4922
rect 27813 4870 27827 4922
rect 27851 4870 27865 4922
rect 27865 4870 27877 4922
rect 27877 4870 27907 4922
rect 27931 4870 27941 4922
rect 27941 4870 27987 4922
rect 27691 4868 27747 4870
rect 27771 4868 27827 4870
rect 27851 4868 27907 4870
rect 27931 4868 27987 4870
rect 11650 4378 11706 4380
rect 11730 4378 11786 4380
rect 11810 4378 11866 4380
rect 11890 4378 11946 4380
rect 11650 4326 11696 4378
rect 11696 4326 11706 4378
rect 11730 4326 11760 4378
rect 11760 4326 11772 4378
rect 11772 4326 11786 4378
rect 11810 4326 11824 4378
rect 11824 4326 11836 4378
rect 11836 4326 11866 4378
rect 11890 4326 11900 4378
rect 11900 4326 11946 4378
rect 11650 4324 11706 4326
rect 11730 4324 11786 4326
rect 11810 4324 11866 4326
rect 11890 4324 11946 4326
rect 6303 3834 6359 3836
rect 6383 3834 6439 3836
rect 6463 3834 6519 3836
rect 6543 3834 6599 3836
rect 6303 3782 6349 3834
rect 6349 3782 6359 3834
rect 6383 3782 6413 3834
rect 6413 3782 6425 3834
rect 6425 3782 6439 3834
rect 6463 3782 6477 3834
rect 6477 3782 6489 3834
rect 6489 3782 6519 3834
rect 6543 3782 6553 3834
rect 6553 3782 6599 3834
rect 6303 3780 6359 3782
rect 6383 3780 6439 3782
rect 6463 3780 6519 3782
rect 6543 3780 6599 3782
rect 6303 2746 6359 2748
rect 6383 2746 6439 2748
rect 6463 2746 6519 2748
rect 6543 2746 6599 2748
rect 6303 2694 6349 2746
rect 6349 2694 6359 2746
rect 6383 2694 6413 2746
rect 6413 2694 6425 2746
rect 6425 2694 6439 2746
rect 6463 2694 6477 2746
rect 6477 2694 6489 2746
rect 6489 2694 6519 2746
rect 6543 2694 6553 2746
rect 6553 2694 6599 2746
rect 6303 2692 6359 2694
rect 6383 2692 6439 2694
rect 6463 2692 6519 2694
rect 6543 2692 6599 2694
rect 6303 1658 6359 1660
rect 6383 1658 6439 1660
rect 6463 1658 6519 1660
rect 6543 1658 6599 1660
rect 6303 1606 6349 1658
rect 6349 1606 6359 1658
rect 6383 1606 6413 1658
rect 6413 1606 6425 1658
rect 6425 1606 6439 1658
rect 6463 1606 6477 1658
rect 6477 1606 6489 1658
rect 6489 1606 6519 1658
rect 6543 1606 6553 1658
rect 6553 1606 6599 1658
rect 6303 1604 6359 1606
rect 6383 1604 6439 1606
rect 6463 1604 6519 1606
rect 6543 1604 6599 1606
rect 16997 3834 17053 3836
rect 17077 3834 17133 3836
rect 17157 3834 17213 3836
rect 17237 3834 17293 3836
rect 16997 3782 17043 3834
rect 17043 3782 17053 3834
rect 17077 3782 17107 3834
rect 17107 3782 17119 3834
rect 17119 3782 17133 3834
rect 17157 3782 17171 3834
rect 17171 3782 17183 3834
rect 17183 3782 17213 3834
rect 17237 3782 17247 3834
rect 17247 3782 17293 3834
rect 16997 3780 17053 3782
rect 17077 3780 17133 3782
rect 17157 3780 17213 3782
rect 17237 3780 17293 3782
rect 11650 3290 11706 3292
rect 11730 3290 11786 3292
rect 11810 3290 11866 3292
rect 11890 3290 11946 3292
rect 11650 3238 11696 3290
rect 11696 3238 11706 3290
rect 11730 3238 11760 3290
rect 11760 3238 11772 3290
rect 11772 3238 11786 3290
rect 11810 3238 11824 3290
rect 11824 3238 11836 3290
rect 11836 3238 11866 3290
rect 11890 3238 11900 3290
rect 11900 3238 11946 3290
rect 11650 3236 11706 3238
rect 11730 3236 11786 3238
rect 11810 3236 11866 3238
rect 11890 3236 11946 3238
rect 16997 2746 17053 2748
rect 17077 2746 17133 2748
rect 17157 2746 17213 2748
rect 17237 2746 17293 2748
rect 16997 2694 17043 2746
rect 17043 2694 17053 2746
rect 17077 2694 17107 2746
rect 17107 2694 17119 2746
rect 17119 2694 17133 2746
rect 17157 2694 17171 2746
rect 17171 2694 17183 2746
rect 17183 2694 17213 2746
rect 17237 2694 17247 2746
rect 17247 2694 17293 2746
rect 16997 2692 17053 2694
rect 17077 2692 17133 2694
rect 17157 2692 17213 2694
rect 17237 2692 17293 2694
rect 11650 2202 11706 2204
rect 11730 2202 11786 2204
rect 11810 2202 11866 2204
rect 11890 2202 11946 2204
rect 11650 2150 11696 2202
rect 11696 2150 11706 2202
rect 11730 2150 11760 2202
rect 11760 2150 11772 2202
rect 11772 2150 11786 2202
rect 11810 2150 11824 2202
rect 11824 2150 11836 2202
rect 11836 2150 11866 2202
rect 11890 2150 11900 2202
rect 11900 2150 11946 2202
rect 11650 2148 11706 2150
rect 11730 2148 11786 2150
rect 11810 2148 11866 2150
rect 11890 2148 11946 2150
rect 16997 1658 17053 1660
rect 17077 1658 17133 1660
rect 17157 1658 17213 1660
rect 17237 1658 17293 1660
rect 16997 1606 17043 1658
rect 17043 1606 17053 1658
rect 17077 1606 17107 1658
rect 17107 1606 17119 1658
rect 17119 1606 17133 1658
rect 17157 1606 17171 1658
rect 17171 1606 17183 1658
rect 17183 1606 17213 1658
rect 17237 1606 17247 1658
rect 17247 1606 17293 1658
rect 16997 1604 17053 1606
rect 17077 1604 17133 1606
rect 17157 1604 17213 1606
rect 17237 1604 17293 1606
rect 11650 1114 11706 1116
rect 11730 1114 11786 1116
rect 11810 1114 11866 1116
rect 11890 1114 11946 1116
rect 11650 1062 11696 1114
rect 11696 1062 11706 1114
rect 11730 1062 11760 1114
rect 11760 1062 11772 1114
rect 11772 1062 11786 1114
rect 11810 1062 11824 1114
rect 11824 1062 11836 1114
rect 11836 1062 11866 1114
rect 11890 1062 11900 1114
rect 11900 1062 11946 1114
rect 11650 1060 11706 1062
rect 11730 1060 11786 1062
rect 11810 1060 11866 1062
rect 11890 1060 11946 1062
rect 22344 4378 22400 4380
rect 22424 4378 22480 4380
rect 22504 4378 22560 4380
rect 22584 4378 22640 4380
rect 22344 4326 22390 4378
rect 22390 4326 22400 4378
rect 22424 4326 22454 4378
rect 22454 4326 22466 4378
rect 22466 4326 22480 4378
rect 22504 4326 22518 4378
rect 22518 4326 22530 4378
rect 22530 4326 22560 4378
rect 22584 4326 22594 4378
rect 22594 4326 22640 4378
rect 22344 4324 22400 4326
rect 22424 4324 22480 4326
rect 22504 4324 22560 4326
rect 22584 4324 22640 4326
rect 22344 3290 22400 3292
rect 22424 3290 22480 3292
rect 22504 3290 22560 3292
rect 22584 3290 22640 3292
rect 22344 3238 22390 3290
rect 22390 3238 22400 3290
rect 22424 3238 22454 3290
rect 22454 3238 22466 3290
rect 22466 3238 22480 3290
rect 22504 3238 22518 3290
rect 22518 3238 22530 3290
rect 22530 3238 22560 3290
rect 22584 3238 22594 3290
rect 22594 3238 22640 3290
rect 22344 3236 22400 3238
rect 22424 3236 22480 3238
rect 22504 3236 22560 3238
rect 22584 3236 22640 3238
rect 22344 2202 22400 2204
rect 22424 2202 22480 2204
rect 22504 2202 22560 2204
rect 22584 2202 22640 2204
rect 22344 2150 22390 2202
rect 22390 2150 22400 2202
rect 22424 2150 22454 2202
rect 22454 2150 22466 2202
rect 22466 2150 22480 2202
rect 22504 2150 22518 2202
rect 22518 2150 22530 2202
rect 22530 2150 22560 2202
rect 22584 2150 22594 2202
rect 22594 2150 22640 2202
rect 22344 2148 22400 2150
rect 22424 2148 22480 2150
rect 22504 2148 22560 2150
rect 22584 2148 22640 2150
rect 22344 1114 22400 1116
rect 22424 1114 22480 1116
rect 22504 1114 22560 1116
rect 22584 1114 22640 1116
rect 22344 1062 22390 1114
rect 22390 1062 22400 1114
rect 22424 1062 22454 1114
rect 22454 1062 22466 1114
rect 22466 1062 22480 1114
rect 22504 1062 22518 1114
rect 22518 1062 22530 1114
rect 22530 1062 22560 1114
rect 22584 1062 22594 1114
rect 22594 1062 22640 1114
rect 22344 1060 22400 1062
rect 22424 1060 22480 1062
rect 22504 1060 22560 1062
rect 22584 1060 22640 1062
rect 27691 3834 27747 3836
rect 27771 3834 27827 3836
rect 27851 3834 27907 3836
rect 27931 3834 27987 3836
rect 27691 3782 27737 3834
rect 27737 3782 27747 3834
rect 27771 3782 27801 3834
rect 27801 3782 27813 3834
rect 27813 3782 27827 3834
rect 27851 3782 27865 3834
rect 27865 3782 27877 3834
rect 27877 3782 27907 3834
rect 27931 3782 27941 3834
rect 27941 3782 27987 3834
rect 27691 3780 27747 3782
rect 27771 3780 27827 3782
rect 27851 3780 27907 3782
rect 27931 3780 27987 3782
rect 31942 8472 31998 8528
rect 32218 8880 32274 8936
rect 33038 8730 33094 8732
rect 33118 8730 33174 8732
rect 33198 8730 33254 8732
rect 33278 8730 33334 8732
rect 33038 8678 33084 8730
rect 33084 8678 33094 8730
rect 33118 8678 33148 8730
rect 33148 8678 33160 8730
rect 33160 8678 33174 8730
rect 33198 8678 33212 8730
rect 33212 8678 33224 8730
rect 33224 8678 33254 8730
rect 33278 8678 33288 8730
rect 33288 8678 33334 8730
rect 33038 8676 33094 8678
rect 33118 8676 33174 8678
rect 33198 8676 33254 8678
rect 33278 8676 33334 8678
rect 27691 2746 27747 2748
rect 27771 2746 27827 2748
rect 27851 2746 27907 2748
rect 27931 2746 27987 2748
rect 27691 2694 27737 2746
rect 27737 2694 27747 2746
rect 27771 2694 27801 2746
rect 27801 2694 27813 2746
rect 27813 2694 27827 2746
rect 27851 2694 27865 2746
rect 27865 2694 27877 2746
rect 27877 2694 27907 2746
rect 27931 2694 27941 2746
rect 27941 2694 27987 2746
rect 27691 2692 27747 2694
rect 27771 2692 27827 2694
rect 27851 2692 27907 2694
rect 27931 2692 27987 2694
rect 27691 1658 27747 1660
rect 27771 1658 27827 1660
rect 27851 1658 27907 1660
rect 27931 1658 27987 1660
rect 27691 1606 27737 1658
rect 27737 1606 27747 1658
rect 27771 1606 27801 1658
rect 27801 1606 27813 1658
rect 27813 1606 27827 1658
rect 27851 1606 27865 1658
rect 27865 1606 27877 1658
rect 27877 1606 27907 1658
rect 27931 1606 27941 1658
rect 27941 1606 27987 1658
rect 27691 1604 27747 1606
rect 27771 1604 27827 1606
rect 27851 1604 27907 1606
rect 27931 1604 27987 1606
rect 33038 7642 33094 7644
rect 33118 7642 33174 7644
rect 33198 7642 33254 7644
rect 33278 7642 33334 7644
rect 33038 7590 33084 7642
rect 33084 7590 33094 7642
rect 33118 7590 33148 7642
rect 33148 7590 33160 7642
rect 33160 7590 33174 7642
rect 33198 7590 33212 7642
rect 33212 7590 33224 7642
rect 33224 7590 33254 7642
rect 33278 7590 33288 7642
rect 33288 7590 33334 7642
rect 33038 7588 33094 7590
rect 33118 7588 33174 7590
rect 33198 7588 33254 7590
rect 33278 7588 33334 7590
rect 33966 7384 34022 7440
rect 33038 6554 33094 6556
rect 33118 6554 33174 6556
rect 33198 6554 33254 6556
rect 33278 6554 33334 6556
rect 33038 6502 33084 6554
rect 33084 6502 33094 6554
rect 33118 6502 33148 6554
rect 33148 6502 33160 6554
rect 33160 6502 33174 6554
rect 33198 6502 33212 6554
rect 33212 6502 33224 6554
rect 33224 6502 33254 6554
rect 33278 6502 33288 6554
rect 33288 6502 33334 6554
rect 33038 6500 33094 6502
rect 33118 6500 33174 6502
rect 33198 6500 33254 6502
rect 33278 6500 33334 6502
rect 33038 5466 33094 5468
rect 33118 5466 33174 5468
rect 33198 5466 33254 5468
rect 33278 5466 33334 5468
rect 33038 5414 33084 5466
rect 33084 5414 33094 5466
rect 33118 5414 33148 5466
rect 33148 5414 33160 5466
rect 33160 5414 33174 5466
rect 33198 5414 33212 5466
rect 33212 5414 33224 5466
rect 33224 5414 33254 5466
rect 33278 5414 33288 5466
rect 33288 5414 33334 5466
rect 33038 5412 33094 5414
rect 33118 5412 33174 5414
rect 33198 5412 33254 5414
rect 33278 5412 33334 5414
rect 33038 4378 33094 4380
rect 33118 4378 33174 4380
rect 33198 4378 33254 4380
rect 33278 4378 33334 4380
rect 33038 4326 33084 4378
rect 33084 4326 33094 4378
rect 33118 4326 33148 4378
rect 33148 4326 33160 4378
rect 33160 4326 33174 4378
rect 33198 4326 33212 4378
rect 33212 4326 33224 4378
rect 33224 4326 33254 4378
rect 33278 4326 33288 4378
rect 33288 4326 33334 4378
rect 33038 4324 33094 4326
rect 33118 4324 33174 4326
rect 33198 4324 33254 4326
rect 33278 4324 33334 4326
rect 33038 3290 33094 3292
rect 33118 3290 33174 3292
rect 33198 3290 33254 3292
rect 33278 3290 33334 3292
rect 33038 3238 33084 3290
rect 33084 3238 33094 3290
rect 33118 3238 33148 3290
rect 33148 3238 33160 3290
rect 33160 3238 33174 3290
rect 33198 3238 33212 3290
rect 33212 3238 33224 3290
rect 33224 3238 33254 3290
rect 33278 3238 33288 3290
rect 33288 3238 33334 3290
rect 33038 3236 33094 3238
rect 33118 3236 33174 3238
rect 33198 3236 33254 3238
rect 33278 3236 33334 3238
rect 33038 2202 33094 2204
rect 33118 2202 33174 2204
rect 33198 2202 33254 2204
rect 33278 2202 33334 2204
rect 33038 2150 33084 2202
rect 33084 2150 33094 2202
rect 33118 2150 33148 2202
rect 33148 2150 33160 2202
rect 33160 2150 33174 2202
rect 33198 2150 33212 2202
rect 33212 2150 33224 2202
rect 33224 2150 33254 2202
rect 33278 2150 33288 2202
rect 33288 2150 33334 2202
rect 33038 2148 33094 2150
rect 33118 2148 33174 2150
rect 33198 2148 33254 2150
rect 33278 2148 33334 2150
rect 38385 8186 38441 8188
rect 38465 8186 38521 8188
rect 38545 8186 38601 8188
rect 38625 8186 38681 8188
rect 38385 8134 38431 8186
rect 38431 8134 38441 8186
rect 38465 8134 38495 8186
rect 38495 8134 38507 8186
rect 38507 8134 38521 8186
rect 38545 8134 38559 8186
rect 38559 8134 38571 8186
rect 38571 8134 38601 8186
rect 38625 8134 38635 8186
rect 38635 8134 38681 8186
rect 38385 8132 38441 8134
rect 38465 8132 38521 8134
rect 38545 8132 38601 8134
rect 38625 8132 38681 8134
rect 38385 7098 38441 7100
rect 38465 7098 38521 7100
rect 38545 7098 38601 7100
rect 38625 7098 38681 7100
rect 38385 7046 38431 7098
rect 38431 7046 38441 7098
rect 38465 7046 38495 7098
rect 38495 7046 38507 7098
rect 38507 7046 38521 7098
rect 38545 7046 38559 7098
rect 38559 7046 38571 7098
rect 38571 7046 38601 7098
rect 38625 7046 38635 7098
rect 38635 7046 38681 7098
rect 38385 7044 38441 7046
rect 38465 7044 38521 7046
rect 38545 7044 38601 7046
rect 38625 7044 38681 7046
rect 38385 6010 38441 6012
rect 38465 6010 38521 6012
rect 38545 6010 38601 6012
rect 38625 6010 38681 6012
rect 38385 5958 38431 6010
rect 38431 5958 38441 6010
rect 38465 5958 38495 6010
rect 38495 5958 38507 6010
rect 38507 5958 38521 6010
rect 38545 5958 38559 6010
rect 38559 5958 38571 6010
rect 38571 5958 38601 6010
rect 38625 5958 38635 6010
rect 38635 5958 38681 6010
rect 38385 5956 38441 5958
rect 38465 5956 38521 5958
rect 38545 5956 38601 5958
rect 38625 5956 38681 5958
rect 38385 4922 38441 4924
rect 38465 4922 38521 4924
rect 38545 4922 38601 4924
rect 38625 4922 38681 4924
rect 38385 4870 38431 4922
rect 38431 4870 38441 4922
rect 38465 4870 38495 4922
rect 38495 4870 38507 4922
rect 38507 4870 38521 4922
rect 38545 4870 38559 4922
rect 38559 4870 38571 4922
rect 38571 4870 38601 4922
rect 38625 4870 38635 4922
rect 38635 4870 38681 4922
rect 38385 4868 38441 4870
rect 38465 4868 38521 4870
rect 38545 4868 38601 4870
rect 38625 4868 38681 4870
rect 43732 8730 43788 8732
rect 43812 8730 43868 8732
rect 43892 8730 43948 8732
rect 43972 8730 44028 8732
rect 43732 8678 43778 8730
rect 43778 8678 43788 8730
rect 43812 8678 43842 8730
rect 43842 8678 43854 8730
rect 43854 8678 43868 8730
rect 43892 8678 43906 8730
rect 43906 8678 43918 8730
rect 43918 8678 43948 8730
rect 43972 8678 43982 8730
rect 43982 8678 44028 8730
rect 43732 8676 43788 8678
rect 43812 8676 43868 8678
rect 43892 8676 43948 8678
rect 43972 8676 44028 8678
rect 33038 1114 33094 1116
rect 33118 1114 33174 1116
rect 33198 1114 33254 1116
rect 33278 1114 33334 1116
rect 33038 1062 33084 1114
rect 33084 1062 33094 1114
rect 33118 1062 33148 1114
rect 33148 1062 33160 1114
rect 33160 1062 33174 1114
rect 33198 1062 33212 1114
rect 33212 1062 33224 1114
rect 33224 1062 33254 1114
rect 33278 1062 33288 1114
rect 33288 1062 33334 1114
rect 33038 1060 33094 1062
rect 33118 1060 33174 1062
rect 33198 1060 33254 1062
rect 33278 1060 33334 1062
rect 38385 3834 38441 3836
rect 38465 3834 38521 3836
rect 38545 3834 38601 3836
rect 38625 3834 38681 3836
rect 38385 3782 38431 3834
rect 38431 3782 38441 3834
rect 38465 3782 38495 3834
rect 38495 3782 38507 3834
rect 38507 3782 38521 3834
rect 38545 3782 38559 3834
rect 38559 3782 38571 3834
rect 38571 3782 38601 3834
rect 38625 3782 38635 3834
rect 38635 3782 38681 3834
rect 38385 3780 38441 3782
rect 38465 3780 38521 3782
rect 38545 3780 38601 3782
rect 38625 3780 38681 3782
rect 38385 2746 38441 2748
rect 38465 2746 38521 2748
rect 38545 2746 38601 2748
rect 38625 2746 38681 2748
rect 38385 2694 38431 2746
rect 38431 2694 38441 2746
rect 38465 2694 38495 2746
rect 38495 2694 38507 2746
rect 38507 2694 38521 2746
rect 38545 2694 38559 2746
rect 38559 2694 38571 2746
rect 38571 2694 38601 2746
rect 38625 2694 38635 2746
rect 38635 2694 38681 2746
rect 38385 2692 38441 2694
rect 38465 2692 38521 2694
rect 38545 2692 38601 2694
rect 38625 2692 38681 2694
rect 43732 7642 43788 7644
rect 43812 7642 43868 7644
rect 43892 7642 43948 7644
rect 43972 7642 44028 7644
rect 43732 7590 43778 7642
rect 43778 7590 43788 7642
rect 43812 7590 43842 7642
rect 43842 7590 43854 7642
rect 43854 7590 43868 7642
rect 43892 7590 43906 7642
rect 43906 7590 43918 7642
rect 43918 7590 43948 7642
rect 43972 7590 43982 7642
rect 43982 7590 44028 7642
rect 43732 7588 43788 7590
rect 43812 7588 43868 7590
rect 43892 7588 43948 7590
rect 43972 7588 44028 7590
rect 43732 6554 43788 6556
rect 43812 6554 43868 6556
rect 43892 6554 43948 6556
rect 43972 6554 44028 6556
rect 43732 6502 43778 6554
rect 43778 6502 43788 6554
rect 43812 6502 43842 6554
rect 43842 6502 43854 6554
rect 43854 6502 43868 6554
rect 43892 6502 43906 6554
rect 43906 6502 43918 6554
rect 43918 6502 43948 6554
rect 43972 6502 43982 6554
rect 43982 6502 44028 6554
rect 43732 6500 43788 6502
rect 43812 6500 43868 6502
rect 43892 6500 43948 6502
rect 43972 6500 44028 6502
rect 43732 5466 43788 5468
rect 43812 5466 43868 5468
rect 43892 5466 43948 5468
rect 43972 5466 44028 5468
rect 43732 5414 43778 5466
rect 43778 5414 43788 5466
rect 43812 5414 43842 5466
rect 43842 5414 43854 5466
rect 43854 5414 43868 5466
rect 43892 5414 43906 5466
rect 43906 5414 43918 5466
rect 43918 5414 43948 5466
rect 43972 5414 43982 5466
rect 43982 5414 44028 5466
rect 43732 5412 43788 5414
rect 43812 5412 43868 5414
rect 43892 5412 43948 5414
rect 43972 5412 44028 5414
rect 43732 4378 43788 4380
rect 43812 4378 43868 4380
rect 43892 4378 43948 4380
rect 43972 4378 44028 4380
rect 43732 4326 43778 4378
rect 43778 4326 43788 4378
rect 43812 4326 43842 4378
rect 43842 4326 43854 4378
rect 43854 4326 43868 4378
rect 43892 4326 43906 4378
rect 43906 4326 43918 4378
rect 43918 4326 43948 4378
rect 43972 4326 43982 4378
rect 43982 4326 44028 4378
rect 43732 4324 43788 4326
rect 43812 4324 43868 4326
rect 43892 4324 43948 4326
rect 43972 4324 44028 4326
rect 43732 3290 43788 3292
rect 43812 3290 43868 3292
rect 43892 3290 43948 3292
rect 43972 3290 44028 3292
rect 43732 3238 43778 3290
rect 43778 3238 43788 3290
rect 43812 3238 43842 3290
rect 43842 3238 43854 3290
rect 43854 3238 43868 3290
rect 43892 3238 43906 3290
rect 43906 3238 43918 3290
rect 43918 3238 43948 3290
rect 43972 3238 43982 3290
rect 43982 3238 44028 3290
rect 43732 3236 43788 3238
rect 43812 3236 43868 3238
rect 43892 3236 43948 3238
rect 43972 3236 44028 3238
rect 38385 1658 38441 1660
rect 38465 1658 38521 1660
rect 38545 1658 38601 1660
rect 38625 1658 38681 1660
rect 38385 1606 38431 1658
rect 38431 1606 38441 1658
rect 38465 1606 38495 1658
rect 38495 1606 38507 1658
rect 38507 1606 38521 1658
rect 38545 1606 38559 1658
rect 38559 1606 38571 1658
rect 38571 1606 38601 1658
rect 38625 1606 38635 1658
rect 38635 1606 38681 1658
rect 38385 1604 38441 1606
rect 38465 1604 38521 1606
rect 38545 1604 38601 1606
rect 38625 1604 38681 1606
rect 43732 2202 43788 2204
rect 43812 2202 43868 2204
rect 43892 2202 43948 2204
rect 43972 2202 44028 2204
rect 43732 2150 43778 2202
rect 43778 2150 43788 2202
rect 43812 2150 43842 2202
rect 43842 2150 43854 2202
rect 43854 2150 43868 2202
rect 43892 2150 43906 2202
rect 43906 2150 43918 2202
rect 43918 2150 43948 2202
rect 43972 2150 43982 2202
rect 43982 2150 44028 2202
rect 43732 2148 43788 2150
rect 43812 2148 43868 2150
rect 43892 2148 43948 2150
rect 43972 2148 44028 2150
rect 43732 1114 43788 1116
rect 43812 1114 43868 1116
rect 43892 1114 43948 1116
rect 43972 1114 44028 1116
rect 43732 1062 43778 1114
rect 43778 1062 43788 1114
rect 43812 1062 43842 1114
rect 43842 1062 43854 1114
rect 43854 1062 43868 1114
rect 43892 1062 43906 1114
rect 43906 1062 43918 1114
rect 43918 1062 43948 1114
rect 43972 1062 43982 1114
rect 43982 1062 44028 1114
rect 43732 1060 43788 1062
rect 43812 1060 43868 1062
rect 43892 1060 43948 1062
rect 43972 1060 44028 1062
<< metal3 >>
rect 20069 9892 20135 9893
rect 20069 9890 20116 9892
rect 20024 9888 20116 9890
rect 20024 9832 20074 9888
rect 20024 9830 20116 9832
rect 20069 9828 20116 9830
rect 20180 9828 20186 9892
rect 20069 9827 20135 9828
rect 17125 9482 17191 9485
rect 21541 9482 21607 9485
rect 17125 9480 21607 9482
rect 17125 9424 17130 9480
rect 17186 9424 21546 9480
rect 21602 9424 21607 9480
rect 17125 9422 21607 9424
rect 17125 9419 17191 9422
rect 21541 9419 21607 9422
rect 19057 9346 19123 9349
rect 20161 9346 20227 9349
rect 19057 9344 20227 9346
rect 19057 9288 19062 9344
rect 19118 9288 20166 9344
rect 20222 9288 20227 9344
rect 19057 9286 20227 9288
rect 19057 9283 19123 9286
rect 20161 9283 20227 9286
rect 12709 9210 12775 9213
rect 27245 9210 27311 9213
rect 12709 9208 27311 9210
rect 12709 9152 12714 9208
rect 12770 9152 27250 9208
rect 27306 9152 27311 9208
rect 12709 9150 27311 9152
rect 12709 9147 12775 9150
rect 27245 9147 27311 9150
rect 4889 9074 4955 9077
rect 19742 9074 19748 9076
rect 4889 9072 19748 9074
rect 4889 9016 4894 9072
rect 4950 9016 19748 9072
rect 4889 9014 19748 9016
rect 4889 9011 4955 9014
rect 19742 9012 19748 9014
rect 19812 9012 19818 9076
rect 21909 9074 21975 9077
rect 26877 9074 26943 9077
rect 21909 9072 26943 9074
rect 21909 9016 21914 9072
rect 21970 9016 26882 9072
rect 26938 9016 26943 9072
rect 21909 9014 26943 9016
rect 21909 9011 21975 9014
rect 26877 9011 26943 9014
rect 32213 8938 32279 8941
rect 18462 8936 32279 8938
rect 18462 8880 32218 8936
rect 32274 8880 32279 8936
rect 18462 8878 32279 8880
rect 11640 8736 11956 8737
rect 11640 8672 11646 8736
rect 11710 8672 11726 8736
rect 11790 8672 11806 8736
rect 11870 8672 11886 8736
rect 11950 8672 11956 8736
rect 11640 8671 11956 8672
rect 18229 8530 18295 8533
rect 18462 8530 18522 8878
rect 32213 8875 32279 8878
rect 18689 8802 18755 8805
rect 20437 8802 20503 8805
rect 18689 8800 20503 8802
rect 18689 8744 18694 8800
rect 18750 8744 20442 8800
rect 20498 8744 20503 8800
rect 18689 8742 20503 8744
rect 18689 8739 18755 8742
rect 20437 8739 20503 8742
rect 22334 8736 22650 8737
rect 22334 8672 22340 8736
rect 22404 8672 22420 8736
rect 22484 8672 22500 8736
rect 22564 8672 22580 8736
rect 22644 8672 22650 8736
rect 22334 8671 22650 8672
rect 33028 8736 33344 8737
rect 33028 8672 33034 8736
rect 33098 8672 33114 8736
rect 33178 8672 33194 8736
rect 33258 8672 33274 8736
rect 33338 8672 33344 8736
rect 33028 8671 33344 8672
rect 43722 8736 44038 8737
rect 43722 8672 43728 8736
rect 43792 8672 43808 8736
rect 43872 8672 43888 8736
rect 43952 8672 43968 8736
rect 44032 8672 44038 8736
rect 43722 8671 44038 8672
rect 31937 8530 32003 8533
rect 18229 8528 18522 8530
rect 18229 8472 18234 8528
rect 18290 8472 18522 8528
rect 18229 8470 18522 8472
rect 18646 8528 32003 8530
rect 18646 8472 31942 8528
rect 31998 8472 32003 8528
rect 18646 8470 32003 8472
rect 18229 8467 18295 8470
rect 18646 8261 18706 8470
rect 31937 8467 32003 8470
rect 18781 8394 18847 8397
rect 22185 8394 22251 8397
rect 18781 8392 22251 8394
rect 18781 8336 18786 8392
rect 18842 8336 22190 8392
rect 22246 8336 22251 8392
rect 18781 8334 22251 8336
rect 18781 8331 18847 8334
rect 22185 8331 22251 8334
rect 18597 8256 18706 8261
rect 18597 8200 18602 8256
rect 18658 8200 18706 8256
rect 18597 8198 18706 8200
rect 19701 8258 19767 8261
rect 19926 8258 19932 8260
rect 19701 8256 19932 8258
rect 19701 8200 19706 8256
rect 19762 8200 19932 8256
rect 19701 8198 19932 8200
rect 18597 8195 18663 8198
rect 19701 8195 19767 8198
rect 19926 8196 19932 8198
rect 19996 8196 20002 8260
rect 20713 8258 20779 8261
rect 24669 8258 24735 8261
rect 20713 8256 24735 8258
rect 20713 8200 20718 8256
rect 20774 8200 24674 8256
rect 24730 8200 24735 8256
rect 20713 8198 24735 8200
rect 20713 8195 20779 8198
rect 24669 8195 24735 8198
rect 6293 8192 6609 8193
rect 6293 8128 6299 8192
rect 6363 8128 6379 8192
rect 6443 8128 6459 8192
rect 6523 8128 6539 8192
rect 6603 8128 6609 8192
rect 6293 8127 6609 8128
rect 16987 8192 17303 8193
rect 16987 8128 16993 8192
rect 17057 8128 17073 8192
rect 17137 8128 17153 8192
rect 17217 8128 17233 8192
rect 17297 8128 17303 8192
rect 16987 8127 17303 8128
rect 27681 8192 27997 8193
rect 27681 8128 27687 8192
rect 27751 8128 27767 8192
rect 27831 8128 27847 8192
rect 27911 8128 27927 8192
rect 27991 8128 27997 8192
rect 27681 8127 27997 8128
rect 38375 8192 38691 8193
rect 38375 8128 38381 8192
rect 38445 8128 38461 8192
rect 38525 8128 38541 8192
rect 38605 8128 38621 8192
rect 38685 8128 38691 8192
rect 38375 8127 38691 8128
rect 19374 8060 19380 8124
rect 19444 8122 19450 8124
rect 25497 8122 25563 8125
rect 19444 8120 25563 8122
rect 19444 8064 25502 8120
rect 25558 8064 25563 8120
rect 19444 8062 25563 8064
rect 19444 8060 19450 8062
rect 25497 8059 25563 8062
rect 12985 7986 13051 7989
rect 27337 7986 27403 7989
rect 12985 7984 27403 7986
rect 12985 7928 12990 7984
rect 13046 7928 27342 7984
rect 27398 7928 27403 7984
rect 12985 7926 27403 7928
rect 12985 7923 13051 7926
rect 27337 7923 27403 7926
rect 6729 7850 6795 7853
rect 17953 7850 18019 7853
rect 24025 7850 24091 7853
rect 6729 7848 12450 7850
rect 6729 7792 6734 7848
rect 6790 7792 12450 7848
rect 6729 7790 12450 7792
rect 6729 7787 6795 7790
rect 11640 7648 11956 7649
rect 11640 7584 11646 7648
rect 11710 7584 11726 7648
rect 11790 7584 11806 7648
rect 11870 7584 11886 7648
rect 11950 7584 11956 7648
rect 11640 7583 11956 7584
rect 12390 7578 12450 7790
rect 17953 7848 24091 7850
rect 17953 7792 17958 7848
rect 18014 7792 24030 7848
rect 24086 7792 24091 7848
rect 17953 7790 24091 7792
rect 17953 7787 18019 7790
rect 24025 7787 24091 7790
rect 15101 7714 15167 7717
rect 19374 7714 19380 7716
rect 15101 7712 19380 7714
rect 15101 7656 15106 7712
rect 15162 7656 19380 7712
rect 15101 7654 19380 7656
rect 15101 7651 15167 7654
rect 19374 7652 19380 7654
rect 19444 7652 19450 7716
rect 20069 7714 20135 7717
rect 20069 7712 20362 7714
rect 20069 7656 20074 7712
rect 20130 7656 20362 7712
rect 20069 7654 20362 7656
rect 20069 7651 20135 7654
rect 20161 7578 20227 7581
rect 12390 7576 20227 7578
rect 12390 7520 20166 7576
rect 20222 7520 20227 7576
rect 12390 7518 20227 7520
rect 20161 7515 20227 7518
rect 9581 7442 9647 7445
rect 20302 7442 20362 7654
rect 22334 7648 22650 7649
rect 22334 7584 22340 7648
rect 22404 7584 22420 7648
rect 22484 7584 22500 7648
rect 22564 7584 22580 7648
rect 22644 7584 22650 7648
rect 22334 7583 22650 7584
rect 33028 7648 33344 7649
rect 33028 7584 33034 7648
rect 33098 7584 33114 7648
rect 33178 7584 33194 7648
rect 33258 7584 33274 7648
rect 33338 7584 33344 7648
rect 33028 7583 33344 7584
rect 43722 7648 44038 7649
rect 43722 7584 43728 7648
rect 43792 7584 43808 7648
rect 43872 7584 43888 7648
rect 43952 7584 43968 7648
rect 44032 7584 44038 7648
rect 43722 7583 44038 7584
rect 9581 7440 20362 7442
rect 9581 7384 9586 7440
rect 9642 7384 20362 7440
rect 9581 7382 20362 7384
rect 22001 7442 22067 7445
rect 33961 7442 34027 7445
rect 22001 7440 34027 7442
rect 22001 7384 22006 7440
rect 22062 7384 33966 7440
rect 34022 7384 34027 7440
rect 22001 7382 34027 7384
rect 9581 7379 9647 7382
rect 22001 7379 22067 7382
rect 33961 7379 34027 7382
rect 6545 7306 6611 7309
rect 19609 7306 19675 7309
rect 6545 7304 19675 7306
rect 6545 7248 6550 7304
rect 6606 7248 19614 7304
rect 19670 7248 19675 7304
rect 6545 7246 19675 7248
rect 6545 7243 6611 7246
rect 19609 7243 19675 7246
rect 19742 7244 19748 7308
rect 19812 7244 19818 7308
rect 20161 7306 20227 7309
rect 24853 7306 24919 7309
rect 20161 7304 24919 7306
rect 20161 7248 20166 7304
rect 20222 7248 24858 7304
rect 24914 7248 24919 7304
rect 20161 7246 24919 7248
rect 19750 7170 19810 7244
rect 20161 7243 20227 7246
rect 24853 7243 24919 7246
rect 20161 7170 20227 7173
rect 19750 7168 20227 7170
rect 19750 7112 20166 7168
rect 20222 7112 20227 7168
rect 19750 7110 20227 7112
rect 20161 7107 20227 7110
rect 6293 7104 6609 7105
rect 6293 7040 6299 7104
rect 6363 7040 6379 7104
rect 6443 7040 6459 7104
rect 6523 7040 6539 7104
rect 6603 7040 6609 7104
rect 6293 7039 6609 7040
rect 16987 7104 17303 7105
rect 16987 7040 16993 7104
rect 17057 7040 17073 7104
rect 17137 7040 17153 7104
rect 17217 7040 17233 7104
rect 17297 7040 17303 7104
rect 16987 7039 17303 7040
rect 27681 7104 27997 7105
rect 27681 7040 27687 7104
rect 27751 7040 27767 7104
rect 27831 7040 27847 7104
rect 27911 7040 27927 7104
rect 27991 7040 27997 7104
rect 27681 7039 27997 7040
rect 38375 7104 38691 7105
rect 38375 7040 38381 7104
rect 38445 7040 38461 7104
rect 38525 7040 38541 7104
rect 38605 7040 38621 7104
rect 38685 7040 38691 7104
rect 38375 7039 38691 7040
rect 19977 7036 20043 7037
rect 19926 7034 19932 7036
rect 19886 6974 19932 7034
rect 19996 7032 20043 7036
rect 20038 6976 20043 7032
rect 19926 6972 19932 6974
rect 19996 6972 20043 6976
rect 20110 6972 20116 7036
rect 20180 7034 20186 7036
rect 20253 7034 20319 7037
rect 20180 7032 20319 7034
rect 20180 6976 20258 7032
rect 20314 6976 20319 7032
rect 20180 6974 20319 6976
rect 20180 6972 20186 6974
rect 19977 6971 20043 6972
rect 20253 6971 20319 6974
rect 15561 6898 15627 6901
rect 22829 6898 22895 6901
rect 15561 6896 22895 6898
rect 15561 6840 15566 6896
rect 15622 6840 22834 6896
rect 22890 6840 22895 6896
rect 15561 6838 22895 6840
rect 15561 6835 15627 6838
rect 22829 6835 22895 6838
rect 7465 6762 7531 6765
rect 21357 6762 21423 6765
rect 7465 6760 21423 6762
rect 7465 6704 7470 6760
rect 7526 6704 21362 6760
rect 21418 6704 21423 6760
rect 7465 6702 21423 6704
rect 7465 6699 7531 6702
rect 21357 6699 21423 6702
rect 14825 6626 14891 6629
rect 21449 6626 21515 6629
rect 14825 6624 21515 6626
rect 14825 6568 14830 6624
rect 14886 6568 21454 6624
rect 21510 6568 21515 6624
rect 14825 6566 21515 6568
rect 14825 6563 14891 6566
rect 21449 6563 21515 6566
rect 11640 6560 11956 6561
rect 11640 6496 11646 6560
rect 11710 6496 11726 6560
rect 11790 6496 11806 6560
rect 11870 6496 11886 6560
rect 11950 6496 11956 6560
rect 11640 6495 11956 6496
rect 22334 6560 22650 6561
rect 22334 6496 22340 6560
rect 22404 6496 22420 6560
rect 22484 6496 22500 6560
rect 22564 6496 22580 6560
rect 22644 6496 22650 6560
rect 22334 6495 22650 6496
rect 33028 6560 33344 6561
rect 33028 6496 33034 6560
rect 33098 6496 33114 6560
rect 33178 6496 33194 6560
rect 33258 6496 33274 6560
rect 33338 6496 33344 6560
rect 33028 6495 33344 6496
rect 43722 6560 44038 6561
rect 43722 6496 43728 6560
rect 43792 6496 43808 6560
rect 43872 6496 43888 6560
rect 43952 6496 43968 6560
rect 44032 6496 44038 6560
rect 43722 6495 44038 6496
rect 7005 6354 7071 6357
rect 23749 6354 23815 6357
rect 7005 6352 23815 6354
rect 7005 6296 7010 6352
rect 7066 6296 23754 6352
rect 23810 6296 23815 6352
rect 7005 6294 23815 6296
rect 7005 6291 7071 6294
rect 23749 6291 23815 6294
rect 8017 6218 8083 6221
rect 22093 6218 22159 6221
rect 8017 6216 22159 6218
rect 8017 6160 8022 6216
rect 8078 6160 22098 6216
rect 22154 6160 22159 6216
rect 8017 6158 22159 6160
rect 8017 6155 8083 6158
rect 22093 6155 22159 6158
rect 6293 6016 6609 6017
rect 6293 5952 6299 6016
rect 6363 5952 6379 6016
rect 6443 5952 6459 6016
rect 6523 5952 6539 6016
rect 6603 5952 6609 6016
rect 6293 5951 6609 5952
rect 16987 6016 17303 6017
rect 16987 5952 16993 6016
rect 17057 5952 17073 6016
rect 17137 5952 17153 6016
rect 17217 5952 17233 6016
rect 17297 5952 17303 6016
rect 16987 5951 17303 5952
rect 27681 6016 27997 6017
rect 27681 5952 27687 6016
rect 27751 5952 27767 6016
rect 27831 5952 27847 6016
rect 27911 5952 27927 6016
rect 27991 5952 27997 6016
rect 27681 5951 27997 5952
rect 38375 6016 38691 6017
rect 38375 5952 38381 6016
rect 38445 5952 38461 6016
rect 38525 5952 38541 6016
rect 38605 5952 38621 6016
rect 38685 5952 38691 6016
rect 38375 5951 38691 5952
rect 8201 5810 8267 5813
rect 23473 5810 23539 5813
rect 8201 5808 23539 5810
rect 8201 5752 8206 5808
rect 8262 5752 23478 5808
rect 23534 5752 23539 5808
rect 8201 5750 23539 5752
rect 8201 5747 8267 5750
rect 23473 5747 23539 5750
rect 11640 5472 11956 5473
rect 11640 5408 11646 5472
rect 11710 5408 11726 5472
rect 11790 5408 11806 5472
rect 11870 5408 11886 5472
rect 11950 5408 11956 5472
rect 11640 5407 11956 5408
rect 22334 5472 22650 5473
rect 22334 5408 22340 5472
rect 22404 5408 22420 5472
rect 22484 5408 22500 5472
rect 22564 5408 22580 5472
rect 22644 5408 22650 5472
rect 22334 5407 22650 5408
rect 33028 5472 33344 5473
rect 33028 5408 33034 5472
rect 33098 5408 33114 5472
rect 33178 5408 33194 5472
rect 33258 5408 33274 5472
rect 33338 5408 33344 5472
rect 33028 5407 33344 5408
rect 43722 5472 44038 5473
rect 43722 5408 43728 5472
rect 43792 5408 43808 5472
rect 43872 5408 43888 5472
rect 43952 5408 43968 5472
rect 44032 5408 44038 5472
rect 43722 5407 44038 5408
rect 6293 4928 6609 4929
rect 6293 4864 6299 4928
rect 6363 4864 6379 4928
rect 6443 4864 6459 4928
rect 6523 4864 6539 4928
rect 6603 4864 6609 4928
rect 6293 4863 6609 4864
rect 16987 4928 17303 4929
rect 16987 4864 16993 4928
rect 17057 4864 17073 4928
rect 17137 4864 17153 4928
rect 17217 4864 17233 4928
rect 17297 4864 17303 4928
rect 16987 4863 17303 4864
rect 27681 4928 27997 4929
rect 27681 4864 27687 4928
rect 27751 4864 27767 4928
rect 27831 4864 27847 4928
rect 27911 4864 27927 4928
rect 27991 4864 27997 4928
rect 27681 4863 27997 4864
rect 38375 4928 38691 4929
rect 38375 4864 38381 4928
rect 38445 4864 38461 4928
rect 38525 4864 38541 4928
rect 38605 4864 38621 4928
rect 38685 4864 38691 4928
rect 38375 4863 38691 4864
rect 11640 4384 11956 4385
rect 11640 4320 11646 4384
rect 11710 4320 11726 4384
rect 11790 4320 11806 4384
rect 11870 4320 11886 4384
rect 11950 4320 11956 4384
rect 11640 4319 11956 4320
rect 22334 4384 22650 4385
rect 22334 4320 22340 4384
rect 22404 4320 22420 4384
rect 22484 4320 22500 4384
rect 22564 4320 22580 4384
rect 22644 4320 22650 4384
rect 22334 4319 22650 4320
rect 33028 4384 33344 4385
rect 33028 4320 33034 4384
rect 33098 4320 33114 4384
rect 33178 4320 33194 4384
rect 33258 4320 33274 4384
rect 33338 4320 33344 4384
rect 33028 4319 33344 4320
rect 43722 4384 44038 4385
rect 43722 4320 43728 4384
rect 43792 4320 43808 4384
rect 43872 4320 43888 4384
rect 43952 4320 43968 4384
rect 44032 4320 44038 4384
rect 43722 4319 44038 4320
rect 6293 3840 6609 3841
rect 6293 3776 6299 3840
rect 6363 3776 6379 3840
rect 6443 3776 6459 3840
rect 6523 3776 6539 3840
rect 6603 3776 6609 3840
rect 6293 3775 6609 3776
rect 16987 3840 17303 3841
rect 16987 3776 16993 3840
rect 17057 3776 17073 3840
rect 17137 3776 17153 3840
rect 17217 3776 17233 3840
rect 17297 3776 17303 3840
rect 16987 3775 17303 3776
rect 27681 3840 27997 3841
rect 27681 3776 27687 3840
rect 27751 3776 27767 3840
rect 27831 3776 27847 3840
rect 27911 3776 27927 3840
rect 27991 3776 27997 3840
rect 27681 3775 27997 3776
rect 38375 3840 38691 3841
rect 38375 3776 38381 3840
rect 38445 3776 38461 3840
rect 38525 3776 38541 3840
rect 38605 3776 38621 3840
rect 38685 3776 38691 3840
rect 38375 3775 38691 3776
rect 11640 3296 11956 3297
rect 11640 3232 11646 3296
rect 11710 3232 11726 3296
rect 11790 3232 11806 3296
rect 11870 3232 11886 3296
rect 11950 3232 11956 3296
rect 11640 3231 11956 3232
rect 22334 3296 22650 3297
rect 22334 3232 22340 3296
rect 22404 3232 22420 3296
rect 22484 3232 22500 3296
rect 22564 3232 22580 3296
rect 22644 3232 22650 3296
rect 22334 3231 22650 3232
rect 33028 3296 33344 3297
rect 33028 3232 33034 3296
rect 33098 3232 33114 3296
rect 33178 3232 33194 3296
rect 33258 3232 33274 3296
rect 33338 3232 33344 3296
rect 33028 3231 33344 3232
rect 43722 3296 44038 3297
rect 43722 3232 43728 3296
rect 43792 3232 43808 3296
rect 43872 3232 43888 3296
rect 43952 3232 43968 3296
rect 44032 3232 44038 3296
rect 43722 3231 44038 3232
rect 6293 2752 6609 2753
rect 6293 2688 6299 2752
rect 6363 2688 6379 2752
rect 6443 2688 6459 2752
rect 6523 2688 6539 2752
rect 6603 2688 6609 2752
rect 6293 2687 6609 2688
rect 16987 2752 17303 2753
rect 16987 2688 16993 2752
rect 17057 2688 17073 2752
rect 17137 2688 17153 2752
rect 17217 2688 17233 2752
rect 17297 2688 17303 2752
rect 16987 2687 17303 2688
rect 27681 2752 27997 2753
rect 27681 2688 27687 2752
rect 27751 2688 27767 2752
rect 27831 2688 27847 2752
rect 27911 2688 27927 2752
rect 27991 2688 27997 2752
rect 27681 2687 27997 2688
rect 38375 2752 38691 2753
rect 38375 2688 38381 2752
rect 38445 2688 38461 2752
rect 38525 2688 38541 2752
rect 38605 2688 38621 2752
rect 38685 2688 38691 2752
rect 38375 2687 38691 2688
rect 11640 2208 11956 2209
rect 11640 2144 11646 2208
rect 11710 2144 11726 2208
rect 11790 2144 11806 2208
rect 11870 2144 11886 2208
rect 11950 2144 11956 2208
rect 11640 2143 11956 2144
rect 22334 2208 22650 2209
rect 22334 2144 22340 2208
rect 22404 2144 22420 2208
rect 22484 2144 22500 2208
rect 22564 2144 22580 2208
rect 22644 2144 22650 2208
rect 22334 2143 22650 2144
rect 33028 2208 33344 2209
rect 33028 2144 33034 2208
rect 33098 2144 33114 2208
rect 33178 2144 33194 2208
rect 33258 2144 33274 2208
rect 33338 2144 33344 2208
rect 33028 2143 33344 2144
rect 43722 2208 44038 2209
rect 43722 2144 43728 2208
rect 43792 2144 43808 2208
rect 43872 2144 43888 2208
rect 43952 2144 43968 2208
rect 44032 2144 44038 2208
rect 43722 2143 44038 2144
rect 6293 1664 6609 1665
rect 6293 1600 6299 1664
rect 6363 1600 6379 1664
rect 6443 1600 6459 1664
rect 6523 1600 6539 1664
rect 6603 1600 6609 1664
rect 6293 1599 6609 1600
rect 16987 1664 17303 1665
rect 16987 1600 16993 1664
rect 17057 1600 17073 1664
rect 17137 1600 17153 1664
rect 17217 1600 17233 1664
rect 17297 1600 17303 1664
rect 16987 1599 17303 1600
rect 27681 1664 27997 1665
rect 27681 1600 27687 1664
rect 27751 1600 27767 1664
rect 27831 1600 27847 1664
rect 27911 1600 27927 1664
rect 27991 1600 27997 1664
rect 27681 1599 27997 1600
rect 38375 1664 38691 1665
rect 38375 1600 38381 1664
rect 38445 1600 38461 1664
rect 38525 1600 38541 1664
rect 38605 1600 38621 1664
rect 38685 1600 38691 1664
rect 38375 1599 38691 1600
rect 11640 1120 11956 1121
rect 11640 1056 11646 1120
rect 11710 1056 11726 1120
rect 11790 1056 11806 1120
rect 11870 1056 11886 1120
rect 11950 1056 11956 1120
rect 11640 1055 11956 1056
rect 22334 1120 22650 1121
rect 22334 1056 22340 1120
rect 22404 1056 22420 1120
rect 22484 1056 22500 1120
rect 22564 1056 22580 1120
rect 22644 1056 22650 1120
rect 22334 1055 22650 1056
rect 33028 1120 33344 1121
rect 33028 1056 33034 1120
rect 33098 1056 33114 1120
rect 33178 1056 33194 1120
rect 33258 1056 33274 1120
rect 33338 1056 33344 1120
rect 33028 1055 33344 1056
rect 43722 1120 44038 1121
rect 43722 1056 43728 1120
rect 43792 1056 43808 1120
rect 43872 1056 43888 1120
rect 43952 1056 43968 1120
rect 44032 1056 44038 1120
rect 43722 1055 44038 1056
<< via3 >>
rect 20116 9888 20180 9892
rect 20116 9832 20130 9888
rect 20130 9832 20180 9888
rect 20116 9828 20180 9832
rect 19748 9012 19812 9076
rect 11646 8732 11710 8736
rect 11646 8676 11650 8732
rect 11650 8676 11706 8732
rect 11706 8676 11710 8732
rect 11646 8672 11710 8676
rect 11726 8732 11790 8736
rect 11726 8676 11730 8732
rect 11730 8676 11786 8732
rect 11786 8676 11790 8732
rect 11726 8672 11790 8676
rect 11806 8732 11870 8736
rect 11806 8676 11810 8732
rect 11810 8676 11866 8732
rect 11866 8676 11870 8732
rect 11806 8672 11870 8676
rect 11886 8732 11950 8736
rect 11886 8676 11890 8732
rect 11890 8676 11946 8732
rect 11946 8676 11950 8732
rect 11886 8672 11950 8676
rect 22340 8732 22404 8736
rect 22340 8676 22344 8732
rect 22344 8676 22400 8732
rect 22400 8676 22404 8732
rect 22340 8672 22404 8676
rect 22420 8732 22484 8736
rect 22420 8676 22424 8732
rect 22424 8676 22480 8732
rect 22480 8676 22484 8732
rect 22420 8672 22484 8676
rect 22500 8732 22564 8736
rect 22500 8676 22504 8732
rect 22504 8676 22560 8732
rect 22560 8676 22564 8732
rect 22500 8672 22564 8676
rect 22580 8732 22644 8736
rect 22580 8676 22584 8732
rect 22584 8676 22640 8732
rect 22640 8676 22644 8732
rect 22580 8672 22644 8676
rect 33034 8732 33098 8736
rect 33034 8676 33038 8732
rect 33038 8676 33094 8732
rect 33094 8676 33098 8732
rect 33034 8672 33098 8676
rect 33114 8732 33178 8736
rect 33114 8676 33118 8732
rect 33118 8676 33174 8732
rect 33174 8676 33178 8732
rect 33114 8672 33178 8676
rect 33194 8732 33258 8736
rect 33194 8676 33198 8732
rect 33198 8676 33254 8732
rect 33254 8676 33258 8732
rect 33194 8672 33258 8676
rect 33274 8732 33338 8736
rect 33274 8676 33278 8732
rect 33278 8676 33334 8732
rect 33334 8676 33338 8732
rect 33274 8672 33338 8676
rect 43728 8732 43792 8736
rect 43728 8676 43732 8732
rect 43732 8676 43788 8732
rect 43788 8676 43792 8732
rect 43728 8672 43792 8676
rect 43808 8732 43872 8736
rect 43808 8676 43812 8732
rect 43812 8676 43868 8732
rect 43868 8676 43872 8732
rect 43808 8672 43872 8676
rect 43888 8732 43952 8736
rect 43888 8676 43892 8732
rect 43892 8676 43948 8732
rect 43948 8676 43952 8732
rect 43888 8672 43952 8676
rect 43968 8732 44032 8736
rect 43968 8676 43972 8732
rect 43972 8676 44028 8732
rect 44028 8676 44032 8732
rect 43968 8672 44032 8676
rect 19932 8196 19996 8260
rect 6299 8188 6363 8192
rect 6299 8132 6303 8188
rect 6303 8132 6359 8188
rect 6359 8132 6363 8188
rect 6299 8128 6363 8132
rect 6379 8188 6443 8192
rect 6379 8132 6383 8188
rect 6383 8132 6439 8188
rect 6439 8132 6443 8188
rect 6379 8128 6443 8132
rect 6459 8188 6523 8192
rect 6459 8132 6463 8188
rect 6463 8132 6519 8188
rect 6519 8132 6523 8188
rect 6459 8128 6523 8132
rect 6539 8188 6603 8192
rect 6539 8132 6543 8188
rect 6543 8132 6599 8188
rect 6599 8132 6603 8188
rect 6539 8128 6603 8132
rect 16993 8188 17057 8192
rect 16993 8132 16997 8188
rect 16997 8132 17053 8188
rect 17053 8132 17057 8188
rect 16993 8128 17057 8132
rect 17073 8188 17137 8192
rect 17073 8132 17077 8188
rect 17077 8132 17133 8188
rect 17133 8132 17137 8188
rect 17073 8128 17137 8132
rect 17153 8188 17217 8192
rect 17153 8132 17157 8188
rect 17157 8132 17213 8188
rect 17213 8132 17217 8188
rect 17153 8128 17217 8132
rect 17233 8188 17297 8192
rect 17233 8132 17237 8188
rect 17237 8132 17293 8188
rect 17293 8132 17297 8188
rect 17233 8128 17297 8132
rect 27687 8188 27751 8192
rect 27687 8132 27691 8188
rect 27691 8132 27747 8188
rect 27747 8132 27751 8188
rect 27687 8128 27751 8132
rect 27767 8188 27831 8192
rect 27767 8132 27771 8188
rect 27771 8132 27827 8188
rect 27827 8132 27831 8188
rect 27767 8128 27831 8132
rect 27847 8188 27911 8192
rect 27847 8132 27851 8188
rect 27851 8132 27907 8188
rect 27907 8132 27911 8188
rect 27847 8128 27911 8132
rect 27927 8188 27991 8192
rect 27927 8132 27931 8188
rect 27931 8132 27987 8188
rect 27987 8132 27991 8188
rect 27927 8128 27991 8132
rect 38381 8188 38445 8192
rect 38381 8132 38385 8188
rect 38385 8132 38441 8188
rect 38441 8132 38445 8188
rect 38381 8128 38445 8132
rect 38461 8188 38525 8192
rect 38461 8132 38465 8188
rect 38465 8132 38521 8188
rect 38521 8132 38525 8188
rect 38461 8128 38525 8132
rect 38541 8188 38605 8192
rect 38541 8132 38545 8188
rect 38545 8132 38601 8188
rect 38601 8132 38605 8188
rect 38541 8128 38605 8132
rect 38621 8188 38685 8192
rect 38621 8132 38625 8188
rect 38625 8132 38681 8188
rect 38681 8132 38685 8188
rect 38621 8128 38685 8132
rect 19380 8060 19444 8124
rect 11646 7644 11710 7648
rect 11646 7588 11650 7644
rect 11650 7588 11706 7644
rect 11706 7588 11710 7644
rect 11646 7584 11710 7588
rect 11726 7644 11790 7648
rect 11726 7588 11730 7644
rect 11730 7588 11786 7644
rect 11786 7588 11790 7644
rect 11726 7584 11790 7588
rect 11806 7644 11870 7648
rect 11806 7588 11810 7644
rect 11810 7588 11866 7644
rect 11866 7588 11870 7644
rect 11806 7584 11870 7588
rect 11886 7644 11950 7648
rect 11886 7588 11890 7644
rect 11890 7588 11946 7644
rect 11946 7588 11950 7644
rect 11886 7584 11950 7588
rect 19380 7652 19444 7716
rect 22340 7644 22404 7648
rect 22340 7588 22344 7644
rect 22344 7588 22400 7644
rect 22400 7588 22404 7644
rect 22340 7584 22404 7588
rect 22420 7644 22484 7648
rect 22420 7588 22424 7644
rect 22424 7588 22480 7644
rect 22480 7588 22484 7644
rect 22420 7584 22484 7588
rect 22500 7644 22564 7648
rect 22500 7588 22504 7644
rect 22504 7588 22560 7644
rect 22560 7588 22564 7644
rect 22500 7584 22564 7588
rect 22580 7644 22644 7648
rect 22580 7588 22584 7644
rect 22584 7588 22640 7644
rect 22640 7588 22644 7644
rect 22580 7584 22644 7588
rect 33034 7644 33098 7648
rect 33034 7588 33038 7644
rect 33038 7588 33094 7644
rect 33094 7588 33098 7644
rect 33034 7584 33098 7588
rect 33114 7644 33178 7648
rect 33114 7588 33118 7644
rect 33118 7588 33174 7644
rect 33174 7588 33178 7644
rect 33114 7584 33178 7588
rect 33194 7644 33258 7648
rect 33194 7588 33198 7644
rect 33198 7588 33254 7644
rect 33254 7588 33258 7644
rect 33194 7584 33258 7588
rect 33274 7644 33338 7648
rect 33274 7588 33278 7644
rect 33278 7588 33334 7644
rect 33334 7588 33338 7644
rect 33274 7584 33338 7588
rect 43728 7644 43792 7648
rect 43728 7588 43732 7644
rect 43732 7588 43788 7644
rect 43788 7588 43792 7644
rect 43728 7584 43792 7588
rect 43808 7644 43872 7648
rect 43808 7588 43812 7644
rect 43812 7588 43868 7644
rect 43868 7588 43872 7644
rect 43808 7584 43872 7588
rect 43888 7644 43952 7648
rect 43888 7588 43892 7644
rect 43892 7588 43948 7644
rect 43948 7588 43952 7644
rect 43888 7584 43952 7588
rect 43968 7644 44032 7648
rect 43968 7588 43972 7644
rect 43972 7588 44028 7644
rect 44028 7588 44032 7644
rect 43968 7584 44032 7588
rect 19748 7244 19812 7308
rect 6299 7100 6363 7104
rect 6299 7044 6303 7100
rect 6303 7044 6359 7100
rect 6359 7044 6363 7100
rect 6299 7040 6363 7044
rect 6379 7100 6443 7104
rect 6379 7044 6383 7100
rect 6383 7044 6439 7100
rect 6439 7044 6443 7100
rect 6379 7040 6443 7044
rect 6459 7100 6523 7104
rect 6459 7044 6463 7100
rect 6463 7044 6519 7100
rect 6519 7044 6523 7100
rect 6459 7040 6523 7044
rect 6539 7100 6603 7104
rect 6539 7044 6543 7100
rect 6543 7044 6599 7100
rect 6599 7044 6603 7100
rect 6539 7040 6603 7044
rect 16993 7100 17057 7104
rect 16993 7044 16997 7100
rect 16997 7044 17053 7100
rect 17053 7044 17057 7100
rect 16993 7040 17057 7044
rect 17073 7100 17137 7104
rect 17073 7044 17077 7100
rect 17077 7044 17133 7100
rect 17133 7044 17137 7100
rect 17073 7040 17137 7044
rect 17153 7100 17217 7104
rect 17153 7044 17157 7100
rect 17157 7044 17213 7100
rect 17213 7044 17217 7100
rect 17153 7040 17217 7044
rect 17233 7100 17297 7104
rect 17233 7044 17237 7100
rect 17237 7044 17293 7100
rect 17293 7044 17297 7100
rect 17233 7040 17297 7044
rect 27687 7100 27751 7104
rect 27687 7044 27691 7100
rect 27691 7044 27747 7100
rect 27747 7044 27751 7100
rect 27687 7040 27751 7044
rect 27767 7100 27831 7104
rect 27767 7044 27771 7100
rect 27771 7044 27827 7100
rect 27827 7044 27831 7100
rect 27767 7040 27831 7044
rect 27847 7100 27911 7104
rect 27847 7044 27851 7100
rect 27851 7044 27907 7100
rect 27907 7044 27911 7100
rect 27847 7040 27911 7044
rect 27927 7100 27991 7104
rect 27927 7044 27931 7100
rect 27931 7044 27987 7100
rect 27987 7044 27991 7100
rect 27927 7040 27991 7044
rect 38381 7100 38445 7104
rect 38381 7044 38385 7100
rect 38385 7044 38441 7100
rect 38441 7044 38445 7100
rect 38381 7040 38445 7044
rect 38461 7100 38525 7104
rect 38461 7044 38465 7100
rect 38465 7044 38521 7100
rect 38521 7044 38525 7100
rect 38461 7040 38525 7044
rect 38541 7100 38605 7104
rect 38541 7044 38545 7100
rect 38545 7044 38601 7100
rect 38601 7044 38605 7100
rect 38541 7040 38605 7044
rect 38621 7100 38685 7104
rect 38621 7044 38625 7100
rect 38625 7044 38681 7100
rect 38681 7044 38685 7100
rect 38621 7040 38685 7044
rect 19932 7032 19996 7036
rect 19932 6976 19982 7032
rect 19982 6976 19996 7032
rect 19932 6972 19996 6976
rect 20116 6972 20180 7036
rect 11646 6556 11710 6560
rect 11646 6500 11650 6556
rect 11650 6500 11706 6556
rect 11706 6500 11710 6556
rect 11646 6496 11710 6500
rect 11726 6556 11790 6560
rect 11726 6500 11730 6556
rect 11730 6500 11786 6556
rect 11786 6500 11790 6556
rect 11726 6496 11790 6500
rect 11806 6556 11870 6560
rect 11806 6500 11810 6556
rect 11810 6500 11866 6556
rect 11866 6500 11870 6556
rect 11806 6496 11870 6500
rect 11886 6556 11950 6560
rect 11886 6500 11890 6556
rect 11890 6500 11946 6556
rect 11946 6500 11950 6556
rect 11886 6496 11950 6500
rect 22340 6556 22404 6560
rect 22340 6500 22344 6556
rect 22344 6500 22400 6556
rect 22400 6500 22404 6556
rect 22340 6496 22404 6500
rect 22420 6556 22484 6560
rect 22420 6500 22424 6556
rect 22424 6500 22480 6556
rect 22480 6500 22484 6556
rect 22420 6496 22484 6500
rect 22500 6556 22564 6560
rect 22500 6500 22504 6556
rect 22504 6500 22560 6556
rect 22560 6500 22564 6556
rect 22500 6496 22564 6500
rect 22580 6556 22644 6560
rect 22580 6500 22584 6556
rect 22584 6500 22640 6556
rect 22640 6500 22644 6556
rect 22580 6496 22644 6500
rect 33034 6556 33098 6560
rect 33034 6500 33038 6556
rect 33038 6500 33094 6556
rect 33094 6500 33098 6556
rect 33034 6496 33098 6500
rect 33114 6556 33178 6560
rect 33114 6500 33118 6556
rect 33118 6500 33174 6556
rect 33174 6500 33178 6556
rect 33114 6496 33178 6500
rect 33194 6556 33258 6560
rect 33194 6500 33198 6556
rect 33198 6500 33254 6556
rect 33254 6500 33258 6556
rect 33194 6496 33258 6500
rect 33274 6556 33338 6560
rect 33274 6500 33278 6556
rect 33278 6500 33334 6556
rect 33334 6500 33338 6556
rect 33274 6496 33338 6500
rect 43728 6556 43792 6560
rect 43728 6500 43732 6556
rect 43732 6500 43788 6556
rect 43788 6500 43792 6556
rect 43728 6496 43792 6500
rect 43808 6556 43872 6560
rect 43808 6500 43812 6556
rect 43812 6500 43868 6556
rect 43868 6500 43872 6556
rect 43808 6496 43872 6500
rect 43888 6556 43952 6560
rect 43888 6500 43892 6556
rect 43892 6500 43948 6556
rect 43948 6500 43952 6556
rect 43888 6496 43952 6500
rect 43968 6556 44032 6560
rect 43968 6500 43972 6556
rect 43972 6500 44028 6556
rect 44028 6500 44032 6556
rect 43968 6496 44032 6500
rect 6299 6012 6363 6016
rect 6299 5956 6303 6012
rect 6303 5956 6359 6012
rect 6359 5956 6363 6012
rect 6299 5952 6363 5956
rect 6379 6012 6443 6016
rect 6379 5956 6383 6012
rect 6383 5956 6439 6012
rect 6439 5956 6443 6012
rect 6379 5952 6443 5956
rect 6459 6012 6523 6016
rect 6459 5956 6463 6012
rect 6463 5956 6519 6012
rect 6519 5956 6523 6012
rect 6459 5952 6523 5956
rect 6539 6012 6603 6016
rect 6539 5956 6543 6012
rect 6543 5956 6599 6012
rect 6599 5956 6603 6012
rect 6539 5952 6603 5956
rect 16993 6012 17057 6016
rect 16993 5956 16997 6012
rect 16997 5956 17053 6012
rect 17053 5956 17057 6012
rect 16993 5952 17057 5956
rect 17073 6012 17137 6016
rect 17073 5956 17077 6012
rect 17077 5956 17133 6012
rect 17133 5956 17137 6012
rect 17073 5952 17137 5956
rect 17153 6012 17217 6016
rect 17153 5956 17157 6012
rect 17157 5956 17213 6012
rect 17213 5956 17217 6012
rect 17153 5952 17217 5956
rect 17233 6012 17297 6016
rect 17233 5956 17237 6012
rect 17237 5956 17293 6012
rect 17293 5956 17297 6012
rect 17233 5952 17297 5956
rect 27687 6012 27751 6016
rect 27687 5956 27691 6012
rect 27691 5956 27747 6012
rect 27747 5956 27751 6012
rect 27687 5952 27751 5956
rect 27767 6012 27831 6016
rect 27767 5956 27771 6012
rect 27771 5956 27827 6012
rect 27827 5956 27831 6012
rect 27767 5952 27831 5956
rect 27847 6012 27911 6016
rect 27847 5956 27851 6012
rect 27851 5956 27907 6012
rect 27907 5956 27911 6012
rect 27847 5952 27911 5956
rect 27927 6012 27991 6016
rect 27927 5956 27931 6012
rect 27931 5956 27987 6012
rect 27987 5956 27991 6012
rect 27927 5952 27991 5956
rect 38381 6012 38445 6016
rect 38381 5956 38385 6012
rect 38385 5956 38441 6012
rect 38441 5956 38445 6012
rect 38381 5952 38445 5956
rect 38461 6012 38525 6016
rect 38461 5956 38465 6012
rect 38465 5956 38521 6012
rect 38521 5956 38525 6012
rect 38461 5952 38525 5956
rect 38541 6012 38605 6016
rect 38541 5956 38545 6012
rect 38545 5956 38601 6012
rect 38601 5956 38605 6012
rect 38541 5952 38605 5956
rect 38621 6012 38685 6016
rect 38621 5956 38625 6012
rect 38625 5956 38681 6012
rect 38681 5956 38685 6012
rect 38621 5952 38685 5956
rect 11646 5468 11710 5472
rect 11646 5412 11650 5468
rect 11650 5412 11706 5468
rect 11706 5412 11710 5468
rect 11646 5408 11710 5412
rect 11726 5468 11790 5472
rect 11726 5412 11730 5468
rect 11730 5412 11786 5468
rect 11786 5412 11790 5468
rect 11726 5408 11790 5412
rect 11806 5468 11870 5472
rect 11806 5412 11810 5468
rect 11810 5412 11866 5468
rect 11866 5412 11870 5468
rect 11806 5408 11870 5412
rect 11886 5468 11950 5472
rect 11886 5412 11890 5468
rect 11890 5412 11946 5468
rect 11946 5412 11950 5468
rect 11886 5408 11950 5412
rect 22340 5468 22404 5472
rect 22340 5412 22344 5468
rect 22344 5412 22400 5468
rect 22400 5412 22404 5468
rect 22340 5408 22404 5412
rect 22420 5468 22484 5472
rect 22420 5412 22424 5468
rect 22424 5412 22480 5468
rect 22480 5412 22484 5468
rect 22420 5408 22484 5412
rect 22500 5468 22564 5472
rect 22500 5412 22504 5468
rect 22504 5412 22560 5468
rect 22560 5412 22564 5468
rect 22500 5408 22564 5412
rect 22580 5468 22644 5472
rect 22580 5412 22584 5468
rect 22584 5412 22640 5468
rect 22640 5412 22644 5468
rect 22580 5408 22644 5412
rect 33034 5468 33098 5472
rect 33034 5412 33038 5468
rect 33038 5412 33094 5468
rect 33094 5412 33098 5468
rect 33034 5408 33098 5412
rect 33114 5468 33178 5472
rect 33114 5412 33118 5468
rect 33118 5412 33174 5468
rect 33174 5412 33178 5468
rect 33114 5408 33178 5412
rect 33194 5468 33258 5472
rect 33194 5412 33198 5468
rect 33198 5412 33254 5468
rect 33254 5412 33258 5468
rect 33194 5408 33258 5412
rect 33274 5468 33338 5472
rect 33274 5412 33278 5468
rect 33278 5412 33334 5468
rect 33334 5412 33338 5468
rect 33274 5408 33338 5412
rect 43728 5468 43792 5472
rect 43728 5412 43732 5468
rect 43732 5412 43788 5468
rect 43788 5412 43792 5468
rect 43728 5408 43792 5412
rect 43808 5468 43872 5472
rect 43808 5412 43812 5468
rect 43812 5412 43868 5468
rect 43868 5412 43872 5468
rect 43808 5408 43872 5412
rect 43888 5468 43952 5472
rect 43888 5412 43892 5468
rect 43892 5412 43948 5468
rect 43948 5412 43952 5468
rect 43888 5408 43952 5412
rect 43968 5468 44032 5472
rect 43968 5412 43972 5468
rect 43972 5412 44028 5468
rect 44028 5412 44032 5468
rect 43968 5408 44032 5412
rect 6299 4924 6363 4928
rect 6299 4868 6303 4924
rect 6303 4868 6359 4924
rect 6359 4868 6363 4924
rect 6299 4864 6363 4868
rect 6379 4924 6443 4928
rect 6379 4868 6383 4924
rect 6383 4868 6439 4924
rect 6439 4868 6443 4924
rect 6379 4864 6443 4868
rect 6459 4924 6523 4928
rect 6459 4868 6463 4924
rect 6463 4868 6519 4924
rect 6519 4868 6523 4924
rect 6459 4864 6523 4868
rect 6539 4924 6603 4928
rect 6539 4868 6543 4924
rect 6543 4868 6599 4924
rect 6599 4868 6603 4924
rect 6539 4864 6603 4868
rect 16993 4924 17057 4928
rect 16993 4868 16997 4924
rect 16997 4868 17053 4924
rect 17053 4868 17057 4924
rect 16993 4864 17057 4868
rect 17073 4924 17137 4928
rect 17073 4868 17077 4924
rect 17077 4868 17133 4924
rect 17133 4868 17137 4924
rect 17073 4864 17137 4868
rect 17153 4924 17217 4928
rect 17153 4868 17157 4924
rect 17157 4868 17213 4924
rect 17213 4868 17217 4924
rect 17153 4864 17217 4868
rect 17233 4924 17297 4928
rect 17233 4868 17237 4924
rect 17237 4868 17293 4924
rect 17293 4868 17297 4924
rect 17233 4864 17297 4868
rect 27687 4924 27751 4928
rect 27687 4868 27691 4924
rect 27691 4868 27747 4924
rect 27747 4868 27751 4924
rect 27687 4864 27751 4868
rect 27767 4924 27831 4928
rect 27767 4868 27771 4924
rect 27771 4868 27827 4924
rect 27827 4868 27831 4924
rect 27767 4864 27831 4868
rect 27847 4924 27911 4928
rect 27847 4868 27851 4924
rect 27851 4868 27907 4924
rect 27907 4868 27911 4924
rect 27847 4864 27911 4868
rect 27927 4924 27991 4928
rect 27927 4868 27931 4924
rect 27931 4868 27987 4924
rect 27987 4868 27991 4924
rect 27927 4864 27991 4868
rect 38381 4924 38445 4928
rect 38381 4868 38385 4924
rect 38385 4868 38441 4924
rect 38441 4868 38445 4924
rect 38381 4864 38445 4868
rect 38461 4924 38525 4928
rect 38461 4868 38465 4924
rect 38465 4868 38521 4924
rect 38521 4868 38525 4924
rect 38461 4864 38525 4868
rect 38541 4924 38605 4928
rect 38541 4868 38545 4924
rect 38545 4868 38601 4924
rect 38601 4868 38605 4924
rect 38541 4864 38605 4868
rect 38621 4924 38685 4928
rect 38621 4868 38625 4924
rect 38625 4868 38681 4924
rect 38681 4868 38685 4924
rect 38621 4864 38685 4868
rect 11646 4380 11710 4384
rect 11646 4324 11650 4380
rect 11650 4324 11706 4380
rect 11706 4324 11710 4380
rect 11646 4320 11710 4324
rect 11726 4380 11790 4384
rect 11726 4324 11730 4380
rect 11730 4324 11786 4380
rect 11786 4324 11790 4380
rect 11726 4320 11790 4324
rect 11806 4380 11870 4384
rect 11806 4324 11810 4380
rect 11810 4324 11866 4380
rect 11866 4324 11870 4380
rect 11806 4320 11870 4324
rect 11886 4380 11950 4384
rect 11886 4324 11890 4380
rect 11890 4324 11946 4380
rect 11946 4324 11950 4380
rect 11886 4320 11950 4324
rect 22340 4380 22404 4384
rect 22340 4324 22344 4380
rect 22344 4324 22400 4380
rect 22400 4324 22404 4380
rect 22340 4320 22404 4324
rect 22420 4380 22484 4384
rect 22420 4324 22424 4380
rect 22424 4324 22480 4380
rect 22480 4324 22484 4380
rect 22420 4320 22484 4324
rect 22500 4380 22564 4384
rect 22500 4324 22504 4380
rect 22504 4324 22560 4380
rect 22560 4324 22564 4380
rect 22500 4320 22564 4324
rect 22580 4380 22644 4384
rect 22580 4324 22584 4380
rect 22584 4324 22640 4380
rect 22640 4324 22644 4380
rect 22580 4320 22644 4324
rect 33034 4380 33098 4384
rect 33034 4324 33038 4380
rect 33038 4324 33094 4380
rect 33094 4324 33098 4380
rect 33034 4320 33098 4324
rect 33114 4380 33178 4384
rect 33114 4324 33118 4380
rect 33118 4324 33174 4380
rect 33174 4324 33178 4380
rect 33114 4320 33178 4324
rect 33194 4380 33258 4384
rect 33194 4324 33198 4380
rect 33198 4324 33254 4380
rect 33254 4324 33258 4380
rect 33194 4320 33258 4324
rect 33274 4380 33338 4384
rect 33274 4324 33278 4380
rect 33278 4324 33334 4380
rect 33334 4324 33338 4380
rect 33274 4320 33338 4324
rect 43728 4380 43792 4384
rect 43728 4324 43732 4380
rect 43732 4324 43788 4380
rect 43788 4324 43792 4380
rect 43728 4320 43792 4324
rect 43808 4380 43872 4384
rect 43808 4324 43812 4380
rect 43812 4324 43868 4380
rect 43868 4324 43872 4380
rect 43808 4320 43872 4324
rect 43888 4380 43952 4384
rect 43888 4324 43892 4380
rect 43892 4324 43948 4380
rect 43948 4324 43952 4380
rect 43888 4320 43952 4324
rect 43968 4380 44032 4384
rect 43968 4324 43972 4380
rect 43972 4324 44028 4380
rect 44028 4324 44032 4380
rect 43968 4320 44032 4324
rect 6299 3836 6363 3840
rect 6299 3780 6303 3836
rect 6303 3780 6359 3836
rect 6359 3780 6363 3836
rect 6299 3776 6363 3780
rect 6379 3836 6443 3840
rect 6379 3780 6383 3836
rect 6383 3780 6439 3836
rect 6439 3780 6443 3836
rect 6379 3776 6443 3780
rect 6459 3836 6523 3840
rect 6459 3780 6463 3836
rect 6463 3780 6519 3836
rect 6519 3780 6523 3836
rect 6459 3776 6523 3780
rect 6539 3836 6603 3840
rect 6539 3780 6543 3836
rect 6543 3780 6599 3836
rect 6599 3780 6603 3836
rect 6539 3776 6603 3780
rect 16993 3836 17057 3840
rect 16993 3780 16997 3836
rect 16997 3780 17053 3836
rect 17053 3780 17057 3836
rect 16993 3776 17057 3780
rect 17073 3836 17137 3840
rect 17073 3780 17077 3836
rect 17077 3780 17133 3836
rect 17133 3780 17137 3836
rect 17073 3776 17137 3780
rect 17153 3836 17217 3840
rect 17153 3780 17157 3836
rect 17157 3780 17213 3836
rect 17213 3780 17217 3836
rect 17153 3776 17217 3780
rect 17233 3836 17297 3840
rect 17233 3780 17237 3836
rect 17237 3780 17293 3836
rect 17293 3780 17297 3836
rect 17233 3776 17297 3780
rect 27687 3836 27751 3840
rect 27687 3780 27691 3836
rect 27691 3780 27747 3836
rect 27747 3780 27751 3836
rect 27687 3776 27751 3780
rect 27767 3836 27831 3840
rect 27767 3780 27771 3836
rect 27771 3780 27827 3836
rect 27827 3780 27831 3836
rect 27767 3776 27831 3780
rect 27847 3836 27911 3840
rect 27847 3780 27851 3836
rect 27851 3780 27907 3836
rect 27907 3780 27911 3836
rect 27847 3776 27911 3780
rect 27927 3836 27991 3840
rect 27927 3780 27931 3836
rect 27931 3780 27987 3836
rect 27987 3780 27991 3836
rect 27927 3776 27991 3780
rect 38381 3836 38445 3840
rect 38381 3780 38385 3836
rect 38385 3780 38441 3836
rect 38441 3780 38445 3836
rect 38381 3776 38445 3780
rect 38461 3836 38525 3840
rect 38461 3780 38465 3836
rect 38465 3780 38521 3836
rect 38521 3780 38525 3836
rect 38461 3776 38525 3780
rect 38541 3836 38605 3840
rect 38541 3780 38545 3836
rect 38545 3780 38601 3836
rect 38601 3780 38605 3836
rect 38541 3776 38605 3780
rect 38621 3836 38685 3840
rect 38621 3780 38625 3836
rect 38625 3780 38681 3836
rect 38681 3780 38685 3836
rect 38621 3776 38685 3780
rect 11646 3292 11710 3296
rect 11646 3236 11650 3292
rect 11650 3236 11706 3292
rect 11706 3236 11710 3292
rect 11646 3232 11710 3236
rect 11726 3292 11790 3296
rect 11726 3236 11730 3292
rect 11730 3236 11786 3292
rect 11786 3236 11790 3292
rect 11726 3232 11790 3236
rect 11806 3292 11870 3296
rect 11806 3236 11810 3292
rect 11810 3236 11866 3292
rect 11866 3236 11870 3292
rect 11806 3232 11870 3236
rect 11886 3292 11950 3296
rect 11886 3236 11890 3292
rect 11890 3236 11946 3292
rect 11946 3236 11950 3292
rect 11886 3232 11950 3236
rect 22340 3292 22404 3296
rect 22340 3236 22344 3292
rect 22344 3236 22400 3292
rect 22400 3236 22404 3292
rect 22340 3232 22404 3236
rect 22420 3292 22484 3296
rect 22420 3236 22424 3292
rect 22424 3236 22480 3292
rect 22480 3236 22484 3292
rect 22420 3232 22484 3236
rect 22500 3292 22564 3296
rect 22500 3236 22504 3292
rect 22504 3236 22560 3292
rect 22560 3236 22564 3292
rect 22500 3232 22564 3236
rect 22580 3292 22644 3296
rect 22580 3236 22584 3292
rect 22584 3236 22640 3292
rect 22640 3236 22644 3292
rect 22580 3232 22644 3236
rect 33034 3292 33098 3296
rect 33034 3236 33038 3292
rect 33038 3236 33094 3292
rect 33094 3236 33098 3292
rect 33034 3232 33098 3236
rect 33114 3292 33178 3296
rect 33114 3236 33118 3292
rect 33118 3236 33174 3292
rect 33174 3236 33178 3292
rect 33114 3232 33178 3236
rect 33194 3292 33258 3296
rect 33194 3236 33198 3292
rect 33198 3236 33254 3292
rect 33254 3236 33258 3292
rect 33194 3232 33258 3236
rect 33274 3292 33338 3296
rect 33274 3236 33278 3292
rect 33278 3236 33334 3292
rect 33334 3236 33338 3292
rect 33274 3232 33338 3236
rect 43728 3292 43792 3296
rect 43728 3236 43732 3292
rect 43732 3236 43788 3292
rect 43788 3236 43792 3292
rect 43728 3232 43792 3236
rect 43808 3292 43872 3296
rect 43808 3236 43812 3292
rect 43812 3236 43868 3292
rect 43868 3236 43872 3292
rect 43808 3232 43872 3236
rect 43888 3292 43952 3296
rect 43888 3236 43892 3292
rect 43892 3236 43948 3292
rect 43948 3236 43952 3292
rect 43888 3232 43952 3236
rect 43968 3292 44032 3296
rect 43968 3236 43972 3292
rect 43972 3236 44028 3292
rect 44028 3236 44032 3292
rect 43968 3232 44032 3236
rect 6299 2748 6363 2752
rect 6299 2692 6303 2748
rect 6303 2692 6359 2748
rect 6359 2692 6363 2748
rect 6299 2688 6363 2692
rect 6379 2748 6443 2752
rect 6379 2692 6383 2748
rect 6383 2692 6439 2748
rect 6439 2692 6443 2748
rect 6379 2688 6443 2692
rect 6459 2748 6523 2752
rect 6459 2692 6463 2748
rect 6463 2692 6519 2748
rect 6519 2692 6523 2748
rect 6459 2688 6523 2692
rect 6539 2748 6603 2752
rect 6539 2692 6543 2748
rect 6543 2692 6599 2748
rect 6599 2692 6603 2748
rect 6539 2688 6603 2692
rect 16993 2748 17057 2752
rect 16993 2692 16997 2748
rect 16997 2692 17053 2748
rect 17053 2692 17057 2748
rect 16993 2688 17057 2692
rect 17073 2748 17137 2752
rect 17073 2692 17077 2748
rect 17077 2692 17133 2748
rect 17133 2692 17137 2748
rect 17073 2688 17137 2692
rect 17153 2748 17217 2752
rect 17153 2692 17157 2748
rect 17157 2692 17213 2748
rect 17213 2692 17217 2748
rect 17153 2688 17217 2692
rect 17233 2748 17297 2752
rect 17233 2692 17237 2748
rect 17237 2692 17293 2748
rect 17293 2692 17297 2748
rect 17233 2688 17297 2692
rect 27687 2748 27751 2752
rect 27687 2692 27691 2748
rect 27691 2692 27747 2748
rect 27747 2692 27751 2748
rect 27687 2688 27751 2692
rect 27767 2748 27831 2752
rect 27767 2692 27771 2748
rect 27771 2692 27827 2748
rect 27827 2692 27831 2748
rect 27767 2688 27831 2692
rect 27847 2748 27911 2752
rect 27847 2692 27851 2748
rect 27851 2692 27907 2748
rect 27907 2692 27911 2748
rect 27847 2688 27911 2692
rect 27927 2748 27991 2752
rect 27927 2692 27931 2748
rect 27931 2692 27987 2748
rect 27987 2692 27991 2748
rect 27927 2688 27991 2692
rect 38381 2748 38445 2752
rect 38381 2692 38385 2748
rect 38385 2692 38441 2748
rect 38441 2692 38445 2748
rect 38381 2688 38445 2692
rect 38461 2748 38525 2752
rect 38461 2692 38465 2748
rect 38465 2692 38521 2748
rect 38521 2692 38525 2748
rect 38461 2688 38525 2692
rect 38541 2748 38605 2752
rect 38541 2692 38545 2748
rect 38545 2692 38601 2748
rect 38601 2692 38605 2748
rect 38541 2688 38605 2692
rect 38621 2748 38685 2752
rect 38621 2692 38625 2748
rect 38625 2692 38681 2748
rect 38681 2692 38685 2748
rect 38621 2688 38685 2692
rect 11646 2204 11710 2208
rect 11646 2148 11650 2204
rect 11650 2148 11706 2204
rect 11706 2148 11710 2204
rect 11646 2144 11710 2148
rect 11726 2204 11790 2208
rect 11726 2148 11730 2204
rect 11730 2148 11786 2204
rect 11786 2148 11790 2204
rect 11726 2144 11790 2148
rect 11806 2204 11870 2208
rect 11806 2148 11810 2204
rect 11810 2148 11866 2204
rect 11866 2148 11870 2204
rect 11806 2144 11870 2148
rect 11886 2204 11950 2208
rect 11886 2148 11890 2204
rect 11890 2148 11946 2204
rect 11946 2148 11950 2204
rect 11886 2144 11950 2148
rect 22340 2204 22404 2208
rect 22340 2148 22344 2204
rect 22344 2148 22400 2204
rect 22400 2148 22404 2204
rect 22340 2144 22404 2148
rect 22420 2204 22484 2208
rect 22420 2148 22424 2204
rect 22424 2148 22480 2204
rect 22480 2148 22484 2204
rect 22420 2144 22484 2148
rect 22500 2204 22564 2208
rect 22500 2148 22504 2204
rect 22504 2148 22560 2204
rect 22560 2148 22564 2204
rect 22500 2144 22564 2148
rect 22580 2204 22644 2208
rect 22580 2148 22584 2204
rect 22584 2148 22640 2204
rect 22640 2148 22644 2204
rect 22580 2144 22644 2148
rect 33034 2204 33098 2208
rect 33034 2148 33038 2204
rect 33038 2148 33094 2204
rect 33094 2148 33098 2204
rect 33034 2144 33098 2148
rect 33114 2204 33178 2208
rect 33114 2148 33118 2204
rect 33118 2148 33174 2204
rect 33174 2148 33178 2204
rect 33114 2144 33178 2148
rect 33194 2204 33258 2208
rect 33194 2148 33198 2204
rect 33198 2148 33254 2204
rect 33254 2148 33258 2204
rect 33194 2144 33258 2148
rect 33274 2204 33338 2208
rect 33274 2148 33278 2204
rect 33278 2148 33334 2204
rect 33334 2148 33338 2204
rect 33274 2144 33338 2148
rect 43728 2204 43792 2208
rect 43728 2148 43732 2204
rect 43732 2148 43788 2204
rect 43788 2148 43792 2204
rect 43728 2144 43792 2148
rect 43808 2204 43872 2208
rect 43808 2148 43812 2204
rect 43812 2148 43868 2204
rect 43868 2148 43872 2204
rect 43808 2144 43872 2148
rect 43888 2204 43952 2208
rect 43888 2148 43892 2204
rect 43892 2148 43948 2204
rect 43948 2148 43952 2204
rect 43888 2144 43952 2148
rect 43968 2204 44032 2208
rect 43968 2148 43972 2204
rect 43972 2148 44028 2204
rect 44028 2148 44032 2204
rect 43968 2144 44032 2148
rect 6299 1660 6363 1664
rect 6299 1604 6303 1660
rect 6303 1604 6359 1660
rect 6359 1604 6363 1660
rect 6299 1600 6363 1604
rect 6379 1660 6443 1664
rect 6379 1604 6383 1660
rect 6383 1604 6439 1660
rect 6439 1604 6443 1660
rect 6379 1600 6443 1604
rect 6459 1660 6523 1664
rect 6459 1604 6463 1660
rect 6463 1604 6519 1660
rect 6519 1604 6523 1660
rect 6459 1600 6523 1604
rect 6539 1660 6603 1664
rect 6539 1604 6543 1660
rect 6543 1604 6599 1660
rect 6599 1604 6603 1660
rect 6539 1600 6603 1604
rect 16993 1660 17057 1664
rect 16993 1604 16997 1660
rect 16997 1604 17053 1660
rect 17053 1604 17057 1660
rect 16993 1600 17057 1604
rect 17073 1660 17137 1664
rect 17073 1604 17077 1660
rect 17077 1604 17133 1660
rect 17133 1604 17137 1660
rect 17073 1600 17137 1604
rect 17153 1660 17217 1664
rect 17153 1604 17157 1660
rect 17157 1604 17213 1660
rect 17213 1604 17217 1660
rect 17153 1600 17217 1604
rect 17233 1660 17297 1664
rect 17233 1604 17237 1660
rect 17237 1604 17293 1660
rect 17293 1604 17297 1660
rect 17233 1600 17297 1604
rect 27687 1660 27751 1664
rect 27687 1604 27691 1660
rect 27691 1604 27747 1660
rect 27747 1604 27751 1660
rect 27687 1600 27751 1604
rect 27767 1660 27831 1664
rect 27767 1604 27771 1660
rect 27771 1604 27827 1660
rect 27827 1604 27831 1660
rect 27767 1600 27831 1604
rect 27847 1660 27911 1664
rect 27847 1604 27851 1660
rect 27851 1604 27907 1660
rect 27907 1604 27911 1660
rect 27847 1600 27911 1604
rect 27927 1660 27991 1664
rect 27927 1604 27931 1660
rect 27931 1604 27987 1660
rect 27987 1604 27991 1660
rect 27927 1600 27991 1604
rect 38381 1660 38445 1664
rect 38381 1604 38385 1660
rect 38385 1604 38441 1660
rect 38441 1604 38445 1660
rect 38381 1600 38445 1604
rect 38461 1660 38525 1664
rect 38461 1604 38465 1660
rect 38465 1604 38521 1660
rect 38521 1604 38525 1660
rect 38461 1600 38525 1604
rect 38541 1660 38605 1664
rect 38541 1604 38545 1660
rect 38545 1604 38601 1660
rect 38601 1604 38605 1660
rect 38541 1600 38605 1604
rect 38621 1660 38685 1664
rect 38621 1604 38625 1660
rect 38625 1604 38681 1660
rect 38681 1604 38685 1660
rect 38621 1600 38685 1604
rect 11646 1116 11710 1120
rect 11646 1060 11650 1116
rect 11650 1060 11706 1116
rect 11706 1060 11710 1116
rect 11646 1056 11710 1060
rect 11726 1116 11790 1120
rect 11726 1060 11730 1116
rect 11730 1060 11786 1116
rect 11786 1060 11790 1116
rect 11726 1056 11790 1060
rect 11806 1116 11870 1120
rect 11806 1060 11810 1116
rect 11810 1060 11866 1116
rect 11866 1060 11870 1116
rect 11806 1056 11870 1060
rect 11886 1116 11950 1120
rect 11886 1060 11890 1116
rect 11890 1060 11946 1116
rect 11946 1060 11950 1116
rect 11886 1056 11950 1060
rect 22340 1116 22404 1120
rect 22340 1060 22344 1116
rect 22344 1060 22400 1116
rect 22400 1060 22404 1116
rect 22340 1056 22404 1060
rect 22420 1116 22484 1120
rect 22420 1060 22424 1116
rect 22424 1060 22480 1116
rect 22480 1060 22484 1116
rect 22420 1056 22484 1060
rect 22500 1116 22564 1120
rect 22500 1060 22504 1116
rect 22504 1060 22560 1116
rect 22560 1060 22564 1116
rect 22500 1056 22564 1060
rect 22580 1116 22644 1120
rect 22580 1060 22584 1116
rect 22584 1060 22640 1116
rect 22640 1060 22644 1116
rect 22580 1056 22644 1060
rect 33034 1116 33098 1120
rect 33034 1060 33038 1116
rect 33038 1060 33094 1116
rect 33094 1060 33098 1116
rect 33034 1056 33098 1060
rect 33114 1116 33178 1120
rect 33114 1060 33118 1116
rect 33118 1060 33174 1116
rect 33174 1060 33178 1116
rect 33114 1056 33178 1060
rect 33194 1116 33258 1120
rect 33194 1060 33198 1116
rect 33198 1060 33254 1116
rect 33254 1060 33258 1116
rect 33194 1056 33258 1060
rect 33274 1116 33338 1120
rect 33274 1060 33278 1116
rect 33278 1060 33334 1116
rect 33334 1060 33338 1116
rect 33274 1056 33338 1060
rect 43728 1116 43792 1120
rect 43728 1060 43732 1116
rect 43732 1060 43788 1116
rect 43788 1060 43792 1116
rect 43728 1056 43792 1060
rect 43808 1116 43872 1120
rect 43808 1060 43812 1116
rect 43812 1060 43868 1116
rect 43868 1060 43872 1116
rect 43808 1056 43872 1060
rect 43888 1116 43952 1120
rect 43888 1060 43892 1116
rect 43892 1060 43948 1116
rect 43948 1060 43952 1116
rect 43888 1056 43952 1060
rect 43968 1116 44032 1120
rect 43968 1060 43972 1116
rect 43972 1060 44028 1116
rect 44028 1060 44032 1116
rect 43968 1056 44032 1060
<< metal4 >>
rect 20115 9892 20181 9893
rect 20115 9828 20116 9892
rect 20180 9828 20181 9892
rect 20115 9827 20181 9828
rect 19747 9076 19813 9077
rect 19747 9012 19748 9076
rect 19812 9012 19813 9076
rect 19747 9011 19813 9012
rect 6291 8192 6611 8752
rect 6291 8128 6299 8192
rect 6363 8128 6379 8192
rect 6443 8128 6459 8192
rect 6523 8128 6539 8192
rect 6603 8128 6611 8192
rect 6291 7104 6611 8128
rect 6291 7040 6299 7104
rect 6363 7040 6379 7104
rect 6443 7040 6459 7104
rect 6523 7040 6539 7104
rect 6603 7040 6611 7104
rect 6291 6016 6611 7040
rect 6291 5952 6299 6016
rect 6363 5952 6379 6016
rect 6443 5952 6459 6016
rect 6523 5952 6539 6016
rect 6603 5952 6611 6016
rect 6291 4928 6611 5952
rect 6291 4864 6299 4928
rect 6363 4864 6379 4928
rect 6443 4864 6459 4928
rect 6523 4864 6539 4928
rect 6603 4864 6611 4928
rect 6291 3840 6611 4864
rect 6291 3776 6299 3840
rect 6363 3776 6379 3840
rect 6443 3776 6459 3840
rect 6523 3776 6539 3840
rect 6603 3776 6611 3840
rect 6291 2752 6611 3776
rect 6291 2688 6299 2752
rect 6363 2688 6379 2752
rect 6443 2688 6459 2752
rect 6523 2688 6539 2752
rect 6603 2688 6611 2752
rect 6291 1664 6611 2688
rect 6291 1600 6299 1664
rect 6363 1600 6379 1664
rect 6443 1600 6459 1664
rect 6523 1600 6539 1664
rect 6603 1600 6611 1664
rect 6291 1040 6611 1600
rect 11638 8736 11958 8752
rect 11638 8672 11646 8736
rect 11710 8672 11726 8736
rect 11790 8672 11806 8736
rect 11870 8672 11886 8736
rect 11950 8672 11958 8736
rect 11638 7648 11958 8672
rect 11638 7584 11646 7648
rect 11710 7584 11726 7648
rect 11790 7584 11806 7648
rect 11870 7584 11886 7648
rect 11950 7584 11958 7648
rect 11638 6560 11958 7584
rect 11638 6496 11646 6560
rect 11710 6496 11726 6560
rect 11790 6496 11806 6560
rect 11870 6496 11886 6560
rect 11950 6496 11958 6560
rect 11638 5472 11958 6496
rect 11638 5408 11646 5472
rect 11710 5408 11726 5472
rect 11790 5408 11806 5472
rect 11870 5408 11886 5472
rect 11950 5408 11958 5472
rect 11638 4384 11958 5408
rect 11638 4320 11646 4384
rect 11710 4320 11726 4384
rect 11790 4320 11806 4384
rect 11870 4320 11886 4384
rect 11950 4320 11958 4384
rect 11638 3296 11958 4320
rect 11638 3232 11646 3296
rect 11710 3232 11726 3296
rect 11790 3232 11806 3296
rect 11870 3232 11886 3296
rect 11950 3232 11958 3296
rect 11638 2208 11958 3232
rect 11638 2144 11646 2208
rect 11710 2144 11726 2208
rect 11790 2144 11806 2208
rect 11870 2144 11886 2208
rect 11950 2144 11958 2208
rect 11638 1120 11958 2144
rect 11638 1056 11646 1120
rect 11710 1056 11726 1120
rect 11790 1056 11806 1120
rect 11870 1056 11886 1120
rect 11950 1056 11958 1120
rect 11638 1040 11958 1056
rect 16985 8192 17305 8752
rect 16985 8128 16993 8192
rect 17057 8128 17073 8192
rect 17137 8128 17153 8192
rect 17217 8128 17233 8192
rect 17297 8128 17305 8192
rect 16985 7104 17305 8128
rect 19379 8124 19445 8125
rect 19379 8060 19380 8124
rect 19444 8060 19445 8124
rect 19379 8059 19445 8060
rect 19382 7717 19442 8059
rect 19379 7716 19445 7717
rect 19379 7652 19380 7716
rect 19444 7652 19445 7716
rect 19379 7651 19445 7652
rect 19750 7309 19810 9011
rect 19931 8260 19997 8261
rect 19931 8196 19932 8260
rect 19996 8196 19997 8260
rect 19931 8195 19997 8196
rect 19747 7308 19813 7309
rect 19747 7244 19748 7308
rect 19812 7244 19813 7308
rect 19747 7243 19813 7244
rect 16985 7040 16993 7104
rect 17057 7040 17073 7104
rect 17137 7040 17153 7104
rect 17217 7040 17233 7104
rect 17297 7040 17305 7104
rect 16985 6016 17305 7040
rect 19934 7037 19994 8195
rect 20118 7037 20178 9827
rect 22332 8736 22652 8752
rect 22332 8672 22340 8736
rect 22404 8672 22420 8736
rect 22484 8672 22500 8736
rect 22564 8672 22580 8736
rect 22644 8672 22652 8736
rect 22332 7648 22652 8672
rect 22332 7584 22340 7648
rect 22404 7584 22420 7648
rect 22484 7584 22500 7648
rect 22564 7584 22580 7648
rect 22644 7584 22652 7648
rect 19931 7036 19997 7037
rect 19931 6972 19932 7036
rect 19996 6972 19997 7036
rect 19931 6971 19997 6972
rect 20115 7036 20181 7037
rect 20115 6972 20116 7036
rect 20180 6972 20181 7036
rect 20115 6971 20181 6972
rect 16985 5952 16993 6016
rect 17057 5952 17073 6016
rect 17137 5952 17153 6016
rect 17217 5952 17233 6016
rect 17297 5952 17305 6016
rect 16985 4928 17305 5952
rect 16985 4864 16993 4928
rect 17057 4864 17073 4928
rect 17137 4864 17153 4928
rect 17217 4864 17233 4928
rect 17297 4864 17305 4928
rect 16985 3840 17305 4864
rect 16985 3776 16993 3840
rect 17057 3776 17073 3840
rect 17137 3776 17153 3840
rect 17217 3776 17233 3840
rect 17297 3776 17305 3840
rect 16985 2752 17305 3776
rect 16985 2688 16993 2752
rect 17057 2688 17073 2752
rect 17137 2688 17153 2752
rect 17217 2688 17233 2752
rect 17297 2688 17305 2752
rect 16985 1664 17305 2688
rect 16985 1600 16993 1664
rect 17057 1600 17073 1664
rect 17137 1600 17153 1664
rect 17217 1600 17233 1664
rect 17297 1600 17305 1664
rect 16985 1040 17305 1600
rect 22332 6560 22652 7584
rect 22332 6496 22340 6560
rect 22404 6496 22420 6560
rect 22484 6496 22500 6560
rect 22564 6496 22580 6560
rect 22644 6496 22652 6560
rect 22332 5472 22652 6496
rect 22332 5408 22340 5472
rect 22404 5408 22420 5472
rect 22484 5408 22500 5472
rect 22564 5408 22580 5472
rect 22644 5408 22652 5472
rect 22332 4384 22652 5408
rect 22332 4320 22340 4384
rect 22404 4320 22420 4384
rect 22484 4320 22500 4384
rect 22564 4320 22580 4384
rect 22644 4320 22652 4384
rect 22332 3296 22652 4320
rect 22332 3232 22340 3296
rect 22404 3232 22420 3296
rect 22484 3232 22500 3296
rect 22564 3232 22580 3296
rect 22644 3232 22652 3296
rect 22332 2208 22652 3232
rect 22332 2144 22340 2208
rect 22404 2144 22420 2208
rect 22484 2144 22500 2208
rect 22564 2144 22580 2208
rect 22644 2144 22652 2208
rect 22332 1120 22652 2144
rect 22332 1056 22340 1120
rect 22404 1056 22420 1120
rect 22484 1056 22500 1120
rect 22564 1056 22580 1120
rect 22644 1056 22652 1120
rect 22332 1040 22652 1056
rect 27679 8192 27999 8752
rect 27679 8128 27687 8192
rect 27751 8128 27767 8192
rect 27831 8128 27847 8192
rect 27911 8128 27927 8192
rect 27991 8128 27999 8192
rect 27679 7104 27999 8128
rect 27679 7040 27687 7104
rect 27751 7040 27767 7104
rect 27831 7040 27847 7104
rect 27911 7040 27927 7104
rect 27991 7040 27999 7104
rect 27679 6016 27999 7040
rect 27679 5952 27687 6016
rect 27751 5952 27767 6016
rect 27831 5952 27847 6016
rect 27911 5952 27927 6016
rect 27991 5952 27999 6016
rect 27679 4928 27999 5952
rect 27679 4864 27687 4928
rect 27751 4864 27767 4928
rect 27831 4864 27847 4928
rect 27911 4864 27927 4928
rect 27991 4864 27999 4928
rect 27679 3840 27999 4864
rect 27679 3776 27687 3840
rect 27751 3776 27767 3840
rect 27831 3776 27847 3840
rect 27911 3776 27927 3840
rect 27991 3776 27999 3840
rect 27679 2752 27999 3776
rect 27679 2688 27687 2752
rect 27751 2688 27767 2752
rect 27831 2688 27847 2752
rect 27911 2688 27927 2752
rect 27991 2688 27999 2752
rect 27679 1664 27999 2688
rect 27679 1600 27687 1664
rect 27751 1600 27767 1664
rect 27831 1600 27847 1664
rect 27911 1600 27927 1664
rect 27991 1600 27999 1664
rect 27679 1040 27999 1600
rect 33026 8736 33346 8752
rect 33026 8672 33034 8736
rect 33098 8672 33114 8736
rect 33178 8672 33194 8736
rect 33258 8672 33274 8736
rect 33338 8672 33346 8736
rect 33026 7648 33346 8672
rect 33026 7584 33034 7648
rect 33098 7584 33114 7648
rect 33178 7584 33194 7648
rect 33258 7584 33274 7648
rect 33338 7584 33346 7648
rect 33026 6560 33346 7584
rect 33026 6496 33034 6560
rect 33098 6496 33114 6560
rect 33178 6496 33194 6560
rect 33258 6496 33274 6560
rect 33338 6496 33346 6560
rect 33026 5472 33346 6496
rect 33026 5408 33034 5472
rect 33098 5408 33114 5472
rect 33178 5408 33194 5472
rect 33258 5408 33274 5472
rect 33338 5408 33346 5472
rect 33026 4384 33346 5408
rect 33026 4320 33034 4384
rect 33098 4320 33114 4384
rect 33178 4320 33194 4384
rect 33258 4320 33274 4384
rect 33338 4320 33346 4384
rect 33026 3296 33346 4320
rect 33026 3232 33034 3296
rect 33098 3232 33114 3296
rect 33178 3232 33194 3296
rect 33258 3232 33274 3296
rect 33338 3232 33346 3296
rect 33026 2208 33346 3232
rect 33026 2144 33034 2208
rect 33098 2144 33114 2208
rect 33178 2144 33194 2208
rect 33258 2144 33274 2208
rect 33338 2144 33346 2208
rect 33026 1120 33346 2144
rect 33026 1056 33034 1120
rect 33098 1056 33114 1120
rect 33178 1056 33194 1120
rect 33258 1056 33274 1120
rect 33338 1056 33346 1120
rect 33026 1040 33346 1056
rect 38373 8192 38693 8752
rect 38373 8128 38381 8192
rect 38445 8128 38461 8192
rect 38525 8128 38541 8192
rect 38605 8128 38621 8192
rect 38685 8128 38693 8192
rect 38373 7104 38693 8128
rect 38373 7040 38381 7104
rect 38445 7040 38461 7104
rect 38525 7040 38541 7104
rect 38605 7040 38621 7104
rect 38685 7040 38693 7104
rect 38373 6016 38693 7040
rect 38373 5952 38381 6016
rect 38445 5952 38461 6016
rect 38525 5952 38541 6016
rect 38605 5952 38621 6016
rect 38685 5952 38693 6016
rect 38373 4928 38693 5952
rect 38373 4864 38381 4928
rect 38445 4864 38461 4928
rect 38525 4864 38541 4928
rect 38605 4864 38621 4928
rect 38685 4864 38693 4928
rect 38373 3840 38693 4864
rect 38373 3776 38381 3840
rect 38445 3776 38461 3840
rect 38525 3776 38541 3840
rect 38605 3776 38621 3840
rect 38685 3776 38693 3840
rect 38373 2752 38693 3776
rect 38373 2688 38381 2752
rect 38445 2688 38461 2752
rect 38525 2688 38541 2752
rect 38605 2688 38621 2752
rect 38685 2688 38693 2752
rect 38373 1664 38693 2688
rect 38373 1600 38381 1664
rect 38445 1600 38461 1664
rect 38525 1600 38541 1664
rect 38605 1600 38621 1664
rect 38685 1600 38693 1664
rect 38373 1040 38693 1600
rect 43720 8736 44040 8752
rect 43720 8672 43728 8736
rect 43792 8672 43808 8736
rect 43872 8672 43888 8736
rect 43952 8672 43968 8736
rect 44032 8672 44040 8736
rect 43720 7648 44040 8672
rect 43720 7584 43728 7648
rect 43792 7584 43808 7648
rect 43872 7584 43888 7648
rect 43952 7584 43968 7648
rect 44032 7584 44040 7648
rect 43720 6560 44040 7584
rect 43720 6496 43728 6560
rect 43792 6496 43808 6560
rect 43872 6496 43888 6560
rect 43952 6496 43968 6560
rect 44032 6496 44040 6560
rect 43720 5472 44040 6496
rect 43720 5408 43728 5472
rect 43792 5408 43808 5472
rect 43872 5408 43888 5472
rect 43952 5408 43968 5472
rect 44032 5408 44040 5472
rect 43720 4384 44040 5408
rect 43720 4320 43728 4384
rect 43792 4320 43808 4384
rect 43872 4320 43888 4384
rect 43952 4320 43968 4384
rect 44032 4320 44040 4384
rect 43720 3296 44040 4320
rect 43720 3232 43728 3296
rect 43792 3232 43808 3296
rect 43872 3232 43888 3296
rect 43952 3232 43968 3296
rect 44032 3232 44040 3296
rect 43720 2208 44040 3232
rect 43720 2144 43728 2208
rect 43792 2144 43808 2208
rect 43872 2144 43888 2208
rect 43952 2144 43968 2208
rect 44032 2144 44040 2208
rect 43720 1120 44040 2144
rect 43720 1056 43728 1120
rect 43792 1056 43808 1120
rect 43872 1056 43888 1120
rect 43952 1056 43968 1120
rect 44032 1056 44040 1120
rect 43720 1040 44040 1056
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 12696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 7912 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 6900 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1688980957
transform 1 0 6716 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_32
timestamp 1688980957
transform 1 0 4048 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_44 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_48 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_52
timestamp 1688980957
transform 1 0 5888 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_69 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_75
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_93
timestamp 1688980957
transform 1 0 9660 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_98
timestamp 1688980957
transform 1 0 10120 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 1688980957
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_117
timestamp 1688980957
transform 1 0 11868 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_121
timestamp 1688980957
transform 1 0 12236 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_133 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_144
timestamp 1688980957
transform 1 0 14352 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_156
timestamp 1688980957
transform 1 0 15456 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1688980957
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_190
timestamp 1688980957
transform 1 0 18584 0 1 1088
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_213
timestamp 1688980957
transform 1 0 20700 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_236
timestamp 1688980957
transform 1 0 22816 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_248
timestamp 1688980957
transform 1 0 23920 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_259
timestamp 1688980957
transform 1 0 24932 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_271
timestamp 1688980957
transform 1 0 26036 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_284
timestamp 1688980957
transform 1 0 27232 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_296
timestamp 1688980957
transform 1 0 28336 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1688980957
transform 1 0 29164 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_328
timestamp 1688980957
transform 1 0 31280 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_345
timestamp 1688980957
transform 1 0 32844 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_351
timestamp 1688980957
transform 1 0 33396 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_363
timestamp 1688980957
transform 1 0 34500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 1088
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_374
timestamp 1688980957
transform 1 0 35512 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_386
timestamp 1688980957
transform 1 0 36616 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_397
timestamp 1688980957
transform 1 0 37628 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_409
timestamp 1688980957
transform 1 0 38732 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_439
timestamp 1688980957
transform 1 0 41492 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_443
timestamp 1688980957
transform 1 0 41860 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_447
timestamp 1688980957
transform 1 0 42228 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_457
timestamp 1688980957
transform 1 0 43148 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_231
timestamp 1688980957
transform 1 0 22356 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_243
timestamp 1688980957
transform 1 0 23460 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_255
timestamp 1688980957
transform 1 0 24564 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_267
timestamp 1688980957
transform 1 0 25668 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_413
timestamp 1688980957
transform 1 0 39100 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_417
timestamp 1688980957
transform 1 0 39468 0 -1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_426
timestamp 1688980957
transform 1 0 40296 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_438
timestamp 1688980957
transform 1 0 41400 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_446
timestamp 1688980957
transform 1 0 42136 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_461
timestamp 1688980957
transform 1 0 43516 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_217
timestamp 1688980957
transform 1 0 21068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_239
timestamp 1688980957
transform 1 0 23092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_409
timestamp 1688980957
transform 1 0 38732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_414
timestamp 1688980957
transform 1 0 39192 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_424
timestamp 1688980957
transform 1 0 40112 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_436
timestamp 1688980957
transform 1 0 41216 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_448
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_460
timestamp 1688980957
transform 1 0 43424 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_189
timestamp 1688980957
transform 1 0 18492 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_195
timestamp 1688980957
transform 1 0 19044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_207
timestamp 1688980957
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_219
timestamp 1688980957
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_230
timestamp 1688980957
transform 1 0 22264 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_234
timestamp 1688980957
transform 1 0 22632 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_246
timestamp 1688980957
transform 1 0 23736 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_258
timestamp 1688980957
transform 1 0 24840 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_270
timestamp 1688980957
transform 1 0 25944 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_278
timestamp 1688980957
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_310
timestamp 1688980957
transform 1 0 29624 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_322
timestamp 1688980957
transform 1 0 30728 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_334
timestamp 1688980957
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_384
timestamp 1688980957
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_433
timestamp 1688980957
transform 1 0 40940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_445
timestamp 1688980957
transform 1 0 42044 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_203
timestamp 1688980957
transform 1 0 19780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_215
timestamp 1688980957
transform 1 0 20884 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_227
timestamp 1688980957
transform 1 0 21988 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_235
timestamp 1688980957
transform 1 0 22724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_241
timestamp 1688980957
transform 1 0 23276 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_249
timestamp 1688980957
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_318
timestamp 1688980957
transform 1 0 30360 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_330
timestamp 1688980957
transform 1 0 31464 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_342
timestamp 1688980957
transform 1 0 32568 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_354
timestamp 1688980957
transform 1 0 33672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_362
timestamp 1688980957
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_396
timestamp 1688980957
transform 1 0 37536 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_408
timestamp 1688980957
transform 1 0 38640 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_425
timestamp 1688980957
transform 1 0 40204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_437
timestamp 1688980957
transform 1 0 41308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_449
timestamp 1688980957
transform 1 0 42412 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_461
timestamp 1688980957
transform 1 0 43516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_213
timestamp 1688980957
transform 1 0 20700 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_218
timestamp 1688980957
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_245
timestamp 1688980957
transform 1 0 23644 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_264
timestamp 1688980957
transform 1 0 25392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_276
timestamp 1688980957
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_287
timestamp 1688980957
transform 1 0 27508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_299
timestamp 1688980957
transform 1 0 28612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_311
timestamp 1688980957
transform 1 0 29716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_323
timestamp 1688980957
transform 1 0 30820 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_333
timestamp 1688980957
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_400
timestamp 1688980957
transform 1 0 37904 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_412
timestamp 1688980957
transform 1 0 39008 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_424
timestamp 1688980957
transform 1 0 40112 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_436
timestamp 1688980957
transform 1 0 41216 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_226
timestamp 1688980957
transform 1 0 21896 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_232
timestamp 1688980957
transform 1 0 22448 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_272
timestamp 1688980957
transform 1 0 26128 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_284
timestamp 1688980957
transform 1 0 27232 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_295
timestamp 1688980957
transform 1 0 28244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_337
timestamp 1688980957
transform 1 0 32108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_341
timestamp 1688980957
transform 1 0 32476 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_353
timestamp 1688980957
transform 1 0 33580 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_361
timestamp 1688980957
transform 1 0 34316 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_385
timestamp 1688980957
transform 1 0 36524 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_406
timestamp 1688980957
transform 1 0 38456 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_418
timestamp 1688980957
transform 1 0 39560 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_461
timestamp 1688980957
transform 1 0 43516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_398
timestamp 1688980957
transform 1 0 37720 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_410
timestamp 1688980957
transform 1 0 38824 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_422
timestamp 1688980957
transform 1 0 39928 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_434
timestamp 1688980957
transform 1 0 41032 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_446
timestamp 1688980957
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_461
timestamp 1688980957
transform 1 0 43516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_61
timestamp 1688980957
transform 1 0 6716 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_193
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_461
timestamp 1688980957
transform 1 0 43516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_61
timestamp 1688980957
transform 1 0 6716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_72
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_76
timestamp 1688980957
transform 1 0 8096 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_88
timestamp 1688980957
transform 1 0 9200 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_100
timestamp 1688980957
transform 1 0 10304 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_120
timestamp 1688980957
transform 1 0 12144 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_130
timestamp 1688980957
transform 1 0 13064 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_142
timestamp 1688980957
transform 1 0 14168 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_154
timestamp 1688980957
transform 1 0 15272 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_177
timestamp 1688980957
transform 1 0 17388 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_184
timestamp 1688980957
transform 1 0 18032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_194
timestamp 1688980957
transform 1 0 18952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_208
timestamp 1688980957
transform 1 0 20240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_212
timestamp 1688980957
transform 1 0 20608 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_231
timestamp 1688980957
transform 1 0 22356 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_238
timestamp 1688980957
transform 1 0 23000 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_244
timestamp 1688980957
transform 1 0 23552 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_256
timestamp 1688980957
transform 1 0 24656 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_268
timestamp 1688980957
transform 1 0 25760 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_274
timestamp 1688980957
transform 1 0 26312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_278
timestamp 1688980957
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_461
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_47
timestamp 1688980957
transform 1 0 5428 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_66
timestamp 1688980957
transform 1 0 7176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_93
timestamp 1688980957
transform 1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_102
timestamp 1688980957
transform 1 0 10488 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_126
timestamp 1688980957
transform 1 0 12696 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_154
timestamp 1688980957
transform 1 0 15272 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_162
timestamp 1688980957
transform 1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_186
timestamp 1688980957
transform 1 0 18216 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1688980957
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_295
timestamp 1688980957
transform 1 0 28244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_359
timestamp 1688980957
transform 1 0 34132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_392
timestamp 1688980957
transform 1 0 37168 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_457
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_461
timestamp 1688980957
transform 1 0 43516 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_35
timestamp 1688980957
transform 1 0 4324 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_38
timestamp 1688980957
transform 1 0 4600 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_63
timestamp 1688980957
transform 1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_71
timestamp 1688980957
transform 1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_124
timestamp 1688980957
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_128
timestamp 1688980957
transform 1 0 12880 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_156
timestamp 1688980957
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_197
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_210
timestamp 1688980957
transform 1 0 20424 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_251
timestamp 1688980957
transform 1 0 24196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_358
timestamp 1688980957
transform 1 0 34040 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_363
timestamp 1688980957
transform 1 0 34500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_375
timestamp 1688980957
transform 1 0 35604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_389
timestamp 1688980957
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_417
timestamp 1688980957
transform 1 0 39468 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_439
timestamp 1688980957
transform 1 0 41492 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1688980957
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_461
timestamp 1688980957
transform 1 0 43516 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24656 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 26956 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 28888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 31004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 33120 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 35236 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 37352 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 39468 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 41584 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 43332 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 5612 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 11960 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 16192 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 20424 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 22540 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 20332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 18308 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 19688 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 21988 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 22264 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 22540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 23092 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 23368 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 23644 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 23920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 24932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 25208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 25484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 28336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 28612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 29532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 29808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 25760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform 1 0 26036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 26312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 27232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 27508 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 27784 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform 1 0 30084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1688980957
transform 1 0 32936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1688980957
transform 1 0 33488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform 1 0 33764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1688980957
transform 1 0 33580 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1688980957
transform 1 0 33856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1688980957
transform 1 0 30360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1688980957
transform 1 0 30636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1688980957
transform 1 0 30912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1688980957
transform 1 0 31188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1688980957
transform 1 0 31464 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1688980957
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1688980957
transform 1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1688980957
transform 1 0 32660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  inst_clk_buf
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__00_
timestamp 1688980957
transform 1 0 24932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__01_
timestamp 1688980957
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__02_
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__03_
timestamp 1688980957
transform 1 0 23552 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__04_
timestamp 1688980957
transform 1 0 23276 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__05_
timestamp 1688980957
transform 1 0 22724 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__06_
timestamp 1688980957
transform 1 0 22724 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__07_
timestamp 1688980957
transform 1 0 22172 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__08_
timestamp 1688980957
transform 1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__09_
timestamp 1688980957
transform 1 0 21620 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__10_
timestamp 1688980957
transform 1 0 21068 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__11_
timestamp 1688980957
transform 1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__12_
timestamp 1688980957
transform 1 0 20516 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__13_
timestamp 1688980957
transform 1 0 20792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__14_
timestamp 1688980957
transform 1 0 20240 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__15_
timestamp 1688980957
transform 1 0 19964 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__16_
timestamp 1688980957
transform 1 0 22448 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__17_
timestamp 1688980957
transform 1 0 23000 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__18_
timestamp 1688980957
transform 1 0 26864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__19_
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__20_
timestamp 1688980957
transform 1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__21_
timestamp 1688980957
transform 1 0 26036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__22_
timestamp 1688980957
transform 1 0 25760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__23_
timestamp 1688980957
transform 1 0 25208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__24_
timestamp 1688980957
transform 1 0 23276 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__25_
timestamp 1688980957
transform 1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__26_
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__27_
timestamp 1688980957
transform 1 0 26404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__28_
timestamp 1688980957
transform 1 0 27968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__29_
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__30_
timestamp 1688980957
transform 1 0 27416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__31_
timestamp 1688980957
transform 1 0 27140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__32_
timestamp 1688980957
transform 1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__33_
timestamp 1688980957
transform 1 0 20792 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__34_
timestamp 1688980957
transform 1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__35_
timestamp 1688980957
transform 1 0 18676 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__36_
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__37_
timestamp 1688980957
transform 1 0 18584 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__38_
timestamp 1688980957
transform 1 0 18584 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__39_
timestamp 1688980957
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__40_
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__41_
timestamp 1688980957
transform 1 0 22080 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__42_
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__43_
timestamp 1688980957
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__44_
timestamp 1688980957
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__45_
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__46_
timestamp 1688980957
transform 1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__47_
timestamp 1688980957
transform 1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__48_
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__49_
timestamp 1688980957
transform 1 0 19688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__50_
timestamp 1688980957
transform 1 0 19412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__51_
timestamp 1688980957
transform 1 0 19136 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 37444 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 38916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 39836 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 38548 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 40388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 40940 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 40388 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1688980957
transform 1 0 35420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 35788 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 36340 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 36064 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 36616 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 37812 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 4784 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 5520 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output96
timestamp 1688980957
transform 1 0 5336 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 6072 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1688980957
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 6624 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 7084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform 1 0 6992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1688980957
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 7728 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1688980957
transform 1 0 7360 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 7912 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1688980957
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 9108 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1688980957
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 9936 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1688980957
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1688980957
transform 1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 10304 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1688980957
transform 1 0 13064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 14352 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1688980957
transform 1 0 14904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1688980957
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 11040 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 11592 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1688980957
transform 1 0 11776 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 12144 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 11960 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1688980957
transform 1 0 11592 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1688980957
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 12880 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 17480 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1688980957
transform 1 0 18032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1688980957
transform 1 0 18400 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1688980957
transform 1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 19872 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 19320 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 15456 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1688980957
transform 1 0 14536 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1688980957
transform 1 0 15640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 16836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1688980957
transform 1 0 16744 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1688980957
transform 1 0 17112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 17664 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1688980957
transform 1 0 34132 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 43884 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 43884 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 43884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 43884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 43884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 43884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 43884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 43884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 43884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 43884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 43884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 22080 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform 1 0 22356 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 21528 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 20884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 27232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 29348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 31464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 36616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 36156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 37628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 39192 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 40664 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 40020 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 23092 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 23368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 21620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 27968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 30084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 32200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 37444 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 37260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 38180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 38916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 39928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 37168 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 3422 0 3478 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 24582 0 24638 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 26698 0 26754 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 28814 0 28870 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 30930 0 30986 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 33046 0 33102 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 35162 0 35218 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 37278 0 37334 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 39394 0 39450 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 41510 0 41566 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 43626 0 43682 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 5538 0 5594 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 7654 0 7710 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 9770 0 9826 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 11886 0 11942 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 14002 0 14058 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 16118 0 16174 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 18234 0 18290 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 20350 0 20406 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 22466 0 22522 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 34334 9840 34390 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 37094 9840 37150 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 37370 9840 37426 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 37646 9840 37702 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 37922 9840 37978 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 38198 9840 38254 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 38474 9840 38530 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 38750 9840 38806 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 39026 9840 39082 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 39302 9840 39358 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 39578 9840 39634 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 34610 9840 34666 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 34886 9840 34942 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 35162 9840 35218 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 35438 9840 35494 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 35714 9840 35770 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 35990 9840 36046 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 36266 9840 36322 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 36542 9840 36598 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 36818 9840 36874 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 5354 9840 5410 10000 0 FreeSans 224 90 0 0 N1BEG[0]
port 40 nsew signal tristate
flabel metal2 s 5630 9840 5686 10000 0 FreeSans 224 90 0 0 N1BEG[1]
port 41 nsew signal tristate
flabel metal2 s 5906 9840 5962 10000 0 FreeSans 224 90 0 0 N1BEG[2]
port 42 nsew signal tristate
flabel metal2 s 6182 9840 6238 10000 0 FreeSans 224 90 0 0 N1BEG[3]
port 43 nsew signal tristate
flabel metal2 s 6458 9840 6514 10000 0 FreeSans 224 90 0 0 N2BEG[0]
port 44 nsew signal tristate
flabel metal2 s 6734 9840 6790 10000 0 FreeSans 224 90 0 0 N2BEG[1]
port 45 nsew signal tristate
flabel metal2 s 7010 9840 7066 10000 0 FreeSans 224 90 0 0 N2BEG[2]
port 46 nsew signal tristate
flabel metal2 s 7286 9840 7342 10000 0 FreeSans 224 90 0 0 N2BEG[3]
port 47 nsew signal tristate
flabel metal2 s 7562 9840 7618 10000 0 FreeSans 224 90 0 0 N2BEG[4]
port 48 nsew signal tristate
flabel metal2 s 7838 9840 7894 10000 0 FreeSans 224 90 0 0 N2BEG[5]
port 49 nsew signal tristate
flabel metal2 s 8114 9840 8170 10000 0 FreeSans 224 90 0 0 N2BEG[6]
port 50 nsew signal tristate
flabel metal2 s 8390 9840 8446 10000 0 FreeSans 224 90 0 0 N2BEG[7]
port 51 nsew signal tristate
flabel metal2 s 8666 9840 8722 10000 0 FreeSans 224 90 0 0 N2BEGb[0]
port 52 nsew signal tristate
flabel metal2 s 8942 9840 8998 10000 0 FreeSans 224 90 0 0 N2BEGb[1]
port 53 nsew signal tristate
flabel metal2 s 9218 9840 9274 10000 0 FreeSans 224 90 0 0 N2BEGb[2]
port 54 nsew signal tristate
flabel metal2 s 9494 9840 9550 10000 0 FreeSans 224 90 0 0 N2BEGb[3]
port 55 nsew signal tristate
flabel metal2 s 9770 9840 9826 10000 0 FreeSans 224 90 0 0 N2BEGb[4]
port 56 nsew signal tristate
flabel metal2 s 10046 9840 10102 10000 0 FreeSans 224 90 0 0 N2BEGb[5]
port 57 nsew signal tristate
flabel metal2 s 10322 9840 10378 10000 0 FreeSans 224 90 0 0 N2BEGb[6]
port 58 nsew signal tristate
flabel metal2 s 10598 9840 10654 10000 0 FreeSans 224 90 0 0 N2BEGb[7]
port 59 nsew signal tristate
flabel metal2 s 10874 9840 10930 10000 0 FreeSans 224 90 0 0 N4BEG[0]
port 60 nsew signal tristate
flabel metal2 s 13634 9840 13690 10000 0 FreeSans 224 90 0 0 N4BEG[10]
port 61 nsew signal tristate
flabel metal2 s 13910 9840 13966 10000 0 FreeSans 224 90 0 0 N4BEG[11]
port 62 nsew signal tristate
flabel metal2 s 14186 9840 14242 10000 0 FreeSans 224 90 0 0 N4BEG[12]
port 63 nsew signal tristate
flabel metal2 s 14462 9840 14518 10000 0 FreeSans 224 90 0 0 N4BEG[13]
port 64 nsew signal tristate
flabel metal2 s 14738 9840 14794 10000 0 FreeSans 224 90 0 0 N4BEG[14]
port 65 nsew signal tristate
flabel metal2 s 15014 9840 15070 10000 0 FreeSans 224 90 0 0 N4BEG[15]
port 66 nsew signal tristate
flabel metal2 s 11150 9840 11206 10000 0 FreeSans 224 90 0 0 N4BEG[1]
port 67 nsew signal tristate
flabel metal2 s 11426 9840 11482 10000 0 FreeSans 224 90 0 0 N4BEG[2]
port 68 nsew signal tristate
flabel metal2 s 11702 9840 11758 10000 0 FreeSans 224 90 0 0 N4BEG[3]
port 69 nsew signal tristate
flabel metal2 s 11978 9840 12034 10000 0 FreeSans 224 90 0 0 N4BEG[4]
port 70 nsew signal tristate
flabel metal2 s 12254 9840 12310 10000 0 FreeSans 224 90 0 0 N4BEG[5]
port 71 nsew signal tristate
flabel metal2 s 12530 9840 12586 10000 0 FreeSans 224 90 0 0 N4BEG[6]
port 72 nsew signal tristate
flabel metal2 s 12806 9840 12862 10000 0 FreeSans 224 90 0 0 N4BEG[7]
port 73 nsew signal tristate
flabel metal2 s 13082 9840 13138 10000 0 FreeSans 224 90 0 0 N4BEG[8]
port 74 nsew signal tristate
flabel metal2 s 13358 9840 13414 10000 0 FreeSans 224 90 0 0 N4BEG[9]
port 75 nsew signal tristate
flabel metal2 s 15290 9840 15346 10000 0 FreeSans 224 90 0 0 NN4BEG[0]
port 76 nsew signal tristate
flabel metal2 s 18050 9840 18106 10000 0 FreeSans 224 90 0 0 NN4BEG[10]
port 77 nsew signal tristate
flabel metal2 s 18326 9840 18382 10000 0 FreeSans 224 90 0 0 NN4BEG[11]
port 78 nsew signal tristate
flabel metal2 s 18602 9840 18658 10000 0 FreeSans 224 90 0 0 NN4BEG[12]
port 79 nsew signal tristate
flabel metal2 s 18878 9840 18934 10000 0 FreeSans 224 90 0 0 NN4BEG[13]
port 80 nsew signal tristate
flabel metal2 s 19154 9840 19210 10000 0 FreeSans 224 90 0 0 NN4BEG[14]
port 81 nsew signal tristate
flabel metal2 s 19430 9840 19486 10000 0 FreeSans 224 90 0 0 NN4BEG[15]
port 82 nsew signal tristate
flabel metal2 s 15566 9840 15622 10000 0 FreeSans 224 90 0 0 NN4BEG[1]
port 83 nsew signal tristate
flabel metal2 s 15842 9840 15898 10000 0 FreeSans 224 90 0 0 NN4BEG[2]
port 84 nsew signal tristate
flabel metal2 s 16118 9840 16174 10000 0 FreeSans 224 90 0 0 NN4BEG[3]
port 85 nsew signal tristate
flabel metal2 s 16394 9840 16450 10000 0 FreeSans 224 90 0 0 NN4BEG[4]
port 86 nsew signal tristate
flabel metal2 s 16670 9840 16726 10000 0 FreeSans 224 90 0 0 NN4BEG[5]
port 87 nsew signal tristate
flabel metal2 s 16946 9840 17002 10000 0 FreeSans 224 90 0 0 NN4BEG[6]
port 88 nsew signal tristate
flabel metal2 s 17222 9840 17278 10000 0 FreeSans 224 90 0 0 NN4BEG[7]
port 89 nsew signal tristate
flabel metal2 s 17498 9840 17554 10000 0 FreeSans 224 90 0 0 NN4BEG[8]
port 90 nsew signal tristate
flabel metal2 s 17774 9840 17830 10000 0 FreeSans 224 90 0 0 NN4BEG[9]
port 91 nsew signal tristate
flabel metal2 s 19706 9840 19762 10000 0 FreeSans 224 90 0 0 S1END[0]
port 92 nsew signal input
flabel metal2 s 19982 9840 20038 10000 0 FreeSans 224 90 0 0 S1END[1]
port 93 nsew signal input
flabel metal2 s 20258 9840 20314 10000 0 FreeSans 224 90 0 0 S1END[2]
port 94 nsew signal input
flabel metal2 s 20534 9840 20590 10000 0 FreeSans 224 90 0 0 S1END[3]
port 95 nsew signal input
flabel metal2 s 20810 9840 20866 10000 0 FreeSans 224 90 0 0 S2END[0]
port 96 nsew signal input
flabel metal2 s 21086 9840 21142 10000 0 FreeSans 224 90 0 0 S2END[1]
port 97 nsew signal input
flabel metal2 s 21362 9840 21418 10000 0 FreeSans 224 90 0 0 S2END[2]
port 98 nsew signal input
flabel metal2 s 21638 9840 21694 10000 0 FreeSans 224 90 0 0 S2END[3]
port 99 nsew signal input
flabel metal2 s 21914 9840 21970 10000 0 FreeSans 224 90 0 0 S2END[4]
port 100 nsew signal input
flabel metal2 s 22190 9840 22246 10000 0 FreeSans 224 90 0 0 S2END[5]
port 101 nsew signal input
flabel metal2 s 22466 9840 22522 10000 0 FreeSans 224 90 0 0 S2END[6]
port 102 nsew signal input
flabel metal2 s 22742 9840 22798 10000 0 FreeSans 224 90 0 0 S2END[7]
port 103 nsew signal input
flabel metal2 s 23018 9840 23074 10000 0 FreeSans 224 90 0 0 S2MID[0]
port 104 nsew signal input
flabel metal2 s 23294 9840 23350 10000 0 FreeSans 224 90 0 0 S2MID[1]
port 105 nsew signal input
flabel metal2 s 23570 9840 23626 10000 0 FreeSans 224 90 0 0 S2MID[2]
port 106 nsew signal input
flabel metal2 s 23846 9840 23902 10000 0 FreeSans 224 90 0 0 S2MID[3]
port 107 nsew signal input
flabel metal2 s 24122 9840 24178 10000 0 FreeSans 224 90 0 0 S2MID[4]
port 108 nsew signal input
flabel metal2 s 24398 9840 24454 10000 0 FreeSans 224 90 0 0 S2MID[5]
port 109 nsew signal input
flabel metal2 s 24674 9840 24730 10000 0 FreeSans 224 90 0 0 S2MID[6]
port 110 nsew signal input
flabel metal2 s 24950 9840 25006 10000 0 FreeSans 224 90 0 0 S2MID[7]
port 111 nsew signal input
flabel metal2 s 25226 9840 25282 10000 0 FreeSans 224 90 0 0 S4END[0]
port 112 nsew signal input
flabel metal2 s 27986 9840 28042 10000 0 FreeSans 224 90 0 0 S4END[10]
port 113 nsew signal input
flabel metal2 s 28262 9840 28318 10000 0 FreeSans 224 90 0 0 S4END[11]
port 114 nsew signal input
flabel metal2 s 28538 9840 28594 10000 0 FreeSans 224 90 0 0 S4END[12]
port 115 nsew signal input
flabel metal2 s 28814 9840 28870 10000 0 FreeSans 224 90 0 0 S4END[13]
port 116 nsew signal input
flabel metal2 s 29090 9840 29146 10000 0 FreeSans 224 90 0 0 S4END[14]
port 117 nsew signal input
flabel metal2 s 29366 9840 29422 10000 0 FreeSans 224 90 0 0 S4END[15]
port 118 nsew signal input
flabel metal2 s 25502 9840 25558 10000 0 FreeSans 224 90 0 0 S4END[1]
port 119 nsew signal input
flabel metal2 s 25778 9840 25834 10000 0 FreeSans 224 90 0 0 S4END[2]
port 120 nsew signal input
flabel metal2 s 26054 9840 26110 10000 0 FreeSans 224 90 0 0 S4END[3]
port 121 nsew signal input
flabel metal2 s 26330 9840 26386 10000 0 FreeSans 224 90 0 0 S4END[4]
port 122 nsew signal input
flabel metal2 s 26606 9840 26662 10000 0 FreeSans 224 90 0 0 S4END[5]
port 123 nsew signal input
flabel metal2 s 26882 9840 26938 10000 0 FreeSans 224 90 0 0 S4END[6]
port 124 nsew signal input
flabel metal2 s 27158 9840 27214 10000 0 FreeSans 224 90 0 0 S4END[7]
port 125 nsew signal input
flabel metal2 s 27434 9840 27490 10000 0 FreeSans 224 90 0 0 S4END[8]
port 126 nsew signal input
flabel metal2 s 27710 9840 27766 10000 0 FreeSans 224 90 0 0 S4END[9]
port 127 nsew signal input
flabel metal2 s 29642 9840 29698 10000 0 FreeSans 224 90 0 0 SS4END[0]
port 128 nsew signal input
flabel metal2 s 32402 9840 32458 10000 0 FreeSans 224 90 0 0 SS4END[10]
port 129 nsew signal input
flabel metal2 s 32678 9840 32734 10000 0 FreeSans 224 90 0 0 SS4END[11]
port 130 nsew signal input
flabel metal2 s 32954 9840 33010 10000 0 FreeSans 224 90 0 0 SS4END[12]
port 131 nsew signal input
flabel metal2 s 33230 9840 33286 10000 0 FreeSans 224 90 0 0 SS4END[13]
port 132 nsew signal input
flabel metal2 s 33506 9840 33562 10000 0 FreeSans 224 90 0 0 SS4END[14]
port 133 nsew signal input
flabel metal2 s 33782 9840 33838 10000 0 FreeSans 224 90 0 0 SS4END[15]
port 134 nsew signal input
flabel metal2 s 29918 9840 29974 10000 0 FreeSans 224 90 0 0 SS4END[1]
port 135 nsew signal input
flabel metal2 s 30194 9840 30250 10000 0 FreeSans 224 90 0 0 SS4END[2]
port 136 nsew signal input
flabel metal2 s 30470 9840 30526 10000 0 FreeSans 224 90 0 0 SS4END[3]
port 137 nsew signal input
flabel metal2 s 30746 9840 30802 10000 0 FreeSans 224 90 0 0 SS4END[4]
port 138 nsew signal input
flabel metal2 s 31022 9840 31078 10000 0 FreeSans 224 90 0 0 SS4END[5]
port 139 nsew signal input
flabel metal2 s 31298 9840 31354 10000 0 FreeSans 224 90 0 0 SS4END[6]
port 140 nsew signal input
flabel metal2 s 31574 9840 31630 10000 0 FreeSans 224 90 0 0 SS4END[7]
port 141 nsew signal input
flabel metal2 s 31850 9840 31906 10000 0 FreeSans 224 90 0 0 SS4END[8]
port 142 nsew signal input
flabel metal2 s 32126 9840 32182 10000 0 FreeSans 224 90 0 0 SS4END[9]
port 143 nsew signal input
flabel metal2 s 1306 0 1362 160 0 FreeSans 224 90 0 0 UserCLK
port 144 nsew signal input
flabel metal2 s 34058 9840 34114 10000 0 FreeSans 224 90 0 0 UserCLKo
port 145 nsew signal tristate
flabel metal4 s 6291 1040 6611 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 16985 1040 17305 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 27679 1040 27999 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 38373 1040 38693 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 11638 1040 11958 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 22332 1040 22652 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 33026 1040 33346 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 43720 1040 44040 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
rlabel metal1 22494 8160 22494 8160 0 vccd1
rlabel via1 22572 8704 22572 8704 0 vssd1
rlabel metal2 3641 68 3641 68 0 FrameStrobe[0]
rlabel metal2 24755 68 24755 68 0 FrameStrobe[10]
rlabel metal2 26726 704 26726 704 0 FrameStrobe[11]
rlabel metal2 28987 68 28987 68 0 FrameStrobe[12]
rlabel metal2 31103 68 31103 68 0 FrameStrobe[13]
rlabel metal2 33265 68 33265 68 0 FrameStrobe[14]
rlabel metal2 35335 68 35335 68 0 FrameStrobe[15]
rlabel metal2 37451 68 37451 68 0 FrameStrobe[16]
rlabel metal2 39422 704 39422 704 0 FrameStrobe[17]
rlabel metal2 41683 68 41683 68 0 FrameStrobe[18]
rlabel metal2 43601 68 43601 68 0 FrameStrobe[19]
rlabel metal2 5619 68 5619 68 0 FrameStrobe[1]
rlabel metal2 7735 68 7735 68 0 FrameStrobe[2]
rlabel metal2 9851 68 9851 68 0 FrameStrobe[3]
rlabel metal2 11967 68 11967 68 0 FrameStrobe[4]
rlabel metal2 14175 68 14175 68 0 FrameStrobe[5]
rlabel metal2 16291 68 16291 68 0 FrameStrobe[6]
rlabel metal2 18407 68 18407 68 0 FrameStrobe[7]
rlabel metal2 20523 68 20523 68 0 FrameStrobe[8]
rlabel metal2 22639 68 22639 68 0 FrameStrobe[9]
rlabel metal2 34362 9462 34362 9462 0 FrameStrobe_O[0]
rlabel metal2 37122 9037 37122 9037 0 FrameStrobe_O[10]
rlabel metal2 37398 8952 37398 8952 0 FrameStrobe_O[11]
rlabel metal2 37674 9156 37674 9156 0 FrameStrobe_O[12]
rlabel metal2 37950 9445 37950 9445 0 FrameStrobe_O[13]
rlabel metal1 38778 6834 38778 6834 0 FrameStrobe_O[14]
rlabel metal2 38502 9088 38502 9088 0 FrameStrobe_O[15]
rlabel metal2 38778 9309 38778 9309 0 FrameStrobe_O[16]
rlabel metal2 39054 9836 39054 9836 0 FrameStrobe_O[17]
rlabel metal2 39330 9224 39330 9224 0 FrameStrobe_O[18]
rlabel metal2 39606 9836 39606 9836 0 FrameStrobe_O[19]
rlabel metal1 35052 8330 35052 8330 0 FrameStrobe_O[1]
rlabel metal1 35282 8058 35282 8058 0 FrameStrobe_O[2]
rlabel metal2 35190 9224 35190 9224 0 FrameStrobe_O[3]
rlabel metal1 36570 8568 36570 8568 0 FrameStrobe_O[4]
rlabel metal2 35742 9088 35742 9088 0 FrameStrobe_O[5]
rlabel metal2 36018 8952 36018 8952 0 FrameStrobe_O[6]
rlabel metal2 36294 9309 36294 9309 0 FrameStrobe_O[7]
rlabel metal2 36570 9122 36570 9122 0 FrameStrobe_O[8]
rlabel metal2 36846 9326 36846 9326 0 FrameStrobe_O[9]
rlabel metal1 22494 2074 22494 2074 0 FrameStrobe_O_i\[0\]
rlabel metal1 25530 4250 25530 4250 0 FrameStrobe_O_i\[10\]
rlabel metal1 27646 3978 27646 3978 0 FrameStrobe_O_i\[11\]
rlabel metal1 29762 3162 29762 3162 0 FrameStrobe_O_i\[12\]
rlabel metal1 32246 4012 32246 4012 0 FrameStrobe_O_i\[13\]
rlabel metal1 37168 4794 37168 4794 0 FrameStrobe_O_i\[14\]
rlabel metal1 36846 3162 36846 3162 0 FrameStrobe_O_i\[15\]
rlabel metal1 38042 4250 38042 4250 0 FrameStrobe_O_i\[16\]
rlabel metal1 39192 2074 39192 2074 0 FrameStrobe_O_i\[17\]
rlabel metal1 40434 3162 40434 3162 0 FrameStrobe_O_i\[18\]
rlabel metal2 40066 2244 40066 2244 0 FrameStrobe_O_i\[19\]
rlabel metal2 22218 4284 22218 4284 0 FrameStrobe_O_i\[1\]
rlabel metal1 22126 4216 22126 4216 0 FrameStrobe_O_i\[2\]
rlabel metal1 22770 3910 22770 3910 0 FrameStrobe_O_i\[3\]
rlabel metal1 23046 4250 23046 4250 0 FrameStrobe_O_i\[4\]
rlabel metal1 21988 2550 21988 2550 0 FrameStrobe_O_i\[5\]
rlabel metal1 21666 2618 21666 2618 0 FrameStrobe_O_i\[6\]
rlabel metal1 19182 3162 19182 3162 0 FrameStrobe_O_i\[7\]
rlabel metal1 21298 4250 21298 4250 0 FrameStrobe_O_i\[8\]
rlabel metal1 23414 3706 23414 3706 0 FrameStrobe_O_i\[9\]
rlabel metal1 5290 8602 5290 8602 0 N1BEG[0]
rlabel metal2 5658 9309 5658 9309 0 N1BEG[1]
rlabel metal1 5842 8602 5842 8602 0 N1BEG[2]
rlabel metal2 6210 8952 6210 8952 0 N1BEG[3]
rlabel metal1 6394 7514 6394 7514 0 N2BEG[0]
rlabel metal2 6762 9037 6762 9037 0 N2BEG[1]
rlabel metal2 7038 9224 7038 9224 0 N2BEG[2]
rlabel metal1 7268 7514 7268 7514 0 N2BEG[3]
rlabel metal2 7590 8952 7590 8952 0 N2BEG[4]
rlabel metal2 7866 8952 7866 8952 0 N2BEG[5]
rlabel metal1 7590 7276 7590 7276 0 N2BEG[6]
rlabel metal2 8418 8952 8418 8952 0 N2BEG[7]
rlabel metal1 8510 8602 8510 8602 0 N2BEGb[0]
rlabel metal2 8970 9173 8970 9173 0 N2BEGb[1]
rlabel metal2 9246 8952 9246 8952 0 N2BEGb[2]
rlabel metal1 8694 8432 8694 8432 0 N2BEGb[3]
rlabel metal2 9798 9224 9798 9224 0 N2BEGb[4]
rlabel metal2 10074 8952 10074 8952 0 N2BEGb[5]
rlabel metal1 9890 6834 9890 6834 0 N2BEGb[6]
rlabel metal1 10396 8602 10396 8602 0 N2BEGb[7]
rlabel metal1 10810 8602 10810 8602 0 N4BEG[0]
rlabel metal1 13478 8602 13478 8602 0 N4BEG[10]
rlabel metal1 13892 8058 13892 8058 0 N4BEG[11]
rlabel metal1 14030 8602 14030 8602 0 N4BEG[12]
rlabel metal2 14490 9309 14490 9309 0 N4BEG[13]
rlabel metal1 14950 8058 14950 8058 0 N4BEG[14]
rlabel metal1 14720 8602 14720 8602 0 N4BEG[15]
rlabel metal2 11178 8952 11178 8952 0 N4BEG[1]
rlabel metal1 11362 8602 11362 8602 0 N4BEG[2]
rlabel metal2 11730 9377 11730 9377 0 N4BEG[3]
rlabel metal2 12006 8680 12006 8680 0 N4BEG[4]
rlabel metal2 12282 8918 12282 8918 0 N4BEG[5]
rlabel metal2 12558 9224 12558 9224 0 N4BEG[6]
rlabel metal2 12834 9836 12834 9836 0 N4BEG[7]
rlabel metal1 13018 7514 13018 7514 0 N4BEG[8]
rlabel metal1 13340 8058 13340 8058 0 N4BEG[9]
rlabel metal2 15318 9224 15318 9224 0 NN4BEG[0]
rlabel metal2 17894 9231 17894 9231 0 NN4BEG[10]
rlabel metal1 18308 8602 18308 8602 0 NN4BEG[11]
rlabel metal2 18630 9224 18630 9224 0 NN4BEG[12]
rlabel metal1 18952 8602 18952 8602 0 NN4BEG[13]
rlabel metal2 19182 9836 19182 9836 0 NN4BEG[14]
rlabel metal2 19458 9224 19458 9224 0 NN4BEG[15]
rlabel metal2 15594 9309 15594 9309 0 NN4BEG[1]
rlabel metal1 14720 8330 14720 8330 0 NN4BEG[2]
rlabel metal1 16008 8602 16008 8602 0 NN4BEG[3]
rlabel metal2 16422 8918 16422 8918 0 NN4BEG[4]
rlabel metal1 16468 8602 16468 8602 0 NN4BEG[5]
rlabel metal2 16974 9309 16974 9309 0 NN4BEG[6]
rlabel metal1 17112 8602 17112 8602 0 NN4BEG[7]
rlabel metal1 17434 8602 17434 8602 0 NN4BEG[8]
rlabel metal2 17802 8918 17802 8918 0 NN4BEG[9]
rlabel metal2 19734 9037 19734 9037 0 S1END[0]
rlabel metal2 20010 9836 20010 9836 0 S1END[1]
rlabel metal2 20286 8884 20286 8884 0 S1END[2]
rlabel metal2 20562 9836 20562 9836 0 S1END[3]
rlabel metal2 20838 9836 20838 9836 0 S2END[0]
rlabel metal2 21114 9836 21114 9836 0 S2END[1]
rlabel metal2 21390 9836 21390 9836 0 S2END[2]
rlabel metal2 21666 9156 21666 9156 0 S2END[3]
rlabel metal2 21942 9513 21942 9513 0 S2END[4]
rlabel metal2 22218 9156 22218 9156 0 S2END[5]
rlabel metal2 22494 9513 22494 9513 0 S2END[6]
rlabel metal2 22770 9581 22770 9581 0 S2END[7]
rlabel metal2 23046 9513 23046 9513 0 S2MID[0]
rlabel metal2 23322 9513 23322 9513 0 S2MID[1]
rlabel metal2 23598 9513 23598 9513 0 S2MID[2]
rlabel metal2 23874 9513 23874 9513 0 S2MID[3]
rlabel metal2 24150 9513 24150 9513 0 S2MID[4]
rlabel metal2 24426 9190 24426 9190 0 S2MID[5]
rlabel metal2 24702 9224 24702 9224 0 S2MID[6]
rlabel metal2 24978 9122 24978 9122 0 S2MID[7]
rlabel metal2 25254 9190 25254 9190 0 S4END[0]
rlabel metal2 28014 9224 28014 9224 0 S4END[10]
rlabel metal2 28290 9224 28290 9224 0 S4END[11]
rlabel metal2 28566 9088 28566 9088 0 S4END[12]
rlabel metal2 28842 9513 28842 9513 0 S4END[13]
rlabel metal2 29118 9224 29118 9224 0 S4END[14]
rlabel metal2 29394 9122 29394 9122 0 S4END[15]
rlabel metal2 25530 9224 25530 9224 0 S4END[1]
rlabel metal2 25806 9156 25806 9156 0 S4END[2]
rlabel metal2 26082 9513 26082 9513 0 S4END[3]
rlabel metal2 26358 9224 26358 9224 0 S4END[4]
rlabel metal2 26634 9156 26634 9156 0 S4END[5]
rlabel metal2 26910 9513 26910 9513 0 S4END[6]
rlabel metal2 27186 9224 27186 9224 0 S4END[7]
rlabel metal2 27462 9122 27462 9122 0 S4END[8]
rlabel metal2 27738 9513 27738 9513 0 S4END[9]
rlabel metal2 29670 9190 29670 9190 0 SS4END[0]
rlabel metal2 32430 9190 32430 9190 0 SS4END[10]
rlabel metal2 32706 9224 32706 9224 0 SS4END[11]
rlabel metal2 32982 9156 32982 9156 0 SS4END[12]
rlabel metal2 33258 9513 33258 9513 0 SS4END[13]
rlabel metal2 33534 8850 33534 8850 0 SS4END[14]
rlabel metal2 33810 8850 33810 8850 0 SS4END[15]
rlabel metal2 29946 9122 29946 9122 0 SS4END[1]
rlabel metal2 30222 9190 30222 9190 0 SS4END[2]
rlabel metal2 30498 9224 30498 9224 0 SS4END[3]
rlabel metal2 30774 9122 30774 9122 0 SS4END[4]
rlabel metal2 31050 9190 31050 9190 0 SS4END[5]
rlabel metal1 31786 8432 31786 8432 0 SS4END[6]
rlabel metal1 32154 8500 32154 8500 0 SS4END[7]
rlabel metal2 31878 9224 31878 9224 0 SS4END[8]
rlabel metal2 32154 9122 32154 9122 0 SS4END[9]
rlabel metal2 1334 704 1334 704 0 UserCLK
rlabel metal1 34224 8602 34224 8602 0 UserCLKo
rlabel metal2 4002 1700 4002 1700 0 net1
rlabel metal1 41262 1190 41262 1190 0 net10
rlabel metal1 7728 8534 7728 8534 0 net100
rlabel metal2 7038 6851 7038 6851 0 net101
rlabel metal1 7820 7854 7820 7854 0 net102
rlabel metal1 11086 7786 11086 7786 0 net103
rlabel metal2 7406 7820 7406 7820 0 net104
rlabel metal2 8418 7514 8418 7514 0 net105
rlabel metal2 8050 7990 8050 7990 0 net106
rlabel metal1 7268 6766 7268 6766 0 net107
rlabel metal2 9246 7548 9246 7548 0 net108
rlabel metal1 8326 9520 8326 9520 0 net109
rlabel metal2 43378 1734 43378 1734 0 net11
rlabel metal2 9890 8636 9890 8636 0 net110
rlabel metal2 10074 7378 10074 7378 0 net111
rlabel metal1 9062 9860 9062 9860 0 net112
rlabel metal1 9982 9282 9982 9282 0 net113
rlabel metal1 10442 9520 10442 9520 0 net114
rlabel metal1 13294 8466 13294 8466 0 net115
rlabel metal2 15502 6970 15502 6970 0 net116
rlabel metal2 16054 8976 16054 8976 0 net117
rlabel metal2 16698 7004 16698 7004 0 net118
rlabel metal2 17618 6834 17618 6834 0 net119
rlabel metal1 5842 1258 5842 1258 0 net12
rlabel metal1 14398 9452 14398 9452 0 net120
rlabel metal1 12374 8024 12374 8024 0 net121
rlabel metal1 10994 8432 10994 8432 0 net122
rlabel metal1 11730 7854 11730 7854 0 net123
rlabel metal1 11822 7412 11822 7412 0 net124
rlabel metal2 12282 7004 12282 7004 0 net125
rlabel metal2 12098 8738 12098 8738 0 net126
rlabel metal1 12029 8466 12029 8466 0 net127
rlabel metal2 12742 8279 12742 8279 0 net128
rlabel metal2 13018 7905 13018 7905 0 net129
rlabel metal2 7958 2618 7958 2618 0 net13
rlabel metal1 15594 8398 15594 8398 0 net130
rlabel metal1 18262 7174 18262 7174 0 net131
rlabel metal1 18584 7514 18584 7514 0 net132
rlabel metal2 17434 8228 17434 8228 0 net133
rlabel metal1 18676 6630 18676 6630 0 net134
rlabel metal1 19090 7718 19090 7718 0 net135
rlabel metal2 18906 8262 18906 8262 0 net136
rlabel metal1 15594 7752 15594 7752 0 net137
rlabel metal1 18630 8466 18630 8466 0 net138
rlabel metal1 17342 8364 17342 8364 0 net139
rlabel metal1 14214 1224 14214 1224 0 net14
rlabel metal1 18262 7378 18262 7378 0 net140
rlabel metal1 16146 8500 16146 8500 0 net141
rlabel metal1 16974 7888 16974 7888 0 net142
rlabel metal1 17296 7174 17296 7174 0 net143
rlabel metal2 17526 7990 17526 7990 0 net144
rlabel metal1 17986 7514 17986 7514 0 net145
rlabel metal1 28106 1802 28106 1802 0 net146
rlabel metal2 18170 1088 18170 1088 0 net15
rlabel metal2 21758 1700 21758 1700 0 net16
rlabel metal1 18446 1292 18446 1292 0 net17
rlabel metal1 18676 1190 18676 1190 0 net18
rlabel metal1 20516 1190 20516 1190 0 net19
rlabel metal1 24748 1190 24748 1190 0 net2
rlabel metal1 22908 1190 22908 1190 0 net20
rlabel metal1 19504 6630 19504 6630 0 net21
rlabel metal1 19826 6970 19826 6970 0 net22
rlabel metal1 19780 7378 19780 7378 0 net23
rlabel metal1 20010 7412 20010 7412 0 net24
rlabel metal1 20010 7820 20010 7820 0 net25
rlabel metal1 20378 7830 20378 7830 0 net26
rlabel metal1 20884 7378 20884 7378 0 net27
rlabel metal1 20562 7888 20562 7888 0 net28
rlabel metal1 21574 7378 21574 7378 0 net29
rlabel metal1 27232 1190 27232 1190 0 net3
rlabel metal2 21114 8058 21114 8058 0 net30
rlabel metal2 21666 8092 21666 8092 0 net31
rlabel metal1 21942 7888 21942 7888 0 net32
rlabel metal1 22218 7820 22218 7820 0 net33
rlabel viali 22770 7380 22770 7380 0 net34
rlabel metal1 22770 7922 22770 7922 0 net35
rlabel metal1 23644 7378 23644 7378 0 net36
rlabel metal1 23598 7888 23598 7888 0 net37
rlabel metal1 24472 7854 24472 7854 0 net38
rlabel metal1 24794 7854 24794 7854 0 net39
rlabel metal1 28934 1258 28934 1258 0 net4
rlabel metal1 25024 7854 25024 7854 0 net40
rlabel metal1 25300 7854 25300 7854 0 net41
rlabel metal1 27416 7378 27416 7378 0 net42
rlabel metal1 25530 7922 25530 7922 0 net43
rlabel metal1 24104 7854 24104 7854 0 net44
rlabel via1 23318 7854 23318 7854 0 net45
rlabel metal1 23046 7888 23046 7888 0 net46
rlabel metal1 22586 7854 22586 7854 0 net47
rlabel metal2 25806 8058 25806 8058 0 net48
rlabel metal2 26082 8058 26082 8058 0 net49
rlabel metal1 31372 1190 31372 1190 0 net5
rlabel metal2 26358 8058 26358 8058 0 net50
rlabel metal2 26634 8058 26634 8058 0 net51
rlabel metal1 26956 7854 26956 7854 0 net52
rlabel metal1 27232 7854 27232 7854 0 net53
rlabel metal1 27508 7854 27508 7854 0 net54
rlabel metal1 27738 7820 27738 7820 0 net55
rlabel metal1 28014 7888 28014 7888 0 net56
rlabel metal2 19090 8398 19090 8398 0 net57
rlabel metal1 33120 8262 33120 8262 0 net58
rlabel metal1 33580 8262 33580 8262 0 net59
rlabel metal1 33856 1190 33856 1190 0 net6
rlabel metal2 33718 8806 33718 8806 0 net60
rlabel metal2 33994 7871 33994 7871 0 net61
rlabel metal1 33810 7412 33810 7412 0 net62
rlabel metal1 34086 7378 34086 7378 0 net63
rlabel metal1 18998 8976 18998 8976 0 net64
rlabel metal2 18814 6324 18814 6324 0 net65
rlabel metal2 17618 8500 17618 8500 0 net66
rlabel metal2 19182 8500 19182 8500 0 net67
rlabel metal2 19090 9843 19090 9843 0 net68
rlabel metal2 31970 8415 31970 8415 0 net69
rlabel metal1 35282 1258 35282 1258 0 net7
rlabel metal1 32246 8262 32246 8262 0 net70
rlabel metal1 32430 8330 32430 8330 0 net71
rlabel metal2 32890 8942 32890 8942 0 net72
rlabel metal2 1610 1734 1610 1734 0 net73
rlabel metal1 28014 2278 28014 2278 0 net74
rlabel metal1 37214 7922 37214 7922 0 net75
rlabel metal1 36846 7752 36846 7752 0 net76
rlabel metal1 37582 8874 37582 8874 0 net77
rlabel metal1 39652 8466 39652 8466 0 net78
rlabel metal1 38410 7718 38410 7718 0 net79
rlabel metal2 37398 2652 37398 2652 0 net8
rlabel metal1 37812 7310 37812 7310 0 net80
rlabel metal1 38732 7854 38732 7854 0 net81
rlabel metal1 39744 2550 39744 2550 0 net82
rlabel metal1 40526 3706 40526 3706 0 net83
rlabel metal1 40204 7854 40204 7854 0 net84
rlabel metal2 35282 8670 35282 8670 0 net85
rlabel metal2 35466 6256 35466 6256 0 net86
rlabel metal1 35926 8432 35926 8432 0 net87
rlabel metal2 36478 6494 36478 6494 0 net88
rlabel metal1 37398 8568 37398 8568 0 net89
rlabel metal1 39468 1530 39468 1530 0 net9
rlabel metal1 36110 7786 36110 7786 0 net90
rlabel metal1 36754 7820 36754 7820 0 net91
rlabel metal1 37720 8534 37720 8534 0 net92
rlabel metal1 38502 8568 38502 8568 0 net93
rlabel metal2 4922 8789 4922 8789 0 net94
rlabel metal1 5658 7752 5658 7752 0 net95
rlabel metal1 6210 7446 6210 7446 0 net96
rlabel metal1 6555 7854 6555 7854 0 net97
rlabel metal2 5934 6902 5934 6902 0 net98
rlabel via2 6762 7803 6762 7803 0 net99
<< properties >>
string FIXED_BBOX 0 0 45000 10000
<< end >>
