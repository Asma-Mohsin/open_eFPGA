magic
tech sky130A
magscale 1 2
timestamp 1733242052
<< viali >>
rect 2053 43401 2087 43435
rect 2421 43401 2455 43435
rect 2973 43401 3007 43435
rect 3525 43401 3559 43435
rect 4813 43401 4847 43435
rect 5365 43401 5399 43435
rect 5733 43401 5767 43435
rect 6377 43401 6411 43435
rect 7021 43401 7055 43435
rect 7573 43401 7607 43435
rect 8125 43401 8159 43435
rect 8677 43401 8711 43435
rect 9137 43401 9171 43435
rect 9781 43401 9815 43435
rect 10517 43401 10551 43435
rect 16865 43401 16899 43435
rect 17325 43401 17359 43435
rect 17601 43401 17635 43435
rect 18429 43401 18463 43435
rect 20453 43401 20487 43435
rect 21005 43401 21039 43435
rect 22201 43401 22235 43435
rect 22569 43401 22603 43435
rect 23673 43401 23707 43435
rect 2329 43333 2363 43367
rect 6745 43333 6779 43367
rect 11621 43333 11655 43367
rect 12449 43333 12483 43367
rect 12817 43333 12851 43367
rect 13737 43333 13771 43367
rect 14197 43333 14231 43367
rect 14749 43333 14783 43367
rect 15117 43333 15151 43367
rect 15577 43333 15611 43367
rect 15945 43333 15979 43367
rect 16313 43333 16347 43367
rect 16773 43333 16807 43367
rect 23029 43333 23063 43367
rect 1593 43265 1627 43299
rect 1777 43265 1811 43299
rect 2881 43265 2915 43299
rect 3341 43265 3375 43299
rect 3985 43265 4019 43299
rect 4169 43265 4203 43299
rect 4537 43265 4571 43299
rect 4629 43265 4663 43299
rect 5089 43265 5123 43299
rect 5641 43265 5675 43299
rect 6561 43265 6595 43299
rect 7389 43265 7423 43299
rect 7849 43265 7883 43299
rect 8401 43265 8435 43299
rect 8953 43265 8987 43299
rect 9505 43265 9539 43299
rect 9965 43265 9999 43299
rect 10333 43265 10367 43299
rect 10701 43265 10735 43299
rect 11069 43265 11103 43299
rect 12081 43265 12115 43299
rect 16497 43265 16531 43299
rect 17233 43265 17267 43299
rect 17509 43265 17543 43299
rect 17785 43265 17819 43299
rect 18061 43265 18095 43299
rect 18337 43265 18371 43299
rect 18613 43265 18647 43299
rect 18889 43265 18923 43299
rect 19441 43265 19475 43299
rect 19809 43265 19843 43299
rect 20177 43265 20211 43299
rect 20361 43265 20395 43299
rect 20913 43265 20947 43299
rect 21373 43265 21407 43299
rect 21925 43265 21959 43299
rect 22477 43265 22511 43299
rect 23581 43265 23615 43299
rect 24225 43265 24259 43299
rect 1409 43129 1443 43163
rect 11805 43129 11839 43163
rect 12633 43129 12667 43163
rect 14933 43129 14967 43163
rect 15301 43129 15335 43163
rect 16129 43129 16163 43163
rect 17049 43129 17083 43163
rect 18153 43129 18187 43163
rect 24041 43129 24075 43163
rect 3801 43061 3835 43095
rect 10149 43061 10183 43095
rect 10885 43061 10919 43095
rect 11253 43061 11287 43095
rect 12265 43061 12299 43095
rect 12909 43061 12943 43095
rect 13829 43061 13863 43095
rect 14289 43061 14323 43095
rect 15669 43061 15703 43095
rect 17877 43061 17911 43095
rect 18705 43061 18739 43095
rect 19257 43061 19291 43095
rect 21557 43061 21591 43095
rect 23121 43061 23155 43095
rect 3341 42857 3375 42891
rect 4353 42857 4387 42891
rect 6101 42857 6135 42891
rect 6653 42857 6687 42891
rect 7205 42857 7239 42891
rect 8953 42857 8987 42891
rect 12081 42857 12115 42891
rect 16957 42857 16991 42891
rect 23305 42857 23339 42891
rect 4721 42789 4755 42823
rect 10333 42789 10367 42823
rect 18613 42789 18647 42823
rect 21189 42789 21223 42823
rect 2973 42721 3007 42755
rect 5365 42721 5399 42755
rect 8677 42721 8711 42755
rect 22937 42721 22971 42755
rect 24041 42721 24075 42755
rect 3801 42653 3835 42687
rect 4905 42653 4939 42687
rect 5549 42653 5583 42687
rect 7573 42653 7607 42687
rect 8125 42653 8159 42687
rect 9137 42653 9171 42687
rect 10241 42653 10275 42687
rect 10517 42653 10551 42687
rect 10885 42653 10919 42687
rect 10977 42653 11011 42687
rect 11621 42653 11655 42687
rect 11897 42653 11931 42687
rect 12357 42653 12391 42687
rect 13001 42653 13035 42687
rect 14105 42653 14139 42687
rect 14381 42653 14415 42687
rect 14657 42653 14691 42687
rect 15117 42653 15151 42687
rect 15393 42653 15427 42687
rect 16589 42653 16623 42687
rect 17141 42653 17175 42687
rect 17417 42653 17451 42687
rect 17693 42653 17727 42687
rect 17969 42653 18003 42687
rect 18245 42653 18279 42687
rect 18521 42653 18555 42687
rect 18797 42653 18831 42687
rect 19073 42653 19107 42687
rect 21373 42653 21407 42687
rect 22109 42653 22143 42687
rect 22477 42653 22511 42687
rect 1409 42585 1443 42619
rect 2145 42585 2179 42619
rect 2697 42585 2731 42619
rect 3249 42585 3283 42619
rect 4261 42585 4295 42619
rect 5089 42585 5123 42619
rect 6009 42585 6043 42619
rect 6561 42585 6595 42619
rect 7113 42585 7147 42619
rect 8401 42585 8435 42619
rect 9505 42585 9539 42619
rect 19257 42585 19291 42619
rect 21005 42585 21039 42619
rect 21557 42585 21591 42619
rect 21925 42585 21959 42619
rect 22661 42585 22695 42619
rect 23213 42585 23247 42619
rect 23765 42585 23799 42619
rect 3985 42517 4019 42551
rect 5733 42517 5767 42551
rect 7757 42517 7791 42551
rect 7941 42517 7975 42551
rect 9781 42517 9815 42551
rect 10057 42517 10091 42551
rect 10701 42517 10735 42551
rect 11161 42517 11195 42551
rect 11805 42517 11839 42551
rect 12541 42517 12575 42551
rect 13185 42517 13219 42551
rect 14289 42517 14323 42551
rect 14565 42517 14599 42551
rect 14841 42517 14875 42551
rect 15301 42517 15335 42551
rect 15577 42517 15611 42551
rect 16773 42517 16807 42551
rect 17233 42517 17267 42551
rect 17509 42517 17543 42551
rect 17785 42517 17819 42551
rect 18061 42517 18095 42551
rect 18337 42517 18371 42551
rect 18889 42517 18923 42551
rect 2605 42313 2639 42347
rect 3157 42313 3191 42347
rect 6469 42313 6503 42347
rect 7573 42313 7607 42347
rect 8493 42313 8527 42347
rect 19625 42313 19659 42347
rect 20545 42313 20579 42347
rect 20821 42313 20855 42347
rect 22753 42313 22787 42347
rect 23305 42313 23339 42347
rect 4721 42245 4755 42279
rect 16773 42245 16807 42279
rect 17141 42245 17175 42279
rect 17509 42245 17543 42279
rect 17877 42245 17911 42279
rect 18245 42245 18279 42279
rect 18981 42245 19015 42279
rect 19349 42245 19383 42279
rect 22293 42245 22327 42279
rect 1409 42177 1443 42211
rect 2513 42177 2547 42211
rect 3065 42177 3099 42211
rect 3617 42177 3651 42211
rect 4169 42177 4203 42211
rect 5457 42177 5491 42211
rect 5917 42177 5951 42211
rect 6193 42177 6227 42211
rect 6653 42177 6687 42211
rect 6929 42177 6963 42211
rect 7389 42177 7423 42211
rect 7941 42177 7975 42211
rect 8217 42177 8251 42211
rect 8401 42177 8435 42211
rect 9287 42187 9321 42221
rect 16221 42177 16255 42211
rect 16497 42177 16531 42211
rect 18613 42177 18647 42211
rect 19809 42177 19843 42211
rect 20177 42177 20211 42211
rect 20453 42177 20487 42211
rect 20729 42177 20763 42211
rect 21005 42177 21039 42211
rect 21281 42177 21315 42211
rect 21925 42177 21959 42211
rect 22477 42177 22511 42211
rect 23029 42177 23063 42211
rect 23581 42177 23615 42211
rect 23949 42177 23983 42211
rect 24133 42177 24167 42211
rect 24501 42177 24535 42211
rect 2237 42109 2271 42143
rect 9045 42109 9079 42143
rect 4353 42041 4387 42075
rect 7757 42041 7791 42075
rect 16037 42041 16071 42075
rect 16957 42041 16991 42075
rect 17325 42041 17359 42075
rect 18429 42041 18463 42075
rect 19993 42041 20027 42075
rect 20269 42041 20303 42075
rect 21557 42041 21591 42075
rect 3709 41973 3743 42007
rect 4813 41973 4847 42007
rect 5733 41973 5767 42007
rect 6009 41973 6043 42007
rect 6745 41973 6779 42007
rect 7297 41973 7331 42007
rect 8033 41973 8067 42007
rect 10057 41973 10091 42007
rect 16313 41973 16347 42007
rect 17601 41973 17635 42007
rect 17969 41973 18003 42007
rect 18705 41973 18739 42007
rect 19073 41973 19107 42007
rect 19441 41973 19475 42007
rect 3433 41769 3467 41803
rect 4537 41769 4571 41803
rect 4997 41769 5031 41803
rect 5457 41769 5491 41803
rect 5825 41769 5859 41803
rect 6193 41769 6227 41803
rect 6561 41769 6595 41803
rect 6837 41769 6871 41803
rect 7297 41769 7331 41803
rect 7757 41769 7791 41803
rect 8401 41769 8435 41803
rect 8953 41769 8987 41803
rect 18889 41769 18923 41803
rect 19809 41769 19843 41803
rect 20085 41769 20119 41803
rect 21281 41769 21315 41803
rect 21741 41769 21775 41803
rect 22293 41769 22327 41803
rect 23581 41769 23615 41803
rect 23949 41769 23983 41803
rect 4721 41701 4755 41735
rect 18613 41701 18647 41735
rect 20729 41701 20763 41735
rect 21833 41701 21867 41735
rect 23029 41701 23063 41735
rect 2237 41633 2271 41667
rect 3249 41633 3283 41667
rect 3617 41565 3651 41599
rect 3893 41565 3927 41599
rect 4353 41565 4387 41599
rect 4905 41565 4939 41599
rect 5181 41565 5215 41599
rect 5641 41565 5675 41599
rect 6009 41565 6043 41599
rect 6377 41565 6411 41599
rect 6745 41565 6779 41599
rect 7021 41565 7055 41599
rect 7481 41565 7515 41599
rect 7941 41565 7975 41599
rect 8309 41565 8343 41599
rect 8577 41565 8611 41599
rect 9137 41565 9171 41599
rect 9781 41565 9815 41599
rect 10039 41535 10073 41569
rect 16129 41565 16163 41599
rect 16497 41565 16531 41599
rect 18521 41565 18555 41599
rect 18797 41565 18831 41599
rect 19073 41565 19107 41599
rect 19441 41565 19475 41599
rect 19717 41565 19751 41599
rect 19993 41565 20027 41599
rect 20269 41565 20303 41599
rect 20545 41565 20579 41599
rect 20913 41565 20947 41599
rect 21189 41565 21223 41599
rect 21465 41565 21499 41599
rect 21557 41565 21591 41599
rect 22017 41565 22051 41599
rect 1409 41497 1443 41531
rect 2421 41497 2455 41531
rect 22201 41497 22235 41531
rect 22753 41497 22787 41531
rect 23305 41497 23339 41531
rect 23857 41497 23891 41531
rect 3985 41429 4019 41463
rect 8125 41429 8159 41463
rect 9413 41429 9447 41463
rect 10793 41429 10827 41463
rect 16221 41429 16255 41463
rect 16589 41429 16623 41463
rect 18337 41429 18371 41463
rect 19257 41429 19291 41463
rect 19533 41429 19567 41463
rect 20361 41429 20395 41463
rect 21005 41429 21039 41463
rect 4721 41225 4755 41259
rect 5273 41225 5307 41259
rect 5549 41225 5583 41259
rect 5825 41225 5859 41259
rect 6377 41225 6411 41259
rect 6929 41225 6963 41259
rect 9505 41225 9539 41259
rect 18613 41225 18647 41259
rect 20453 41225 20487 41259
rect 21189 41225 21223 41259
rect 21833 41225 21867 41259
rect 22109 41225 22143 41259
rect 22477 41225 22511 41259
rect 23121 41225 23155 41259
rect 24225 41225 24259 41259
rect 1869 41157 1903 41191
rect 18981 41157 19015 41191
rect 22845 41157 22879 41191
rect 1501 41089 1535 41123
rect 2237 41089 2271 41123
rect 2329 41089 2363 41123
rect 3065 41089 3099 41123
rect 3615 41089 3649 41123
rect 4905 41089 4939 41123
rect 5181 41089 5215 41123
rect 5457 41089 5491 41123
rect 5733 41089 5767 41123
rect 6009 41089 6043 41123
rect 6561 41089 6595 41123
rect 6837 41089 6871 41123
rect 7113 41089 7147 41123
rect 7941 41089 7975 41123
rect 8217 41089 8251 41123
rect 9689 41089 9723 41123
rect 10057 41089 10091 41123
rect 10331 41089 10365 41123
rect 18797 41089 18831 41123
rect 19625 41089 19659 41123
rect 20085 41089 20119 41123
rect 20361 41089 20395 41123
rect 20637 41089 20671 41123
rect 21005 41089 21039 41123
rect 21373 41089 21407 41123
rect 21649 41089 21683 41123
rect 22017 41089 22051 41123
rect 22293 41089 22327 41123
rect 22661 41089 22695 41123
rect 23397 41089 23431 41123
rect 23949 41089 23983 41123
rect 3341 41021 3375 41055
rect 1685 40953 1719 40987
rect 4353 40953 4387 40987
rect 4997 40953 5031 40987
rect 6653 40953 6687 40987
rect 7757 40953 7791 40987
rect 11713 40953 11747 40987
rect 19165 40953 19199 40987
rect 19901 40953 19935 40987
rect 8033 40885 8067 40919
rect 11069 40885 11103 40919
rect 19441 40885 19475 40919
rect 20177 40885 20211 40919
rect 20821 40885 20855 40919
rect 21465 40885 21499 40919
rect 23673 40885 23707 40919
rect 3801 40681 3835 40715
rect 4077 40681 4111 40715
rect 20453 40681 20487 40715
rect 20729 40681 20763 40715
rect 22109 40681 22143 40715
rect 22569 40681 22603 40715
rect 22937 40681 22971 40715
rect 23581 40681 23615 40715
rect 10517 40613 10551 40647
rect 19625 40613 19659 40647
rect 21005 40613 21039 40647
rect 21281 40613 21315 40647
rect 21557 40613 21591 40647
rect 1409 40545 1443 40579
rect 10057 40545 10091 40579
rect 10793 40545 10827 40579
rect 11069 40545 11103 40579
rect 1685 40477 1719 40511
rect 2329 40477 2363 40511
rect 2603 40477 2637 40511
rect 3985 40477 4019 40511
rect 4261 40477 4295 40511
rect 4353 40477 4387 40511
rect 4627 40477 4661 40511
rect 5733 40477 5767 40511
rect 6007 40477 6041 40511
rect 7481 40477 7515 40511
rect 7755 40477 7789 40511
rect 9873 40477 9907 40511
rect 10910 40477 10944 40511
rect 19349 40477 19383 40511
rect 19809 40477 19843 40511
rect 20085 40477 20119 40511
rect 20361 40477 20395 40511
rect 20637 40477 20671 40511
rect 20913 40477 20947 40511
rect 21189 40477 21223 40511
rect 21465 40477 21499 40511
rect 21741 40477 21775 40511
rect 22017 40477 22051 40511
rect 22293 40477 22327 40511
rect 22753 40477 22787 40511
rect 23121 40477 23155 40511
rect 23305 40409 23339 40443
rect 23857 40409 23891 40443
rect 24225 40409 24259 40443
rect 3341 40341 3375 40375
rect 5365 40341 5399 40375
rect 6745 40341 6779 40375
rect 8493 40341 8527 40375
rect 11713 40341 11747 40375
rect 19441 40341 19475 40375
rect 19901 40341 19935 40375
rect 20177 40341 20211 40375
rect 21833 40341 21867 40375
rect 2789 40137 2823 40171
rect 4353 40137 4387 40171
rect 19993 40137 20027 40171
rect 20269 40137 20303 40171
rect 20545 40137 20579 40171
rect 21465 40137 21499 40171
rect 22109 40137 22143 40171
rect 22385 40137 22419 40171
rect 22845 40137 22879 40171
rect 23397 40137 23431 40171
rect 23765 40137 23799 40171
rect 3249 40069 3283 40103
rect 3617 40069 3651 40103
rect 8677 40069 8711 40103
rect 9045 40069 9079 40103
rect 1683 40001 1717 40035
rect 2973 40001 3007 40035
rect 3525 40001 3559 40035
rect 3985 40001 4019 40035
rect 5147 40001 5181 40035
rect 6835 40001 6869 40035
rect 8953 40001 8987 40035
rect 9413 40001 9447 40035
rect 9795 40001 9829 40035
rect 20177 40001 20211 40035
rect 20453 40001 20487 40035
rect 20729 40001 20763 40035
rect 21097 40001 21131 40035
rect 21373 40001 21407 40035
rect 21649 40001 21683 40035
rect 22017 40001 22051 40035
rect 22293 40001 22327 40035
rect 22569 40001 22603 40035
rect 23029 40001 23063 40035
rect 23305 40001 23339 40035
rect 23581 40001 23615 40035
rect 23949 40001 23983 40035
rect 24133 40001 24167 40035
rect 1409 39933 1443 39967
rect 4905 39933 4939 39967
rect 6561 39933 6595 39967
rect 20913 39865 20947 39899
rect 21189 39865 21223 39899
rect 23121 39865 23155 39899
rect 2421 39797 2455 39831
rect 4537 39797 4571 39831
rect 5917 39797 5951 39831
rect 7573 39797 7607 39831
rect 9965 39797 9999 39831
rect 21833 39797 21867 39831
rect 24409 39797 24443 39831
rect 3801 39593 3835 39627
rect 7941 39593 7975 39627
rect 21097 39593 21131 39627
rect 21649 39593 21683 39627
rect 21925 39593 21959 39627
rect 22477 39593 22511 39627
rect 22753 39593 22787 39627
rect 3433 39525 3467 39559
rect 4813 39525 4847 39559
rect 6745 39525 6779 39559
rect 20821 39525 20855 39559
rect 21373 39525 21407 39559
rect 22201 39525 22235 39559
rect 23489 39525 23523 39559
rect 2053 39457 2087 39491
rect 4169 39457 4203 39491
rect 5089 39457 5123 39491
rect 5365 39457 5399 39491
rect 6101 39457 6135 39491
rect 7297 39457 7331 39491
rect 9229 39457 9263 39491
rect 12265 39457 12299 39491
rect 1409 39389 1443 39423
rect 2295 39389 2329 39423
rect 3617 39389 3651 39423
rect 3985 39389 4019 39423
rect 4353 39389 4387 39423
rect 5206 39389 5240 39423
rect 6285 39389 6319 39423
rect 7021 39389 7055 39423
rect 7159 39389 7193 39423
rect 9503 39389 9537 39423
rect 10885 39389 10919 39423
rect 11159 39389 11193 39423
rect 12507 39389 12541 39423
rect 21005 39389 21039 39423
rect 21281 39389 21315 39423
rect 21557 39389 21591 39423
rect 21833 39389 21867 39423
rect 22109 39389 22143 39423
rect 22385 39389 22419 39423
rect 22661 39389 22695 39423
rect 22937 39389 22971 39423
rect 23213 39389 23247 39423
rect 23673 39389 23707 39423
rect 23949 39389 23983 39423
rect 1685 39321 1719 39355
rect 3065 39253 3099 39287
rect 6009 39253 6043 39287
rect 10241 39253 10275 39287
rect 11897 39253 11931 39287
rect 13277 39253 13311 39287
rect 23029 39253 23063 39287
rect 24133 39253 24167 39287
rect 3157 39049 3191 39083
rect 13369 39049 13403 39083
rect 20177 39049 20211 39083
rect 20453 39049 20487 39083
rect 21097 39049 21131 39083
rect 22293 39049 22327 39083
rect 22937 39049 22971 39083
rect 23213 39049 23247 39083
rect 23765 39049 23799 39083
rect 3525 38981 3559 39015
rect 4261 38981 4295 39015
rect 8585 38981 8619 39015
rect 1409 38913 1443 38947
rect 2421 38913 2455 38947
rect 3433 38913 3467 38947
rect 3893 38913 3927 38947
rect 7021 38913 7055 38947
rect 7295 38913 7329 38947
rect 8861 38913 8895 38947
rect 8953 38913 8987 38947
rect 9321 38913 9355 38947
rect 9703 38913 9737 38947
rect 10057 38913 10091 38947
rect 10331 38913 10365 38947
rect 12449 38913 12483 38947
rect 12725 38913 12759 38947
rect 19441 38913 19475 38947
rect 20361 38913 20395 38947
rect 20637 38913 20671 38947
rect 21281 38913 21315 38947
rect 21833 38913 21867 38947
rect 22477 38913 22511 38947
rect 22569 38913 22603 38947
rect 22761 38919 22795 38953
rect 23121 38913 23155 38947
rect 23397 38913 23431 38947
rect 23673 38913 23707 38947
rect 23949 38913 23983 38947
rect 24133 38913 24167 38947
rect 2237 38845 2271 38879
rect 2605 38845 2639 38879
rect 11529 38845 11563 38879
rect 11713 38845 11747 38879
rect 12566 38845 12600 38879
rect 8033 38777 8067 38811
rect 9873 38777 9907 38811
rect 11069 38777 11103 38811
rect 12173 38777 12207 38811
rect 19257 38777 19291 38811
rect 23489 38777 23523 38811
rect 4445 38709 4479 38743
rect 13645 38709 13679 38743
rect 21925 38709 21959 38743
rect 22661 38709 22695 38743
rect 24409 38709 24443 38743
rect 4813 38505 4847 38539
rect 18705 38505 18739 38539
rect 22017 38505 22051 38539
rect 23489 38505 23523 38539
rect 12725 38437 12759 38471
rect 2237 38369 2271 38403
rect 3157 38369 3191 38403
rect 12265 38369 12299 38403
rect 13001 38369 13035 38403
rect 20637 38369 20671 38403
rect 1409 38301 1443 38335
rect 2421 38301 2455 38335
rect 2973 38301 3007 38335
rect 3801 38301 3835 38335
rect 4075 38301 4109 38335
rect 7481 38301 7515 38335
rect 7739 38271 7773 38305
rect 10241 38301 10275 38335
rect 10499 38271 10533 38305
rect 12081 38301 12115 38335
rect 13118 38301 13152 38335
rect 13277 38301 13311 38335
rect 18889 38301 18923 38335
rect 19625 38301 19659 38335
rect 22109 38301 22143 38335
rect 22351 38301 22385 38335
rect 23673 38301 23707 38335
rect 23949 38301 23983 38335
rect 2697 38233 2731 38267
rect 13921 38233 13955 38267
rect 20882 38233 20916 38267
rect 8493 38165 8527 38199
rect 11253 38165 11287 38199
rect 19441 38165 19475 38199
rect 23121 38165 23155 38199
rect 24133 38165 24167 38199
rect 13737 37961 13771 37995
rect 18153 37961 18187 37995
rect 20913 37961 20947 37995
rect 21925 37961 21959 37995
rect 23397 37961 23431 37995
rect 8493 37893 8527 37927
rect 8769 37893 8803 37927
rect 8861 37893 8895 37927
rect 9597 37893 9631 37927
rect 22845 37893 22879 37927
rect 2605 37825 2639 37859
rect 3341 37825 3375 37859
rect 3893 37825 3927 37859
rect 4871 37825 4905 37859
rect 7389 37825 7423 37859
rect 7573 37825 7607 37859
rect 9229 37825 9263 37859
rect 12967 37825 13001 37859
rect 18337 37825 18371 37859
rect 21097 37825 21131 37859
rect 22109 37825 22143 37859
rect 22477 37825 22511 37859
rect 23121 37825 23155 37859
rect 23581 37825 23615 37859
rect 23857 37825 23891 37859
rect 24133 37825 24167 37859
rect 1409 37757 1443 37791
rect 1593 37757 1627 37791
rect 2329 37757 2363 37791
rect 2467 37757 2501 37791
rect 3525 37757 3559 37791
rect 4169 37757 4203 37791
rect 4629 37757 4663 37791
rect 12725 37757 12759 37791
rect 22293 37757 22327 37791
rect 2053 37689 2087 37723
rect 22937 37689 22971 37723
rect 3249 37621 3283 37655
rect 5641 37621 5675 37655
rect 7481 37621 7515 37655
rect 9781 37621 9815 37655
rect 22753 37621 22787 37655
rect 23673 37621 23707 37655
rect 24409 37621 24443 37655
rect 2421 37417 2455 37451
rect 7573 37417 7607 37451
rect 9965 37417 9999 37451
rect 22477 37417 22511 37451
rect 23121 37417 23155 37451
rect 23673 37417 23707 37451
rect 5089 37281 5123 37315
rect 8217 37281 8251 37315
rect 1409 37213 1443 37247
rect 1683 37213 1717 37247
rect 2789 37213 2823 37247
rect 3801 37213 3835 37247
rect 4353 37213 4387 37247
rect 5363 37213 5397 37247
rect 6561 37213 6595 37247
rect 6835 37203 6869 37237
rect 7941 37213 7975 37247
rect 8033 37213 8067 37247
rect 8953 37213 8987 37247
rect 9227 37203 9261 37237
rect 19441 37213 19475 37247
rect 19993 37213 20027 37247
rect 20361 37213 20395 37247
rect 21925 37213 21959 37247
rect 22661 37213 22695 37247
rect 23397 37213 23431 37247
rect 23857 37213 23891 37247
rect 23949 37213 23983 37247
rect 3065 37145 3099 37179
rect 4077 37145 4111 37179
rect 4629 37145 4663 37179
rect 8217 37145 8251 37179
rect 6101 37077 6135 37111
rect 19257 37077 19291 37111
rect 19809 37077 19843 37111
rect 20177 37077 20211 37111
rect 21741 37077 21775 37111
rect 23213 37077 23247 37111
rect 24133 37077 24167 37111
rect 3157 36873 3191 36907
rect 5641 36873 5675 36907
rect 7481 36873 7515 36907
rect 18613 36873 18647 36907
rect 19533 36873 19567 36907
rect 22385 36873 22419 36907
rect 23397 36873 23431 36907
rect 23673 36873 23707 36907
rect 3525 36805 3559 36839
rect 4261 36805 4295 36839
rect 7297 36805 7331 36839
rect 24133 36805 24167 36839
rect 1409 36737 1443 36771
rect 1961 36737 1995 36771
rect 3433 36737 3467 36771
rect 3893 36737 3927 36771
rect 4903 36737 4937 36771
rect 7205 36737 7239 36771
rect 7665 36737 7699 36771
rect 9873 36737 9907 36771
rect 10147 36737 10181 36771
rect 18797 36737 18831 36771
rect 19717 36737 19751 36771
rect 22569 36737 22603 36771
rect 23581 36737 23615 36771
rect 23857 36737 23891 36771
rect 1685 36669 1719 36703
rect 2145 36669 2179 36703
rect 4629 36669 4663 36703
rect 2697 36601 2731 36635
rect 4445 36533 4479 36567
rect 10885 36533 10919 36567
rect 23029 36533 23063 36567
rect 24409 36533 24443 36567
rect 3341 36329 3375 36363
rect 6929 36329 6963 36363
rect 21557 36329 21591 36363
rect 22845 36329 22879 36363
rect 5641 36261 5675 36295
rect 6837 36261 6871 36295
rect 22569 36261 22603 36295
rect 23213 36261 23247 36295
rect 2329 36193 2363 36227
rect 5181 36193 5215 36227
rect 6034 36193 6068 36227
rect 6193 36193 6227 36227
rect 10793 36193 10827 36227
rect 1409 36125 1443 36159
rect 2571 36125 2605 36159
rect 3801 36125 3835 36159
rect 4353 36125 4387 36159
rect 4997 36125 5031 36159
rect 5917 36125 5951 36159
rect 7113 36125 7147 36159
rect 9413 36125 9447 36159
rect 9687 36125 9721 36159
rect 11035 36125 11069 36159
rect 12265 36125 12299 36159
rect 12539 36125 12573 36159
rect 18337 36125 18371 36159
rect 18705 36125 18739 36159
rect 18797 36125 18831 36159
rect 19441 36125 19475 36159
rect 20269 36125 20303 36159
rect 21741 36125 21775 36159
rect 22753 36125 22787 36159
rect 23029 36125 23063 36159
rect 23397 36125 23431 36159
rect 23673 36125 23707 36159
rect 23857 36125 23891 36159
rect 1685 36057 1719 36091
rect 4077 36057 4111 36091
rect 4629 36057 4663 36091
rect 10425 35989 10459 36023
rect 11805 35989 11839 36023
rect 13277 35989 13311 36023
rect 18153 35989 18187 36023
rect 19257 35989 19291 36023
rect 20085 35989 20119 36023
rect 23489 35989 23523 36023
rect 24133 35989 24167 36023
rect 6193 35785 6227 35819
rect 11805 35785 11839 35819
rect 19073 35785 19107 35819
rect 21005 35785 21039 35819
rect 22661 35785 22695 35819
rect 22937 35785 22971 35819
rect 23305 35785 23339 35819
rect 23581 35785 23615 35819
rect 8033 35717 8067 35751
rect 8309 35717 8343 35751
rect 9137 35717 9171 35751
rect 12541 35717 12575 35751
rect 12909 35717 12943 35751
rect 19870 35717 19904 35751
rect 21373 35717 21407 35751
rect 1409 35649 1443 35683
rect 2695 35649 2729 35683
rect 3801 35649 3835 35683
rect 8401 35649 8435 35683
rect 8769 35649 8803 35683
rect 9689 35649 9723 35683
rect 10425 35649 10459 35683
rect 10542 35649 10576 35683
rect 11345 35649 11379 35683
rect 12081 35649 12115 35683
rect 12173 35649 12207 35683
rect 14363 35679 14397 35713
rect 17960 35649 17994 35683
rect 19165 35649 19199 35683
rect 19257 35649 19291 35683
rect 19625 35649 19659 35683
rect 21097 35649 21131 35683
rect 21465 35649 21499 35683
rect 22009 35653 22043 35687
rect 22109 35649 22143 35683
rect 22293 35649 22327 35683
rect 22569 35649 22603 35683
rect 22845 35649 22879 35683
rect 23121 35649 23155 35683
rect 23489 35649 23523 35683
rect 23765 35649 23799 35683
rect 24133 35649 24167 35683
rect 1685 35581 1719 35615
rect 2421 35581 2455 35615
rect 3985 35581 4019 35615
rect 4353 35581 4387 35615
rect 4537 35581 4571 35615
rect 5273 35581 5307 35615
rect 5390 35581 5424 35615
rect 5549 35581 5583 35615
rect 9505 35581 9539 35615
rect 10711 35581 10745 35615
rect 14105 35581 14139 35615
rect 17693 35581 17727 35615
rect 19441 35581 19475 35615
rect 21373 35581 21407 35615
rect 22201 35581 22235 35615
rect 4997 35513 5031 35547
rect 10149 35513 10183 35547
rect 21189 35513 21223 35547
rect 21557 35513 21591 35547
rect 21833 35513 21867 35547
rect 22385 35513 22419 35547
rect 3433 35445 3467 35479
rect 9321 35445 9355 35479
rect 13093 35445 13127 35479
rect 15117 35445 15151 35479
rect 19349 35445 19383 35479
rect 24409 35445 24443 35479
rect 3433 35241 3467 35275
rect 8309 35241 8343 35275
rect 13093 35241 13127 35275
rect 19349 35241 19383 35275
rect 21281 35241 21315 35275
rect 23213 35241 23247 35275
rect 10793 35173 10827 35207
rect 18797 35173 18831 35207
rect 22201 35173 22235 35207
rect 1593 35105 1627 35139
rect 2237 35105 2271 35139
rect 2513 35105 2547 35139
rect 2651 35105 2685 35139
rect 5733 35105 5767 35139
rect 7297 35105 7331 35139
rect 10333 35105 10367 35139
rect 12081 35105 12115 35139
rect 1777 35037 1811 35071
rect 2789 35037 2823 35071
rect 4261 35037 4295 35071
rect 6007 35037 6041 35071
rect 7571 35037 7605 35071
rect 10149 35037 10183 35071
rect 11069 35037 11103 35071
rect 11186 35037 11220 35071
rect 11345 35037 11379 35071
rect 12355 35037 12389 35071
rect 17785 35037 17819 35071
rect 18059 35037 18093 35071
rect 19257 35037 19291 35071
rect 19441 35037 19475 35071
rect 20269 35037 20303 35071
rect 20543 35037 20577 35071
rect 22385 35037 22419 35071
rect 23397 35037 23431 35071
rect 23673 35037 23707 35071
rect 4353 34969 4387 35003
rect 4721 34969 4755 35003
rect 23857 34969 23891 35003
rect 24225 34969 24259 35003
rect 3985 34901 4019 34935
rect 5089 34901 5123 34935
rect 5273 34901 5307 34935
rect 6745 34901 6779 34935
rect 11989 34901 12023 34935
rect 23489 34901 23523 34935
rect 2513 34697 2547 34731
rect 4261 34697 4295 34731
rect 7389 34697 7423 34731
rect 9045 34697 9079 34731
rect 17693 34697 17727 34731
rect 20637 34697 20671 34731
rect 21465 34697 21499 34731
rect 21833 34697 21867 34731
rect 22753 34697 22787 34731
rect 23305 34697 23339 34731
rect 23673 34697 23707 34731
rect 4813 34629 4847 34663
rect 5089 34629 5123 34663
rect 5181 34629 5215 34663
rect 5917 34629 5951 34663
rect 24133 34629 24167 34663
rect 1775 34561 1809 34595
rect 3523 34561 3557 34595
rect 5549 34561 5583 34595
rect 6377 34561 6411 34595
rect 6635 34591 6669 34625
rect 8275 34561 8309 34595
rect 14363 34591 14397 34625
rect 16221 34561 16255 34595
rect 16681 34561 16715 34595
rect 16955 34571 16989 34605
rect 20821 34561 20855 34595
rect 21649 34561 21683 34595
rect 22017 34561 22051 34595
rect 22661 34561 22695 34595
rect 22937 34561 22971 34595
rect 23213 34561 23247 34595
rect 23489 34561 23523 34595
rect 23857 34561 23891 34595
rect 1501 34493 1535 34527
rect 3249 34493 3283 34527
rect 8033 34493 8067 34527
rect 14105 34493 14139 34527
rect 16497 34493 16531 34527
rect 24409 34493 24443 34527
rect 22477 34425 22511 34459
rect 23029 34425 23063 34459
rect 6101 34357 6135 34391
rect 15117 34357 15151 34391
rect 16313 34357 16347 34391
rect 16405 34357 16439 34391
rect 2421 34153 2455 34187
rect 10333 34153 10367 34187
rect 17233 34153 17267 34187
rect 17509 34153 17543 34187
rect 23857 34153 23891 34187
rect 9413 34085 9447 34119
rect 21465 34085 21499 34119
rect 22477 34085 22511 34119
rect 3065 34017 3099 34051
rect 4629 34017 4663 34051
rect 7021 34017 7055 34051
rect 9321 34017 9355 34051
rect 9505 34017 9539 34051
rect 10057 34017 10091 34051
rect 12173 34017 12207 34051
rect 14105 34017 14139 34051
rect 15485 34017 15519 34051
rect 1409 33949 1443 33983
rect 1683 33949 1717 33983
rect 2789 33949 2823 33983
rect 3801 33949 3835 33983
rect 4353 33949 4387 33983
rect 5549 33949 5583 33983
rect 5823 33949 5857 33983
rect 7295 33939 7329 33973
rect 9229 33949 9263 33983
rect 9781 33949 9815 33983
rect 9965 33949 9999 33983
rect 10149 33949 10183 33983
rect 10241 33949 10275 33983
rect 12447 33949 12481 33983
rect 14379 33949 14413 33983
rect 15727 33949 15761 33983
rect 17141 33949 17175 33983
rect 17407 33949 17441 33983
rect 17601 33949 17635 33983
rect 21649 33949 21683 33983
rect 22385 33949 22419 33983
rect 22661 33949 22695 33983
rect 23213 33949 23247 33983
rect 23581 33949 23615 33983
rect 23673 33949 23707 33983
rect 23949 33949 23983 33983
rect 4077 33881 4111 33915
rect 6561 33813 6595 33847
rect 8033 33813 8067 33847
rect 9597 33813 9631 33847
rect 13185 33813 13219 33847
rect 15117 33813 15151 33847
rect 16497 33813 16531 33847
rect 22201 33813 22235 33847
rect 23029 33813 23063 33847
rect 23397 33813 23431 33847
rect 24133 33813 24167 33847
rect 9413 33609 9447 33643
rect 10517 33609 10551 33643
rect 15761 33609 15795 33643
rect 17141 33609 17175 33643
rect 19717 33609 19751 33643
rect 22753 33609 22787 33643
rect 23029 33609 23063 33643
rect 23765 33609 23799 33643
rect 2789 33541 2823 33575
rect 24133 33541 24167 33575
rect 1409 33473 1443 33507
rect 1685 33473 1719 33507
rect 1961 33473 1995 33507
rect 2513 33473 2547 33507
rect 3399 33473 3433 33507
rect 7573 33473 7607 33507
rect 8631 33473 8665 33507
rect 8769 33473 8803 33507
rect 9763 33473 9797 33507
rect 11805 33473 11839 33507
rect 15117 33473 15151 33507
rect 17325 33473 17359 33507
rect 18337 33473 18371 33507
rect 18705 33473 18739 33507
rect 19073 33473 19107 33507
rect 19441 33473 19475 33507
rect 19625 33473 19659 33507
rect 19901 33473 19935 33507
rect 20177 33473 20211 33507
rect 22293 33473 22327 33507
rect 22937 33473 22971 33507
rect 23213 33473 23247 33507
rect 23581 33473 23615 33507
rect 23949 33473 23983 33507
rect 2237 33405 2271 33439
rect 3157 33405 3191 33439
rect 7757 33405 7791 33439
rect 8217 33405 8251 33439
rect 8493 33405 8527 33439
rect 9505 33405 9539 33439
rect 11621 33405 11655 33439
rect 12541 33405 12575 33439
rect 12658 33405 12692 33439
rect 12817 33405 12851 33439
rect 13921 33405 13955 33439
rect 14105 33405 14139 33439
rect 14565 33405 14599 33439
rect 14841 33405 14875 33439
rect 14958 33405 14992 33439
rect 19349 33405 19383 33439
rect 19533 33405 19567 33439
rect 12265 33337 12299 33371
rect 18153 33337 18187 33371
rect 4169 33269 4203 33303
rect 4721 33269 4755 33303
rect 13461 33269 13495 33303
rect 18797 33269 18831 33303
rect 19165 33269 19199 33303
rect 19257 33269 19291 33303
rect 20269 33269 20303 33303
rect 22109 33269 22143 33303
rect 23397 33269 23431 33303
rect 24409 33269 24443 33303
rect 9321 33065 9355 33099
rect 12265 33065 12299 33099
rect 17325 33065 17359 33099
rect 20821 33065 20855 33099
rect 23029 33065 23063 33099
rect 16037 32997 16071 33031
rect 20637 32997 20671 33031
rect 21373 32997 21407 33031
rect 22661 32997 22695 33031
rect 9781 32929 9815 32963
rect 11253 32929 11287 32963
rect 12633 32929 12667 32963
rect 16430 32929 16464 32963
rect 16589 32929 16623 32963
rect 21005 32929 21039 32963
rect 21189 32929 21223 32963
rect 1409 32861 1443 32895
rect 1683 32861 1717 32895
rect 2789 32861 2823 32895
rect 3617 32861 3651 32895
rect 4261 32861 4295 32895
rect 4353 32861 4387 32895
rect 9505 32861 9539 32895
rect 10055 32861 10089 32895
rect 11527 32861 11561 32895
rect 12907 32861 12941 32895
rect 15393 32861 15427 32895
rect 15577 32861 15611 32895
rect 16313 32861 16347 32895
rect 17233 32861 17267 32895
rect 17509 32861 17543 32895
rect 17693 32861 17727 32895
rect 19257 32861 19291 32895
rect 20729 32861 20763 32895
rect 21097 32861 21131 32895
rect 21281 32861 21315 32895
rect 21557 32861 21591 32895
rect 22017 32861 22051 32895
rect 22845 32861 22879 32895
rect 23213 32861 23247 32895
rect 23489 32861 23523 32895
rect 23765 32861 23799 32895
rect 23949 32861 23983 32895
rect 3065 32793 3099 32827
rect 4721 32793 4755 32827
rect 5733 32793 5767 32827
rect 6469 32793 6503 32827
rect 6561 32793 6595 32827
rect 6929 32793 6963 32827
rect 7297 32793 7331 32827
rect 17938 32793 17972 32827
rect 19524 32793 19558 32827
rect 2421 32725 2455 32759
rect 3433 32725 3467 32759
rect 3985 32725 4019 32759
rect 5089 32725 5123 32759
rect 5273 32725 5307 32759
rect 6193 32725 6227 32759
rect 7481 32725 7515 32759
rect 10793 32725 10827 32759
rect 13645 32725 13679 32759
rect 19073 32725 19107 32759
rect 21005 32725 21039 32759
rect 21833 32725 21867 32759
rect 23305 32725 23339 32759
rect 23581 32725 23615 32759
rect 24133 32725 24167 32759
rect 3249 32521 3283 32555
rect 4813 32521 4847 32555
rect 9413 32521 9447 32555
rect 19073 32521 19107 32555
rect 19441 32521 19475 32555
rect 20729 32521 20763 32555
rect 23213 32521 23247 32555
rect 11713 32453 11747 32487
rect 14105 32453 14139 32487
rect 14473 32453 14507 32487
rect 14841 32453 14875 32487
rect 15209 32453 15243 32487
rect 22078 32453 22112 32487
rect 24133 32453 24167 32487
rect 2329 32385 2363 32419
rect 3801 32385 3835 32419
rect 4075 32385 4109 32419
rect 8769 32385 8803 32419
rect 10057 32385 10091 32419
rect 10331 32385 10365 32419
rect 14381 32385 14415 32419
rect 16681 32385 16715 32419
rect 16923 32385 16957 32419
rect 18319 32415 18353 32449
rect 19625 32385 19659 32419
rect 19717 32385 19751 32419
rect 19991 32385 20025 32419
rect 21649 32385 21683 32419
rect 23673 32385 23707 32419
rect 23949 32385 23983 32419
rect 1409 32317 1443 32351
rect 1593 32317 1627 32351
rect 2053 32317 2087 32351
rect 2446 32317 2480 32351
rect 2605 32317 2639 32351
rect 7573 32317 7607 32351
rect 7757 32317 7791 32351
rect 8493 32317 8527 32351
rect 8631 32317 8665 32351
rect 18061 32317 18095 32351
rect 21833 32317 21867 32351
rect 8217 32249 8251 32283
rect 11897 32249 11931 32283
rect 11069 32181 11103 32215
rect 15393 32181 15427 32215
rect 17693 32181 17727 32215
rect 21465 32181 21499 32215
rect 23489 32181 23523 32215
rect 23765 32181 23799 32215
rect 24409 32181 24443 32215
rect 2421 31977 2455 32011
rect 7113 31977 7147 32011
rect 8493 31977 8527 32011
rect 11529 31977 11563 32011
rect 17509 31977 17543 32011
rect 10333 31909 10367 31943
rect 16313 31909 16347 31943
rect 23029 31909 23063 31943
rect 2973 31841 3007 31875
rect 6101 31841 6135 31875
rect 7481 31841 7515 31875
rect 9689 31841 9723 31875
rect 9873 31841 9907 31875
rect 10726 31841 10760 31875
rect 10885 31841 10919 31875
rect 11897 31841 11931 31875
rect 12173 31841 12207 31875
rect 16589 31841 16623 31875
rect 16865 31841 16899 31875
rect 22385 31841 22419 31875
rect 23305 31841 23339 31875
rect 1409 31773 1443 31807
rect 1667 31743 1701 31777
rect 2789 31773 2823 31807
rect 4169 31773 4203 31807
rect 4443 31773 4477 31807
rect 6343 31773 6377 31807
rect 7755 31773 7789 31807
rect 10609 31773 10643 31807
rect 12415 31763 12449 31797
rect 15669 31773 15703 31807
rect 15853 31773 15887 31807
rect 16706 31773 16740 31807
rect 22293 31773 22327 31807
rect 22753 31773 22787 31807
rect 22937 31773 22971 31807
rect 23121 31773 23155 31807
rect 23213 31773 23247 31807
rect 23397 31773 23431 31807
rect 23673 31773 23707 31807
rect 23857 31773 23891 31807
rect 24225 31773 24259 31807
rect 5181 31637 5215 31671
rect 13185 31637 13219 31671
rect 23489 31637 23523 31671
rect 3985 31433 4019 31467
rect 12817 31433 12851 31467
rect 22845 31433 22879 31467
rect 23673 31433 23707 31467
rect 13921 31365 13955 31399
rect 24133 31365 24167 31399
rect 1501 31297 1535 31331
rect 2143 31297 2177 31331
rect 3249 31297 3283 31331
rect 3525 31297 3559 31331
rect 3801 31297 3835 31331
rect 4905 31297 4939 31331
rect 5179 31297 5213 31331
rect 8125 31297 8159 31331
rect 8399 31297 8433 31331
rect 13093 31297 13127 31331
rect 13185 31297 13219 31331
rect 13553 31297 13587 31331
rect 15467 31327 15501 31361
rect 18153 31297 18187 31331
rect 22075 31297 22109 31331
rect 23397 31297 23431 31331
rect 23857 31297 23891 31331
rect 1869 31229 1903 31263
rect 15209 31229 15243 31263
rect 21833 31229 21867 31263
rect 1685 31161 1719 31195
rect 3709 31161 3743 31195
rect 2881 31093 2915 31127
rect 3433 31093 3467 31127
rect 5917 31093 5951 31127
rect 9137 31093 9171 31127
rect 14105 31093 14139 31127
rect 16221 31093 16255 31127
rect 17969 31093 18003 31127
rect 23213 31093 23247 31127
rect 24409 31093 24443 31127
rect 3985 30889 4019 30923
rect 6101 30889 6135 30923
rect 12265 30889 12299 30923
rect 13645 30889 13679 30923
rect 23029 30889 23063 30923
rect 23305 30889 23339 30923
rect 18889 30821 18923 30855
rect 7481 30753 7515 30787
rect 10057 30753 10091 30787
rect 12633 30753 12667 30787
rect 15945 30753 15979 30787
rect 16221 30753 16255 30787
rect 16338 30753 16372 30787
rect 16497 30753 16531 30787
rect 17509 30753 17543 30787
rect 1409 30685 1443 30719
rect 1685 30685 1719 30719
rect 2329 30685 2363 30719
rect 2603 30685 2637 30719
rect 3801 30685 3835 30719
rect 5181 30685 5215 30719
rect 7723 30685 7757 30719
rect 10331 30685 10365 30719
rect 12875 30685 12909 30719
rect 15301 30685 15335 30719
rect 15485 30685 15519 30719
rect 17141 30685 17175 30719
rect 17776 30685 17810 30719
rect 19257 30685 19291 30719
rect 19533 30685 19567 30719
rect 19717 30685 19751 30719
rect 19993 30685 20027 30719
rect 20913 30685 20947 30719
rect 21097 30685 21131 30719
rect 23213 30685 23247 30719
rect 23489 30685 23523 30719
rect 5089 30617 5123 30651
rect 5549 30617 5583 30651
rect 11529 30617 11563 30651
rect 23857 30617 23891 30651
rect 24225 30617 24259 30651
rect 3341 30549 3375 30583
rect 4813 30549 4847 30583
rect 5917 30549 5951 30583
rect 8493 30549 8527 30583
rect 11069 30549 11103 30583
rect 11621 30549 11655 30583
rect 19349 30549 19383 30583
rect 19625 30549 19659 30583
rect 19809 30549 19843 30583
rect 21097 30549 21131 30583
rect 3985 30345 4019 30379
rect 15577 30345 15611 30379
rect 18981 30345 19015 30379
rect 20729 30345 20763 30379
rect 21465 30345 21499 30379
rect 23581 30345 23615 30379
rect 2697 30277 2731 30311
rect 3065 30277 3099 30311
rect 3801 30277 3835 30311
rect 7941 30277 7975 30311
rect 8217 30277 8251 30311
rect 8309 30277 8343 30311
rect 9045 30277 9079 30311
rect 12725 30277 12759 30311
rect 24133 30277 24167 30311
rect 1409 30209 1443 30243
rect 2053 30209 2087 30243
rect 2973 30209 3007 30243
rect 3433 30209 3467 30243
rect 4629 30209 4663 30243
rect 5147 30209 5181 30243
rect 6619 30209 6653 30243
rect 8677 30209 8711 30243
rect 9505 30209 9539 30243
rect 10425 30209 10459 30243
rect 12081 30209 12115 30243
rect 12265 30209 12299 30243
rect 14839 30209 14873 30243
rect 17969 30209 18003 30243
rect 18243 30209 18277 30243
rect 19605 30209 19639 30243
rect 20821 30209 20855 30243
rect 21189 30209 21223 30243
rect 21649 30209 21683 30243
rect 22661 30209 22695 30243
rect 22937 30209 22971 30243
rect 23213 30209 23247 30243
rect 23489 30209 23523 30243
rect 23765 30209 23799 30243
rect 1593 30141 1627 30175
rect 4905 30141 4939 30175
rect 6377 30141 6411 30175
rect 9689 30141 9723 30175
rect 10542 30141 10576 30175
rect 10701 30141 10735 30175
rect 14565 30141 14599 30175
rect 19349 30141 19383 30175
rect 21097 30171 21131 30205
rect 4813 30073 4847 30107
rect 10149 30073 10183 30107
rect 11897 30073 11931 30107
rect 12909 30073 12943 30107
rect 20913 30073 20947 30107
rect 21281 30073 21315 30107
rect 23029 30073 23063 30107
rect 2145 30005 2179 30039
rect 5917 30005 5951 30039
rect 7389 30005 7423 30039
rect 9229 30005 9263 30039
rect 11345 30005 11379 30039
rect 12357 30005 12391 30039
rect 21005 30005 21039 30039
rect 22477 30005 22511 30039
rect 22753 30005 22787 30039
rect 23305 30005 23339 30039
rect 24409 30005 24443 30039
rect 3525 29801 3559 29835
rect 11621 29801 11655 29835
rect 13553 29801 13587 29835
rect 19349 29801 19383 29835
rect 20913 29801 20947 29835
rect 23121 29801 23155 29835
rect 3985 29733 4019 29767
rect 5089 29733 5123 29767
rect 7849 29733 7883 29767
rect 12725 29733 12759 29767
rect 16497 29733 16531 29767
rect 4077 29665 4111 29699
rect 10425 29665 10459 29699
rect 10701 29665 10735 29699
rect 10839 29665 10873 29699
rect 13093 29665 13127 29699
rect 19533 29665 19567 29699
rect 19901 29665 19935 29699
rect 21373 29665 21407 29699
rect 1501 29597 1535 29631
rect 1775 29597 1809 29631
rect 3341 29597 3375 29631
rect 3801 29597 3835 29631
rect 4351 29597 4385 29631
rect 5457 29597 5491 29631
rect 5733 29597 5767 29631
rect 6837 29597 6871 29631
rect 6929 29597 6963 29631
rect 9781 29597 9815 29631
rect 9965 29597 9999 29631
rect 10977 29597 11011 29631
rect 11713 29597 11747 29631
rect 11987 29597 12021 29631
rect 13277 29597 13311 29631
rect 14105 29597 14139 29631
rect 14363 29567 14397 29601
rect 15485 29597 15519 29631
rect 15759 29597 15793 29631
rect 19257 29597 19291 29631
rect 19809 29597 19843 29631
rect 20175 29597 20209 29631
rect 21647 29597 21681 29631
rect 23305 29597 23339 29631
rect 23673 29597 23707 29631
rect 7297 29529 7331 29563
rect 13645 29529 13679 29563
rect 23857 29529 23891 29563
rect 24225 29529 24259 29563
rect 2513 29461 2547 29495
rect 6561 29461 6595 29495
rect 7665 29461 7699 29495
rect 15117 29461 15151 29495
rect 19533 29461 19567 29495
rect 19625 29461 19659 29495
rect 22385 29461 22419 29495
rect 23489 29461 23523 29495
rect 10149 29257 10183 29291
rect 11989 29257 12023 29291
rect 12633 29257 12667 29291
rect 2329 29121 2363 29155
rect 2605 29121 2639 29155
rect 3433 29121 3467 29155
rect 4995 29121 5029 29155
rect 9395 29151 9429 29185
rect 12173 29121 12207 29155
rect 12449 29121 12483 29155
rect 12633 29121 12667 29155
rect 12999 29121 13033 29155
rect 14379 29121 14413 29155
rect 17291 29121 17325 29155
rect 21373 29121 21407 29155
rect 22385 29121 22419 29155
rect 22569 29121 22603 29155
rect 23121 29121 23155 29155
rect 23397 29121 23431 29155
rect 23857 29121 23891 29155
rect 24133 29121 24167 29155
rect 1409 29053 1443 29087
rect 1593 29053 1627 29087
rect 2467 29053 2501 29087
rect 3709 29053 3743 29087
rect 4721 29053 4755 29087
rect 9137 29053 9171 29087
rect 12725 29053 12759 29087
rect 14105 29053 14139 29087
rect 17049 29053 17083 29087
rect 2053 28985 2087 29019
rect 3249 28985 3283 29019
rect 13737 28985 13771 29019
rect 15117 28985 15151 29019
rect 21189 28985 21223 29019
rect 22937 28985 22971 29019
rect 23213 28985 23247 29019
rect 24409 28985 24443 29019
rect 5733 28917 5767 28951
rect 18061 28917 18095 28951
rect 22477 28917 22511 28951
rect 23673 28917 23707 28951
rect 19073 28713 19107 28747
rect 20361 28713 20395 28747
rect 22845 28713 22879 28747
rect 23397 28713 23431 28747
rect 3341 28645 3375 28679
rect 5273 28645 5307 28679
rect 17877 28645 17911 28679
rect 22385 28645 22419 28679
rect 12633 28577 12667 28611
rect 15945 28577 15979 28611
rect 16338 28577 16372 28611
rect 16497 28577 16531 28611
rect 18153 28577 18187 28611
rect 22477 28577 22511 28611
rect 1869 28509 1903 28543
rect 2329 28509 2363 28543
rect 2603 28509 2637 28543
rect 4261 28509 4295 28543
rect 6285 28509 6319 28543
rect 6527 28509 6561 28543
rect 12891 28479 12925 28513
rect 15301 28509 15335 28543
rect 15485 28509 15519 28543
rect 16221 28509 16255 28543
rect 17233 28509 17267 28543
rect 17417 28509 17451 28543
rect 18270 28509 18304 28543
rect 18429 28509 18463 28543
rect 19901 28509 19935 28543
rect 19993 28509 20027 28543
rect 20177 28509 20211 28543
rect 20545 28509 20579 28543
rect 20637 28509 20671 28543
rect 22201 28509 22235 28543
rect 22293 28509 22327 28543
rect 22569 28509 22603 28543
rect 23029 28509 23063 28543
rect 23305 28509 23339 28543
rect 23581 28509 23615 28543
rect 23857 28509 23891 28543
rect 23949 28509 23983 28543
rect 1501 28441 1535 28475
rect 1685 28441 1719 28475
rect 4353 28441 4387 28475
rect 4721 28441 4755 28475
rect 20904 28441 20938 28475
rect 22661 28441 22695 28475
rect 1961 28373 1995 28407
rect 3985 28373 4019 28407
rect 5089 28373 5123 28407
rect 7297 28373 7331 28407
rect 13645 28373 13679 28407
rect 17141 28373 17175 28407
rect 19717 28373 19751 28407
rect 20085 28373 20119 28407
rect 22017 28373 22051 28407
rect 23121 28373 23155 28407
rect 23673 28373 23707 28407
rect 24133 28373 24167 28407
rect 2421 28169 2455 28203
rect 4077 28169 4111 28203
rect 4629 28169 4663 28203
rect 5733 28169 5767 28203
rect 11069 28169 11103 28203
rect 11805 28169 11839 28203
rect 17693 28169 17727 28203
rect 19441 28169 19475 28203
rect 21925 28169 21959 28203
rect 23213 28169 23247 28203
rect 5365 28101 5399 28135
rect 18306 28101 18340 28135
rect 24133 28101 24167 28135
rect 1683 28033 1717 28067
rect 2789 28033 2823 28067
rect 3307 28033 3341 28067
rect 4905 28033 4939 28067
rect 4997 28033 5031 28067
rect 7555 28033 7589 28067
rect 8919 28033 8953 28067
rect 10331 28033 10365 28067
rect 11529 28033 11563 28067
rect 15083 28033 15117 28067
rect 16681 28033 16715 28067
rect 16955 28033 16989 28067
rect 19807 28033 19841 28067
rect 21373 28033 21407 28067
rect 22109 28033 22143 28067
rect 22661 28033 22695 28067
rect 23397 28033 23431 28067
rect 23857 28033 23891 28067
rect 1409 27965 1443 27999
rect 3065 27965 3099 27999
rect 7297 27965 7331 27999
rect 8677 27965 8711 27999
rect 10057 27965 10091 27999
rect 11805 27965 11839 27999
rect 14841 27965 14875 27999
rect 18061 27965 18095 27999
rect 19533 27965 19567 27999
rect 5917 27897 5951 27931
rect 15853 27897 15887 27931
rect 21189 27897 21223 27931
rect 22477 27897 22511 27931
rect 2973 27829 3007 27863
rect 8309 27829 8343 27863
rect 9689 27829 9723 27863
rect 11621 27829 11655 27863
rect 20545 27829 20579 27863
rect 23673 27829 23707 27863
rect 24409 27829 24443 27863
rect 11253 27625 11287 27659
rect 11529 27625 11563 27659
rect 2973 27557 3007 27591
rect 3525 27557 3559 27591
rect 5641 27557 5675 27591
rect 10609 27557 10643 27591
rect 23121 27557 23155 27591
rect 11897 27489 11931 27523
rect 19441 27489 19475 27523
rect 19901 27489 19935 27523
rect 20085 27489 20119 27523
rect 1409 27421 1443 27455
rect 1683 27421 1717 27455
rect 2781 27417 2815 27451
rect 3065 27421 3099 27455
rect 3341 27421 3375 27455
rect 3801 27421 3835 27455
rect 4629 27421 4663 27455
rect 4903 27421 4937 27455
rect 6469 27421 6503 27455
rect 6561 27421 6595 27455
rect 11161 27421 11195 27455
rect 11437 27421 11471 27455
rect 11621 27421 11655 27455
rect 12171 27421 12205 27455
rect 14197 27421 14231 27455
rect 14471 27421 14505 27455
rect 18797 27421 18831 27455
rect 19349 27421 19383 27455
rect 19809 27421 19843 27455
rect 22661 27421 22695 27455
rect 23029 27421 23063 27455
rect 23305 27421 23339 27455
rect 23397 27421 23431 27455
rect 23857 27421 23891 27455
rect 6193 27353 6227 27387
rect 6929 27353 6963 27387
rect 9597 27353 9631 27387
rect 9689 27353 9723 27387
rect 10057 27353 10091 27387
rect 24225 27353 24259 27387
rect 2421 27285 2455 27319
rect 3249 27285 3283 27319
rect 3985 27285 4019 27319
rect 7297 27285 7331 27319
rect 7481 27285 7515 27319
rect 9321 27285 9355 27319
rect 10425 27285 10459 27319
rect 12909 27285 12943 27319
rect 15209 27285 15243 27319
rect 18613 27285 18647 27319
rect 20085 27285 20119 27319
rect 22477 27285 22511 27319
rect 22845 27285 22879 27319
rect 23581 27285 23615 27319
rect 1777 27081 1811 27115
rect 3065 27081 3099 27115
rect 3709 27081 3743 27115
rect 10333 27081 10367 27115
rect 11621 27081 11655 27115
rect 11897 27081 11931 27115
rect 15393 27081 15427 27115
rect 21833 27081 21867 27115
rect 2881 27013 2915 27047
rect 7757 27013 7791 27047
rect 8033 27013 8067 27047
rect 8125 27013 8159 27047
rect 8493 27013 8527 27047
rect 22652 27013 22686 27047
rect 23949 27013 23983 27047
rect 2053 26945 2087 26979
rect 2145 26945 2179 26979
rect 2513 26945 2547 26979
rect 3525 26945 3559 26979
rect 3801 26945 3835 26979
rect 4075 26945 4109 26979
rect 8875 26945 8909 26979
rect 9563 26945 9597 26979
rect 11805 26945 11839 26979
rect 12081 26945 12115 26979
rect 12447 26945 12481 26979
rect 13737 26945 13771 26979
rect 14590 26945 14624 26979
rect 14749 26945 14783 26979
rect 16955 26945 16989 26979
rect 22017 26945 22051 26979
rect 22109 26945 22143 26979
rect 22293 26945 22327 26979
rect 9321 26877 9355 26911
rect 12173 26877 12207 26911
rect 13553 26877 13587 26911
rect 14197 26877 14231 26911
rect 14473 26877 14507 26911
rect 16681 26877 16715 26911
rect 22385 26877 22419 26911
rect 4813 26741 4847 26775
rect 9045 26741 9079 26775
rect 13185 26741 13219 26775
rect 17693 26741 17727 26775
rect 22201 26741 22235 26775
rect 23765 26741 23799 26775
rect 24225 26741 24259 26775
rect 2789 26537 2823 26571
rect 8309 26537 8343 26571
rect 21373 26537 21407 26571
rect 22477 26537 22511 26571
rect 1593 26469 1627 26503
rect 14749 26469 14783 26503
rect 18061 26469 18095 26503
rect 1777 26401 1811 26435
rect 7297 26401 7331 26435
rect 14289 26401 14323 26435
rect 15301 26401 15335 26435
rect 16037 26401 16071 26435
rect 16221 26401 16255 26435
rect 16681 26401 16715 26435
rect 16957 26401 16991 26435
rect 17233 26401 17267 26435
rect 21465 26401 21499 26435
rect 22845 26401 22879 26435
rect 1409 26333 1443 26367
rect 2035 26303 2069 26337
rect 4261 26333 4295 26367
rect 4535 26323 4569 26357
rect 7571 26333 7605 26367
rect 11529 26333 11563 26367
rect 11803 26333 11837 26367
rect 14105 26333 14139 26367
rect 15025 26333 15059 26367
rect 15142 26333 15176 26367
rect 17074 26333 17108 26367
rect 17877 26333 17911 26367
rect 18245 26333 18279 26367
rect 18429 26333 18463 26367
rect 19993 26333 20027 26367
rect 21707 26333 21741 26367
rect 23119 26333 23153 26367
rect 15945 26265 15979 26299
rect 20238 26265 20272 26299
rect 5273 26197 5307 26231
rect 12541 26197 12575 26231
rect 18521 26197 18555 26231
rect 23857 26197 23891 26231
rect 2145 25993 2179 26027
rect 2697 25993 2731 26027
rect 5457 25993 5491 26027
rect 16221 25993 16255 26027
rect 18981 25993 19015 26027
rect 4169 25925 4203 25959
rect 4537 25925 4571 25959
rect 4905 25925 4939 25959
rect 5273 25925 5307 25959
rect 17868 25925 17902 25959
rect 24133 25925 24167 25959
rect 1409 25857 1443 25891
rect 1869 25857 1903 25891
rect 1961 25857 1995 25891
rect 2237 25857 2271 25891
rect 2513 25857 2547 25891
rect 4445 25857 4479 25891
rect 7847 25857 7881 25891
rect 10239 25857 10273 25891
rect 15483 25857 15517 25891
rect 19073 25857 19107 25891
rect 19165 25857 19199 25891
rect 19441 25857 19475 25891
rect 19625 25857 19659 25891
rect 19901 25857 19935 25891
rect 20637 25857 20671 25891
rect 21097 25857 21131 25891
rect 21833 25857 21867 25891
rect 22937 25857 22971 25891
rect 23213 25857 23247 25891
rect 23397 25857 23431 25891
rect 23673 25857 23707 25891
rect 7573 25789 7607 25823
rect 9965 25789 9999 25823
rect 15209 25789 15243 25823
rect 17601 25789 17635 25823
rect 19349 25789 19383 25823
rect 19533 25789 19567 25823
rect 22109 25789 22143 25823
rect 23305 25789 23339 25823
rect 23949 25789 23983 25823
rect 2421 25721 2455 25755
rect 19717 25721 19751 25755
rect 20453 25721 20487 25755
rect 23029 25721 23063 25755
rect 23765 25721 23799 25755
rect 1593 25653 1627 25687
rect 1685 25653 1719 25687
rect 6745 25653 6779 25687
rect 8585 25653 8619 25687
rect 10977 25653 11011 25687
rect 19257 25653 19291 25687
rect 21189 25653 21223 25687
rect 21925 25653 21959 25687
rect 22017 25653 22051 25687
rect 23857 25653 23891 25687
rect 24409 25653 24443 25687
rect 11529 25449 11563 25483
rect 18613 25449 18647 25483
rect 23489 25449 23523 25483
rect 2145 25381 2179 25415
rect 5733 25381 5767 25415
rect 12541 25381 12575 25415
rect 4721 25313 4755 25347
rect 9873 25313 9907 25347
rect 10333 25313 10367 25347
rect 10726 25313 10760 25347
rect 10885 25313 10919 25347
rect 11897 25313 11931 25347
rect 12817 25313 12851 25347
rect 14105 25313 14139 25347
rect 14749 25313 14783 25347
rect 15025 25313 15059 25347
rect 15142 25313 15176 25347
rect 15301 25313 15335 25347
rect 1409 25245 1443 25279
rect 1685 25245 1719 25279
rect 1961 25245 1995 25279
rect 2329 25245 2363 25279
rect 2603 25245 2637 25279
rect 4963 25245 4997 25279
rect 9689 25245 9723 25279
rect 10609 25245 10643 25279
rect 12081 25245 12115 25279
rect 12934 25245 12968 25279
rect 13093 25245 13127 25279
rect 14289 25245 14323 25279
rect 17601 25245 17635 25279
rect 17875 25245 17909 25279
rect 20269 25245 20303 25279
rect 20361 25245 20395 25279
rect 20545 25245 20579 25279
rect 23673 25245 23707 25279
rect 6561 25177 6595 25211
rect 6653 25177 6687 25211
rect 7021 25177 7055 25211
rect 7389 25177 7423 25211
rect 23857 25177 23891 25211
rect 1593 25109 1627 25143
rect 1869 25109 1903 25143
rect 3341 25109 3375 25143
rect 6285 25109 6319 25143
rect 7573 25109 7607 25143
rect 13737 25109 13771 25143
rect 15945 25109 15979 25143
rect 20085 25109 20119 25143
rect 20453 25109 20487 25143
rect 24133 25109 24167 25143
rect 4537 24905 4571 24939
rect 7389 24905 7423 24939
rect 9321 24905 9355 24939
rect 13185 24905 13219 24939
rect 19901 24905 19935 24939
rect 3433 24837 3467 24871
rect 4169 24837 4203 24871
rect 8033 24837 8067 24871
rect 8309 24837 8343 24871
rect 9137 24837 9171 24871
rect 1409 24769 1443 24803
rect 1683 24769 1717 24803
rect 2789 24769 2823 24803
rect 3709 24769 3743 24803
rect 3801 24769 3835 24803
rect 6619 24769 6653 24803
rect 8401 24769 8435 24803
rect 8769 24769 8803 24803
rect 10542 24769 10576 24803
rect 10701 24769 10735 24803
rect 11345 24769 11379 24803
rect 12447 24769 12481 24803
rect 16405 24769 16439 24803
rect 17509 24769 17543 24803
rect 18777 24769 18811 24803
rect 19993 24769 20027 24803
rect 20267 24769 20301 24803
rect 22109 24769 22143 24803
rect 22753 24769 22787 24803
rect 23213 24769 23247 24803
rect 23305 24769 23339 24803
rect 23581 24769 23615 24803
rect 23765 24769 23799 24803
rect 24133 24769 24167 24803
rect 6377 24701 6411 24735
rect 9505 24701 9539 24735
rect 9689 24701 9723 24735
rect 10149 24701 10183 24735
rect 10425 24701 10459 24735
rect 12173 24701 12207 24735
rect 18521 24701 18555 24735
rect 2973 24633 3007 24667
rect 4721 24633 4755 24667
rect 23029 24633 23063 24667
rect 2421 24565 2455 24599
rect 16221 24565 16255 24599
rect 17325 24565 17359 24599
rect 21005 24565 21039 24599
rect 21925 24565 21959 24599
rect 22569 24565 22603 24599
rect 23489 24565 23523 24599
rect 23673 24565 23707 24599
rect 24409 24565 24443 24599
rect 3065 24361 3099 24395
rect 4813 24361 4847 24395
rect 10241 24361 10275 24395
rect 15945 24361 15979 24395
rect 21741 24361 21775 24395
rect 23397 24361 23431 24395
rect 14749 24293 14783 24327
rect 3801 24225 3835 24259
rect 9229 24225 9263 24259
rect 11621 24225 11655 24259
rect 11805 24225 11839 24259
rect 12265 24225 12299 24259
rect 12679 24225 12713 24259
rect 14105 24225 14139 24259
rect 14289 24225 14323 24259
rect 15025 24225 15059 24259
rect 15142 24225 15176 24259
rect 15301 24225 15335 24259
rect 17049 24225 17083 24259
rect 19809 24225 19843 24259
rect 20085 24225 20119 24259
rect 20269 24225 20303 24259
rect 4075 24157 4109 24191
rect 9503 24157 9537 24191
rect 12541 24157 12575 24191
rect 12817 24157 12851 24191
rect 16589 24157 16623 24191
rect 16773 24157 16807 24191
rect 17323 24157 17357 24191
rect 19441 24157 19475 24191
rect 19717 24157 19751 24191
rect 19993 24157 20027 24191
rect 20361 24157 20395 24191
rect 22017 24157 22051 24191
rect 22273 24157 22307 24191
rect 23489 24157 23523 24191
rect 23949 24157 23983 24191
rect 1777 24089 1811 24123
rect 2053 24089 2087 24123
rect 2145 24089 2179 24123
rect 2513 24089 2547 24123
rect 20606 24089 20640 24123
rect 2881 24021 2915 24055
rect 13461 24021 13495 24055
rect 16865 24021 16899 24055
rect 18061 24021 18095 24055
rect 19257 24021 19291 24055
rect 20269 24021 20303 24055
rect 23581 24021 23615 24055
rect 24133 24021 24167 24055
rect 2789 23817 2823 23851
rect 3617 23817 3651 23851
rect 9137 23817 9171 23851
rect 12541 23817 12575 23851
rect 20821 23817 20855 23851
rect 23489 23817 23523 23851
rect 1501 23681 1535 23715
rect 1777 23681 1811 23715
rect 2051 23681 2085 23715
rect 3157 23681 3191 23715
rect 3433 23681 3467 23715
rect 4353 23681 4387 23715
rect 4537 23681 4571 23715
rect 5273 23681 5307 23715
rect 8399 23681 8433 23715
rect 11529 23681 11563 23715
rect 11803 23681 11837 23715
rect 15267 23681 15301 23715
rect 16939 23711 16973 23745
rect 18061 23681 18095 23715
rect 18245 23681 18279 23715
rect 18613 23681 18647 23715
rect 21005 23681 21039 23715
rect 21465 23681 21499 23715
rect 21833 23681 21867 23715
rect 22201 23681 22235 23715
rect 22385 23681 22419 23715
rect 22477 23681 22511 23715
rect 22751 23681 22785 23715
rect 24133 23681 24167 23715
rect 5390 23613 5424 23647
rect 5549 23613 5583 23647
rect 8125 23613 8159 23647
rect 15025 23613 15059 23647
rect 16681 23613 16715 23647
rect 22109 23613 22143 23647
rect 22293 23613 22327 23647
rect 1685 23545 1719 23579
rect 4997 23545 5031 23579
rect 18337 23545 18371 23579
rect 3341 23477 3375 23511
rect 6193 23477 6227 23511
rect 16037 23477 16071 23511
rect 17693 23477 17727 23511
rect 21557 23477 21591 23511
rect 21925 23477 21959 23511
rect 22017 23477 22051 23511
rect 24409 23477 24443 23511
rect 5825 23273 5859 23307
rect 6929 23273 6963 23307
rect 17785 23273 17819 23307
rect 21925 23273 21959 23307
rect 23949 23273 23983 23307
rect 24041 23273 24075 23307
rect 16037 23205 16071 23239
rect 1409 23137 1443 23171
rect 3065 23137 3099 23171
rect 7389 23137 7423 23171
rect 15393 23137 15427 23171
rect 16430 23137 16464 23171
rect 20913 23137 20947 23171
rect 24133 23137 24167 23171
rect 1683 23069 1717 23103
rect 2789 23069 2823 23103
rect 4813 23069 4847 23103
rect 5087 23069 5121 23103
rect 6653 23069 6687 23103
rect 6837 23069 6871 23103
rect 7113 23069 7147 23103
rect 7297 23069 7331 23103
rect 7663 23069 7697 23103
rect 9137 23069 9171 23103
rect 9965 23069 9999 23103
rect 10239 23069 10273 23103
rect 15577 23069 15611 23103
rect 16313 23069 16347 23103
rect 16589 23069 16623 23103
rect 17693 23069 17727 23103
rect 17877 23069 17911 23103
rect 21155 23069 21189 23103
rect 23397 23069 23431 23103
rect 23489 23069 23523 23103
rect 23857 23069 23891 23103
rect 2421 22933 2455 22967
rect 6469 22933 6503 22967
rect 7297 22933 7331 22967
rect 8401 22933 8435 22967
rect 10977 22933 11011 22967
rect 17233 22933 17267 22967
rect 23213 22933 23247 22967
rect 23673 22933 23707 22967
rect 9045 22729 9079 22763
rect 9229 22729 9263 22763
rect 9965 22729 9999 22763
rect 19901 22729 19935 22763
rect 23673 22729 23707 22763
rect 7941 22661 7975 22695
rect 8217 22661 8251 22695
rect 10241 22661 10275 22695
rect 10333 22661 10367 22695
rect 11069 22661 11103 22695
rect 18398 22661 18432 22695
rect 1409 22593 1443 22627
rect 1683 22603 1717 22637
rect 2789 22593 2823 22627
rect 3801 22593 3835 22627
rect 4353 22593 4387 22627
rect 5390 22593 5424 22627
rect 6651 22593 6685 22627
rect 8309 22593 8343 22627
rect 8677 22593 8711 22627
rect 10701 22593 10735 22627
rect 11713 22593 11747 22627
rect 12967 22593 13001 22627
rect 14439 22593 14473 22627
rect 19625 22593 19659 22627
rect 20085 22593 20119 22627
rect 20177 22593 20211 22627
rect 20361 22593 20395 22627
rect 23397 22593 23431 22627
rect 23581 22593 23615 22627
rect 23857 22593 23891 22627
rect 24133 22593 24167 22627
rect 4537 22525 4571 22559
rect 4997 22525 5031 22559
rect 5273 22525 5307 22559
rect 5549 22525 5583 22559
rect 6377 22525 6411 22559
rect 12725 22525 12759 22559
rect 14197 22525 14231 22559
rect 18153 22525 18187 22559
rect 2973 22457 3007 22491
rect 11253 22457 11287 22491
rect 19533 22457 19567 22491
rect 2421 22389 2455 22423
rect 3985 22389 4019 22423
rect 6193 22389 6227 22423
rect 7389 22389 7423 22423
rect 11897 22389 11931 22423
rect 13737 22389 13771 22423
rect 15209 22389 15243 22423
rect 15761 22389 15795 22423
rect 19717 22389 19751 22423
rect 20269 22389 20303 22423
rect 23489 22389 23523 22423
rect 24409 22389 24443 22423
rect 2881 22185 2915 22219
rect 4905 22185 4939 22219
rect 7573 22185 7607 22219
rect 10517 22185 10551 22219
rect 19809 22185 19843 22219
rect 7389 22117 7423 22151
rect 15117 22117 15151 22151
rect 21649 22117 21683 22151
rect 21833 22117 21867 22151
rect 3893 22049 3927 22083
rect 7205 22049 7239 22083
rect 9505 22049 9539 22083
rect 11253 22049 11287 22083
rect 12633 22049 12667 22083
rect 15393 22049 15427 22083
rect 15531 22049 15565 22083
rect 19993 22049 20027 22083
rect 20269 22049 20303 22083
rect 1961 21981 1995 22015
rect 4151 21951 4185 21985
rect 7113 21981 7147 22015
rect 7481 21981 7515 22015
rect 7757 21981 7791 22015
rect 9779 21981 9813 22015
rect 11511 21951 11545 21985
rect 12875 21981 12909 22015
rect 14473 21981 14507 22015
rect 14657 21981 14691 22015
rect 15669 21981 15703 22015
rect 18889 21981 18923 22015
rect 19717 21981 19751 22015
rect 22017 21981 22051 22015
rect 22385 21981 22419 22015
rect 23949 21981 23983 22015
rect 1869 21913 1903 21947
rect 2329 21913 2363 21947
rect 2697 21913 2731 21947
rect 20536 21913 20570 21947
rect 22630 21913 22664 21947
rect 1593 21845 1627 21879
rect 12265 21845 12299 21879
rect 13645 21845 13679 21879
rect 16313 21845 16347 21879
rect 18705 21845 18739 21879
rect 19993 21845 20027 21879
rect 23765 21845 23799 21879
rect 24133 21845 24167 21879
rect 1869 21641 1903 21675
rect 9229 21641 9263 21675
rect 13185 21641 13219 21675
rect 14289 21641 14323 21675
rect 15761 21641 15795 21675
rect 19901 21641 19935 21675
rect 23765 21641 23799 21675
rect 13553 21573 13587 21607
rect 1409 21505 1443 21539
rect 1685 21505 1719 21539
rect 1961 21505 1995 21539
rect 2237 21505 2271 21539
rect 2511 21505 2545 21539
rect 3891 21505 3925 21539
rect 6895 21505 6929 21539
rect 8217 21505 8251 21539
rect 8491 21515 8525 21549
rect 11803 21505 11837 21539
rect 13461 21505 13495 21539
rect 13921 21505 13955 21539
rect 15023 21505 15057 21539
rect 16681 21505 16715 21539
rect 17718 21505 17752 21539
rect 19131 21505 19165 21539
rect 21005 21505 21039 21539
rect 21465 21505 21499 21539
rect 21833 21505 21867 21539
rect 22201 21505 22235 21539
rect 22385 21505 22419 21539
rect 22661 21505 22695 21539
rect 23011 21535 23045 21569
rect 24133 21505 24167 21539
rect 3617 21437 3651 21471
rect 6653 21437 6687 21471
rect 11529 21437 11563 21471
rect 14749 21437 14783 21471
rect 16865 21437 16899 21471
rect 17601 21437 17635 21471
rect 17877 21437 17911 21471
rect 18889 21437 18923 21471
rect 22109 21437 22143 21471
rect 22293 21437 22327 21471
rect 22753 21437 22787 21471
rect 24409 21437 24443 21471
rect 1593 21369 1627 21403
rect 17325 21369 17359 21403
rect 20821 21369 20855 21403
rect 22017 21369 22051 21403
rect 24317 21369 24351 21403
rect 2145 21301 2179 21335
rect 3249 21301 3283 21335
rect 4629 21301 4663 21335
rect 7665 21301 7699 21335
rect 12541 21301 12575 21335
rect 14473 21301 14507 21335
rect 18521 21301 18555 21335
rect 21557 21301 21591 21335
rect 21925 21301 21959 21335
rect 22477 21301 22511 21335
rect 24225 21301 24259 21335
rect 1593 21097 1627 21131
rect 1961 21097 1995 21131
rect 7113 21097 7147 21131
rect 18981 21097 19015 21131
rect 22201 21097 22235 21131
rect 23397 21097 23431 21131
rect 12173 21029 12207 21063
rect 16037 21029 16071 21063
rect 17049 21029 17083 21063
rect 18337 21029 18371 21063
rect 2145 20961 2179 20995
rect 4721 20961 4755 20995
rect 9413 20961 9447 20995
rect 11529 20961 11563 20995
rect 11713 20961 11747 20995
rect 15025 20961 15059 20995
rect 21189 20961 21223 20995
rect 1777 20893 1811 20927
rect 2419 20893 2453 20927
rect 4995 20893 5029 20927
rect 8125 20893 8159 20927
rect 9655 20893 9689 20927
rect 12449 20893 12483 20927
rect 12566 20893 12600 20927
rect 12725 20893 12759 20927
rect 15283 20863 15317 20897
rect 16405 20893 16439 20927
rect 16589 20893 16623 20927
rect 17325 20893 17359 20927
rect 17442 20893 17476 20927
rect 17601 20893 17635 20927
rect 18529 20889 18563 20923
rect 18797 20893 18831 20927
rect 18889 20893 18923 20927
rect 19901 20893 19935 20927
rect 21431 20893 21465 20927
rect 23305 20893 23339 20927
rect 23673 20893 23707 20927
rect 1501 20825 1535 20859
rect 7389 20825 7423 20859
rect 7665 20825 7699 20859
rect 7757 20825 7791 20859
rect 18245 20825 18279 20859
rect 3157 20757 3191 20791
rect 5733 20757 5767 20791
rect 8493 20757 8527 20791
rect 8677 20757 8711 20791
rect 10425 20757 10459 20791
rect 13369 20757 13403 20791
rect 18613 20757 18647 20791
rect 19717 20757 19751 20791
rect 23949 20757 23983 20791
rect 1639 20553 1673 20587
rect 2513 20553 2547 20587
rect 4813 20553 4847 20587
rect 8585 20553 8619 20587
rect 9413 20553 9447 20587
rect 18061 20553 18095 20587
rect 23121 20553 23155 20587
rect 24317 20553 24351 20587
rect 2881 20485 2915 20519
rect 3617 20485 3651 20519
rect 3985 20485 4019 20519
rect 5917 20485 5951 20519
rect 9781 20485 9815 20519
rect 10517 20485 10551 20519
rect 19421 20485 19455 20519
rect 24041 20485 24075 20519
rect 1409 20417 1443 20451
rect 2329 20417 2363 20451
rect 3157 20417 3191 20451
rect 3249 20417 3283 20451
rect 5089 20417 5123 20451
rect 5181 20417 5215 20451
rect 5549 20417 5583 20451
rect 7815 20417 7849 20451
rect 9689 20417 9723 20451
rect 10149 20417 10183 20451
rect 12725 20417 12759 20451
rect 17049 20417 17083 20451
rect 17291 20417 17325 20451
rect 18521 20417 18555 20451
rect 18613 20417 18647 20451
rect 19165 20417 19199 20451
rect 20637 20417 20671 20451
rect 21097 20417 21131 20451
rect 22845 20417 22879 20451
rect 23305 20417 23339 20451
rect 23489 20417 23523 20451
rect 7573 20349 7607 20383
rect 18797 20349 18831 20383
rect 20545 20281 20579 20315
rect 4169 20213 4203 20247
rect 6101 20213 6135 20247
rect 10701 20213 10735 20247
rect 18705 20213 18739 20247
rect 20729 20213 20763 20247
rect 20913 20213 20947 20247
rect 22661 20213 22695 20247
rect 23765 20213 23799 20247
rect 1593 20009 1627 20043
rect 3525 20009 3559 20043
rect 6285 20009 6319 20043
rect 18705 20009 18739 20043
rect 19349 20009 19383 20043
rect 21281 20009 21315 20043
rect 22017 20009 22051 20043
rect 2697 19941 2731 19975
rect 10701 19941 10735 19975
rect 11713 19941 11747 19975
rect 20821 19941 20855 19975
rect 9689 19873 9723 19907
rect 11069 19873 11103 19907
rect 11253 19873 11287 19907
rect 12106 19873 12140 19907
rect 14473 19873 14507 19907
rect 17693 19873 17727 19907
rect 19809 19873 19843 19907
rect 21465 19873 21499 19907
rect 21649 19873 21683 19907
rect 1409 19805 1443 19839
rect 1685 19805 1719 19839
rect 1959 19805 1993 19839
rect 3065 19805 3099 19839
rect 3341 19805 3375 19839
rect 3801 19805 3835 19839
rect 5273 19805 5307 19839
rect 5547 19805 5581 19839
rect 9947 19775 9981 19809
rect 11989 19805 12023 19839
rect 12263 19805 12297 19839
rect 13921 19805 13955 19839
rect 14747 19805 14781 19839
rect 17951 19775 17985 19809
rect 19257 19805 19291 19839
rect 19441 19805 19475 19839
rect 20067 19775 20101 19809
rect 21189 19805 21223 19839
rect 21557 19805 21591 19839
rect 21741 19805 21775 19839
rect 21833 19805 21867 19839
rect 22201 19805 22235 19839
rect 23857 19805 23891 19839
rect 22468 19737 22502 19771
rect 24225 19737 24259 19771
rect 3249 19669 3283 19703
rect 3985 19669 4019 19703
rect 12909 19669 12943 19703
rect 15485 19669 15519 19703
rect 21465 19669 21499 19703
rect 23581 19669 23615 19703
rect 8493 19465 8527 19499
rect 9965 19465 9999 19499
rect 12541 19465 12575 19499
rect 24133 19397 24167 19431
rect 1409 19329 1443 19363
rect 1683 19329 1717 19363
rect 2881 19329 2915 19363
rect 3431 19329 3465 19363
rect 7739 19329 7773 19363
rect 8953 19329 8987 19363
rect 9211 19329 9245 19363
rect 11529 19329 11563 19363
rect 11787 19359 11821 19393
rect 12909 19329 12943 19363
rect 13183 19329 13217 19363
rect 14289 19329 14323 19363
rect 15485 19329 15519 19363
rect 16939 19359 16973 19393
rect 22477 19329 22511 19363
rect 22751 19329 22785 19363
rect 3152 19261 3186 19295
rect 7481 19261 7515 19295
rect 14473 19261 14507 19295
rect 15209 19261 15243 19295
rect 15326 19261 15360 19295
rect 16681 19261 16715 19295
rect 14933 19193 14967 19227
rect 2421 19125 2455 19159
rect 2973 19125 3007 19159
rect 4169 19125 4203 19159
rect 13921 19125 13955 19159
rect 16129 19125 16163 19159
rect 16497 19125 16531 19159
rect 17693 19125 17727 19159
rect 23489 19125 23523 19159
rect 24409 19125 24443 19159
rect 15117 18921 15151 18955
rect 1961 18853 1995 18887
rect 6837 18853 6871 18887
rect 20545 18853 20579 18887
rect 22937 18853 22971 18887
rect 23489 18853 23523 18887
rect 2329 18785 2363 18819
rect 4261 18785 4295 18819
rect 12449 18785 12483 18819
rect 15761 18785 15795 18819
rect 16405 18785 16439 18819
rect 16681 18785 16715 18819
rect 16957 18785 16991 18819
rect 23673 18785 23707 18819
rect 1409 18717 1443 18751
rect 1777 18717 1811 18751
rect 2587 18687 2621 18721
rect 4535 18717 4569 18751
rect 5825 18717 5859 18751
rect 6083 18687 6117 18721
rect 7665 18717 7699 18751
rect 7757 18717 7791 18751
rect 8125 18717 8159 18751
rect 12691 18717 12725 18751
rect 14105 18717 14139 18751
rect 14379 18717 14413 18751
rect 15945 18717 15979 18751
rect 16819 18717 16853 18751
rect 19625 18717 19659 18751
rect 19809 18717 19843 18751
rect 20729 18717 20763 18751
rect 21281 18717 21315 18751
rect 22845 18717 22879 18751
rect 23305 18717 23339 18751
rect 23397 18717 23431 18751
rect 23857 18717 23891 18751
rect 1593 18581 1627 18615
rect 3341 18581 3375 18615
rect 5273 18581 5307 18615
rect 7389 18581 7423 18615
rect 8493 18581 8527 18615
rect 8677 18581 8711 18615
rect 13461 18581 13495 18615
rect 17601 18581 17635 18615
rect 19717 18581 19751 18615
rect 21373 18581 21407 18615
rect 23121 18581 23155 18615
rect 23673 18581 23707 18615
rect 24133 18581 24167 18615
rect 5825 18377 5859 18411
rect 6561 18377 6595 18411
rect 7849 18377 7883 18411
rect 9689 18377 9723 18411
rect 16221 18377 16255 18411
rect 19349 18377 19383 18411
rect 19717 18377 19751 18411
rect 23581 18377 23615 18411
rect 24409 18377 24443 18411
rect 1501 18309 1535 18343
rect 1685 18309 1719 18343
rect 7665 18309 7699 18343
rect 20341 18309 20375 18343
rect 22109 18309 22143 18343
rect 1961 18241 1995 18275
rect 3249 18241 3283 18275
rect 5022 18241 5056 18275
rect 5181 18241 5215 18275
rect 6193 18241 6227 18275
rect 6837 18241 6871 18275
rect 6929 18241 6963 18275
rect 7297 18241 7331 18275
rect 8951 18241 8985 18275
rect 10609 18241 10643 18275
rect 12817 18241 12851 18275
rect 13001 18241 13035 18275
rect 13737 18241 13771 18275
rect 14013 18241 14047 18275
rect 15209 18241 15243 18275
rect 15467 18271 15501 18305
rect 17969 18241 18003 18275
rect 18225 18241 18259 18275
rect 19441 18241 19475 18275
rect 19901 18241 19935 18275
rect 21833 18241 21867 18275
rect 21925 18241 21959 18275
rect 22385 18241 22419 18275
rect 22477 18241 22511 18275
rect 22661 18241 22695 18275
rect 22845 18241 22879 18275
rect 23305 18241 23339 18275
rect 23397 18241 23431 18275
rect 23581 18241 23615 18275
rect 23765 18241 23799 18275
rect 24225 18241 24259 18275
rect 2053 18173 2087 18207
rect 2237 18173 2271 18207
rect 2973 18173 3007 18207
rect 3111 18173 3145 18207
rect 3985 18173 4019 18207
rect 4169 18173 4203 18207
rect 4629 18173 4663 18207
rect 4905 18173 4939 18207
rect 8677 18173 8711 18207
rect 13461 18173 13495 18207
rect 13854 18173 13888 18207
rect 20085 18173 20119 18207
rect 22109 18173 22143 18207
rect 22569 18173 22603 18207
rect 2697 18105 2731 18139
rect 14657 18105 14691 18139
rect 21465 18105 21499 18139
rect 22201 18105 22235 18139
rect 23121 18105 23155 18139
rect 1777 18037 1811 18071
rect 3893 18037 3927 18071
rect 10425 18037 10459 18071
rect 11989 18037 12023 18071
rect 19533 18037 19567 18071
rect 22937 18037 22971 18071
rect 24041 18037 24075 18071
rect 5457 17833 5491 17867
rect 6837 17833 6871 17867
rect 10885 17833 10919 17867
rect 12817 17833 12851 17867
rect 18429 17833 18463 17867
rect 20269 17833 20303 17867
rect 21741 17833 21775 17867
rect 2329 17765 2363 17799
rect 9689 17765 9723 17799
rect 2605 17697 2639 17731
rect 2881 17697 2915 17731
rect 9965 17697 9999 17731
rect 19257 17697 19291 17731
rect 1593 17629 1627 17663
rect 1685 17629 1719 17663
rect 1869 17629 1903 17663
rect 2743 17629 2777 17663
rect 4445 17629 4479 17663
rect 4719 17629 4753 17663
rect 5825 17629 5859 17663
rect 6099 17629 6133 17663
rect 9045 17629 9079 17663
rect 9229 17629 9263 17663
rect 10103 17629 10137 17663
rect 10241 17629 10275 17663
rect 11805 17629 11839 17663
rect 12265 17629 12299 17663
rect 16957 17629 16991 17663
rect 18245 17629 18279 17663
rect 18613 17629 18647 17663
rect 19531 17629 19565 17663
rect 20729 17629 20763 17663
rect 20971 17629 21005 17663
rect 22569 17629 22603 17663
rect 22661 17629 22695 17663
rect 22917 17629 22951 17663
rect 11529 17561 11563 17595
rect 11897 17561 11931 17595
rect 1409 17493 1443 17527
rect 3525 17493 3559 17527
rect 12633 17493 12667 17527
rect 17141 17493 17175 17527
rect 22385 17493 22419 17527
rect 24041 17493 24075 17527
rect 1777 17289 1811 17323
rect 2329 17289 2363 17323
rect 3801 17289 3835 17323
rect 10517 17289 10551 17323
rect 12725 17289 12759 17323
rect 24501 17289 24535 17323
rect 1685 17221 1719 17255
rect 3341 17221 3375 17255
rect 2237 17153 2271 17187
rect 2789 17153 2823 17187
rect 3985 17153 4019 17187
rect 8275 17153 8309 17187
rect 9505 17153 9539 17187
rect 9779 17153 9813 17187
rect 11987 17153 12021 17187
rect 15025 17153 15059 17187
rect 15299 17153 15333 17187
rect 16681 17153 16715 17187
rect 16955 17153 16989 17187
rect 18303 17153 18337 17187
rect 19441 17153 19475 17187
rect 19533 17153 19567 17187
rect 22017 17153 22051 17187
rect 23087 17153 23121 17187
rect 24225 17153 24259 17187
rect 8033 17085 8067 17119
rect 11713 17085 11747 17119
rect 18061 17085 18095 17119
rect 19717 17085 19751 17119
rect 22845 17085 22879 17119
rect 24317 17085 24351 17119
rect 24501 17085 24535 17119
rect 19625 17017 19659 17051
rect 2881 16949 2915 16983
rect 3433 16949 3467 16983
rect 9045 16949 9079 16983
rect 14197 16949 14231 16983
rect 16037 16949 16071 16983
rect 17693 16949 17727 16983
rect 19073 16949 19107 16983
rect 21833 16949 21867 16983
rect 23857 16949 23891 16983
rect 3249 16745 3283 16779
rect 11805 16745 11839 16779
rect 17325 16745 17359 16779
rect 23397 16745 23431 16779
rect 8217 16677 8251 16711
rect 4077 16609 4111 16643
rect 7205 16609 7239 16643
rect 10793 16609 10827 16643
rect 12633 16609 12667 16643
rect 15485 16609 15519 16643
rect 15669 16609 15703 16643
rect 16129 16609 16163 16643
rect 16522 16609 16556 16643
rect 16681 16609 16715 16643
rect 21005 16609 21039 16643
rect 23949 16609 23983 16643
rect 1593 16541 1627 16575
rect 1685 16541 1719 16575
rect 1959 16541 1993 16575
rect 4351 16541 4385 16575
rect 7447 16541 7481 16575
rect 11051 16511 11085 16545
rect 12907 16541 12941 16575
rect 14105 16541 14139 16575
rect 14379 16541 14413 16575
rect 16405 16541 16439 16575
rect 17417 16541 17451 16575
rect 17675 16511 17709 16545
rect 21272 16541 21306 16575
rect 22477 16541 22511 16575
rect 22937 16541 22971 16575
rect 23029 16541 23063 16575
rect 23213 16541 23247 16575
rect 23305 16541 23339 16575
rect 23489 16541 23523 16575
rect 23673 16541 23707 16575
rect 3157 16473 3191 16507
rect 1409 16405 1443 16439
rect 2697 16405 2731 16439
rect 5089 16405 5123 16439
rect 13645 16405 13679 16439
rect 15117 16405 15151 16439
rect 18429 16405 18463 16439
rect 22385 16405 22419 16439
rect 22569 16405 22603 16439
rect 22753 16405 22787 16439
rect 23213 16405 23247 16439
rect 5641 16201 5675 16235
rect 9505 16201 9539 16235
rect 10977 16201 11011 16235
rect 13645 16201 13679 16235
rect 14933 16201 14967 16235
rect 20453 16201 20487 16235
rect 24317 16201 24351 16235
rect 1501 16133 1535 16167
rect 13921 16133 13955 16167
rect 14749 16133 14783 16167
rect 18889 16133 18923 16167
rect 19340 16133 19374 16167
rect 24041 16133 24075 16167
rect 2329 16065 2363 16099
rect 2421 16065 2455 16099
rect 2695 16065 2729 16099
rect 3801 16065 3835 16099
rect 4838 16065 4872 16099
rect 4997 16065 5031 16099
rect 7665 16065 7699 16099
rect 8861 16065 8895 16099
rect 9871 16065 9905 16099
rect 11161 16065 11195 16099
rect 14013 16065 14047 16099
rect 14381 16065 14415 16099
rect 17049 16065 17083 16099
rect 17969 16065 18003 16099
rect 19073 16065 19107 16099
rect 20545 16065 20579 16099
rect 21005 16065 21039 16099
rect 22091 16095 22125 16129
rect 23489 16065 23523 16099
rect 3985 15997 4019 16031
rect 4721 15997 4755 16031
rect 7849 15997 7883 16031
rect 8309 15997 8343 16031
rect 8585 15997 8619 16031
rect 8723 15997 8757 16031
rect 9597 15997 9631 16031
rect 17233 15997 17267 16031
rect 18086 15997 18120 16031
rect 18245 15997 18279 16031
rect 21833 15997 21867 16031
rect 3433 15929 3467 15963
rect 4445 15929 4479 15963
rect 17693 15929 17727 15963
rect 1593 15861 1627 15895
rect 2145 15861 2179 15895
rect 10609 15861 10643 15895
rect 20637 15861 20671 15895
rect 20821 15861 20855 15895
rect 22845 15861 22879 15895
rect 23765 15861 23799 15895
rect 4629 15657 4663 15691
rect 11253 15657 11287 15691
rect 19533 15657 19567 15691
rect 21281 15657 21315 15691
rect 23305 15657 23339 15691
rect 2421 15589 2455 15623
rect 3801 15589 3835 15623
rect 10057 15589 10091 15623
rect 20821 15589 20855 15623
rect 1777 15521 1811 15555
rect 2697 15521 2731 15555
rect 2835 15521 2869 15555
rect 7021 15521 7055 15555
rect 9413 15521 9447 15555
rect 10333 15521 10367 15555
rect 19809 15521 19843 15555
rect 21465 15521 21499 15555
rect 21649 15521 21683 15555
rect 23489 15521 23523 15555
rect 1961 15453 1995 15487
rect 2973 15453 3007 15487
rect 3617 15453 3651 15487
rect 3985 15453 4019 15487
rect 5917 15453 5951 15487
rect 7295 15453 7329 15487
rect 9597 15453 9631 15487
rect 10450 15453 10484 15487
rect 10609 15453 10643 15487
rect 11805 15453 11839 15487
rect 12079 15453 12113 15487
rect 13185 15453 13219 15487
rect 13553 15453 13587 15487
rect 19717 15453 19751 15487
rect 20067 15423 20101 15457
rect 21189 15453 21223 15487
rect 21557 15453 21591 15487
rect 21741 15453 21775 15487
rect 22661 15453 22695 15487
rect 22937 15453 22971 15487
rect 23121 15453 23155 15487
rect 23213 15453 23247 15487
rect 23857 15453 23891 15487
rect 4537 15385 4571 15419
rect 5089 15385 5123 15419
rect 5825 15385 5859 15419
rect 6285 15385 6319 15419
rect 22753 15385 22787 15419
rect 5549 15317 5583 15351
rect 6653 15317 6687 15351
rect 6837 15317 6871 15351
rect 8033 15317 8067 15351
rect 12817 15317 12851 15351
rect 13369 15317 13403 15351
rect 13737 15317 13771 15351
rect 21465 15317 21499 15351
rect 23121 15317 23155 15351
rect 23489 15317 23523 15351
rect 24133 15317 24167 15351
rect 1777 15113 1811 15147
rect 3157 15113 3191 15147
rect 3709 15113 3743 15147
rect 5917 15113 5951 15147
rect 10701 15113 10735 15147
rect 11713 15113 11747 15147
rect 12817 15113 12851 15147
rect 13001 15113 13035 15147
rect 22385 15113 22419 15147
rect 23673 15113 23707 15147
rect 1685 15045 1719 15079
rect 3617 15045 3651 15079
rect 12081 15045 12115 15079
rect 24133 15045 24167 15079
rect 2387 14977 2421 15011
rect 5147 14977 5181 15011
rect 6929 14977 6963 15011
rect 7782 14977 7816 15011
rect 9689 14977 9723 15011
rect 9963 14977 9997 15011
rect 11989 14977 12023 15011
rect 12495 14977 12529 15011
rect 14381 14977 14415 15011
rect 18245 14977 18279 15011
rect 18501 14977 18535 15011
rect 22569 14977 22603 15011
rect 22919 15007 22953 15041
rect 2145 14909 2179 14943
rect 4905 14909 4939 14943
rect 6745 14909 6779 14943
rect 7389 14909 7423 14943
rect 7665 14909 7699 14943
rect 7941 14909 7975 14943
rect 14197 14909 14231 14943
rect 15117 14909 15151 14943
rect 15234 14909 15268 14943
rect 15393 14909 15427 14943
rect 22661 14909 22695 14943
rect 14841 14841 14875 14875
rect 8585 14773 8619 14807
rect 16037 14773 16071 14807
rect 19625 14773 19659 14807
rect 24409 14773 24443 14807
rect 1593 14569 1627 14603
rect 3065 14569 3099 14603
rect 6561 14569 6595 14603
rect 8033 14569 8067 14603
rect 11805 14569 11839 14603
rect 15117 14569 15151 14603
rect 16497 14569 16531 14603
rect 24225 14569 24259 14603
rect 4169 14501 4203 14535
rect 5549 14433 5583 14467
rect 7021 14433 7055 14467
rect 14105 14433 14139 14467
rect 15485 14433 15519 14467
rect 20729 14433 20763 14467
rect 22845 14433 22879 14467
rect 1501 14365 1535 14399
rect 2237 14365 2271 14399
rect 3617 14365 3651 14399
rect 5791 14365 5825 14399
rect 7263 14365 7297 14399
rect 10793 14365 10827 14399
rect 11067 14365 11101 14399
rect 14347 14365 14381 14399
rect 15743 14335 15777 14369
rect 18889 14365 18923 14399
rect 19349 14365 19383 14399
rect 19993 14365 20027 14399
rect 20996 14365 21030 14399
rect 22201 14365 22235 14399
rect 22661 14365 22695 14399
rect 2421 14297 2455 14331
rect 2973 14297 3007 14331
rect 3893 14297 3927 14331
rect 23112 14297 23146 14331
rect 2053 14229 2087 14263
rect 2513 14229 2547 14263
rect 3433 14229 3467 14263
rect 4537 14229 4571 14263
rect 18705 14229 18739 14263
rect 19441 14229 19475 14263
rect 19809 14229 19843 14263
rect 22109 14229 22143 14263
rect 22293 14229 22327 14263
rect 22477 14229 22511 14263
rect 1777 14025 1811 14059
rect 9413 14025 9447 14059
rect 9965 14025 9999 14059
rect 21281 14025 21315 14059
rect 1685 13957 1719 13991
rect 2237 13957 2271 13991
rect 2697 13889 2731 13923
rect 2971 13889 3005 13923
rect 4335 13919 4369 13953
rect 8401 13889 8435 13923
rect 8675 13889 8709 13923
rect 9781 13889 9815 13923
rect 12999 13889 13033 13923
rect 15209 13889 15243 13923
rect 15451 13889 15485 13923
rect 16681 13889 16715 13923
rect 16955 13889 16989 13923
rect 18061 13889 18095 13923
rect 18335 13889 18369 13923
rect 19683 13889 19717 13923
rect 21465 13889 21499 13923
rect 22107 13889 22141 13923
rect 23397 13889 23431 13923
rect 23673 13889 23707 13923
rect 24133 13889 24167 13923
rect 4077 13821 4111 13855
rect 12725 13821 12759 13855
rect 19441 13821 19475 13855
rect 21833 13821 21867 13855
rect 24041 13753 24075 13787
rect 2329 13685 2363 13719
rect 3709 13685 3743 13719
rect 5089 13685 5123 13719
rect 13737 13685 13771 13719
rect 16221 13685 16255 13719
rect 17693 13685 17727 13719
rect 19073 13685 19107 13719
rect 20453 13685 20487 13719
rect 22845 13685 22879 13719
rect 1777 13481 1811 13515
rect 5917 13481 5951 13515
rect 10793 13481 10827 13515
rect 17509 13481 17543 13515
rect 19809 13481 19843 13515
rect 22293 13481 22327 13515
rect 23029 13481 23063 13515
rect 4445 13413 4479 13447
rect 8493 13413 8527 13447
rect 9597 13413 9631 13447
rect 16313 13413 16347 13447
rect 23397 13413 23431 13447
rect 2237 13345 2271 13379
rect 3801 13345 3835 13379
rect 4721 13345 4755 13379
rect 4838 13345 4872 13379
rect 4997 13345 5031 13379
rect 7481 13345 7515 13379
rect 9137 13345 9171 13379
rect 9990 13345 10024 13379
rect 10149 13345 10183 13379
rect 10885 13345 10919 13379
rect 12265 13345 12299 13379
rect 15669 13345 15703 13379
rect 16706 13345 16740 13379
rect 16865 13345 16899 13379
rect 18061 13345 18095 13379
rect 18705 13345 18739 13379
rect 19993 13345 20027 13379
rect 20177 13345 20211 13379
rect 22477 13345 22511 13379
rect 1685 13277 1719 13311
rect 2511 13277 2545 13311
rect 3985 13277 4019 13311
rect 5825 13277 5859 13311
rect 7755 13277 7789 13311
rect 8953 13277 8987 13311
rect 9873 13277 9907 13311
rect 11159 13267 11193 13301
rect 12539 13277 12573 13311
rect 15853 13277 15887 13311
rect 16589 13277 16623 13311
rect 18153 13277 18187 13311
rect 18613 13277 18647 13311
rect 18889 13277 18923 13311
rect 19073 13277 19107 13311
rect 19717 13277 19751 13311
rect 20085 13277 20119 13311
rect 20269 13277 20303 13311
rect 22201 13277 22235 13311
rect 22845 13253 22879 13287
rect 22943 13277 22977 13311
rect 23121 13277 23155 13311
rect 23213 13277 23247 13311
rect 23673 13277 23707 13311
rect 18429 13209 18463 13243
rect 18521 13209 18555 13243
rect 18981 13209 19015 13243
rect 24041 13209 24075 13243
rect 3249 13141 3283 13175
rect 5641 13141 5675 13175
rect 11897 13141 11931 13175
rect 13277 13141 13311 13175
rect 19993 13141 20027 13175
rect 22477 13141 22511 13175
rect 22661 13141 22695 13175
rect 1685 12937 1719 12971
rect 4169 12937 4203 12971
rect 19441 12937 19475 12971
rect 24409 12937 24443 12971
rect 14473 12869 14507 12903
rect 24133 12869 24167 12903
rect 1593 12801 1627 12835
rect 3090 12801 3124 12835
rect 4077 12801 4111 12835
rect 5147 12801 5181 12835
rect 6651 12801 6685 12835
rect 9597 12801 9631 12835
rect 11253 12801 11287 12835
rect 11529 12801 11563 12835
rect 13553 12801 13587 12835
rect 13670 12801 13704 12835
rect 13829 12801 13863 12835
rect 14565 12801 14599 12835
rect 14807 12801 14841 12835
rect 17877 12801 17911 12835
rect 18236 12801 18270 12835
rect 19625 12801 19659 12835
rect 20913 12801 20947 12835
rect 21189 12801 21223 12835
rect 21373 12801 21407 12835
rect 21649 12801 21683 12835
rect 23581 12801 23615 12835
rect 2053 12733 2087 12767
rect 2237 12733 2271 12767
rect 2973 12733 3007 12767
rect 3249 12733 3283 12767
rect 4905 12733 4939 12767
rect 6377 12733 6411 12767
rect 9413 12733 9447 12767
rect 10333 12733 10367 12767
rect 10450 12733 10484 12767
rect 10609 12733 10643 12767
rect 12633 12733 12667 12767
rect 12817 12733 12851 12767
rect 13277 12733 13311 12767
rect 17969 12733 18003 12767
rect 2697 12665 2731 12699
rect 10057 12665 10091 12699
rect 17693 12665 17727 12699
rect 19349 12665 19383 12699
rect 21465 12665 21499 12699
rect 3893 12597 3927 12631
rect 5917 12597 5951 12631
rect 7389 12597 7423 12631
rect 11713 12597 11747 12631
rect 15577 12597 15611 12631
rect 21005 12597 21039 12631
rect 21281 12597 21315 12631
rect 23857 12597 23891 12631
rect 1409 12393 1443 12427
rect 2697 12393 2731 12427
rect 8769 12393 8803 12427
rect 15577 12393 15611 12427
rect 20453 12393 20487 12427
rect 22661 12393 22695 12427
rect 5641 12325 5675 12359
rect 7573 12325 7607 12359
rect 10793 12325 10827 12359
rect 17049 12325 17083 12359
rect 1685 12257 1719 12291
rect 5181 12257 5215 12291
rect 6034 12257 6068 12291
rect 6193 12257 6227 12291
rect 7113 12257 7147 12291
rect 9781 12257 9815 12291
rect 16589 12257 16623 12291
rect 17325 12257 17359 12291
rect 17601 12257 17635 12291
rect 20821 12257 20855 12291
rect 1593 12189 1627 12223
rect 1959 12189 1993 12223
rect 3893 12189 3927 12223
rect 4997 12189 5031 12223
rect 5917 12189 5951 12223
rect 6929 12189 6963 12223
rect 7849 12189 7883 12223
rect 7966 12189 8000 12223
rect 8125 12189 8159 12223
rect 10055 12189 10089 12223
rect 11713 12189 11747 12223
rect 12081 12189 12115 12223
rect 14657 12189 14691 12223
rect 16405 12189 16439 12223
rect 17463 12189 17497 12223
rect 19441 12189 19475 12223
rect 19715 12189 19749 12223
rect 22845 12189 22879 12223
rect 23103 12159 23137 12193
rect 3157 12121 3191 12155
rect 11621 12121 11655 12155
rect 14565 12121 14599 12155
rect 15025 12121 15059 12155
rect 21088 12121 21122 12155
rect 22569 12121 22603 12155
rect 3249 12053 3283 12087
rect 3985 12053 4019 12087
rect 6837 12053 6871 12087
rect 11345 12053 11379 12087
rect 12449 12053 12483 12087
rect 12633 12053 12667 12087
rect 14289 12053 14323 12087
rect 15393 12053 15427 12087
rect 18245 12053 18279 12087
rect 22201 12053 22235 12087
rect 23857 12053 23891 12087
rect 3433 11849 3467 11883
rect 7849 11849 7883 11883
rect 9229 11849 9263 11883
rect 10701 11849 10735 11883
rect 14381 11849 14415 11883
rect 21833 11849 21867 11883
rect 22385 11849 22419 11883
rect 24409 11849 24443 11883
rect 1501 11713 1535 11747
rect 2295 11713 2329 11747
rect 3617 11713 3651 11747
rect 3983 11713 4017 11747
rect 7095 11743 7129 11777
rect 8459 11713 8493 11747
rect 9931 11713 9965 11747
rect 13369 11713 13403 11747
rect 13643 11713 13677 11747
rect 16923 11713 16957 11747
rect 18335 11713 18369 11747
rect 20729 11713 20763 11747
rect 21005 11713 21039 11747
rect 21373 11713 21407 11747
rect 22017 11713 22051 11747
rect 22569 11713 22603 11747
rect 22935 11713 22969 11747
rect 24225 11713 24259 11747
rect 1777 11645 1811 11679
rect 2053 11645 2087 11679
rect 3709 11645 3743 11679
rect 6837 11645 6871 11679
rect 8217 11645 8251 11679
rect 9689 11645 9723 11679
rect 16681 11645 16715 11679
rect 18061 11645 18095 11679
rect 22661 11645 22695 11679
rect 17693 11577 17727 11611
rect 19073 11577 19107 11611
rect 21373 11577 21407 11611
rect 3065 11509 3099 11543
rect 4721 11509 4755 11543
rect 23673 11509 23707 11543
rect 10149 11305 10183 11339
rect 17049 11305 17083 11339
rect 18153 11305 18187 11339
rect 22201 11305 22235 11339
rect 2421 11237 2455 11271
rect 4537 11237 4571 11271
rect 2835 11169 2869 11203
rect 3617 11169 3651 11203
rect 4813 11169 4847 11203
rect 4951 11169 4985 11203
rect 11713 11169 11747 11203
rect 15853 11169 15887 11203
rect 16405 11169 16439 11203
rect 1593 11101 1627 11135
rect 1777 11101 1811 11135
rect 1961 11101 1995 11135
rect 2697 11101 2731 11135
rect 2973 11101 3007 11135
rect 3893 11101 3927 11135
rect 4077 11101 4111 11135
rect 5089 11101 5123 11135
rect 9137 11101 9171 11135
rect 9395 11071 9429 11105
rect 11987 11101 12021 11135
rect 15209 11101 15243 11135
rect 15393 11101 15427 11135
rect 16129 11101 16163 11135
rect 16246 11101 16280 11135
rect 17141 11101 17175 11135
rect 17383 11101 17417 11135
rect 19257 11101 19291 11135
rect 19531 11101 19565 11135
rect 22385 11101 22419 11135
rect 22661 11101 22695 11135
rect 22753 11101 22787 11135
rect 23027 11101 23061 11135
rect 5733 11033 5767 11067
rect 1409 10965 1443 10999
rect 12725 10965 12759 10999
rect 20269 10965 20303 10999
rect 22477 10965 22511 10999
rect 23765 10965 23799 10999
rect 1961 10761 1995 10795
rect 3433 10761 3467 10795
rect 5273 10761 5307 10795
rect 5641 10761 5675 10795
rect 13001 10761 13035 10795
rect 15025 10761 15059 10795
rect 16221 10761 16255 10795
rect 1501 10693 1535 10727
rect 11713 10693 11747 10727
rect 11989 10693 12023 10727
rect 12081 10693 12115 10727
rect 12449 10693 12483 10727
rect 12817 10693 12851 10727
rect 13737 10693 13771 10727
rect 14841 10693 14875 10727
rect 19165 10693 19199 10727
rect 19257 10693 19291 10727
rect 19441 10693 19475 10727
rect 23581 10693 23615 10727
rect 24133 10693 24167 10727
rect 2145 10625 2179 10659
rect 2695 10625 2729 10659
rect 3985 10625 4019 10659
rect 4261 10625 4295 10659
rect 4519 10655 4553 10689
rect 5825 10625 5859 10659
rect 6377 10625 6411 10659
rect 7435 10625 7469 10659
rect 7573 10625 7607 10659
rect 10057 10625 10091 10659
rect 10331 10625 10365 10659
rect 14013 10625 14047 10659
rect 14105 10625 14139 10659
rect 14473 10625 14507 10659
rect 15467 10625 15501 10659
rect 18889 10625 18923 10659
rect 19073 10625 19107 10659
rect 19349 10625 19383 10659
rect 19533 10625 19567 10659
rect 19625 10625 19659 10659
rect 19883 10655 19917 10689
rect 22385 10625 22419 10659
rect 22661 10625 22695 10659
rect 23213 10625 23247 10659
rect 24501 10625 24535 10659
rect 2421 10557 2455 10591
rect 6561 10557 6595 10591
rect 7297 10557 7331 10591
rect 15209 10557 15243 10591
rect 22017 10557 22051 10591
rect 7021 10489 7055 10523
rect 11069 10489 11103 10523
rect 22661 10489 22695 10523
rect 1593 10421 1627 10455
rect 3801 10421 3835 10455
rect 8217 10421 8251 10455
rect 20637 10421 20671 10455
rect 23029 10421 23063 10455
rect 23857 10421 23891 10455
rect 3249 10217 3283 10251
rect 5549 10217 5583 10251
rect 6929 10217 6963 10251
rect 10793 10217 10827 10251
rect 13645 10217 13679 10251
rect 15117 10217 15151 10251
rect 18797 10217 18831 10251
rect 19533 10217 19567 10251
rect 22385 10217 22419 10251
rect 22661 10217 22695 10251
rect 1685 10149 1719 10183
rect 19257 10149 19291 10183
rect 21925 10149 21959 10183
rect 2329 10081 2363 10115
rect 4537 10081 4571 10115
rect 9137 10081 9171 10115
rect 9597 10081 9631 10115
rect 9873 10081 9907 10115
rect 10011 10081 10045 10115
rect 12633 10081 12667 10115
rect 14105 10081 14139 10115
rect 1501 10013 1535 10047
rect 3157 10013 3191 10047
rect 4811 10013 4845 10047
rect 5917 10013 5951 10047
rect 6175 9983 6209 10017
rect 8953 10013 8987 10047
rect 10149 10013 10183 10047
rect 10977 10013 11011 10047
rect 11251 10013 11285 10047
rect 12875 10013 12909 10047
rect 14363 10013 14397 10047
rect 18705 10013 18739 10047
rect 19441 10013 19475 10047
rect 19717 10013 19751 10047
rect 20913 10013 20947 10047
rect 21155 10013 21189 10047
rect 22293 10013 22327 10047
rect 22569 10013 22603 10047
rect 22753 10013 22787 10047
rect 22845 10013 22879 10047
rect 23103 9983 23137 10017
rect 2053 9945 2087 9979
rect 2605 9945 2639 9979
rect 3893 9945 3927 9979
rect 2881 9877 2915 9911
rect 3985 9877 4019 9911
rect 11989 9877 12023 9911
rect 23857 9877 23891 9911
rect 1777 9673 1811 9707
rect 2329 9673 2363 9707
rect 3249 9673 3283 9707
rect 8309 9673 8343 9707
rect 9689 9673 9723 9707
rect 13001 9673 13035 9707
rect 19441 9673 19475 9707
rect 21465 9673 21499 9707
rect 23213 9673 23247 9707
rect 2789 9605 2823 9639
rect 3157 9605 3191 9639
rect 11713 9605 11747 9639
rect 11989 9605 12023 9639
rect 12817 9605 12851 9639
rect 18328 9605 18362 9639
rect 24133 9605 24167 9639
rect 24501 9605 24535 9639
rect 1685 9537 1719 9571
rect 2237 9537 2271 9571
rect 3433 9537 3467 9571
rect 3525 9537 3559 9571
rect 3799 9537 3833 9571
rect 5089 9537 5123 9571
rect 5365 9537 5399 9571
rect 5641 9537 5675 9571
rect 5917 9537 5951 9571
rect 7555 9567 7589 9601
rect 8951 9537 8985 9571
rect 12081 9537 12115 9571
rect 12449 9537 12483 9571
rect 16955 9537 16989 9571
rect 19775 9537 19809 9571
rect 21649 9537 21683 9571
rect 22100 9537 22134 9571
rect 23581 9537 23615 9571
rect 23949 9537 23983 9571
rect 7297 9469 7331 9503
rect 8677 9469 8711 9503
rect 16681 9469 16715 9503
rect 18061 9469 18095 9503
rect 19533 9469 19567 9503
rect 21833 9469 21867 9503
rect 4905 9401 4939 9435
rect 5457 9401 5491 9435
rect 4537 9333 4571 9367
rect 5181 9333 5215 9367
rect 5733 9333 5767 9367
rect 17693 9333 17727 9367
rect 20545 9333 20579 9367
rect 1501 9129 1535 9163
rect 5641 9129 5675 9163
rect 12909 9129 12943 9163
rect 4445 9061 4479 9095
rect 7389 9061 7423 9095
rect 9965 9061 9999 9095
rect 21005 9061 21039 9095
rect 23949 9061 23983 9095
rect 1777 8993 1811 9027
rect 4859 8993 4893 9027
rect 6929 8993 6963 9027
rect 7665 8993 7699 9027
rect 7803 8993 7837 9027
rect 9321 8993 9355 9027
rect 10241 8993 10275 9027
rect 16681 8993 16715 9027
rect 17141 8993 17175 9027
rect 18337 8993 18371 9027
rect 19993 8993 20027 9027
rect 21465 8993 21499 9027
rect 1685 8925 1719 8959
rect 2051 8925 2085 8959
rect 3249 8925 3283 8959
rect 3801 8925 3835 8959
rect 3985 8925 4019 8959
rect 4721 8925 4755 8959
rect 4997 8925 5031 8959
rect 6745 8925 6779 8959
rect 7941 8925 7975 8959
rect 9505 8925 9539 8959
rect 10379 8925 10413 8959
rect 10517 8925 10551 8959
rect 11897 8925 11931 8959
rect 12171 8925 12205 8959
rect 15117 8925 15151 8959
rect 15375 8925 15409 8959
rect 16497 8925 16531 8959
rect 17417 8925 17451 8959
rect 17534 8925 17568 8959
rect 17693 8925 17727 8959
rect 19901 8925 19935 8959
rect 20361 8925 20395 8959
rect 20545 8925 20579 8959
rect 21097 8925 21131 8959
rect 21373 8925 21407 8959
rect 21557 8925 21591 8959
rect 21833 8925 21867 8959
rect 23029 8925 23063 8959
rect 23305 8925 23339 8959
rect 23489 8925 23523 8959
rect 24041 8925 24075 8959
rect 2789 8789 2823 8823
rect 3341 8789 3375 8823
rect 8585 8789 8619 8823
rect 11161 8789 11195 8823
rect 16129 8789 16163 8823
rect 21649 8789 21683 8823
rect 22845 8789 22879 8823
rect 3893 8585 3927 8619
rect 5089 8585 5123 8619
rect 8125 8585 8159 8619
rect 10517 8585 10551 8619
rect 12173 8585 12207 8619
rect 17693 8585 17727 8619
rect 21465 8585 21499 8619
rect 22937 8585 22971 8619
rect 1961 8517 1995 8551
rect 12449 8517 12483 8551
rect 12909 8517 12943 8551
rect 13277 8517 13311 8551
rect 13829 8517 13863 8551
rect 14565 8517 14599 8551
rect 14933 8517 14967 8551
rect 1593 8449 1627 8483
rect 3249 8449 3283 8483
rect 4319 8449 4353 8483
rect 7371 8479 7405 8513
rect 9747 8449 9781 8483
rect 12541 8449 12575 8483
rect 14105 8449 14139 8483
rect 14197 8449 14231 8483
rect 16681 8449 16715 8483
rect 16939 8449 16973 8483
rect 20085 8449 20119 8483
rect 20352 8449 20386 8483
rect 22845 8449 22879 8483
rect 23377 8449 23411 8483
rect 2053 8381 2087 8415
rect 2237 8381 2271 8415
rect 2697 8381 2731 8415
rect 2973 8381 3007 8415
rect 3111 8381 3145 8415
rect 4077 8381 4111 8415
rect 7113 8381 7147 8415
rect 9505 8381 9539 8415
rect 23121 8381 23155 8415
rect 13461 8313 13495 8347
rect 15117 8313 15151 8347
rect 24501 8245 24535 8279
rect 1593 8041 1627 8075
rect 1961 8041 1995 8075
rect 3249 8041 3283 8075
rect 8401 8041 8435 8075
rect 9965 8041 9999 8075
rect 23305 8041 23339 8075
rect 23949 8041 23983 8075
rect 3801 7973 3835 8007
rect 5089 7973 5123 8007
rect 6101 7973 6135 8007
rect 7297 7973 7331 8007
rect 16037 7973 16071 8007
rect 20177 7973 20211 8007
rect 23673 7973 23707 8007
rect 2237 7905 2271 7939
rect 4077 7905 4111 7939
rect 6377 7905 6411 7939
rect 6494 7905 6528 7939
rect 6653 7905 6687 7939
rect 15577 7905 15611 7939
rect 16313 7905 16347 7939
rect 16430 7905 16464 7939
rect 20637 7905 20671 7939
rect 20913 7905 20947 7939
rect 22293 7905 22327 7939
rect 2145 7837 2179 7871
rect 2511 7837 2545 7871
rect 3985 7837 4019 7871
rect 4351 7837 4385 7871
rect 5457 7837 5491 7871
rect 5641 7837 5675 7871
rect 7389 7837 7423 7871
rect 7663 7837 7697 7871
rect 8953 7837 8987 7871
rect 9227 7837 9261 7871
rect 10793 7837 10827 7871
rect 11067 7837 11101 7871
rect 15393 7837 15427 7871
rect 16589 7837 16623 7871
rect 19533 7837 19567 7871
rect 19717 7837 19751 7871
rect 20269 7837 20303 7871
rect 20545 7837 20579 7871
rect 20729 7837 20763 7871
rect 21155 7837 21189 7871
rect 22567 7837 22601 7871
rect 23857 7837 23891 7871
rect 24133 7837 24167 7871
rect 1501 7769 1535 7803
rect 11805 7701 11839 7735
rect 17233 7701 17267 7735
rect 21925 7701 21959 7735
rect 3249 7497 3283 7531
rect 3801 7497 3835 7531
rect 7481 7497 7515 7531
rect 9413 7497 9447 7531
rect 13737 7497 13771 7531
rect 15117 7497 15151 7531
rect 17693 7497 17727 7531
rect 18705 7497 18739 7531
rect 19073 7497 19107 7531
rect 20637 7497 20671 7531
rect 21005 7497 21039 7531
rect 23305 7497 23339 7531
rect 23673 7497 23707 7531
rect 24041 7497 24075 7531
rect 24409 7497 24443 7531
rect 1869 7429 1903 7463
rect 2421 7429 2455 7463
rect 3157 7429 3191 7463
rect 19524 7429 19558 7463
rect 1501 7361 1535 7395
rect 2053 7361 2087 7395
rect 2605 7361 2639 7395
rect 3985 7361 4019 7395
rect 4261 7361 4295 7395
rect 4537 7361 4571 7395
rect 6711 7361 6745 7395
rect 9229 7361 9263 7395
rect 9781 7361 9815 7395
rect 10039 7391 10073 7425
rect 12983 7391 13017 7425
rect 14347 7361 14381 7395
rect 16939 7371 16973 7405
rect 18245 7361 18279 7395
rect 18613 7361 18647 7395
rect 18889 7361 18923 7395
rect 18981 7361 19015 7395
rect 19257 7361 19291 7395
rect 20913 7361 20947 7395
rect 21189 7361 21223 7395
rect 21649 7361 21683 7395
rect 21925 7361 21959 7395
rect 22201 7361 22235 7395
rect 22385 7361 22419 7395
rect 22753 7361 22787 7395
rect 23213 7361 23247 7395
rect 23489 7361 23523 7395
rect 23857 7361 23891 7395
rect 23949 7361 23983 7395
rect 24133 7361 24167 7395
rect 24225 7361 24259 7395
rect 6469 7293 6503 7327
rect 12725 7293 12759 7327
rect 14105 7293 14139 7327
rect 16681 7293 16715 7327
rect 18337 7293 18371 7327
rect 4077 7225 4111 7259
rect 4353 7225 4387 7259
rect 18245 7225 18279 7259
rect 21465 7225 21499 7259
rect 22569 7225 22603 7259
rect 2697 7157 2731 7191
rect 10793 7157 10827 7191
rect 20729 7157 20763 7191
rect 22017 7157 22051 7191
rect 22293 7157 22327 7191
rect 23029 7157 23063 7191
rect 1777 6953 1811 6987
rect 18705 6953 18739 6987
rect 18981 6953 19015 6987
rect 20269 6953 20303 6987
rect 21281 6953 21315 6987
rect 22937 6953 22971 6987
rect 24041 6885 24075 6919
rect 2513 6817 2547 6851
rect 3065 6817 3099 6851
rect 4169 6817 4203 6851
rect 8953 6817 8987 6851
rect 10701 6817 10735 6851
rect 11161 6817 11195 6851
rect 11437 6817 11471 6851
rect 12633 6817 12667 6851
rect 17233 6817 17267 6851
rect 21557 6817 21591 6851
rect 3433 6749 3467 6783
rect 3893 6749 3927 6783
rect 4537 6749 4571 6783
rect 4813 6749 4847 6783
rect 7205 6749 7239 6783
rect 7479 6749 7513 6783
rect 9211 6719 9245 6753
rect 10517 6749 10551 6783
rect 11554 6749 11588 6783
rect 11713 6749 11747 6783
rect 12875 6749 12909 6783
rect 17475 6749 17509 6783
rect 18613 6749 18647 6783
rect 18889 6749 18923 6783
rect 19073 6749 19107 6783
rect 19257 6749 19291 6783
rect 19531 6749 19565 6783
rect 21465 6749 21499 6783
rect 21813 6749 21847 6783
rect 23121 6749 23155 6783
rect 23489 6749 23523 6783
rect 23949 6749 23983 6783
rect 1685 6681 1719 6715
rect 2237 6681 2271 6715
rect 2789 6681 2823 6715
rect 3249 6613 3283 6647
rect 4353 6613 4387 6647
rect 4629 6613 4663 6647
rect 8217 6613 8251 6647
rect 9965 6613 9999 6647
rect 12357 6613 12391 6647
rect 13645 6613 13679 6647
rect 18245 6613 18279 6647
rect 1593 6409 1627 6443
rect 3433 6409 3467 6443
rect 9689 6409 9723 6443
rect 17325 6409 17359 6443
rect 19073 6409 19107 6443
rect 20729 6409 20763 6443
rect 24501 6409 24535 6443
rect 1501 6341 1535 6375
rect 2327 6273 2361 6307
rect 3617 6273 3651 6307
rect 3709 6273 3743 6307
rect 4629 6273 4663 6307
rect 4905 6273 4939 6307
rect 5549 6273 5583 6307
rect 5825 6273 5859 6307
rect 8907 6273 8941 6307
rect 9045 6273 9079 6307
rect 11529 6273 11563 6307
rect 12449 6273 12483 6307
rect 15007 6303 15041 6337
rect 17509 6273 17543 6307
rect 17601 6273 17635 6307
rect 17868 6273 17902 6307
rect 19257 6273 19291 6307
rect 20637 6273 20671 6307
rect 21097 6273 21131 6307
rect 21189 6273 21223 6307
rect 21465 6273 21499 6307
rect 22017 6273 22051 6307
rect 22201 6273 22235 6307
rect 22661 6273 22695 6307
rect 23377 6273 23411 6307
rect 2053 6205 2087 6239
rect 3893 6205 3927 6239
rect 4767 6205 4801 6239
rect 7849 6205 7883 6239
rect 8033 6205 8067 6239
rect 8493 6205 8527 6239
rect 8769 6205 8803 6239
rect 11713 6205 11747 6239
rect 12566 6205 12600 6239
rect 12725 6205 12759 6239
rect 14749 6205 14783 6239
rect 23121 6205 23155 6239
rect 4353 6137 4387 6171
rect 12173 6137 12207 6171
rect 18981 6137 19015 6171
rect 20913 6137 20947 6171
rect 21649 6137 21683 6171
rect 22661 6137 22695 6171
rect 3065 6069 3099 6103
rect 5641 6069 5675 6103
rect 13369 6069 13403 6103
rect 15761 6069 15795 6103
rect 21373 6069 21407 6103
rect 1501 5865 1535 5899
rect 3617 5865 3651 5899
rect 5089 5865 5123 5899
rect 7389 5865 7423 5899
rect 11897 5865 11931 5899
rect 13277 5865 13311 5899
rect 18153 5865 18187 5899
rect 20269 5865 20303 5899
rect 21189 5865 21223 5899
rect 21557 5865 21591 5899
rect 22293 5865 22327 5899
rect 23765 5865 23799 5899
rect 24225 5865 24259 5899
rect 15853 5797 15887 5831
rect 20729 5797 20763 5831
rect 21833 5797 21867 5831
rect 1777 5729 1811 5763
rect 1961 5729 1995 5763
rect 2421 5729 2455 5763
rect 2697 5729 2731 5763
rect 2835 5729 2869 5763
rect 2973 5729 3007 5763
rect 5733 5729 5767 5763
rect 6193 5729 6227 5763
rect 6586 5729 6620 5763
rect 6745 5729 6779 5763
rect 10885 5729 10919 5763
rect 12265 5729 12299 5763
rect 16129 5729 16163 5763
rect 16267 5729 16301 5763
rect 16405 5729 16439 5763
rect 17141 5729 17175 5763
rect 20913 5729 20947 5763
rect 1685 5661 1719 5695
rect 3985 5661 4019 5695
rect 4077 5661 4111 5695
rect 4351 5661 4385 5695
rect 5549 5661 5583 5695
rect 6469 5661 6503 5695
rect 9137 5661 9171 5695
rect 9379 5661 9413 5695
rect 11159 5661 11193 5695
rect 12523 5631 12557 5665
rect 15209 5661 15243 5695
rect 15393 5661 15427 5695
rect 17415 5661 17449 5695
rect 20453 5661 20487 5695
rect 20729 5661 20763 5695
rect 21373 5661 21407 5695
rect 21465 5661 21499 5695
rect 21649 5661 21683 5695
rect 21741 5661 21775 5695
rect 22109 5661 22143 5695
rect 22385 5661 22419 5695
rect 22659 5661 22693 5695
rect 23949 5661 23983 5695
rect 24041 5661 24075 5695
rect 21097 5593 21131 5627
rect 3801 5525 3835 5559
rect 10149 5525 10183 5559
rect 17049 5525 17083 5559
rect 23397 5525 23431 5559
rect 1593 5321 1627 5355
rect 2145 5321 2179 5355
rect 2881 5321 2915 5355
rect 4353 5321 4387 5355
rect 5917 5321 5951 5355
rect 7389 5321 7423 5355
rect 21373 5321 21407 5355
rect 21833 5321 21867 5355
rect 22293 5321 22327 5355
rect 22569 5321 22603 5355
rect 22661 5321 22695 5355
rect 24409 5321 24443 5355
rect 2053 5253 2087 5287
rect 23765 5253 23799 5287
rect 1501 5185 1535 5219
rect 2605 5185 2639 5219
rect 3249 5185 3283 5219
rect 3615 5185 3649 5219
rect 5147 5185 5181 5219
rect 6619 5185 6653 5219
rect 9505 5185 9539 5219
rect 10563 5185 10597 5219
rect 12523 5215 12557 5249
rect 13645 5185 13679 5219
rect 14841 5185 14875 5219
rect 19039 5185 19073 5219
rect 20361 5185 20395 5219
rect 20729 5185 20763 5219
rect 21005 5185 21039 5219
rect 21189 5185 21223 5219
rect 21281 5185 21315 5219
rect 22017 5185 22051 5219
rect 22109 5185 22143 5219
rect 22385 5185 22419 5219
rect 22845 5185 22879 5219
rect 23121 5185 23155 5219
rect 23397 5185 23431 5219
rect 24041 5185 24075 5219
rect 24317 5185 24351 5219
rect 3341 5117 3375 5151
rect 4905 5117 4939 5151
rect 6377 5117 6411 5151
rect 9689 5117 9723 5151
rect 10149 5117 10183 5151
rect 10425 5117 10459 5151
rect 10701 5117 10735 5151
rect 12265 5117 12299 5151
rect 13829 5117 13863 5151
rect 14565 5117 14599 5151
rect 14703 5117 14737 5151
rect 18797 5117 18831 5151
rect 20177 5117 20211 5151
rect 21097 5117 21131 5151
rect 23213 5117 23247 5151
rect 13277 5049 13311 5083
rect 14289 5049 14323 5083
rect 19809 5049 19843 5083
rect 20361 5049 20395 5083
rect 23489 5049 23523 5083
rect 3065 4981 3099 5015
rect 11345 4981 11379 5015
rect 15485 4981 15519 5015
rect 22937 4981 22971 5015
rect 23857 4981 23891 5015
rect 1593 4777 1627 4811
rect 2513 4777 2547 4811
rect 2789 4777 2823 4811
rect 4721 4777 4755 4811
rect 11161 4777 11195 4811
rect 15117 4777 15151 4811
rect 18705 4777 18739 4811
rect 18889 4777 18923 4811
rect 19809 4777 19843 4811
rect 20085 4777 20119 4811
rect 22477 4777 22511 4811
rect 24041 4777 24075 4811
rect 19441 4709 19475 4743
rect 21925 4709 21959 4743
rect 10149 4641 10183 4675
rect 11621 4641 11655 4675
rect 14105 4641 14139 4675
rect 20545 4641 20579 4675
rect 23213 4641 23247 4675
rect 1501 4573 1535 4607
rect 2053 4573 2087 4607
rect 2697 4573 2731 4607
rect 2973 4573 3007 4607
rect 3249 4573 3283 4607
rect 3525 4573 3559 4607
rect 4905 4573 4939 4607
rect 7481 4573 7515 4607
rect 7755 4573 7789 4607
rect 10423 4573 10457 4607
rect 11879 4543 11913 4577
rect 14379 4573 14413 4607
rect 17233 4573 17267 4607
rect 17491 4543 17525 4577
rect 18613 4573 18647 4607
rect 19073 4573 19107 4607
rect 19625 4573 19659 4607
rect 19717 4573 19751 4607
rect 19993 4573 20027 4607
rect 20177 4573 20211 4607
rect 20453 4573 20487 4607
rect 22201 4573 22235 4607
rect 22293 4573 22327 4607
rect 22661 4573 22695 4607
rect 20812 4505 20846 4539
rect 23949 4505 23983 4539
rect 2145 4437 2179 4471
rect 3065 4437 3099 4471
rect 3341 4437 3375 4471
rect 8493 4437 8527 4471
rect 12633 4437 12667 4471
rect 18245 4437 18279 4471
rect 20269 4437 20303 4471
rect 22017 4437 22051 4471
rect 1593 4233 1627 4267
rect 5181 4233 5215 4267
rect 9413 4233 9447 4267
rect 12173 4233 12207 4267
rect 13277 4233 13311 4267
rect 13461 4233 13495 4267
rect 20545 4233 20579 4267
rect 1501 4165 1535 4199
rect 5365 4165 5399 4199
rect 12449 4165 12483 4199
rect 12541 4165 12575 4199
rect 12909 4165 12943 4199
rect 19432 4165 19466 4199
rect 21005 4165 21039 4199
rect 1961 4097 1995 4131
rect 2235 4097 2269 4131
rect 3341 4097 3375 4131
rect 3525 4097 3559 4131
rect 4399 4097 4433 4131
rect 7573 4097 7607 4131
rect 8769 4097 8803 4131
rect 14657 4097 14691 4131
rect 15694 4097 15728 4131
rect 17693 4097 17727 4131
rect 17877 4097 17911 4131
rect 18061 4097 18095 4131
rect 18521 4097 18555 4131
rect 19073 4097 19107 4131
rect 19165 4097 19199 4131
rect 20821 4097 20855 4131
rect 21465 4097 21499 4131
rect 22107 4097 22141 4131
rect 23213 4097 23247 4131
rect 23487 4097 23521 4131
rect 4261 4029 4295 4063
rect 4537 4029 4571 4063
rect 7757 4029 7791 4063
rect 8493 4029 8527 4063
rect 8631 4029 8665 4063
rect 14841 4029 14875 4063
rect 15577 4029 15611 4063
rect 15853 4029 15887 4063
rect 21833 4029 21867 4063
rect 2973 3961 3007 3995
rect 3985 3961 4019 3995
rect 5549 3961 5583 3995
rect 8217 3961 8251 3995
rect 13921 3961 13955 3995
rect 15301 3961 15335 3995
rect 17693 3961 17727 3995
rect 20637 3961 20671 3995
rect 16497 3893 16531 3927
rect 18889 3893 18923 3927
rect 21097 3893 21131 3927
rect 21557 3893 21591 3927
rect 22845 3893 22879 3927
rect 24225 3893 24259 3927
rect 1409 3689 1443 3723
rect 2697 3689 2731 3723
rect 4813 3689 4847 3723
rect 7113 3689 7147 3723
rect 15669 3689 15703 3723
rect 17049 3689 17083 3723
rect 18337 3689 18371 3723
rect 23949 3621 23983 3655
rect 6101 3553 6135 3587
rect 7481 3553 7515 3587
rect 9781 3553 9815 3587
rect 12449 3553 12483 3587
rect 14657 3553 14691 3587
rect 16037 3553 16071 3587
rect 18613 3553 18647 3587
rect 22201 3553 22235 3587
rect 23029 3553 23063 3587
rect 1593 3485 1627 3519
rect 1685 3485 1719 3519
rect 1959 3485 1993 3519
rect 3801 3485 3835 3519
rect 4075 3485 4109 3519
rect 6375 3485 6409 3519
rect 7755 3485 7789 3519
rect 9137 3485 9171 3519
rect 10055 3485 10089 3519
rect 11713 3485 11747 3519
rect 13369 3485 13403 3519
rect 13829 3485 13863 3519
rect 14931 3485 14965 3519
rect 16295 3455 16329 3489
rect 17693 3485 17727 3519
rect 17785 3485 17819 3519
rect 17969 3485 18003 3519
rect 18245 3485 18279 3519
rect 18429 3485 18463 3519
rect 18521 3485 18555 3519
rect 18981 3485 19015 3519
rect 19441 3485 19475 3519
rect 20269 3485 20303 3519
rect 21465 3485 21499 3519
rect 21649 3485 21683 3519
rect 22109 3485 22143 3519
rect 22661 3485 22695 3519
rect 23765 3485 23799 3519
rect 17877 3417 17911 3451
rect 19717 3417 19751 3451
rect 20821 3417 20855 3451
rect 8493 3349 8527 3383
rect 8953 3349 8987 3383
rect 10793 3349 10827 3383
rect 11529 3349 11563 3383
rect 13645 3349 13679 3383
rect 17509 3349 17543 3383
rect 18797 3349 18831 3383
rect 19257 3349 19291 3383
rect 19809 3349 19843 3383
rect 20361 3349 20395 3383
rect 20913 3349 20947 3383
rect 9413 3145 9447 3179
rect 9873 3145 9907 3179
rect 13277 3145 13311 3179
rect 17785 3145 17819 3179
rect 19441 3145 19475 3179
rect 19717 3145 19751 3179
rect 2973 3077 3007 3111
rect 4445 3077 4479 3111
rect 10149 3077 10183 3111
rect 10241 3077 10275 3111
rect 10609 3077 10643 3111
rect 10977 3077 11011 3111
rect 19625 3077 19659 3111
rect 20177 3077 20211 3111
rect 22845 3077 22879 3111
rect 23388 3077 23422 3111
rect 5163 3039 5197 3073
rect 6653 3009 6687 3043
rect 6929 3009 6963 3043
rect 7205 3009 7239 3043
rect 7481 3009 7515 3043
rect 7573 3009 7607 3043
rect 8493 3009 8527 3043
rect 8631 3009 8665 3043
rect 8769 3009 8803 3043
rect 11897 3009 11931 3043
rect 12173 3009 12207 3043
rect 12539 3009 12573 3043
rect 16313 3009 16347 3043
rect 16497 3009 16531 3043
rect 16865 3009 16899 3043
rect 17141 3009 17175 3043
rect 17417 3009 17451 3043
rect 17693 3009 17727 3043
rect 17969 3009 18003 3043
rect 18328 3009 18362 3043
rect 20821 3009 20855 3043
rect 22201 3009 22235 3043
rect 3157 2941 3191 2975
rect 4629 2941 4663 2975
rect 4905 2941 4939 2975
rect 7757 2941 7791 2975
rect 12265 2941 12299 2975
rect 18061 2941 18095 2975
rect 21005 2941 21039 2975
rect 23121 2941 23155 2975
rect 8217 2873 8251 2907
rect 11161 2873 11195 2907
rect 5917 2805 5951 2839
rect 6469 2805 6503 2839
rect 6745 2805 6779 2839
rect 7021 2805 7055 2839
rect 7297 2805 7331 2839
rect 11713 2805 11747 2839
rect 11989 2805 12023 2839
rect 16405 2805 16439 2839
rect 16681 2805 16715 2839
rect 16957 2805 16991 2839
rect 17233 2805 17267 2839
rect 17509 2805 17543 2839
rect 20269 2805 20303 2839
rect 24501 2805 24535 2839
rect 1961 2601 1995 2635
rect 2697 2601 2731 2635
rect 4905 2601 4939 2635
rect 5181 2601 5215 2635
rect 6745 2601 6779 2635
rect 7941 2601 7975 2635
rect 9413 2601 9447 2635
rect 11253 2601 11287 2635
rect 17141 2601 17175 2635
rect 18337 2601 18371 2635
rect 19257 2601 19291 2635
rect 19947 2601 19981 2635
rect 21925 2601 21959 2635
rect 24133 2601 24167 2635
rect 1593 2533 1627 2567
rect 8953 2533 8987 2567
rect 15301 2533 15335 2567
rect 23857 2533 23891 2567
rect 10241 2465 10275 2499
rect 19763 2465 19797 2499
rect 22477 2465 22511 2499
rect 1409 2397 1443 2431
rect 1777 2397 1811 2431
rect 2513 2397 2547 2431
rect 4629 2397 4663 2431
rect 4721 2397 4755 2431
rect 4997 2397 5031 2431
rect 5733 2397 5767 2431
rect 6929 2397 6963 2431
rect 7203 2397 7237 2431
rect 8493 2397 8527 2431
rect 8769 2397 8803 2431
rect 9137 2397 9171 2431
rect 9781 2397 9815 2431
rect 9873 2397 9907 2431
rect 10483 2397 10517 2431
rect 11989 2397 12023 2431
rect 12265 2397 12299 2431
rect 12541 2397 12575 2431
rect 12909 2397 12943 2431
rect 13277 2397 13311 2431
rect 13553 2397 13587 2431
rect 13829 2397 13863 2431
rect 14841 2397 14875 2431
rect 15117 2397 15151 2431
rect 15485 2397 15519 2431
rect 15761 2397 15795 2431
rect 16037 2397 16071 2431
rect 16405 2397 16439 2431
rect 16865 2397 16899 2431
rect 17509 2397 17543 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 24041 2397 24075 2431
rect 5825 2329 5859 2363
rect 6193 2329 6227 2363
rect 6561 2329 6595 2363
rect 9321 2329 9355 2363
rect 17049 2329 17083 2363
rect 17693 2329 17727 2363
rect 18245 2329 18279 2363
rect 20637 2329 20671 2363
rect 22722 2329 22756 2363
rect 4445 2261 4479 2295
rect 5457 2261 5491 2295
rect 8309 2261 8343 2295
rect 8585 2261 8619 2295
rect 9597 2261 9631 2295
rect 10057 2261 10091 2295
rect 11805 2261 11839 2295
rect 12081 2261 12115 2295
rect 12357 2261 12391 2295
rect 12725 2261 12759 2295
rect 13093 2261 13127 2295
rect 13369 2261 13403 2295
rect 13645 2261 13679 2295
rect 14657 2261 14691 2295
rect 14933 2261 14967 2295
rect 15577 2261 15611 2295
rect 15853 2261 15887 2295
rect 16681 2261 16715 2295
rect 17325 2261 17359 2295
rect 17785 2261 17819 2295
rect 18705 2261 18739 2295
rect 2145 2057 2179 2091
rect 3249 2057 3283 2091
rect 3801 2057 3835 2091
rect 4077 2057 4111 2091
rect 4445 2057 4479 2091
rect 4721 2057 4755 2091
rect 5917 2057 5951 2091
rect 6653 2057 6687 2091
rect 7021 2057 7055 2091
rect 7757 2057 7791 2091
rect 8125 2057 8159 2091
rect 8493 2057 8527 2091
rect 8861 2057 8895 2091
rect 10057 2057 10091 2091
rect 19441 2057 19475 2091
rect 23121 2057 23155 2091
rect 23857 2057 23891 2091
rect 1685 1989 1719 2023
rect 6561 1989 6595 2023
rect 6929 1989 6963 2023
rect 7665 1989 7699 2023
rect 8033 1989 8067 2023
rect 8769 1989 8803 2023
rect 10977 1989 11011 2023
rect 11805 1989 11839 2023
rect 15669 1989 15703 2023
rect 16773 1989 16807 2023
rect 17877 1989 17911 2023
rect 18429 1989 18463 2023
rect 18981 1989 19015 2023
rect 1501 1921 1535 1955
rect 1869 1921 1903 1955
rect 2421 1921 2455 1955
rect 2789 1921 2823 1955
rect 3065 1921 3099 1955
rect 3525 1921 3559 1955
rect 3617 1921 3651 1955
rect 3985 1921 4019 1955
rect 4261 1921 4295 1955
rect 4629 1921 4663 1955
rect 4905 1921 4939 1955
rect 5179 1921 5213 1955
rect 7205 1921 7239 1955
rect 8401 1921 8435 1955
rect 9045 1921 9079 1955
rect 9303 1951 9337 1985
rect 10517 1921 10551 1955
rect 12357 1921 12391 1955
rect 13093 1921 13127 1955
rect 13553 1921 13587 1955
rect 13829 1921 13863 1955
rect 14289 1921 14323 1955
rect 14473 1921 14507 1955
rect 14841 1921 14875 1955
rect 15393 1921 15427 1955
rect 16129 1921 16163 1955
rect 17325 1921 17359 1955
rect 17693 1921 17727 1955
rect 19625 1921 19659 1955
rect 19993 1921 20027 1955
rect 20729 1921 20763 1955
rect 21833 1921 21867 1955
rect 24041 1921 24075 1955
rect 24317 1921 24351 1955
rect 19717 1853 19751 1887
rect 21005 1853 21039 1887
rect 2605 1785 2639 1819
rect 2973 1785 3007 1819
rect 7389 1785 7423 1819
rect 10701 1785 10735 1819
rect 11161 1785 11195 1819
rect 11989 1785 12023 1819
rect 15209 1785 15243 1819
rect 24133 1785 24167 1819
rect 3341 1717 3375 1751
rect 12633 1717 12667 1751
rect 13369 1717 13403 1751
rect 13645 1717 13679 1751
rect 14105 1717 14139 1751
rect 14657 1717 14691 1751
rect 15025 1717 15059 1751
rect 15761 1717 15795 1751
rect 16313 1717 16347 1751
rect 16865 1717 16899 1751
rect 17969 1717 18003 1751
rect 18521 1717 18555 1751
rect 19073 1717 19107 1751
rect 10701 1513 10735 1547
rect 12725 1513 12759 1547
rect 14289 1513 14323 1547
rect 15393 1513 15427 1547
rect 15945 1513 15979 1547
rect 16313 1513 16347 1547
rect 16865 1513 16899 1547
rect 17417 1513 17451 1547
rect 23765 1445 23799 1479
rect 10333 1377 10367 1411
rect 1777 1309 1811 1343
rect 2145 1309 2179 1343
rect 2237 1309 2271 1343
rect 2513 1309 2547 1343
rect 3433 1309 3467 1343
rect 4077 1309 4111 1343
rect 4169 1309 4203 1343
rect 4445 1309 4479 1343
rect 5273 1309 5307 1343
rect 5917 1309 5951 1343
rect 6561 1309 6595 1343
rect 6745 1309 6779 1343
rect 7021 1309 7055 1343
rect 8493 1309 8527 1343
rect 8769 1309 8803 1343
rect 9137 1309 9171 1343
rect 9597 1309 9631 1343
rect 10609 1309 10643 1343
rect 11069 1309 11103 1343
rect 11529 1309 11563 1343
rect 12081 1309 12115 1343
rect 12357 1309 12391 1343
rect 12633 1309 12667 1343
rect 13277 1309 13311 1343
rect 13645 1309 13679 1343
rect 14657 1309 14691 1343
rect 15301 1309 15335 1343
rect 16497 1309 16531 1343
rect 16773 1309 16807 1343
rect 17325 1309 17359 1343
rect 17877 1309 17911 1343
rect 18521 1309 18555 1343
rect 19073 1309 19107 1343
rect 19441 1309 19475 1343
rect 20177 1309 20211 1343
rect 20453 1309 20487 1343
rect 22017 1309 22051 1343
rect 22109 1309 22143 1343
rect 1593 1241 1627 1275
rect 1961 1241 1995 1275
rect 3249 1241 3283 1275
rect 5457 1241 5491 1275
rect 7481 1241 7515 1275
rect 7849 1241 7883 1275
rect 9321 1241 9355 1275
rect 9505 1241 9539 1275
rect 10057 1241 10091 1275
rect 14197 1241 14231 1275
rect 15853 1241 15887 1275
rect 21281 1241 21315 1275
rect 22477 1241 22511 1275
rect 3893 1173 3927 1207
rect 5089 1173 5123 1207
rect 5549 1173 5583 1207
rect 6101 1173 6135 1207
rect 6377 1173 6411 1207
rect 6837 1173 6871 1207
rect 7205 1173 7239 1207
rect 7573 1173 7607 1207
rect 7941 1173 7975 1207
rect 8309 1173 8343 1207
rect 8585 1173 8619 1207
rect 8953 1173 8987 1207
rect 9781 1173 9815 1207
rect 11253 1173 11287 1207
rect 11713 1173 11747 1207
rect 11897 1173 11931 1207
rect 13461 1173 13495 1207
rect 13829 1173 13863 1207
rect 14841 1173 14875 1207
rect 17969 1173 18003 1207
rect 18889 1173 18923 1207
rect 21833 1173 21867 1207
rect 22293 1173 22327 1207
<< metal1 >>
rect 17218 44888 17224 44940
rect 17276 44928 17282 44940
rect 18506 44928 18512 44940
rect 17276 44900 18512 44928
rect 17276 44888 17282 44900
rect 18506 44888 18512 44900
rect 18564 44888 18570 44940
rect 8938 44752 8944 44804
rect 8996 44792 9002 44804
rect 9582 44792 9588 44804
rect 8996 44764 9588 44792
rect 8996 44752 9002 44764
rect 9582 44752 9588 44764
rect 9640 44752 9646 44804
rect 3510 44004 3516 44056
rect 3568 44044 3574 44056
rect 4614 44044 4620 44056
rect 3568 44016 4620 44044
rect 3568 44004 3574 44016
rect 4614 44004 4620 44016
rect 4672 44004 4678 44056
rect 3602 43800 3608 43852
rect 3660 43840 3666 43852
rect 6362 43840 6368 43852
rect 3660 43812 6368 43840
rect 3660 43800 3666 43812
rect 6362 43800 6368 43812
rect 6420 43800 6426 43852
rect 4798 43772 4804 43784
rect 1780 43744 4804 43772
rect 1780 43648 1808 43744
rect 4798 43732 4804 43744
rect 4856 43732 4862 43784
rect 17034 43732 17040 43784
rect 17092 43772 17098 43784
rect 18046 43772 18052 43784
rect 17092 43744 18052 43772
rect 17092 43732 17098 43744
rect 18046 43732 18052 43744
rect 18104 43732 18110 43784
rect 3418 43664 3424 43716
rect 3476 43704 3482 43716
rect 10502 43704 10508 43716
rect 3476 43676 10508 43704
rect 3476 43664 3482 43676
rect 10502 43664 10508 43676
rect 10560 43664 10566 43716
rect 17586 43664 17592 43716
rect 17644 43704 17650 43716
rect 18598 43704 18604 43716
rect 17644 43676 18604 43704
rect 17644 43664 17650 43676
rect 18598 43664 18604 43676
rect 18656 43664 18662 43716
rect 1762 43596 1768 43648
rect 1820 43596 1826 43648
rect 3970 43596 3976 43648
rect 4028 43636 4034 43648
rect 5258 43636 5264 43648
rect 4028 43608 5264 43636
rect 4028 43596 4034 43608
rect 5258 43596 5264 43608
rect 5316 43596 5322 43648
rect 9122 43596 9128 43648
rect 9180 43636 9186 43648
rect 16850 43636 16856 43648
rect 9180 43608 16856 43636
rect 9180 43596 9186 43608
rect 16850 43596 16856 43608
rect 16908 43596 16914 43648
rect 17310 43596 17316 43648
rect 17368 43636 17374 43648
rect 18322 43636 18328 43648
rect 17368 43608 18328 43636
rect 17368 43596 17374 43608
rect 18322 43596 18328 43608
rect 18380 43596 18386 43648
rect 19978 43596 19984 43648
rect 20036 43636 20042 43648
rect 22646 43636 22652 43648
rect 20036 43608 22652 43636
rect 20036 43596 20042 43608
rect 22646 43596 22652 43608
rect 22704 43596 22710 43648
rect 1104 43546 25000 43568
rect 1104 43494 6884 43546
rect 6936 43494 6948 43546
rect 7000 43494 7012 43546
rect 7064 43494 7076 43546
rect 7128 43494 7140 43546
rect 7192 43494 12818 43546
rect 12870 43494 12882 43546
rect 12934 43494 12946 43546
rect 12998 43494 13010 43546
rect 13062 43494 13074 43546
rect 13126 43494 18752 43546
rect 18804 43494 18816 43546
rect 18868 43494 18880 43546
rect 18932 43494 18944 43546
rect 18996 43494 19008 43546
rect 19060 43494 24686 43546
rect 24738 43494 24750 43546
rect 24802 43494 24814 43546
rect 24866 43494 24878 43546
rect 24930 43494 24942 43546
rect 24994 43494 25000 43546
rect 1104 43472 25000 43494
rect 2041 43435 2099 43441
rect 2041 43401 2053 43435
rect 2087 43432 2099 43435
rect 2130 43432 2136 43444
rect 2087 43404 2136 43432
rect 2087 43401 2099 43404
rect 2041 43395 2099 43401
rect 2130 43392 2136 43404
rect 2188 43392 2194 43444
rect 2406 43392 2412 43444
rect 2464 43392 2470 43444
rect 2958 43392 2964 43444
rect 3016 43392 3022 43444
rect 3510 43392 3516 43444
rect 3568 43392 3574 43444
rect 3970 43432 3976 43444
rect 3620 43404 3976 43432
rect 2317 43367 2375 43373
rect 2317 43333 2329 43367
rect 2363 43364 2375 43367
rect 3620 43364 3648 43404
rect 3970 43392 3976 43404
rect 4028 43392 4034 43444
rect 4801 43435 4859 43441
rect 4801 43401 4813 43435
rect 4847 43432 4859 43435
rect 5166 43432 5172 43444
rect 4847 43404 5172 43432
rect 4847 43401 4859 43404
rect 4801 43395 4859 43401
rect 5166 43392 5172 43404
rect 5224 43392 5230 43444
rect 5353 43435 5411 43441
rect 5353 43401 5365 43435
rect 5399 43432 5411 43435
rect 5442 43432 5448 43444
rect 5399 43404 5448 43432
rect 5399 43401 5411 43404
rect 5353 43395 5411 43401
rect 5442 43392 5448 43404
rect 5500 43392 5506 43444
rect 5718 43392 5724 43444
rect 5776 43392 5782 43444
rect 6365 43435 6423 43441
rect 6365 43401 6377 43435
rect 6411 43432 6423 43435
rect 6411 43404 6776 43432
rect 6411 43401 6423 43404
rect 6365 43395 6423 43401
rect 6748 43373 6776 43404
rect 6822 43392 6828 43444
rect 6880 43432 6886 43444
rect 7009 43435 7067 43441
rect 7009 43432 7021 43435
rect 6880 43404 7021 43432
rect 6880 43392 6886 43404
rect 7009 43401 7021 43404
rect 7055 43401 7067 43435
rect 7009 43395 7067 43401
rect 7561 43435 7619 43441
rect 7561 43401 7573 43435
rect 7607 43432 7619 43435
rect 7926 43432 7932 43444
rect 7607 43404 7932 43432
rect 7607 43401 7619 43404
rect 7561 43395 7619 43401
rect 7926 43392 7932 43404
rect 7984 43392 7990 43444
rect 8113 43435 8171 43441
rect 8113 43401 8125 43435
rect 8159 43432 8171 43435
rect 8202 43432 8208 43444
rect 8159 43404 8208 43432
rect 8159 43401 8171 43404
rect 8113 43395 8171 43401
rect 8202 43392 8208 43404
rect 8260 43392 8266 43444
rect 8665 43435 8723 43441
rect 8665 43401 8677 43435
rect 8711 43432 8723 43435
rect 8938 43432 8944 43444
rect 8711 43404 8944 43432
rect 8711 43401 8723 43404
rect 8665 43395 8723 43401
rect 8938 43392 8944 43404
rect 8996 43392 9002 43444
rect 9030 43392 9036 43444
rect 9088 43432 9094 43444
rect 9125 43435 9183 43441
rect 9125 43432 9137 43435
rect 9088 43404 9137 43432
rect 9088 43392 9094 43404
rect 9125 43401 9137 43404
rect 9171 43401 9183 43435
rect 9125 43395 9183 43401
rect 9769 43435 9827 43441
rect 9769 43401 9781 43435
rect 9815 43432 9827 43435
rect 9858 43432 9864 43444
rect 9815 43404 9864 43432
rect 9815 43401 9827 43404
rect 9769 43395 9827 43401
rect 9858 43392 9864 43404
rect 9916 43392 9922 43444
rect 10502 43392 10508 43444
rect 10560 43392 10566 43444
rect 13170 43392 13176 43444
rect 13228 43432 13234 43444
rect 13228 43404 14228 43432
rect 13228 43392 13234 43404
rect 6733 43367 6791 43373
rect 2363 43336 3648 43364
rect 3988 43336 6408 43364
rect 2363 43333 2375 43336
rect 2317 43327 2375 43333
rect 1581 43299 1639 43305
rect 1581 43265 1593 43299
rect 1627 43296 1639 43299
rect 1670 43296 1676 43308
rect 1627 43268 1676 43296
rect 1627 43265 1639 43268
rect 1581 43259 1639 43265
rect 1670 43256 1676 43268
rect 1728 43256 1734 43308
rect 1762 43256 1768 43308
rect 1820 43256 1826 43308
rect 2866 43256 2872 43308
rect 2924 43256 2930 43308
rect 3329 43299 3387 43305
rect 3329 43265 3341 43299
rect 3375 43296 3387 43299
rect 3602 43296 3608 43308
rect 3375 43268 3608 43296
rect 3375 43265 3387 43268
rect 3329 43259 3387 43265
rect 3602 43256 3608 43268
rect 3660 43256 3666 43308
rect 3988 43305 4016 43336
rect 3973 43299 4031 43305
rect 3973 43265 3985 43299
rect 4019 43265 4031 43299
rect 3973 43259 4031 43265
rect 4154 43256 4160 43308
rect 4212 43256 4218 43308
rect 4522 43256 4528 43308
rect 4580 43256 4586 43308
rect 4614 43256 4620 43308
rect 4672 43256 4678 43308
rect 5077 43299 5135 43305
rect 5077 43265 5089 43299
rect 5123 43265 5135 43299
rect 5077 43259 5135 43265
rect 1397 43163 1455 43169
rect 1397 43129 1409 43163
rect 1443 43160 1455 43163
rect 5092 43160 5120 43259
rect 5442 43256 5448 43308
rect 5500 43296 5506 43308
rect 5629 43299 5687 43305
rect 5629 43296 5641 43299
rect 5500 43268 5641 43296
rect 5500 43256 5506 43268
rect 5629 43265 5641 43268
rect 5675 43265 5687 43299
rect 5629 43259 5687 43265
rect 6380 43240 6408 43336
rect 6733 43333 6745 43367
rect 6779 43333 6791 43367
rect 6733 43327 6791 43333
rect 11238 43324 11244 43376
rect 11296 43364 11302 43376
rect 11609 43367 11667 43373
rect 11609 43364 11621 43367
rect 11296 43336 11621 43364
rect 11296 43324 11302 43336
rect 11609 43333 11621 43336
rect 11655 43333 11667 43367
rect 11609 43327 11667 43333
rect 12434 43324 12440 43376
rect 12492 43324 12498 43376
rect 12618 43324 12624 43376
rect 12676 43364 12682 43376
rect 12805 43367 12863 43373
rect 12805 43364 12817 43367
rect 12676 43336 12817 43364
rect 12676 43324 12682 43336
rect 12805 43333 12817 43336
rect 12851 43333 12863 43367
rect 12805 43327 12863 43333
rect 13446 43324 13452 43376
rect 13504 43364 13510 43376
rect 14200 43373 14228 43404
rect 16850 43392 16856 43444
rect 16908 43392 16914 43444
rect 17313 43435 17371 43441
rect 17313 43401 17325 43435
rect 17359 43401 17371 43435
rect 17313 43395 17371 43401
rect 17589 43435 17647 43441
rect 17589 43401 17601 43435
rect 17635 43432 17647 43435
rect 17678 43432 17684 43444
rect 17635 43404 17684 43432
rect 17635 43401 17647 43404
rect 17589 43395 17647 43401
rect 13725 43367 13783 43373
rect 13725 43364 13737 43367
rect 13504 43336 13737 43364
rect 13504 43324 13510 43336
rect 13725 43333 13737 43336
rect 13771 43333 13783 43367
rect 13725 43327 13783 43333
rect 14185 43367 14243 43373
rect 14185 43333 14197 43367
rect 14231 43333 14243 43367
rect 14185 43327 14243 43333
rect 14734 43324 14740 43376
rect 14792 43324 14798 43376
rect 14826 43324 14832 43376
rect 14884 43364 14890 43376
rect 15105 43367 15163 43373
rect 15105 43364 15117 43367
rect 14884 43336 15117 43364
rect 14884 43324 14890 43336
rect 15105 43333 15117 43336
rect 15151 43333 15163 43367
rect 15105 43327 15163 43333
rect 15562 43324 15568 43376
rect 15620 43324 15626 43376
rect 15654 43324 15660 43376
rect 15712 43364 15718 43376
rect 15933 43367 15991 43373
rect 15933 43364 15945 43367
rect 15712 43336 15945 43364
rect 15712 43324 15718 43336
rect 15933 43333 15945 43336
rect 15979 43333 15991 43367
rect 15933 43327 15991 43333
rect 16114 43324 16120 43376
rect 16172 43364 16178 43376
rect 16301 43367 16359 43373
rect 16301 43364 16313 43367
rect 16172 43336 16313 43364
rect 16172 43324 16178 43336
rect 16301 43333 16313 43336
rect 16347 43333 16359 43367
rect 16301 43327 16359 43333
rect 16390 43324 16396 43376
rect 16448 43364 16454 43376
rect 16761 43367 16819 43373
rect 16761 43364 16773 43367
rect 16448 43336 16773 43364
rect 16448 43324 16454 43336
rect 16761 43333 16773 43336
rect 16807 43333 16819 43367
rect 16761 43327 16819 43333
rect 17328 43308 17356 43395
rect 17678 43392 17684 43404
rect 17736 43392 17742 43444
rect 17862 43392 17868 43444
rect 17920 43432 17926 43444
rect 18417 43435 18475 43441
rect 18417 43432 18429 43435
rect 17920 43404 18429 43432
rect 17920 43392 17926 43404
rect 18417 43401 18429 43404
rect 18463 43401 18475 43435
rect 18417 43395 18475 43401
rect 20438 43392 20444 43444
rect 20496 43392 20502 43444
rect 20622 43392 20628 43444
rect 20680 43432 20686 43444
rect 20993 43435 21051 43441
rect 20993 43432 21005 43435
rect 20680 43404 21005 43432
rect 20680 43392 20686 43404
rect 20993 43401 21005 43404
rect 21039 43401 21051 43435
rect 20993 43395 21051 43401
rect 21358 43392 21364 43444
rect 21416 43432 21422 43444
rect 22189 43435 22247 43441
rect 22189 43432 22201 43435
rect 21416 43404 22201 43432
rect 21416 43392 21422 43404
rect 22189 43401 22201 43404
rect 22235 43401 22247 43435
rect 22189 43395 22247 43401
rect 22557 43435 22615 43441
rect 22557 43401 22569 43435
rect 22603 43401 22615 43435
rect 22557 43395 22615 43401
rect 18230 43364 18236 43376
rect 17512 43336 18236 43364
rect 6546 43256 6552 43308
rect 6604 43256 6610 43308
rect 7377 43299 7435 43305
rect 7377 43265 7389 43299
rect 7423 43296 7435 43299
rect 7466 43296 7472 43308
rect 7423 43268 7472 43296
rect 7423 43265 7435 43268
rect 7377 43259 7435 43265
rect 7466 43256 7472 43268
rect 7524 43256 7530 43308
rect 7837 43299 7895 43305
rect 7837 43265 7849 43299
rect 7883 43296 7895 43299
rect 8294 43296 8300 43308
rect 7883 43268 8300 43296
rect 7883 43265 7895 43268
rect 7837 43259 7895 43265
rect 8294 43256 8300 43268
rect 8352 43256 8358 43308
rect 8389 43299 8447 43305
rect 8389 43265 8401 43299
rect 8435 43265 8447 43299
rect 8389 43259 8447 43265
rect 8941 43299 8999 43305
rect 8941 43265 8953 43299
rect 8987 43265 8999 43299
rect 8941 43259 8999 43265
rect 9493 43299 9551 43305
rect 9493 43265 9505 43299
rect 9539 43265 9551 43299
rect 9493 43259 9551 43265
rect 6362 43188 6368 43240
rect 6420 43188 6426 43240
rect 1443 43132 5120 43160
rect 1443 43129 1455 43132
rect 1397 43123 1455 43129
rect 3789 43095 3847 43101
rect 3789 43061 3801 43095
rect 3835 43092 3847 43095
rect 5534 43092 5540 43104
rect 3835 43064 5540 43092
rect 3835 43061 3847 43064
rect 3789 43055 3847 43061
rect 5534 43052 5540 43064
rect 5592 43052 5598 43104
rect 8404 43092 8432 43259
rect 8956 43160 8984 43259
rect 9508 43228 9536 43259
rect 9950 43256 9956 43308
rect 10008 43256 10014 43308
rect 10318 43256 10324 43308
rect 10376 43256 10382 43308
rect 10686 43256 10692 43308
rect 10744 43256 10750 43308
rect 11054 43256 11060 43308
rect 11112 43256 11118 43308
rect 12066 43256 12072 43308
rect 12124 43256 12130 43308
rect 12158 43256 12164 43308
rect 12216 43296 12222 43308
rect 16485 43299 16543 43305
rect 16485 43296 16497 43299
rect 12216 43268 16497 43296
rect 12216 43256 12222 43268
rect 16485 43265 16497 43268
rect 16531 43265 16543 43299
rect 16485 43259 16543 43265
rect 17218 43256 17224 43308
rect 17276 43256 17282 43308
rect 17310 43256 17316 43308
rect 17368 43256 17374 43308
rect 17512 43305 17540 43336
rect 18230 43324 18236 43336
rect 18288 43324 18294 43376
rect 21266 43364 21272 43376
rect 18432 43336 18920 43364
rect 17497 43299 17555 43305
rect 17497 43265 17509 43299
rect 17543 43265 17555 43299
rect 17773 43299 17831 43305
rect 17773 43296 17785 43299
rect 17497 43259 17555 43265
rect 17604 43268 17785 43296
rect 13630 43228 13636 43240
rect 9508 43200 13636 43228
rect 13630 43188 13636 43200
rect 13688 43188 13694 43240
rect 16758 43188 16764 43240
rect 16816 43228 16822 43240
rect 17604 43228 17632 43268
rect 17773 43265 17785 43268
rect 17819 43265 17831 43299
rect 17773 43259 17831 43265
rect 18046 43256 18052 43308
rect 18104 43256 18110 43308
rect 18322 43256 18328 43308
rect 18380 43256 18386 43308
rect 16816 43200 17632 43228
rect 16816 43188 16822 43200
rect 17954 43188 17960 43240
rect 18012 43228 18018 43240
rect 18432 43228 18460 43336
rect 18598 43256 18604 43308
rect 18656 43256 18662 43308
rect 18892 43305 18920 43336
rect 19812 43336 21272 43364
rect 18877 43299 18935 43305
rect 18877 43265 18889 43299
rect 18923 43265 18935 43299
rect 18877 43259 18935 43265
rect 19426 43256 19432 43308
rect 19484 43256 19490 43308
rect 19812 43305 19840 43336
rect 21266 43324 21272 43336
rect 21324 43324 21330 43376
rect 21450 43324 21456 43376
rect 21508 43364 21514 43376
rect 22572 43364 22600 43395
rect 22646 43392 22652 43444
rect 22704 43432 22710 43444
rect 22704 43404 23060 43432
rect 22704 43392 22710 43404
rect 23032 43373 23060 43404
rect 23382 43392 23388 43444
rect 23440 43432 23446 43444
rect 23661 43435 23719 43441
rect 23661 43432 23673 43435
rect 23440 43404 23673 43432
rect 23440 43392 23446 43404
rect 23661 43401 23673 43404
rect 23707 43401 23719 43435
rect 23661 43395 23719 43401
rect 21508 43336 22600 43364
rect 23017 43367 23075 43373
rect 21508 43324 21514 43336
rect 23017 43333 23029 43367
rect 23063 43333 23075 43367
rect 23017 43327 23075 43333
rect 19797 43299 19855 43305
rect 19797 43265 19809 43299
rect 19843 43265 19855 43299
rect 19797 43259 19855 43265
rect 20165 43299 20223 43305
rect 20165 43265 20177 43299
rect 20211 43265 20223 43299
rect 20165 43259 20223 43265
rect 18012 43200 18460 43228
rect 18012 43188 18018 43200
rect 18506 43188 18512 43240
rect 18564 43228 18570 43240
rect 19242 43228 19248 43240
rect 18564 43200 19248 43228
rect 18564 43188 18570 43200
rect 19242 43188 19248 43200
rect 19300 43188 19306 43240
rect 20180 43228 20208 43259
rect 20346 43256 20352 43308
rect 20404 43256 20410 43308
rect 20898 43256 20904 43308
rect 20956 43256 20962 43308
rect 21082 43256 21088 43308
rect 21140 43296 21146 43308
rect 21361 43299 21419 43305
rect 21361 43296 21373 43299
rect 21140 43268 21373 43296
rect 21140 43256 21146 43268
rect 21361 43265 21373 43268
rect 21407 43265 21419 43299
rect 21361 43259 21419 43265
rect 21542 43256 21548 43308
rect 21600 43296 21606 43308
rect 21913 43299 21971 43305
rect 21913 43296 21925 43299
rect 21600 43268 21925 43296
rect 21600 43256 21606 43268
rect 21913 43265 21925 43268
rect 21959 43265 21971 43299
rect 21913 43259 21971 43265
rect 22094 43256 22100 43308
rect 22152 43296 22158 43308
rect 22465 43299 22523 43305
rect 22465 43296 22477 43299
rect 22152 43268 22477 43296
rect 22152 43256 22158 43268
rect 22465 43265 22477 43268
rect 22511 43265 22523 43299
rect 22465 43259 22523 43265
rect 22554 43256 22560 43308
rect 22612 43256 22618 43308
rect 23382 43256 23388 43308
rect 23440 43296 23446 43308
rect 23569 43299 23627 43305
rect 23569 43296 23581 43299
rect 23440 43268 23581 43296
rect 23440 43256 23446 43268
rect 23569 43265 23581 43268
rect 23615 43265 23627 43299
rect 23569 43259 23627 43265
rect 24213 43299 24271 43305
rect 24213 43265 24225 43299
rect 24259 43265 24271 43299
rect 24213 43259 24271 43265
rect 22572 43228 22600 43256
rect 20180 43200 22600 43228
rect 23106 43188 23112 43240
rect 23164 43228 23170 43240
rect 24228 43228 24256 43259
rect 23164 43200 24256 43228
rect 23164 43188 23170 43200
rect 10318 43160 10324 43172
rect 8956 43132 10324 43160
rect 10318 43120 10324 43132
rect 10376 43120 10382 43172
rect 11790 43120 11796 43172
rect 11848 43120 11854 43172
rect 12621 43163 12679 43169
rect 12621 43129 12633 43163
rect 12667 43160 12679 43163
rect 13078 43160 13084 43172
rect 12667 43132 13084 43160
rect 12667 43129 12679 43132
rect 12621 43123 12679 43129
rect 13078 43120 13084 43132
rect 13136 43120 13142 43172
rect 14918 43120 14924 43172
rect 14976 43120 14982 43172
rect 15286 43120 15292 43172
rect 15344 43120 15350 43172
rect 16114 43120 16120 43172
rect 16172 43120 16178 43172
rect 17037 43163 17095 43169
rect 17037 43129 17049 43163
rect 17083 43160 17095 43163
rect 17402 43160 17408 43172
rect 17083 43132 17408 43160
rect 17083 43129 17095 43132
rect 17037 43123 17095 43129
rect 17402 43120 17408 43132
rect 17460 43120 17466 43172
rect 17494 43120 17500 43172
rect 17552 43160 17558 43172
rect 18141 43163 18199 43169
rect 18141 43160 18153 43163
rect 17552 43132 18153 43160
rect 17552 43120 17558 43132
rect 18141 43129 18153 43132
rect 18187 43129 18199 43163
rect 18141 43123 18199 43129
rect 20070 43120 20076 43172
rect 20128 43160 20134 43172
rect 24029 43163 24087 43169
rect 24029 43160 24041 43163
rect 20128 43132 24041 43160
rect 20128 43120 20134 43132
rect 24029 43129 24041 43132
rect 24075 43129 24087 43163
rect 24029 43123 24087 43129
rect 9766 43092 9772 43104
rect 8404 43064 9772 43092
rect 9766 43052 9772 43064
rect 9824 43052 9830 43104
rect 10137 43095 10195 43101
rect 10137 43061 10149 43095
rect 10183 43092 10195 43095
rect 10410 43092 10416 43104
rect 10183 43064 10416 43092
rect 10183 43061 10195 43064
rect 10137 43055 10195 43061
rect 10410 43052 10416 43064
rect 10468 43052 10474 43104
rect 10870 43052 10876 43104
rect 10928 43052 10934 43104
rect 11238 43052 11244 43104
rect 11296 43052 11302 43104
rect 12250 43052 12256 43104
rect 12308 43052 12314 43104
rect 12894 43052 12900 43104
rect 12952 43052 12958 43104
rect 13814 43052 13820 43104
rect 13872 43052 13878 43104
rect 14274 43052 14280 43104
rect 14332 43052 14338 43104
rect 15654 43052 15660 43104
rect 15712 43052 15718 43104
rect 17586 43052 17592 43104
rect 17644 43092 17650 43104
rect 17865 43095 17923 43101
rect 17865 43092 17877 43095
rect 17644 43064 17877 43092
rect 17644 43052 17650 43064
rect 17865 43061 17877 43064
rect 17911 43061 17923 43095
rect 17865 43055 17923 43061
rect 18046 43052 18052 43104
rect 18104 43092 18110 43104
rect 18693 43095 18751 43101
rect 18693 43092 18705 43095
rect 18104 43064 18705 43092
rect 18104 43052 18110 43064
rect 18693 43061 18705 43064
rect 18739 43061 18751 43095
rect 18693 43055 18751 43061
rect 19245 43095 19303 43101
rect 19245 43061 19257 43095
rect 19291 43092 19303 43095
rect 19334 43092 19340 43104
rect 19291 43064 19340 43092
rect 19291 43061 19303 43064
rect 19245 43055 19303 43061
rect 19334 43052 19340 43064
rect 19392 43052 19398 43104
rect 20990 43052 20996 43104
rect 21048 43092 21054 43104
rect 21545 43095 21603 43101
rect 21545 43092 21557 43095
rect 21048 43064 21557 43092
rect 21048 43052 21054 43064
rect 21545 43061 21557 43064
rect 21591 43061 21603 43095
rect 21545 43055 21603 43061
rect 21910 43052 21916 43104
rect 21968 43092 21974 43104
rect 23109 43095 23167 43101
rect 23109 43092 23121 43095
rect 21968 43064 23121 43092
rect 21968 43052 21974 43064
rect 23109 43061 23121 43064
rect 23155 43061 23167 43095
rect 23109 43055 23167 43061
rect 1104 43002 24840 43024
rect 1104 42950 3917 43002
rect 3969 42950 3981 43002
rect 4033 42950 4045 43002
rect 4097 42950 4109 43002
rect 4161 42950 4173 43002
rect 4225 42950 9851 43002
rect 9903 42950 9915 43002
rect 9967 42950 9979 43002
rect 10031 42950 10043 43002
rect 10095 42950 10107 43002
rect 10159 42950 15785 43002
rect 15837 42950 15849 43002
rect 15901 42950 15913 43002
rect 15965 42950 15977 43002
rect 16029 42950 16041 43002
rect 16093 42950 21719 43002
rect 21771 42950 21783 43002
rect 21835 42950 21847 43002
rect 21899 42950 21911 43002
rect 21963 42950 21975 43002
rect 22027 42950 24840 43002
rect 1104 42928 24840 42950
rect 3326 42848 3332 42900
rect 3384 42848 3390 42900
rect 4338 42848 4344 42900
rect 4396 42848 4402 42900
rect 6086 42848 6092 42900
rect 6144 42848 6150 42900
rect 6638 42848 6644 42900
rect 6696 42848 6702 42900
rect 7190 42848 7196 42900
rect 7248 42848 7254 42900
rect 8294 42848 8300 42900
rect 8352 42888 8358 42900
rect 8941 42891 8999 42897
rect 8941 42888 8953 42891
rect 8352 42860 8953 42888
rect 8352 42848 8358 42860
rect 8941 42857 8953 42860
rect 8987 42857 8999 42891
rect 12069 42891 12127 42897
rect 12069 42888 12081 42891
rect 8941 42851 8999 42857
rect 9232 42860 12081 42888
rect 4709 42823 4767 42829
rect 4709 42820 4721 42823
rect 4630 42792 4721 42820
rect 2682 42712 2688 42764
rect 2740 42752 2746 42764
rect 2961 42755 3019 42761
rect 2961 42752 2973 42755
rect 2740 42724 2973 42752
rect 2740 42712 2746 42724
rect 2961 42721 2973 42724
rect 3007 42721 3019 42755
rect 2961 42715 3019 42721
rect 3789 42687 3847 42693
rect 3789 42653 3801 42687
rect 3835 42684 3847 42687
rect 4522 42684 4528 42696
rect 3835 42656 4528 42684
rect 3835 42653 3847 42656
rect 3789 42647 3847 42653
rect 4522 42644 4528 42656
rect 4580 42644 4586 42696
rect 1394 42576 1400 42628
rect 1452 42576 1458 42628
rect 2038 42576 2044 42628
rect 2096 42616 2102 42628
rect 2133 42619 2191 42625
rect 2133 42616 2145 42619
rect 2096 42588 2145 42616
rect 2096 42576 2102 42588
rect 2133 42585 2145 42588
rect 2179 42585 2191 42619
rect 2133 42579 2191 42585
rect 2685 42619 2743 42625
rect 2685 42585 2697 42619
rect 2731 42616 2743 42619
rect 3050 42616 3056 42628
rect 2731 42588 3056 42616
rect 2731 42585 2743 42588
rect 2685 42579 2743 42585
rect 3050 42576 3056 42588
rect 3108 42576 3114 42628
rect 3234 42576 3240 42628
rect 3292 42576 3298 42628
rect 4249 42619 4307 42625
rect 4249 42585 4261 42619
rect 4295 42585 4307 42619
rect 4630 42616 4658 42792
rect 4709 42789 4721 42792
rect 4755 42789 4767 42823
rect 4709 42783 4767 42789
rect 4982 42712 4988 42764
rect 5040 42752 5046 42764
rect 5353 42755 5411 42761
rect 5353 42752 5365 42755
rect 5040 42724 5365 42752
rect 5040 42712 5046 42724
rect 5353 42721 5365 42724
rect 5399 42721 5411 42755
rect 5353 42715 5411 42721
rect 8665 42755 8723 42761
rect 8665 42721 8677 42755
rect 8711 42752 8723 42755
rect 8754 42752 8760 42764
rect 8711 42724 8760 42752
rect 8711 42721 8723 42724
rect 8665 42715 8723 42721
rect 8754 42712 8760 42724
rect 8812 42712 8818 42764
rect 9232 42752 9260 42860
rect 12069 42857 12081 42860
rect 12115 42857 12127 42891
rect 12069 42851 12127 42857
rect 13630 42848 13636 42900
rect 13688 42848 13694 42900
rect 16945 42891 17003 42897
rect 16945 42857 16957 42891
rect 16991 42857 17003 42891
rect 16945 42851 17003 42857
rect 9766 42780 9772 42832
rect 9824 42820 9830 42832
rect 10321 42823 10379 42829
rect 10321 42820 10333 42823
rect 9824 42792 10333 42820
rect 9824 42780 9830 42792
rect 10321 42789 10333 42792
rect 10367 42789 10379 42823
rect 13648 42820 13676 42848
rect 13648 42792 14780 42820
rect 10321 42783 10379 42789
rect 8864 42724 9260 42752
rect 4706 42644 4712 42696
rect 4764 42684 4770 42696
rect 4893 42687 4951 42693
rect 4893 42684 4905 42687
rect 4764 42656 4905 42684
rect 4764 42644 4770 42656
rect 4893 42653 4905 42656
rect 4939 42653 4951 42687
rect 4893 42647 4951 42653
rect 5534 42644 5540 42696
rect 5592 42644 5598 42696
rect 7558 42644 7564 42696
rect 7616 42644 7622 42696
rect 8110 42644 8116 42696
rect 8168 42644 8174 42696
rect 8864 42684 8892 42724
rect 9306 42712 9312 42764
rect 9364 42752 9370 42764
rect 13538 42752 13544 42764
rect 9364 42724 10272 42752
rect 9364 42712 9370 42724
rect 8220 42656 8892 42684
rect 5077 42619 5135 42625
rect 5077 42616 5089 42619
rect 4630 42588 5089 42616
rect 4249 42579 4307 42585
rect 5077 42585 5089 42588
rect 5123 42585 5135 42619
rect 5077 42579 5135 42585
rect 3786 42508 3792 42560
rect 3844 42548 3850 42560
rect 3973 42551 4031 42557
rect 3973 42548 3985 42551
rect 3844 42520 3985 42548
rect 3844 42508 3850 42520
rect 3973 42517 3985 42520
rect 4019 42517 4031 42551
rect 4264 42548 4292 42579
rect 5994 42576 6000 42628
rect 6052 42576 6058 42628
rect 6549 42619 6607 42625
rect 6549 42585 6561 42619
rect 6595 42616 6607 42619
rect 6730 42616 6736 42628
rect 6595 42588 6736 42616
rect 6595 42585 6607 42588
rect 6549 42579 6607 42585
rect 6730 42576 6736 42588
rect 6788 42576 6794 42628
rect 7101 42619 7159 42625
rect 7101 42585 7113 42619
rect 7147 42616 7159 42619
rect 7282 42616 7288 42628
rect 7147 42588 7288 42616
rect 7147 42585 7159 42588
rect 7101 42579 7159 42585
rect 7282 42576 7288 42588
rect 7340 42576 7346 42628
rect 7650 42576 7656 42628
rect 7708 42576 7714 42628
rect 7834 42576 7840 42628
rect 7892 42616 7898 42628
rect 8220 42616 8248 42656
rect 9122 42644 9128 42696
rect 9180 42644 9186 42696
rect 10244 42693 10272 42724
rect 10980 42724 13544 42752
rect 10229 42687 10287 42693
rect 9232 42656 9904 42684
rect 7892 42588 8248 42616
rect 8389 42619 8447 42625
rect 7892 42576 7898 42588
rect 8389 42585 8401 42619
rect 8435 42616 8447 42619
rect 9232 42616 9260 42656
rect 8435 42588 9260 42616
rect 8435 42585 8447 42588
rect 8389 42579 8447 42585
rect 9490 42576 9496 42628
rect 9548 42576 9554 42628
rect 9674 42576 9680 42628
rect 9732 42616 9738 42628
rect 9732 42588 9812 42616
rect 9732 42576 9738 42588
rect 5534 42548 5540 42560
rect 4264 42520 5540 42548
rect 3973 42511 4031 42517
rect 5534 42508 5540 42520
rect 5592 42508 5598 42560
rect 5721 42551 5779 42557
rect 5721 42517 5733 42551
rect 5767 42548 5779 42551
rect 6270 42548 6276 42560
rect 5767 42520 6276 42548
rect 5767 42517 5779 42520
rect 5721 42511 5779 42517
rect 6270 42508 6276 42520
rect 6328 42508 6334 42560
rect 7668 42548 7696 42576
rect 7745 42551 7803 42557
rect 7745 42548 7757 42551
rect 7668 42520 7757 42548
rect 7745 42517 7757 42520
rect 7791 42517 7803 42551
rect 7745 42511 7803 42517
rect 7926 42508 7932 42560
rect 7984 42508 7990 42560
rect 8294 42508 8300 42560
rect 8352 42548 8358 42560
rect 9582 42548 9588 42560
rect 8352 42520 9588 42548
rect 8352 42508 8358 42520
rect 9582 42508 9588 42520
rect 9640 42508 9646 42560
rect 9784 42557 9812 42588
rect 9769 42551 9827 42557
rect 9769 42517 9781 42551
rect 9815 42517 9827 42551
rect 9876 42548 9904 42656
rect 10229 42653 10241 42687
rect 10275 42653 10287 42687
rect 10229 42647 10287 42653
rect 10318 42644 10324 42696
rect 10376 42644 10382 42696
rect 10502 42644 10508 42696
rect 10560 42644 10566 42696
rect 10870 42644 10876 42696
rect 10928 42644 10934 42696
rect 10980 42693 11008 42724
rect 13538 42712 13544 42724
rect 13596 42712 13602 42764
rect 13814 42712 13820 42764
rect 13872 42752 13878 42764
rect 14752 42752 14780 42792
rect 16960 42752 16988 42851
rect 17310 42848 17316 42900
rect 17368 42848 17374 42900
rect 17402 42848 17408 42900
rect 17460 42888 17466 42900
rect 17460 42860 18828 42888
rect 17460 42848 17466 42860
rect 13872 42724 14688 42752
rect 14752 42724 16988 42752
rect 17328 42752 17356 42848
rect 18598 42780 18604 42832
rect 18656 42780 18662 42832
rect 17328 42724 18552 42752
rect 13872 42712 13878 42724
rect 10965 42687 11023 42693
rect 10965 42653 10977 42687
rect 11011 42653 11023 42687
rect 10965 42647 11023 42653
rect 11606 42644 11612 42696
rect 11664 42644 11670 42696
rect 11882 42644 11888 42696
rect 11940 42644 11946 42696
rect 12342 42644 12348 42696
rect 12400 42644 12406 42696
rect 12710 42644 12716 42696
rect 12768 42684 12774 42696
rect 12989 42687 13047 42693
rect 12989 42684 13001 42687
rect 12768 42656 13001 42684
rect 12768 42644 12774 42656
rect 12989 42653 13001 42656
rect 13035 42653 13047 42687
rect 12989 42647 13047 42653
rect 14090 42644 14096 42696
rect 14148 42644 14154 42696
rect 14366 42644 14372 42696
rect 14424 42644 14430 42696
rect 14660 42693 14688 42724
rect 14645 42687 14703 42693
rect 14645 42653 14657 42687
rect 14691 42653 14703 42687
rect 14645 42647 14703 42653
rect 15102 42644 15108 42696
rect 15160 42644 15166 42696
rect 15378 42644 15384 42696
rect 15436 42644 15442 42696
rect 16482 42644 16488 42696
rect 16540 42684 16546 42696
rect 16577 42687 16635 42693
rect 16577 42684 16589 42687
rect 16540 42656 16589 42684
rect 16540 42644 16546 42656
rect 16577 42653 16589 42656
rect 16623 42653 16635 42687
rect 16577 42647 16635 42653
rect 17129 42687 17187 42693
rect 17129 42653 17141 42687
rect 17175 42653 17187 42687
rect 17129 42647 17187 42653
rect 17405 42687 17463 42693
rect 17405 42653 17417 42687
rect 17451 42684 17463 42687
rect 17494 42684 17500 42696
rect 17451 42656 17500 42684
rect 17451 42653 17463 42656
rect 17405 42647 17463 42653
rect 10045 42551 10103 42557
rect 10045 42548 10057 42551
rect 9876 42520 10057 42548
rect 9769 42511 9827 42517
rect 10045 42517 10057 42520
rect 10091 42517 10103 42551
rect 10336 42548 10364 42644
rect 10778 42576 10784 42628
rect 10836 42616 10842 42628
rect 10836 42588 13216 42616
rect 10836 42576 10842 42588
rect 10689 42551 10747 42557
rect 10689 42548 10701 42551
rect 10336 42520 10701 42548
rect 10045 42511 10103 42517
rect 10689 42517 10701 42520
rect 10735 42517 10747 42551
rect 10689 42511 10747 42517
rect 11146 42508 11152 42560
rect 11204 42508 11210 42560
rect 11330 42508 11336 42560
rect 11388 42548 11394 42560
rect 11793 42551 11851 42557
rect 11793 42548 11805 42551
rect 11388 42520 11805 42548
rect 11388 42508 11394 42520
rect 11793 42517 11805 42520
rect 11839 42517 11851 42551
rect 11793 42511 11851 42517
rect 12526 42508 12532 42560
rect 12584 42508 12590 42560
rect 13188 42557 13216 42588
rect 13354 42576 13360 42628
rect 13412 42616 13418 42628
rect 13412 42588 14596 42616
rect 13412 42576 13418 42588
rect 13173 42551 13231 42557
rect 13173 42517 13185 42551
rect 13219 42517 13231 42551
rect 13173 42511 13231 42517
rect 13262 42508 13268 42560
rect 13320 42548 13326 42560
rect 14568 42557 14596 42588
rect 15120 42588 15608 42616
rect 15120 42560 15148 42588
rect 14277 42551 14335 42557
rect 14277 42548 14289 42551
rect 13320 42520 14289 42548
rect 13320 42508 13326 42520
rect 14277 42517 14289 42520
rect 14323 42517 14335 42551
rect 14277 42511 14335 42517
rect 14553 42551 14611 42557
rect 14553 42517 14565 42551
rect 14599 42517 14611 42551
rect 14553 42511 14611 42517
rect 14826 42508 14832 42560
rect 14884 42508 14890 42560
rect 15102 42508 15108 42560
rect 15160 42508 15166 42560
rect 15286 42508 15292 42560
rect 15344 42508 15350 42560
rect 15580 42557 15608 42588
rect 16390 42576 16396 42628
rect 16448 42616 16454 42628
rect 17144 42616 17172 42647
rect 17494 42644 17500 42656
rect 17552 42644 17558 42696
rect 17681 42687 17739 42693
rect 17681 42653 17693 42687
rect 17727 42684 17739 42687
rect 17862 42684 17868 42696
rect 17727 42656 17868 42684
rect 17727 42653 17739 42656
rect 17681 42647 17739 42653
rect 17862 42644 17868 42656
rect 17920 42644 17926 42696
rect 17957 42687 18015 42693
rect 17957 42653 17969 42687
rect 18003 42684 18015 42687
rect 18046 42684 18052 42696
rect 18003 42656 18052 42684
rect 18003 42653 18015 42656
rect 17957 42647 18015 42653
rect 18046 42644 18052 42656
rect 18104 42644 18110 42696
rect 18524 42693 18552 42724
rect 18800 42693 18828 42860
rect 20254 42848 20260 42900
rect 20312 42888 20318 42900
rect 21542 42888 21548 42900
rect 20312 42860 21548 42888
rect 20312 42848 20318 42860
rect 21542 42848 21548 42860
rect 21600 42848 21606 42900
rect 22922 42848 22928 42900
rect 22980 42888 22986 42900
rect 23293 42891 23351 42897
rect 23293 42888 23305 42891
rect 22980 42860 23305 42888
rect 22980 42848 22986 42860
rect 23293 42857 23305 42860
rect 23339 42857 23351 42891
rect 23293 42851 23351 42857
rect 19702 42780 19708 42832
rect 19760 42820 19766 42832
rect 21177 42823 21235 42829
rect 21177 42820 21189 42823
rect 19760 42792 21189 42820
rect 19760 42780 19766 42792
rect 21177 42789 21189 42792
rect 21223 42789 21235 42823
rect 21177 42783 21235 42789
rect 20070 42752 20076 42764
rect 18984 42724 20076 42752
rect 18233 42687 18291 42693
rect 18233 42653 18245 42687
rect 18279 42653 18291 42687
rect 18233 42647 18291 42653
rect 18509 42687 18567 42693
rect 18509 42653 18521 42687
rect 18555 42653 18567 42687
rect 18509 42647 18567 42653
rect 18785 42687 18843 42693
rect 18785 42653 18797 42687
rect 18831 42653 18843 42687
rect 18785 42647 18843 42653
rect 16448 42588 17172 42616
rect 18248 42616 18276 42647
rect 18984 42616 19012 42724
rect 20070 42712 20076 42724
rect 20128 42712 20134 42764
rect 20162 42712 20168 42764
rect 20220 42752 20226 42764
rect 20220 42724 22140 42752
rect 20220 42712 20226 42724
rect 19061 42687 19119 42693
rect 19061 42653 19073 42687
rect 19107 42684 19119 42687
rect 19610 42684 19616 42696
rect 19107 42656 19616 42684
rect 19107 42653 19119 42656
rect 19061 42647 19119 42653
rect 19610 42644 19616 42656
rect 19668 42644 19674 42696
rect 21358 42644 21364 42696
rect 21416 42644 21422 42696
rect 22112 42693 22140 42724
rect 22278 42712 22284 42764
rect 22336 42752 22342 42764
rect 22925 42755 22983 42761
rect 22925 42752 22937 42755
rect 22336 42724 22937 42752
rect 22336 42712 22342 42724
rect 22925 42721 22937 42724
rect 22971 42721 22983 42755
rect 22925 42715 22983 42721
rect 23566 42712 23572 42764
rect 23624 42752 23630 42764
rect 24029 42755 24087 42761
rect 24029 42752 24041 42755
rect 23624 42724 24041 42752
rect 23624 42712 23630 42724
rect 24029 42721 24041 42724
rect 24075 42721 24087 42755
rect 24029 42715 24087 42721
rect 22097 42687 22155 42693
rect 22097 42653 22109 42687
rect 22143 42653 22155 42687
rect 22097 42647 22155 42653
rect 22465 42687 22523 42693
rect 22465 42653 22477 42687
rect 22511 42684 22523 42687
rect 24118 42684 24124 42696
rect 22511 42656 24124 42684
rect 22511 42653 22523 42656
rect 22465 42647 22523 42653
rect 24118 42644 24124 42656
rect 24176 42644 24182 42696
rect 18248 42588 19012 42616
rect 16448 42576 16454 42588
rect 19242 42576 19248 42628
rect 19300 42576 19306 42628
rect 20990 42576 20996 42628
rect 21048 42576 21054 42628
rect 21545 42619 21603 42625
rect 21545 42616 21557 42619
rect 21100 42588 21557 42616
rect 15565 42551 15623 42557
rect 15565 42517 15577 42551
rect 15611 42517 15623 42551
rect 15565 42511 15623 42517
rect 16758 42508 16764 42560
rect 16816 42508 16822 42560
rect 17218 42508 17224 42560
rect 17276 42508 17282 42560
rect 17310 42508 17316 42560
rect 17368 42548 17374 42560
rect 17497 42551 17555 42557
rect 17497 42548 17509 42551
rect 17368 42520 17509 42548
rect 17368 42508 17374 42520
rect 17497 42517 17509 42520
rect 17543 42517 17555 42551
rect 17497 42511 17555 42517
rect 17770 42508 17776 42560
rect 17828 42508 17834 42560
rect 18046 42508 18052 42560
rect 18104 42508 18110 42560
rect 18322 42508 18328 42560
rect 18380 42508 18386 42560
rect 18414 42508 18420 42560
rect 18472 42548 18478 42560
rect 18877 42551 18935 42557
rect 18877 42548 18889 42551
rect 18472 42520 18889 42548
rect 18472 42508 18478 42520
rect 18877 42517 18889 42520
rect 18923 42517 18935 42551
rect 18877 42511 18935 42517
rect 20714 42508 20720 42560
rect 20772 42548 20778 42560
rect 21100 42548 21128 42588
rect 21545 42585 21557 42588
rect 21591 42585 21603 42619
rect 21545 42579 21603 42585
rect 21913 42619 21971 42625
rect 21913 42585 21925 42619
rect 21959 42616 21971 42619
rect 21959 42588 22094 42616
rect 21959 42585 21971 42588
rect 21913 42579 21971 42585
rect 20772 42520 21128 42548
rect 22066 42548 22094 42588
rect 22370 42576 22376 42628
rect 22428 42616 22434 42628
rect 22649 42619 22707 42625
rect 22649 42616 22661 42619
rect 22428 42588 22661 42616
rect 22428 42576 22434 42588
rect 22649 42585 22661 42588
rect 22695 42585 22707 42619
rect 22649 42579 22707 42585
rect 22830 42576 22836 42628
rect 22888 42616 22894 42628
rect 23201 42619 23259 42625
rect 23201 42616 23213 42619
rect 22888 42588 23213 42616
rect 22888 42576 22894 42588
rect 23201 42585 23213 42588
rect 23247 42585 23259 42619
rect 23201 42579 23259 42585
rect 23753 42619 23811 42625
rect 23753 42585 23765 42619
rect 23799 42616 23811 42619
rect 23842 42616 23848 42628
rect 23799 42588 23848 42616
rect 23799 42585 23811 42588
rect 23753 42579 23811 42585
rect 23842 42576 23848 42588
rect 23900 42576 23906 42628
rect 25038 42548 25044 42560
rect 22066 42520 25044 42548
rect 20772 42508 20778 42520
rect 25038 42508 25044 42520
rect 25096 42508 25102 42560
rect 1104 42458 25000 42480
rect 1104 42406 6884 42458
rect 6936 42406 6948 42458
rect 7000 42406 7012 42458
rect 7064 42406 7076 42458
rect 7128 42406 7140 42458
rect 7192 42406 12818 42458
rect 12870 42406 12882 42458
rect 12934 42406 12946 42458
rect 12998 42406 13010 42458
rect 13062 42406 13074 42458
rect 13126 42406 18752 42458
rect 18804 42406 18816 42458
rect 18868 42406 18880 42458
rect 18932 42406 18944 42458
rect 18996 42406 19008 42458
rect 19060 42406 24686 42458
rect 24738 42406 24750 42458
rect 24802 42406 24814 42458
rect 24866 42406 24878 42458
rect 24930 42406 24942 42458
rect 24994 42406 25000 42458
rect 1104 42384 25000 42406
rect 1026 42304 1032 42356
rect 1084 42344 1090 42356
rect 2593 42347 2651 42353
rect 2593 42344 2605 42347
rect 1084 42316 2605 42344
rect 1084 42304 1090 42316
rect 2593 42313 2605 42316
rect 2639 42313 2651 42347
rect 3145 42347 3203 42353
rect 3145 42344 3157 42347
rect 2593 42307 2651 42313
rect 2746 42316 3157 42344
rect 1578 42236 1584 42288
rect 1636 42276 1642 42288
rect 2746 42276 2774 42316
rect 3145 42313 3157 42316
rect 3191 42313 3203 42347
rect 3145 42307 3203 42313
rect 3234 42304 3240 42356
rect 3292 42344 3298 42356
rect 5626 42344 5632 42356
rect 3292 42316 5632 42344
rect 3292 42304 3298 42316
rect 5626 42304 5632 42316
rect 5684 42304 5690 42356
rect 6457 42347 6515 42353
rect 6457 42313 6469 42347
rect 6503 42344 6515 42347
rect 6546 42344 6552 42356
rect 6503 42316 6552 42344
rect 6503 42313 6515 42316
rect 6457 42307 6515 42313
rect 6546 42304 6552 42316
rect 6604 42304 6610 42356
rect 7374 42304 7380 42356
rect 7432 42344 7438 42356
rect 7561 42347 7619 42353
rect 7561 42344 7573 42347
rect 7432 42316 7573 42344
rect 7432 42304 7438 42316
rect 7561 42313 7573 42316
rect 7607 42313 7619 42347
rect 7561 42307 7619 42313
rect 8202 42304 8208 42356
rect 8260 42344 8266 42356
rect 8481 42347 8539 42353
rect 8481 42344 8493 42347
rect 8260 42316 8493 42344
rect 8260 42304 8266 42316
rect 8481 42313 8493 42316
rect 8527 42313 8539 42347
rect 8481 42307 8539 42313
rect 8846 42304 8852 42356
rect 8904 42344 8910 42356
rect 10778 42344 10784 42356
rect 8904 42316 10784 42344
rect 8904 42304 8910 42316
rect 10778 42304 10784 42316
rect 10836 42304 10842 42356
rect 11146 42304 11152 42356
rect 11204 42304 11210 42356
rect 12526 42344 12532 42356
rect 12406 42316 12532 42344
rect 4709 42279 4767 42285
rect 1636 42248 2774 42276
rect 3068 42248 4476 42276
rect 1636 42236 1642 42248
rect 1394 42168 1400 42220
rect 1452 42168 1458 42220
rect 2498 42168 2504 42220
rect 2556 42168 2562 42220
rect 3068 42217 3096 42248
rect 4448 42220 4476 42248
rect 4709 42245 4721 42279
rect 4755 42245 4767 42279
rect 4709 42239 4767 42245
rect 3053 42211 3111 42217
rect 3053 42177 3065 42211
rect 3099 42177 3111 42211
rect 3053 42171 3111 42177
rect 3602 42168 3608 42220
rect 3660 42168 3666 42220
rect 3786 42168 3792 42220
rect 3844 42208 3850 42220
rect 4157 42211 4215 42217
rect 4157 42208 4169 42211
rect 3844 42180 4169 42208
rect 3844 42168 3850 42180
rect 4157 42177 4169 42180
rect 4203 42177 4215 42211
rect 4157 42171 4215 42177
rect 4430 42168 4436 42220
rect 4488 42168 4494 42220
rect 2222 42100 2228 42152
rect 2280 42100 2286 42152
rect 4724 42140 4752 42239
rect 5810 42236 5816 42288
rect 5868 42276 5874 42288
rect 8294 42276 8300 42288
rect 5868 42248 7420 42276
rect 5868 42236 5874 42248
rect 5445 42211 5503 42217
rect 5445 42177 5457 42211
rect 5491 42208 5503 42211
rect 5905 42211 5963 42217
rect 5905 42208 5917 42211
rect 5491 42180 5917 42208
rect 5491 42177 5503 42180
rect 5445 42171 5503 42177
rect 5905 42177 5917 42180
rect 5951 42208 5963 42211
rect 6086 42208 6092 42220
rect 5951 42180 6092 42208
rect 5951 42177 5963 42180
rect 5905 42171 5963 42177
rect 6086 42168 6092 42180
rect 6144 42168 6150 42220
rect 6178 42168 6184 42220
rect 6236 42168 6242 42220
rect 6638 42168 6644 42220
rect 6696 42168 6702 42220
rect 6917 42211 6975 42217
rect 6917 42177 6929 42211
rect 6963 42208 6975 42211
rect 7190 42208 7196 42220
rect 6963 42180 7196 42208
rect 6963 42177 6975 42180
rect 6917 42171 6975 42177
rect 7190 42168 7196 42180
rect 7248 42168 7254 42220
rect 7392 42217 7420 42248
rect 7484 42248 8300 42276
rect 7377 42211 7435 42217
rect 7377 42177 7389 42211
rect 7423 42177 7435 42211
rect 7377 42171 7435 42177
rect 7484 42140 7512 42248
rect 8294 42236 8300 42248
rect 8352 42236 8358 42288
rect 9398 42236 9404 42288
rect 9456 42236 9462 42288
rect 9582 42236 9588 42288
rect 9640 42276 9646 42288
rect 11164 42276 11192 42304
rect 9640 42248 11192 42276
rect 9640 42236 9646 42248
rect 9275 42221 9333 42227
rect 7742 42168 7748 42220
rect 7800 42208 7806 42220
rect 7929 42211 7987 42217
rect 7929 42208 7941 42211
rect 7800 42180 7941 42208
rect 7800 42168 7806 42180
rect 7929 42177 7941 42180
rect 7975 42177 7987 42211
rect 7929 42171 7987 42177
rect 8018 42168 8024 42220
rect 8076 42208 8082 42220
rect 8205 42211 8263 42217
rect 8205 42208 8217 42211
rect 8076 42180 8217 42208
rect 8076 42168 8082 42180
rect 8205 42177 8217 42180
rect 8251 42177 8263 42211
rect 8205 42171 8263 42177
rect 8386 42168 8392 42220
rect 8444 42168 8450 42220
rect 8662 42168 8668 42220
rect 8720 42208 8726 42220
rect 9275 42218 9287 42221
rect 9048 42208 9287 42218
rect 8720 42190 9287 42208
rect 8720 42180 9076 42190
rect 9275 42187 9287 42190
rect 9321 42187 9333 42221
rect 9275 42181 9333 42187
rect 9416 42208 9444 42236
rect 12406 42208 12434 42316
rect 12526 42304 12532 42316
rect 12584 42304 12590 42356
rect 17218 42344 17224 42356
rect 16776 42316 17224 42344
rect 16776 42285 16804 42316
rect 17218 42304 17224 42316
rect 17276 42304 17282 42356
rect 17310 42304 17316 42356
rect 17368 42304 17374 42356
rect 17678 42344 17684 42356
rect 17420 42316 17684 42344
rect 16761 42279 16819 42285
rect 16761 42245 16773 42279
rect 16807 42245 16819 42279
rect 16761 42239 16819 42245
rect 17129 42279 17187 42285
rect 17129 42245 17141 42279
rect 17175 42276 17187 42279
rect 17328 42276 17356 42304
rect 17175 42248 17356 42276
rect 17175 42245 17187 42248
rect 17129 42239 17187 42245
rect 9416 42180 12434 42208
rect 8720 42168 8726 42180
rect 16206 42168 16212 42220
rect 16264 42168 16270 42220
rect 16485 42211 16543 42217
rect 16485 42177 16497 42211
rect 16531 42208 16543 42211
rect 17420 42208 17448 42316
rect 17678 42304 17684 42316
rect 17736 42304 17742 42356
rect 17770 42304 17776 42356
rect 17828 42304 17834 42356
rect 18046 42304 18052 42356
rect 18104 42304 18110 42356
rect 18322 42344 18328 42356
rect 18248 42316 18328 42344
rect 17497 42279 17555 42285
rect 17497 42245 17509 42279
rect 17543 42276 17555 42279
rect 17788 42276 17816 42304
rect 17543 42248 17816 42276
rect 17865 42279 17923 42285
rect 17543 42245 17555 42248
rect 17497 42239 17555 42245
rect 17865 42245 17877 42279
rect 17911 42276 17923 42279
rect 18064 42276 18092 42304
rect 18248 42285 18276 42316
rect 18322 42304 18328 42316
rect 18380 42304 18386 42356
rect 19076 42316 19472 42344
rect 17911 42248 18092 42276
rect 18233 42279 18291 42285
rect 17911 42245 17923 42248
rect 17865 42239 17923 42245
rect 18233 42245 18245 42279
rect 18279 42245 18291 42279
rect 18233 42239 18291 42245
rect 18414 42236 18420 42288
rect 18472 42276 18478 42288
rect 18969 42279 19027 42285
rect 18969 42276 18981 42279
rect 18472 42248 18981 42276
rect 18472 42236 18478 42248
rect 18969 42245 18981 42248
rect 19015 42245 19027 42279
rect 18969 42239 19027 42245
rect 16531 42180 17448 42208
rect 16531 42177 16543 42180
rect 16485 42171 16543 42177
rect 18598 42168 18604 42220
rect 18656 42168 18662 42220
rect 18874 42168 18880 42220
rect 18932 42208 18938 42220
rect 19076 42208 19104 42316
rect 19334 42236 19340 42288
rect 19392 42236 19398 42288
rect 19444 42276 19472 42316
rect 19610 42304 19616 42356
rect 19668 42304 19674 42356
rect 19978 42304 19984 42356
rect 20036 42304 20042 42356
rect 20346 42304 20352 42356
rect 20404 42344 20410 42356
rect 20533 42347 20591 42353
rect 20533 42344 20545 42347
rect 20404 42316 20545 42344
rect 20404 42304 20410 42316
rect 20533 42313 20545 42316
rect 20579 42313 20591 42347
rect 20533 42307 20591 42313
rect 20809 42347 20867 42353
rect 20809 42313 20821 42347
rect 20855 42344 20867 42347
rect 20898 42344 20904 42356
rect 20855 42316 20904 42344
rect 20855 42313 20867 42316
rect 20809 42307 20867 42313
rect 20898 42304 20904 42316
rect 20956 42304 20962 42356
rect 22741 42347 22799 42353
rect 22741 42313 22753 42347
rect 22787 42344 22799 42347
rect 23014 42344 23020 42356
rect 22787 42316 23020 42344
rect 22787 42313 22799 42316
rect 22741 42307 22799 42313
rect 23014 42304 23020 42316
rect 23072 42304 23078 42356
rect 23293 42347 23351 42353
rect 23293 42313 23305 42347
rect 23339 42344 23351 42347
rect 24210 42344 24216 42356
rect 23339 42316 24216 42344
rect 23339 42313 23351 42316
rect 23293 42307 23351 42313
rect 24210 42304 24216 42316
rect 24268 42304 24274 42356
rect 19996 42276 20024 42304
rect 19444 42248 20024 42276
rect 20254 42236 20260 42288
rect 20312 42276 20318 42288
rect 22094 42276 22100 42288
rect 20312 42248 22100 42276
rect 20312 42236 20318 42248
rect 22094 42236 22100 42248
rect 22152 42236 22158 42288
rect 22281 42279 22339 42285
rect 22281 42245 22293 42279
rect 22327 42276 22339 42279
rect 23750 42276 23756 42288
rect 22327 42248 23756 42276
rect 22327 42245 22339 42248
rect 22281 42239 22339 42245
rect 23750 42236 23756 42248
rect 23808 42236 23814 42288
rect 18932 42180 19104 42208
rect 18932 42168 18938 42180
rect 19150 42168 19156 42220
rect 19208 42208 19214 42220
rect 19797 42211 19855 42217
rect 19797 42208 19809 42211
rect 19208 42180 19809 42208
rect 19208 42168 19214 42180
rect 19797 42177 19809 42180
rect 19843 42177 19855 42211
rect 19797 42171 19855 42177
rect 19978 42168 19984 42220
rect 20036 42208 20042 42220
rect 20165 42211 20223 42217
rect 20165 42208 20177 42211
rect 20036 42180 20177 42208
rect 20036 42168 20042 42180
rect 20165 42177 20177 42180
rect 20211 42177 20223 42211
rect 20165 42171 20223 42177
rect 20438 42168 20444 42220
rect 20496 42168 20502 42220
rect 20717 42211 20775 42217
rect 20717 42177 20729 42211
rect 20763 42177 20775 42211
rect 20717 42171 20775 42177
rect 20993 42211 21051 42217
rect 20993 42177 21005 42211
rect 21039 42177 21051 42211
rect 20993 42171 21051 42177
rect 21269 42211 21327 42217
rect 21269 42177 21281 42211
rect 21315 42177 21327 42211
rect 21269 42171 21327 42177
rect 21913 42211 21971 42217
rect 21913 42177 21925 42211
rect 21959 42208 21971 42211
rect 21959 42180 22094 42208
rect 21959 42177 21971 42180
rect 21913 42171 21971 42177
rect 2746 42112 4384 42140
rect 4724 42112 7512 42140
rect 474 42032 480 42084
rect 532 42072 538 42084
rect 2746 42072 2774 42112
rect 4356 42081 4384 42112
rect 7834 42100 7840 42152
rect 7892 42140 7898 42152
rect 9033 42143 9091 42149
rect 9033 42140 9045 42143
rect 7892 42112 9045 42140
rect 7892 42100 7898 42112
rect 9033 42109 9045 42112
rect 9079 42109 9091 42143
rect 9033 42103 9091 42109
rect 9766 42100 9772 42152
rect 9824 42140 9830 42152
rect 20732 42140 20760 42171
rect 9824 42112 19932 42140
rect 9824 42100 9830 42112
rect 4341 42075 4399 42081
rect 532 42044 2774 42072
rect 3068 42044 3740 42072
rect 532 42032 538 42044
rect 1302 41964 1308 42016
rect 1360 42004 1366 42016
rect 3068 42004 3096 42044
rect 3712 42013 3740 42044
rect 4341 42041 4353 42075
rect 4387 42041 4399 42075
rect 4341 42035 4399 42041
rect 4522 42032 4528 42084
rect 4580 42072 4586 42084
rect 5902 42072 5908 42084
rect 4580 42044 5908 42072
rect 4580 42032 4586 42044
rect 5902 42032 5908 42044
rect 5960 42032 5966 42084
rect 7745 42075 7803 42081
rect 7745 42041 7757 42075
rect 7791 42072 7803 42075
rect 8202 42072 8208 42084
rect 7791 42044 8208 42072
rect 7791 42041 7803 42044
rect 7745 42035 7803 42041
rect 8202 42032 8208 42044
rect 8260 42032 8266 42084
rect 16025 42075 16083 42081
rect 16025 42041 16037 42075
rect 16071 42072 16083 42075
rect 16390 42072 16396 42084
rect 16071 42044 16396 42072
rect 16071 42041 16083 42044
rect 16025 42035 16083 42041
rect 16390 42032 16396 42044
rect 16448 42032 16454 42084
rect 16942 42032 16948 42084
rect 17000 42032 17006 42084
rect 17310 42032 17316 42084
rect 17368 42032 17374 42084
rect 18414 42032 18420 42084
rect 18472 42032 18478 42084
rect 19904 42016 19932 42112
rect 19996 42112 20760 42140
rect 19996 42081 20024 42112
rect 19981 42075 20039 42081
rect 19981 42041 19993 42075
rect 20027 42041 20039 42075
rect 19981 42035 20039 42041
rect 20257 42075 20315 42081
rect 20257 42041 20269 42075
rect 20303 42072 20315 42075
rect 21008 42072 21036 42171
rect 20303 42044 21036 42072
rect 20303 42041 20315 42044
rect 20257 42035 20315 42041
rect 1360 41976 3096 42004
rect 3697 42007 3755 42013
rect 1360 41964 1366 41976
rect 3697 41973 3709 42007
rect 3743 41973 3755 42007
rect 3697 41967 3755 41973
rect 4798 41964 4804 42016
rect 4856 41964 4862 42016
rect 5718 41964 5724 42016
rect 5776 41964 5782 42016
rect 5997 42007 6055 42013
rect 5997 41973 6009 42007
rect 6043 42004 6055 42007
rect 6270 42004 6276 42016
rect 6043 41976 6276 42004
rect 6043 41973 6055 41976
rect 5997 41967 6055 41973
rect 6270 41964 6276 41976
rect 6328 41964 6334 42016
rect 6730 41964 6736 42016
rect 6788 41964 6794 42016
rect 7190 41964 7196 42016
rect 7248 42004 7254 42016
rect 7285 42007 7343 42013
rect 7285 42004 7297 42007
rect 7248 41976 7297 42004
rect 7248 41964 7254 41976
rect 7285 41973 7297 41976
rect 7331 42004 7343 42007
rect 7374 42004 7380 42016
rect 7331 41976 7380 42004
rect 7331 41973 7343 41976
rect 7285 41967 7343 41973
rect 7374 41964 7380 41976
rect 7432 41964 7438 42016
rect 8021 42007 8079 42013
rect 8021 41973 8033 42007
rect 8067 42004 8079 42007
rect 8294 42004 8300 42016
rect 8067 41976 8300 42004
rect 8067 41973 8079 41976
rect 8021 41967 8079 41973
rect 8294 41964 8300 41976
rect 8352 41964 8358 42016
rect 9030 41964 9036 42016
rect 9088 42004 9094 42016
rect 10045 42007 10103 42013
rect 10045 42004 10057 42007
rect 9088 41976 10057 42004
rect 9088 41964 9094 41976
rect 10045 41973 10057 41976
rect 10091 41973 10103 42007
rect 10045 41967 10103 41973
rect 16298 41964 16304 42016
rect 16356 41964 16362 42016
rect 17586 41964 17592 42016
rect 17644 41964 17650 42016
rect 17954 41964 17960 42016
rect 18012 41964 18018 42016
rect 18690 41964 18696 42016
rect 18748 41964 18754 42016
rect 19058 41964 19064 42016
rect 19116 41964 19122 42016
rect 19334 41964 19340 42016
rect 19392 42004 19398 42016
rect 19429 42007 19487 42013
rect 19429 42004 19441 42007
rect 19392 41976 19441 42004
rect 19392 41964 19398 41976
rect 19429 41973 19441 41976
rect 19475 41973 19487 42007
rect 19429 41967 19487 41973
rect 19886 41964 19892 42016
rect 19944 41964 19950 42016
rect 21284 42004 21312 42171
rect 22066 42140 22094 42180
rect 22462 42168 22468 42220
rect 22520 42168 22526 42220
rect 22554 42168 22560 42220
rect 22612 42208 22618 42220
rect 23017 42211 23075 42217
rect 23017 42208 23029 42211
rect 22612 42180 23029 42208
rect 22612 42168 22618 42180
rect 23017 42177 23029 42180
rect 23063 42177 23075 42211
rect 23017 42171 23075 42177
rect 23566 42168 23572 42220
rect 23624 42168 23630 42220
rect 23937 42211 23995 42217
rect 23937 42177 23949 42211
rect 23983 42208 23995 42211
rect 24026 42208 24032 42220
rect 23983 42180 24032 42208
rect 23983 42177 23995 42180
rect 23937 42171 23995 42177
rect 24026 42168 24032 42180
rect 24084 42168 24090 42220
rect 24118 42168 24124 42220
rect 24176 42168 24182 42220
rect 24489 42211 24547 42217
rect 24489 42177 24501 42211
rect 24535 42208 24547 42211
rect 25038 42208 25044 42220
rect 24535 42180 25044 42208
rect 24535 42177 24547 42180
rect 24489 42171 24547 42177
rect 25038 42168 25044 42180
rect 25096 42168 25102 42220
rect 23750 42140 23756 42152
rect 22066 42112 23756 42140
rect 23750 42100 23756 42112
rect 23808 42100 23814 42152
rect 25590 42100 25596 42152
rect 25648 42100 25654 42152
rect 21545 42075 21603 42081
rect 21545 42041 21557 42075
rect 21591 42072 21603 42075
rect 25608 42072 25636 42100
rect 21591 42044 25636 42072
rect 21591 42041 21603 42044
rect 21545 42035 21603 42041
rect 25682 42004 25688 42016
rect 21284 41976 25688 42004
rect 25682 41964 25688 41976
rect 25740 41964 25746 42016
rect 1104 41914 24840 41936
rect 1104 41862 3917 41914
rect 3969 41862 3981 41914
rect 4033 41862 4045 41914
rect 4097 41862 4109 41914
rect 4161 41862 4173 41914
rect 4225 41862 9851 41914
rect 9903 41862 9915 41914
rect 9967 41862 9979 41914
rect 10031 41862 10043 41914
rect 10095 41862 10107 41914
rect 10159 41862 15785 41914
rect 15837 41862 15849 41914
rect 15901 41862 15913 41914
rect 15965 41862 15977 41914
rect 16029 41862 16041 41914
rect 16093 41862 21719 41914
rect 21771 41862 21783 41914
rect 21835 41862 21847 41914
rect 21899 41862 21911 41914
rect 21963 41862 21975 41914
rect 22027 41862 24840 41914
rect 1104 41840 24840 41862
rect 3421 41803 3479 41809
rect 3421 41769 3433 41803
rect 3467 41800 3479 41803
rect 3786 41800 3792 41812
rect 3467 41772 3792 41800
rect 3467 41769 3479 41772
rect 3421 41763 3479 41769
rect 3786 41760 3792 41772
rect 3844 41760 3850 41812
rect 3878 41760 3884 41812
rect 3936 41800 3942 41812
rect 4525 41803 4583 41809
rect 4525 41800 4537 41803
rect 3936 41772 4537 41800
rect 3936 41760 3942 41772
rect 4525 41769 4537 41772
rect 4571 41769 4583 41803
rect 4525 41763 4583 41769
rect 4614 41760 4620 41812
rect 4672 41800 4678 41812
rect 4985 41803 5043 41809
rect 4985 41800 4997 41803
rect 4672 41772 4997 41800
rect 4672 41760 4678 41772
rect 4985 41769 4997 41772
rect 5031 41769 5043 41803
rect 4985 41763 5043 41769
rect 5442 41760 5448 41812
rect 5500 41760 5506 41812
rect 5718 41760 5724 41812
rect 5776 41760 5782 41812
rect 5810 41760 5816 41812
rect 5868 41760 5874 41812
rect 5994 41760 6000 41812
rect 6052 41800 6058 41812
rect 6181 41803 6239 41809
rect 6181 41800 6193 41803
rect 6052 41772 6193 41800
rect 6052 41760 6058 41772
rect 6181 41769 6193 41772
rect 6227 41769 6239 41803
rect 6181 41763 6239 41769
rect 6362 41760 6368 41812
rect 6420 41800 6426 41812
rect 6549 41803 6607 41809
rect 6549 41800 6561 41803
rect 6420 41772 6561 41800
rect 6420 41760 6426 41772
rect 6549 41769 6561 41772
rect 6595 41769 6607 41803
rect 6549 41763 6607 41769
rect 6730 41760 6736 41812
rect 6788 41760 6794 41812
rect 6822 41760 6828 41812
rect 6880 41760 6886 41812
rect 7282 41760 7288 41812
rect 7340 41760 7346 41812
rect 7558 41760 7564 41812
rect 7616 41800 7622 41812
rect 7745 41803 7803 41809
rect 7745 41800 7757 41803
rect 7616 41772 7757 41800
rect 7616 41760 7622 41772
rect 7745 41769 7757 41772
rect 7791 41769 7803 41803
rect 7745 41763 7803 41769
rect 7926 41760 7932 41812
rect 7984 41760 7990 41812
rect 8202 41760 8208 41812
rect 8260 41760 8266 41812
rect 8294 41760 8300 41812
rect 8352 41760 8358 41812
rect 8386 41760 8392 41812
rect 8444 41760 8450 41812
rect 8941 41803 8999 41809
rect 8941 41769 8953 41803
rect 8987 41800 8999 41803
rect 9122 41800 9128 41812
rect 8987 41772 9128 41800
rect 8987 41769 8999 41772
rect 8941 41763 8999 41769
rect 9122 41760 9128 41772
rect 9180 41760 9186 41812
rect 11330 41800 11336 41812
rect 9232 41772 11336 41800
rect 4709 41735 4767 41741
rect 2746 41704 4660 41732
rect 2225 41667 2283 41673
rect 2225 41633 2237 41667
rect 2271 41664 2283 41667
rect 2746 41664 2774 41704
rect 2271 41636 2774 41664
rect 3237 41667 3295 41673
rect 2271 41633 2283 41636
rect 2225 41627 2283 41633
rect 3237 41633 3249 41667
rect 3283 41664 3295 41667
rect 3283 41636 4108 41664
rect 3283 41633 3295 41636
rect 3237 41627 3295 41633
rect 750 41556 756 41608
rect 808 41596 814 41608
rect 3605 41599 3663 41605
rect 808 41568 3372 41596
rect 808 41556 814 41568
rect 1397 41531 1455 41537
rect 1397 41497 1409 41531
rect 1443 41497 1455 41531
rect 1397 41491 1455 41497
rect 1412 41460 1440 41491
rect 2406 41488 2412 41540
rect 2464 41488 2470 41540
rect 2774 41460 2780 41472
rect 1412 41432 2780 41460
rect 2774 41420 2780 41432
rect 2832 41420 2838 41472
rect 3344 41460 3372 41568
rect 3605 41565 3617 41599
rect 3651 41596 3663 41599
rect 3694 41596 3700 41608
rect 3651 41568 3700 41596
rect 3651 41565 3663 41568
rect 3605 41559 3663 41565
rect 3694 41556 3700 41568
rect 3752 41556 3758 41608
rect 3878 41556 3884 41608
rect 3936 41556 3942 41608
rect 3973 41463 4031 41469
rect 3973 41460 3985 41463
rect 3344 41432 3985 41460
rect 3973 41429 3985 41432
rect 4019 41429 4031 41463
rect 4080 41460 4108 41636
rect 4522 41624 4528 41676
rect 4580 41664 4586 41676
rect 4632 41664 4660 41704
rect 4709 41701 4721 41735
rect 4755 41732 4767 41735
rect 4755 41704 5672 41732
rect 4755 41701 4767 41704
rect 4709 41695 4767 41701
rect 4580 41636 4660 41664
rect 4580 41624 4586 41636
rect 4338 41556 4344 41608
rect 4396 41556 4402 41608
rect 4614 41556 4620 41608
rect 4672 41596 4678 41608
rect 4893 41599 4951 41605
rect 4893 41596 4905 41599
rect 4672 41568 4905 41596
rect 4672 41556 4678 41568
rect 4893 41565 4905 41568
rect 4939 41565 4951 41599
rect 4893 41559 4951 41565
rect 5166 41556 5172 41608
rect 5224 41556 5230 41608
rect 5644 41605 5672 41704
rect 5736 41664 5764 41760
rect 6748 41664 6776 41760
rect 5736 41636 6408 41664
rect 6748 41636 7512 41664
rect 5629 41599 5687 41605
rect 5629 41565 5641 41599
rect 5675 41565 5687 41599
rect 5629 41559 5687 41565
rect 5994 41556 6000 41608
rect 6052 41556 6058 41608
rect 6270 41556 6276 41608
rect 6328 41556 6334 41608
rect 6380 41605 6408 41636
rect 6365 41599 6423 41605
rect 6365 41565 6377 41599
rect 6411 41565 6423 41599
rect 6365 41559 6423 41565
rect 6730 41556 6736 41608
rect 6788 41556 6794 41608
rect 7484 41605 7512 41636
rect 7944 41605 7972 41760
rect 7009 41599 7067 41605
rect 7009 41565 7021 41599
rect 7055 41565 7067 41599
rect 7009 41559 7067 41565
rect 7469 41599 7527 41605
rect 7469 41565 7481 41599
rect 7515 41565 7527 41599
rect 7469 41559 7527 41565
rect 7929 41599 7987 41605
rect 7929 41565 7941 41599
rect 7975 41565 7987 41599
rect 8220 41596 8248 41760
rect 8312 41664 8340 41760
rect 8570 41692 8576 41744
rect 8628 41732 8634 41744
rect 9232 41732 9260 41772
rect 11330 41760 11336 41772
rect 11388 41760 11394 41812
rect 16298 41760 16304 41812
rect 16356 41760 16362 41812
rect 16390 41760 16396 41812
rect 16448 41760 16454 41812
rect 16666 41760 16672 41812
rect 16724 41800 16730 41812
rect 16724 41772 18736 41800
rect 16724 41760 16730 41772
rect 8628 41704 9260 41732
rect 8628 41692 8634 41704
rect 8312 41636 8524 41664
rect 8297 41599 8355 41605
rect 8297 41596 8309 41599
rect 8220 41568 8309 41596
rect 7929 41559 7987 41565
rect 8297 41565 8309 41568
rect 8343 41565 8355 41599
rect 8496 41596 8524 41636
rect 9048 41636 9674 41664
rect 8565 41599 8623 41605
rect 8565 41596 8577 41599
rect 8496 41568 8577 41596
rect 8297 41559 8355 41565
rect 8565 41565 8577 41568
rect 8611 41565 8623 41599
rect 8565 41559 8623 41565
rect 4154 41488 4160 41540
rect 4212 41528 4218 41540
rect 4798 41528 4804 41540
rect 4212 41500 4804 41528
rect 4212 41488 4218 41500
rect 4798 41488 4804 41500
rect 4856 41488 4862 41540
rect 5902 41488 5908 41540
rect 5960 41528 5966 41540
rect 6178 41528 6184 41540
rect 5960 41500 6184 41528
rect 5960 41488 5966 41500
rect 6178 41488 6184 41500
rect 6236 41488 6242 41540
rect 6288 41528 6316 41556
rect 7024 41528 7052 41559
rect 9048 41528 9076 41636
rect 9125 41599 9183 41605
rect 9125 41565 9137 41599
rect 9171 41596 9183 41599
rect 9171 41568 9444 41596
rect 9171 41565 9183 41568
rect 9125 41559 9183 41565
rect 6288 41500 7052 41528
rect 7392 41500 9076 41528
rect 7392 41460 7420 41500
rect 9416 41472 9444 41568
rect 4080 41432 7420 41460
rect 3973 41423 4031 41429
rect 7466 41420 7472 41472
rect 7524 41460 7530 41472
rect 8113 41463 8171 41469
rect 8113 41460 8125 41463
rect 7524 41432 8125 41460
rect 7524 41420 7530 41432
rect 8113 41429 8125 41432
rect 8159 41429 8171 41463
rect 8113 41423 8171 41429
rect 9398 41420 9404 41472
rect 9456 41420 9462 41472
rect 9646 41460 9674 41636
rect 9766 41556 9772 41608
rect 9824 41556 9830 41608
rect 16117 41599 16175 41605
rect 10027 41569 10085 41575
rect 10027 41535 10039 41569
rect 10073 41566 10085 41569
rect 10073 41540 10088 41566
rect 16117 41565 16129 41599
rect 16163 41596 16175 41599
rect 16316 41596 16344 41760
rect 16163 41568 16344 41596
rect 16408 41596 16436 41760
rect 18601 41735 18659 41741
rect 18601 41701 18613 41735
rect 18647 41701 18659 41735
rect 18708 41732 18736 41772
rect 18874 41760 18880 41812
rect 18932 41760 18938 41812
rect 19334 41760 19340 41812
rect 19392 41800 19398 41812
rect 19702 41800 19708 41812
rect 19392 41772 19708 41800
rect 19392 41760 19398 41772
rect 19702 41760 19708 41772
rect 19760 41760 19766 41812
rect 19797 41803 19855 41809
rect 19797 41769 19809 41803
rect 19843 41800 19855 41803
rect 19978 41800 19984 41812
rect 19843 41772 19984 41800
rect 19843 41769 19855 41772
rect 19797 41763 19855 41769
rect 19978 41760 19984 41772
rect 20036 41760 20042 41812
rect 20073 41803 20131 41809
rect 20073 41769 20085 41803
rect 20119 41800 20131 41803
rect 20438 41800 20444 41812
rect 20119 41772 20444 41800
rect 20119 41769 20131 41772
rect 20073 41763 20131 41769
rect 20438 41760 20444 41772
rect 20496 41760 20502 41812
rect 20990 41760 20996 41812
rect 21048 41800 21054 41812
rect 21269 41803 21327 41809
rect 21048 41772 21220 41800
rect 21048 41760 21054 41772
rect 20717 41735 20775 41741
rect 18708 41704 19656 41732
rect 18601 41695 18659 41701
rect 18616 41664 18644 41695
rect 18616 41636 19472 41664
rect 16485 41599 16543 41605
rect 16485 41596 16497 41599
rect 16408 41568 16497 41596
rect 16163 41565 16175 41568
rect 16117 41559 16175 41565
rect 16485 41565 16497 41568
rect 16531 41565 16543 41599
rect 16485 41559 16543 41565
rect 18509 41599 18567 41605
rect 18509 41565 18521 41599
rect 18555 41596 18567 41599
rect 18690 41596 18696 41608
rect 18555 41568 18696 41596
rect 18555 41565 18567 41568
rect 18509 41559 18567 41565
rect 18690 41556 18696 41568
rect 18748 41556 18754 41608
rect 18785 41599 18843 41605
rect 18785 41565 18797 41599
rect 18831 41565 18843 41599
rect 18785 41559 18843 41565
rect 19061 41599 19119 41605
rect 19061 41565 19073 41599
rect 19107 41596 19119 41599
rect 19334 41596 19340 41608
rect 19107 41568 19340 41596
rect 19107 41565 19119 41568
rect 19061 41559 19119 41565
rect 10027 41529 10048 41535
rect 10042 41488 10048 41529
rect 10100 41488 10106 41540
rect 10704 41500 12434 41528
rect 10704 41460 10732 41500
rect 9646 41432 10732 41460
rect 10778 41420 10784 41472
rect 10836 41420 10842 41472
rect 12406 41460 12434 41500
rect 15102 41488 15108 41540
rect 15160 41528 15166 41540
rect 18800 41528 18828 41559
rect 19334 41556 19340 41568
rect 19392 41556 19398 41608
rect 19444 41605 19472 41636
rect 19429 41599 19487 41605
rect 19429 41565 19441 41599
rect 19475 41565 19487 41599
rect 19429 41559 19487 41565
rect 19518 41556 19524 41608
rect 19576 41556 19582 41608
rect 19536 41528 19564 41556
rect 15160 41500 16620 41528
rect 18800 41500 19564 41528
rect 19628 41528 19656 41704
rect 19720 41704 20668 41732
rect 19720 41605 19748 41704
rect 19794 41624 19800 41676
rect 19852 41664 19858 41676
rect 20640 41664 20668 41704
rect 20717 41701 20729 41735
rect 20763 41732 20775 41735
rect 21192 41732 21220 41772
rect 21269 41769 21281 41803
rect 21315 41800 21327 41803
rect 21450 41800 21456 41812
rect 21315 41772 21456 41800
rect 21315 41769 21327 41772
rect 21269 41763 21327 41769
rect 21450 41760 21456 41772
rect 21508 41760 21514 41812
rect 21726 41760 21732 41812
rect 21784 41760 21790 41812
rect 22278 41760 22284 41812
rect 22336 41760 22342 41812
rect 23569 41803 23627 41809
rect 23569 41769 23581 41803
rect 23615 41800 23627 41803
rect 23658 41800 23664 41812
rect 23615 41772 23664 41800
rect 23615 41769 23627 41772
rect 23569 41763 23627 41769
rect 23658 41760 23664 41772
rect 23716 41760 23722 41812
rect 23934 41760 23940 41812
rect 23992 41760 23998 41812
rect 24578 41760 24584 41812
rect 24636 41760 24642 41812
rect 20763 41704 21128 41732
rect 21192 41704 21404 41732
rect 20763 41701 20775 41704
rect 20717 41695 20775 41701
rect 21100 41664 21128 41704
rect 21376 41664 21404 41704
rect 21542 41692 21548 41744
rect 21600 41732 21606 41744
rect 21821 41735 21879 41741
rect 21821 41732 21833 41735
rect 21600 41704 21833 41732
rect 21600 41692 21606 41704
rect 21821 41701 21833 41704
rect 21867 41701 21879 41735
rect 21821 41695 21879 41701
rect 23017 41735 23075 41741
rect 23017 41701 23029 41735
rect 23063 41732 23075 41735
rect 24596 41732 24624 41760
rect 23063 41704 24624 41732
rect 23063 41701 23075 41704
rect 23017 41695 23075 41701
rect 19852 41636 20576 41664
rect 20640 41636 21036 41664
rect 21100 41636 21312 41664
rect 21376 41636 21588 41664
rect 19852 41624 19858 41636
rect 19705 41599 19763 41605
rect 19705 41565 19717 41599
rect 19751 41565 19763 41599
rect 19705 41559 19763 41565
rect 19886 41556 19892 41608
rect 19944 41596 19950 41608
rect 20548 41605 20576 41636
rect 19981 41599 20039 41605
rect 19981 41596 19993 41599
rect 19944 41568 19993 41596
rect 19944 41556 19950 41568
rect 19981 41565 19993 41568
rect 20027 41565 20039 41599
rect 19981 41559 20039 41565
rect 20257 41599 20315 41605
rect 20257 41565 20269 41599
rect 20303 41565 20315 41599
rect 20257 41559 20315 41565
rect 20533 41599 20591 41605
rect 20533 41565 20545 41599
rect 20579 41565 20591 41599
rect 20533 41559 20591 41565
rect 20272 41528 20300 41559
rect 20622 41556 20628 41608
rect 20680 41596 20686 41608
rect 20901 41599 20959 41605
rect 20901 41596 20913 41599
rect 20680 41568 20913 41596
rect 20680 41556 20686 41568
rect 20901 41565 20913 41568
rect 20947 41565 20959 41599
rect 20901 41559 20959 41565
rect 19628 41500 20300 41528
rect 21008 41528 21036 41636
rect 21174 41556 21180 41608
rect 21232 41556 21238 41608
rect 21284 41596 21312 41636
rect 21560 41605 21588 41636
rect 21453 41599 21511 41605
rect 21453 41596 21465 41599
rect 21284 41568 21465 41596
rect 21453 41565 21465 41568
rect 21499 41565 21511 41599
rect 21453 41559 21511 41565
rect 21545 41599 21603 41605
rect 21545 41565 21557 41599
rect 21591 41565 21603 41599
rect 21545 41559 21603 41565
rect 22002 41556 22008 41608
rect 22060 41556 22066 41608
rect 21008 41500 21128 41528
rect 15160 41488 15166 41500
rect 15194 41460 15200 41472
rect 12406 41432 15200 41460
rect 15194 41420 15200 41432
rect 15252 41420 15258 41472
rect 16206 41420 16212 41472
rect 16264 41420 16270 41472
rect 16592 41469 16620 41500
rect 16577 41463 16635 41469
rect 16577 41429 16589 41463
rect 16623 41429 16635 41463
rect 16577 41423 16635 41429
rect 18322 41420 18328 41472
rect 18380 41420 18386 41472
rect 19150 41420 19156 41472
rect 19208 41460 19214 41472
rect 19245 41463 19303 41469
rect 19245 41460 19257 41463
rect 19208 41432 19257 41460
rect 19208 41420 19214 41432
rect 19245 41429 19257 41432
rect 19291 41429 19303 41463
rect 19245 41423 19303 41429
rect 19521 41463 19579 41469
rect 19521 41429 19533 41463
rect 19567 41460 19579 41463
rect 20254 41460 20260 41472
rect 19567 41432 20260 41460
rect 19567 41429 19579 41432
rect 19521 41423 19579 41429
rect 20254 41420 20260 41432
rect 20312 41420 20318 41472
rect 20346 41420 20352 41472
rect 20404 41420 20410 41472
rect 20438 41420 20444 41472
rect 20496 41460 20502 41472
rect 20993 41463 21051 41469
rect 20993 41460 21005 41463
rect 20496 41432 21005 41460
rect 20496 41420 20502 41432
rect 20993 41429 21005 41432
rect 21039 41429 21051 41463
rect 21100 41460 21128 41500
rect 21634 41488 21640 41540
rect 21692 41528 21698 41540
rect 22189 41531 22247 41537
rect 22189 41528 22201 41531
rect 21692 41500 22201 41528
rect 21692 41488 21698 41500
rect 22189 41497 22201 41500
rect 22235 41497 22247 41531
rect 22189 41491 22247 41497
rect 22741 41531 22799 41537
rect 22741 41497 22753 41531
rect 22787 41497 22799 41531
rect 22741 41491 22799 41497
rect 22278 41460 22284 41472
rect 21100 41432 22284 41460
rect 20993 41423 21051 41429
rect 22278 41420 22284 41432
rect 22336 41420 22342 41472
rect 22756 41460 22784 41491
rect 23290 41488 23296 41540
rect 23348 41488 23354 41540
rect 23842 41488 23848 41540
rect 23900 41488 23906 41540
rect 24486 41460 24492 41472
rect 22756 41432 24492 41460
rect 24486 41420 24492 41432
rect 24544 41420 24550 41472
rect 1104 41370 25000 41392
rect 1104 41318 6884 41370
rect 6936 41318 6948 41370
rect 7000 41318 7012 41370
rect 7064 41318 7076 41370
rect 7128 41318 7140 41370
rect 7192 41318 12818 41370
rect 12870 41318 12882 41370
rect 12934 41318 12946 41370
rect 12998 41318 13010 41370
rect 13062 41318 13074 41370
rect 13126 41318 18752 41370
rect 18804 41318 18816 41370
rect 18868 41318 18880 41370
rect 18932 41318 18944 41370
rect 18996 41318 19008 41370
rect 19060 41318 24686 41370
rect 24738 41318 24750 41370
rect 24802 41318 24814 41370
rect 24866 41318 24878 41370
rect 24930 41318 24942 41370
rect 24994 41318 25000 41370
rect 1104 41296 25000 41318
rect 198 41216 204 41268
rect 256 41256 262 41268
rect 4154 41256 4160 41268
rect 256 41228 4160 41256
rect 256 41216 262 41228
rect 4154 41216 4160 41228
rect 4212 41216 4218 41268
rect 4709 41259 4767 41265
rect 4709 41225 4721 41259
rect 4755 41256 4767 41259
rect 4798 41256 4804 41268
rect 4755 41228 4804 41256
rect 4755 41225 4767 41228
rect 4709 41219 4767 41225
rect 4798 41216 4804 41228
rect 4856 41216 4862 41268
rect 5258 41216 5264 41268
rect 5316 41216 5322 41268
rect 5534 41216 5540 41268
rect 5592 41216 5598 41268
rect 5810 41216 5816 41268
rect 5868 41216 5874 41268
rect 6365 41259 6423 41265
rect 6365 41256 6377 41259
rect 5920 41228 6377 41256
rect 1857 41191 1915 41197
rect 1857 41157 1869 41191
rect 1903 41188 1915 41191
rect 5920 41188 5948 41228
rect 6365 41225 6377 41228
rect 6411 41225 6423 41259
rect 6365 41219 6423 41225
rect 6546 41216 6552 41268
rect 6604 41256 6610 41268
rect 6917 41259 6975 41265
rect 6917 41256 6929 41259
rect 6604 41228 6929 41256
rect 6604 41216 6610 41228
rect 6917 41225 6929 41228
rect 6963 41225 6975 41259
rect 6917 41219 6975 41225
rect 7834 41216 7840 41268
rect 7892 41256 7898 41268
rect 8202 41256 8208 41268
rect 7892 41228 8208 41256
rect 7892 41216 7898 41228
rect 8202 41216 8208 41228
rect 8260 41216 8266 41268
rect 9214 41216 9220 41268
rect 9272 41256 9278 41268
rect 9493 41259 9551 41265
rect 9493 41256 9505 41259
rect 9272 41228 9505 41256
rect 9272 41216 9278 41228
rect 9493 41225 9505 41228
rect 9539 41225 9551 41259
rect 9493 41219 9551 41225
rect 9766 41216 9772 41268
rect 9824 41256 9830 41268
rect 18601 41259 18659 41265
rect 9824 41228 12434 41256
rect 9824 41216 9830 41228
rect 1903 41160 4182 41188
rect 1903 41157 1915 41160
rect 1857 41151 1915 41157
rect 1489 41123 1547 41129
rect 1489 41089 1501 41123
rect 1535 41089 1547 41123
rect 1489 41083 1547 41089
rect 1504 41052 1532 41083
rect 2130 41080 2136 41132
rect 2188 41120 2194 41132
rect 2225 41123 2283 41129
rect 2225 41120 2237 41123
rect 2188 41092 2237 41120
rect 2188 41080 2194 41092
rect 2225 41089 2237 41092
rect 2271 41089 2283 41123
rect 2225 41083 2283 41089
rect 2314 41080 2320 41132
rect 2372 41080 2378 41132
rect 2682 41080 2688 41132
rect 2740 41120 2746 41132
rect 3053 41123 3111 41129
rect 3053 41120 3065 41123
rect 2740 41092 3065 41120
rect 2740 41080 2746 41092
rect 3053 41089 3065 41092
rect 3099 41089 3111 41123
rect 3053 41083 3111 41089
rect 3510 41080 3516 41132
rect 3568 41120 3574 41132
rect 3603 41123 3661 41129
rect 3603 41120 3615 41123
rect 3568 41092 3615 41120
rect 3568 41080 3574 41092
rect 3603 41089 3615 41092
rect 3649 41089 3661 41123
rect 4154 41120 4182 41160
rect 4356 41160 5948 41188
rect 6012 41160 12112 41188
rect 4356 41120 4384 41160
rect 4154 41092 4384 41120
rect 4893 41123 4951 41129
rect 3603 41083 3661 41089
rect 4893 41089 4905 41123
rect 4939 41120 4951 41123
rect 5074 41120 5080 41132
rect 4939 41092 5080 41120
rect 4939 41089 4951 41092
rect 4893 41083 4951 41089
rect 5074 41080 5080 41092
rect 5132 41080 5138 41132
rect 5169 41123 5227 41129
rect 5169 41089 5181 41123
rect 5215 41089 5227 41123
rect 5169 41083 5227 41089
rect 2958 41052 2964 41064
rect 1504 41024 2964 41052
rect 2958 41012 2964 41024
rect 3016 41012 3022 41064
rect 3329 41055 3387 41061
rect 3329 41052 3341 41055
rect 3252 41024 3341 41052
rect 3252 40996 3280 41024
rect 3329 41021 3341 41024
rect 3375 41021 3387 41055
rect 3329 41015 3387 41021
rect 4430 41012 4436 41064
rect 4488 41012 4494 41064
rect 4706 41012 4712 41064
rect 4764 41052 4770 41064
rect 5184 41052 5212 41083
rect 5442 41080 5448 41132
rect 5500 41080 5506 41132
rect 5534 41080 5540 41132
rect 5592 41120 5598 41132
rect 6012 41129 6040 41160
rect 5721 41123 5779 41129
rect 5721 41120 5733 41123
rect 5592 41092 5733 41120
rect 5592 41080 5598 41092
rect 5721 41089 5733 41092
rect 5767 41089 5779 41123
rect 5721 41083 5779 41089
rect 5997 41123 6055 41129
rect 5997 41089 6009 41123
rect 6043 41089 6055 41123
rect 5997 41083 6055 41089
rect 6546 41080 6552 41132
rect 6604 41080 6610 41132
rect 6825 41123 6883 41129
rect 6825 41089 6837 41123
rect 6871 41089 6883 41123
rect 6825 41083 6883 41089
rect 7101 41123 7159 41129
rect 7101 41089 7113 41123
rect 7147 41120 7159 41123
rect 7374 41120 7380 41132
rect 7147 41092 7380 41120
rect 7147 41089 7159 41092
rect 7101 41083 7159 41089
rect 4764 41024 5212 41052
rect 4764 41012 4770 41024
rect 6270 41012 6276 41064
rect 6328 41012 6334 41064
rect 6362 41012 6368 41064
rect 6420 41052 6426 41064
rect 6840 41052 6868 41083
rect 7374 41080 7380 41092
rect 7432 41080 7438 41132
rect 7929 41123 7987 41129
rect 7929 41089 7941 41123
rect 7975 41120 7987 41123
rect 8110 41120 8116 41132
rect 7975 41092 8116 41120
rect 7975 41089 7987 41092
rect 7929 41083 7987 41089
rect 8110 41080 8116 41092
rect 8168 41080 8174 41132
rect 8202 41080 8208 41132
rect 8260 41080 8266 41132
rect 9582 41080 9588 41132
rect 9640 41080 9646 41132
rect 9674 41080 9680 41132
rect 9732 41080 9738 41132
rect 9858 41080 9864 41132
rect 9916 41120 9922 41132
rect 10045 41123 10103 41129
rect 10045 41120 10057 41123
rect 9916 41092 10057 41120
rect 9916 41080 9922 41092
rect 10045 41089 10057 41092
rect 10091 41089 10103 41123
rect 10318 41120 10324 41132
rect 10279 41092 10324 41120
rect 10045 41083 10103 41089
rect 10318 41080 10324 41092
rect 10376 41080 10382 41132
rect 6420 41024 6868 41052
rect 6420 41012 6426 41024
rect 1670 40944 1676 40996
rect 1728 40944 1734 40996
rect 3234 40944 3240 40996
rect 3292 40944 3298 40996
rect 4341 40987 4399 40993
rect 4341 40984 4353 40987
rect 3988 40956 4353 40984
rect 3786 40876 3792 40928
rect 3844 40916 3850 40928
rect 3988 40916 4016 40956
rect 4341 40953 4353 40956
rect 4387 40953 4399 40987
rect 4448 40984 4476 41012
rect 4985 40987 5043 40993
rect 4985 40984 4997 40987
rect 4448 40956 4997 40984
rect 4341 40947 4399 40953
rect 4985 40953 4997 40956
rect 5031 40953 5043 40987
rect 4985 40947 5043 40953
rect 5994 40944 6000 40996
rect 6052 40944 6058 40996
rect 6288 40984 6316 41012
rect 6641 40987 6699 40993
rect 6641 40984 6653 40987
rect 6288 40956 6653 40984
rect 6641 40953 6653 40956
rect 6687 40953 6699 40987
rect 6641 40947 6699 40953
rect 7745 40987 7803 40993
rect 7745 40953 7757 40987
rect 7791 40984 7803 40987
rect 9600 40984 9628 41080
rect 7791 40956 9628 40984
rect 7791 40953 7803 40956
rect 7745 40947 7803 40953
rect 3844 40888 4016 40916
rect 6012 40916 6040 40944
rect 8021 40919 8079 40925
rect 8021 40916 8033 40919
rect 6012 40888 8033 40916
rect 3844 40876 3850 40888
rect 8021 40885 8033 40888
rect 8067 40885 8079 40919
rect 8021 40879 8079 40885
rect 9122 40876 9128 40928
rect 9180 40916 9186 40928
rect 9876 40916 9904 41080
rect 10870 40944 10876 40996
rect 10928 40984 10934 40996
rect 11701 40987 11759 40993
rect 11701 40984 11713 40987
rect 10928 40956 11713 40984
rect 10928 40944 10934 40956
rect 11701 40953 11713 40956
rect 11747 40953 11759 40987
rect 12084 40984 12112 41160
rect 12406 41052 12434 41228
rect 18601 41225 18613 41259
rect 18647 41256 18659 41259
rect 19610 41256 19616 41268
rect 18647 41228 19616 41256
rect 18647 41225 18659 41228
rect 18601 41219 18659 41225
rect 19610 41216 19616 41228
rect 19668 41216 19674 41268
rect 20346 41256 20352 41268
rect 19996 41228 20352 41256
rect 18969 41191 19027 41197
rect 18969 41157 18981 41191
rect 19015 41188 19027 41191
rect 19150 41188 19156 41200
rect 19015 41160 19156 41188
rect 19015 41157 19027 41160
rect 18969 41151 19027 41157
rect 19150 41148 19156 41160
rect 19208 41148 19214 41200
rect 18506 41080 18512 41132
rect 18564 41120 18570 41132
rect 18785 41123 18843 41129
rect 18785 41120 18797 41123
rect 18564 41092 18797 41120
rect 18564 41080 18570 41092
rect 18785 41089 18797 41092
rect 18831 41089 18843 41123
rect 18785 41083 18843 41089
rect 19613 41123 19671 41129
rect 19613 41089 19625 41123
rect 19659 41120 19671 41123
rect 19996 41120 20024 41228
rect 20346 41216 20352 41228
rect 20404 41216 20410 41268
rect 20441 41259 20499 41265
rect 20441 41225 20453 41259
rect 20487 41256 20499 41259
rect 20622 41256 20628 41268
rect 20487 41228 20628 41256
rect 20487 41225 20499 41228
rect 20441 41219 20499 41225
rect 20622 41216 20628 41228
rect 20680 41216 20686 41268
rect 21177 41259 21235 41265
rect 21177 41225 21189 41259
rect 21223 41256 21235 41259
rect 21266 41256 21272 41268
rect 21223 41228 21272 41256
rect 21223 41225 21235 41228
rect 21177 41219 21235 41225
rect 21266 41216 21272 41228
rect 21324 41216 21330 41268
rect 21821 41259 21879 41265
rect 21821 41225 21833 41259
rect 21867 41225 21879 41259
rect 21821 41219 21879 41225
rect 22097 41259 22155 41265
rect 22097 41225 22109 41259
rect 22143 41256 22155 41259
rect 22186 41256 22192 41268
rect 22143 41228 22192 41256
rect 22143 41225 22155 41228
rect 22097 41219 22155 41225
rect 21836 41188 21864 41219
rect 22186 41216 22192 41228
rect 22244 41216 22250 41268
rect 22278 41216 22284 41268
rect 22336 41256 22342 41268
rect 22465 41259 22523 41265
rect 22465 41256 22477 41259
rect 22336 41228 22477 41256
rect 22336 41216 22342 41228
rect 22465 41225 22477 41228
rect 22511 41225 22523 41259
rect 22465 41219 22523 41225
rect 23109 41259 23167 41265
rect 23109 41225 23121 41259
rect 23155 41256 23167 41259
rect 23198 41256 23204 41268
rect 23155 41228 23204 41256
rect 23155 41225 23167 41228
rect 23109 41219 23167 41225
rect 23198 41216 23204 41228
rect 23256 41216 23262 41268
rect 24213 41259 24271 41265
rect 24213 41225 24225 41259
rect 24259 41256 24271 41259
rect 24302 41256 24308 41268
rect 24259 41228 24308 41256
rect 24259 41225 24271 41228
rect 24213 41219 24271 41225
rect 24302 41216 24308 41228
rect 24360 41216 24366 41268
rect 22833 41191 22891 41197
rect 22833 41188 22845 41191
rect 20272 41160 21864 41188
rect 22112 41160 22845 41188
rect 19659 41092 20024 41120
rect 20073 41123 20131 41129
rect 19659 41089 19671 41092
rect 19613 41083 19671 41089
rect 20073 41089 20085 41123
rect 20119 41120 20131 41123
rect 20272 41120 20300 41160
rect 22112 41132 22140 41160
rect 22833 41157 22845 41160
rect 22879 41157 22891 41191
rect 22833 41151 22891 41157
rect 20119 41092 20300 41120
rect 20119 41089 20131 41092
rect 20073 41083 20131 41089
rect 20346 41080 20352 41132
rect 20404 41080 20410 41132
rect 20625 41123 20683 41129
rect 20625 41089 20637 41123
rect 20671 41120 20683 41123
rect 20806 41120 20812 41132
rect 20671 41092 20812 41120
rect 20671 41089 20683 41092
rect 20625 41083 20683 41089
rect 20806 41080 20812 41092
rect 20864 41080 20870 41132
rect 20993 41123 21051 41129
rect 20993 41089 21005 41123
rect 21039 41089 21051 41123
rect 20993 41083 21051 41089
rect 21361 41123 21419 41129
rect 21361 41089 21373 41123
rect 21407 41089 21419 41123
rect 21361 41083 21419 41089
rect 21008 41052 21036 41083
rect 12406 41024 21036 41052
rect 21376 41052 21404 41083
rect 21450 41080 21456 41132
rect 21508 41120 21514 41132
rect 21637 41123 21695 41129
rect 21637 41120 21649 41123
rect 21508 41092 21649 41120
rect 21508 41080 21514 41092
rect 21637 41089 21649 41092
rect 21683 41089 21695 41123
rect 21637 41083 21695 41089
rect 22002 41080 22008 41132
rect 22060 41080 22066 41132
rect 22094 41080 22100 41132
rect 22152 41080 22158 41132
rect 22278 41080 22284 41132
rect 22336 41080 22342 41132
rect 22646 41080 22652 41132
rect 22704 41080 22710 41132
rect 23106 41080 23112 41132
rect 23164 41120 23170 41132
rect 23385 41123 23443 41129
rect 23385 41120 23397 41123
rect 23164 41092 23397 41120
rect 23164 41080 23170 41092
rect 23385 41089 23397 41092
rect 23431 41089 23443 41123
rect 23385 41083 23443 41089
rect 23937 41123 23995 41129
rect 23937 41089 23949 41123
rect 23983 41089 23995 41123
rect 23937 41083 23995 41089
rect 22186 41052 22192 41064
rect 21376 41024 22192 41052
rect 22186 41012 22192 41024
rect 22244 41012 22250 41064
rect 17310 40984 17316 40996
rect 12084 40956 17316 40984
rect 11701 40947 11759 40953
rect 17310 40944 17316 40956
rect 17368 40944 17374 40996
rect 19150 40944 19156 40996
rect 19208 40944 19214 40996
rect 19889 40987 19947 40993
rect 19889 40953 19901 40987
rect 19935 40984 19947 40987
rect 21358 40984 21364 40996
rect 19935 40956 21364 40984
rect 19935 40953 19947 40956
rect 19889 40947 19947 40953
rect 21358 40944 21364 40956
rect 21416 40944 21422 40996
rect 23382 40944 23388 40996
rect 23440 40984 23446 40996
rect 23952 40984 23980 41083
rect 23440 40956 23980 40984
rect 23440 40944 23446 40956
rect 9180 40888 9904 40916
rect 9180 40876 9186 40888
rect 11054 40876 11060 40928
rect 11112 40876 11118 40928
rect 19426 40876 19432 40928
rect 19484 40876 19490 40928
rect 20165 40919 20223 40925
rect 20165 40885 20177 40919
rect 20211 40916 20223 40919
rect 20530 40916 20536 40928
rect 20211 40888 20536 40916
rect 20211 40885 20223 40888
rect 20165 40879 20223 40885
rect 20530 40876 20536 40888
rect 20588 40876 20594 40928
rect 20809 40919 20867 40925
rect 20809 40885 20821 40919
rect 20855 40916 20867 40919
rect 21174 40916 21180 40928
rect 20855 40888 21180 40916
rect 20855 40885 20867 40888
rect 20809 40879 20867 40885
rect 21174 40876 21180 40888
rect 21232 40876 21238 40928
rect 21450 40876 21456 40928
rect 21508 40876 21514 40928
rect 23658 40876 23664 40928
rect 23716 40876 23722 40928
rect 1104 40826 24840 40848
rect 1104 40774 3917 40826
rect 3969 40774 3981 40826
rect 4033 40774 4045 40826
rect 4097 40774 4109 40826
rect 4161 40774 4173 40826
rect 4225 40774 9851 40826
rect 9903 40774 9915 40826
rect 9967 40774 9979 40826
rect 10031 40774 10043 40826
rect 10095 40774 10107 40826
rect 10159 40774 15785 40826
rect 15837 40774 15849 40826
rect 15901 40774 15913 40826
rect 15965 40774 15977 40826
rect 16029 40774 16041 40826
rect 16093 40774 21719 40826
rect 21771 40774 21783 40826
rect 21835 40774 21847 40826
rect 21899 40774 21911 40826
rect 21963 40774 21975 40826
rect 22027 40774 24840 40826
rect 1104 40752 24840 40774
rect 1412 40684 3556 40712
rect 1412 40585 1440 40684
rect 3528 40644 3556 40684
rect 3602 40672 3608 40724
rect 3660 40712 3666 40724
rect 3789 40715 3847 40721
rect 3789 40712 3801 40715
rect 3660 40684 3801 40712
rect 3660 40672 3666 40684
rect 3789 40681 3801 40684
rect 3835 40681 3847 40715
rect 3789 40675 3847 40681
rect 4065 40715 4123 40721
rect 4065 40681 4077 40715
rect 4111 40712 4123 40715
rect 4246 40712 4252 40724
rect 4111 40684 4252 40712
rect 4111 40681 4123 40684
rect 4065 40675 4123 40681
rect 4246 40672 4252 40684
rect 4304 40672 4310 40724
rect 5994 40712 6000 40724
rect 4448 40684 6000 40712
rect 4448 40644 4476 40684
rect 5994 40672 6000 40684
rect 6052 40672 6058 40724
rect 7926 40712 7932 40724
rect 7484 40684 7932 40712
rect 3528 40616 4476 40644
rect 1397 40579 1455 40585
rect 1397 40545 1409 40579
rect 1443 40545 1455 40579
rect 1397 40539 1455 40545
rect 3234 40536 3240 40588
rect 3292 40576 3298 40588
rect 3292 40548 4200 40576
rect 3292 40536 3298 40548
rect 1670 40468 1676 40520
rect 1728 40468 1734 40520
rect 2317 40511 2375 40517
rect 2317 40477 2329 40511
rect 2363 40477 2375 40511
rect 2590 40508 2596 40520
rect 2551 40480 2596 40508
rect 2317 40471 2375 40477
rect 2332 40440 2360 40471
rect 2590 40468 2596 40480
rect 2648 40468 2654 40520
rect 3252 40440 3280 40536
rect 3970 40468 3976 40520
rect 4028 40468 4034 40520
rect 4172 40452 4200 40548
rect 7484 40520 7512 40684
rect 7926 40672 7932 40684
rect 7984 40672 7990 40724
rect 8570 40672 8576 40724
rect 8628 40712 8634 40724
rect 10318 40712 10324 40724
rect 8628 40684 10324 40712
rect 8628 40672 8634 40684
rect 10318 40672 10324 40684
rect 10376 40672 10382 40724
rect 10778 40712 10784 40724
rect 10520 40684 10784 40712
rect 9766 40644 9772 40656
rect 9692 40616 9772 40644
rect 4246 40468 4252 40520
rect 4304 40468 4310 40520
rect 4341 40511 4399 40517
rect 4341 40477 4353 40511
rect 4387 40477 4399 40511
rect 4341 40471 4399 40477
rect 4615 40511 4673 40517
rect 4615 40477 4627 40511
rect 4661 40508 4673 40511
rect 5258 40508 5264 40520
rect 4661 40480 5264 40508
rect 4661 40477 4673 40480
rect 4615 40471 4673 40477
rect 2332 40412 3280 40440
rect 4154 40400 4160 40452
rect 4212 40400 4218 40452
rect 4356 40440 4384 40471
rect 5258 40468 5264 40480
rect 5316 40468 5322 40520
rect 5721 40511 5779 40517
rect 5721 40477 5733 40511
rect 5767 40477 5779 40511
rect 5721 40471 5779 40477
rect 5995 40511 6053 40517
rect 5995 40477 6007 40511
rect 6041 40508 6053 40511
rect 6822 40508 6828 40520
rect 6041 40480 6828 40508
rect 6041 40477 6053 40480
rect 5995 40471 6053 40477
rect 4798 40440 4804 40452
rect 4356 40412 4804 40440
rect 4798 40400 4804 40412
rect 4856 40440 4862 40452
rect 5736 40440 5764 40471
rect 6822 40468 6828 40480
rect 6880 40468 6886 40520
rect 6914 40468 6920 40520
rect 6972 40508 6978 40520
rect 7466 40508 7472 40520
rect 6972 40480 7472 40508
rect 6972 40468 6978 40480
rect 7466 40468 7472 40480
rect 7524 40468 7530 40520
rect 7743 40511 7801 40517
rect 7743 40477 7755 40511
rect 7789 40508 7801 40511
rect 8294 40508 8300 40520
rect 7789 40480 8300 40508
rect 7789 40477 7801 40480
rect 7743 40471 7801 40477
rect 8294 40468 8300 40480
rect 8352 40468 8358 40520
rect 9692 40440 9720 40616
rect 9766 40604 9772 40616
rect 9824 40604 9830 40656
rect 10520 40653 10548 40684
rect 10778 40672 10784 40684
rect 10836 40672 10842 40724
rect 20162 40672 20168 40724
rect 20220 40712 20226 40724
rect 20441 40715 20499 40721
rect 20441 40712 20453 40715
rect 20220 40684 20453 40712
rect 20220 40672 20226 40684
rect 20441 40681 20453 40684
rect 20487 40681 20499 40715
rect 20441 40675 20499 40681
rect 20717 40715 20775 40721
rect 20717 40681 20729 40715
rect 20763 40712 20775 40715
rect 21082 40712 21088 40724
rect 20763 40684 21088 40712
rect 20763 40681 20775 40684
rect 20717 40675 20775 40681
rect 21082 40672 21088 40684
rect 21140 40672 21146 40724
rect 22097 40715 22155 40721
rect 22097 40681 22109 40715
rect 22143 40712 22155 40715
rect 22370 40712 22376 40724
rect 22143 40684 22376 40712
rect 22143 40681 22155 40684
rect 22097 40675 22155 40681
rect 22370 40672 22376 40684
rect 22428 40672 22434 40724
rect 22554 40672 22560 40724
rect 22612 40672 22618 40724
rect 22925 40715 22983 40721
rect 22925 40681 22937 40715
rect 22971 40712 22983 40715
rect 23290 40712 23296 40724
rect 22971 40684 23296 40712
rect 22971 40681 22983 40684
rect 22925 40675 22983 40681
rect 23290 40672 23296 40684
rect 23348 40672 23354 40724
rect 23569 40715 23627 40721
rect 23569 40681 23581 40715
rect 23615 40712 23627 40715
rect 25314 40712 25320 40724
rect 23615 40684 25320 40712
rect 23615 40681 23627 40684
rect 23569 40675 23627 40681
rect 25314 40672 25320 40684
rect 25372 40672 25378 40724
rect 10505 40647 10563 40653
rect 10505 40613 10517 40647
rect 10551 40613 10563 40647
rect 10505 40607 10563 40613
rect 19613 40647 19671 40653
rect 19613 40613 19625 40647
rect 19659 40644 19671 40647
rect 20898 40644 20904 40656
rect 19659 40616 20904 40644
rect 19659 40613 19671 40616
rect 19613 40607 19671 40613
rect 20898 40604 20904 40616
rect 20956 40604 20962 40656
rect 20990 40604 20996 40656
rect 21048 40604 21054 40656
rect 21266 40604 21272 40656
rect 21324 40604 21330 40656
rect 21545 40647 21603 40653
rect 21545 40613 21557 40647
rect 21591 40644 21603 40647
rect 21591 40616 21680 40644
rect 21591 40613 21603 40616
rect 21545 40607 21603 40613
rect 10045 40579 10103 40585
rect 10045 40576 10057 40579
rect 9784 40548 10057 40576
rect 9784 40520 9812 40548
rect 10045 40545 10057 40548
rect 10091 40545 10103 40579
rect 10045 40539 10103 40545
rect 10778 40536 10784 40588
rect 10836 40536 10842 40588
rect 11054 40536 11060 40588
rect 11112 40536 11118 40588
rect 16574 40536 16580 40588
rect 16632 40576 16638 40588
rect 16632 40548 19932 40576
rect 16632 40536 16638 40548
rect 9766 40468 9772 40520
rect 9824 40468 9830 40520
rect 9861 40511 9919 40517
rect 9861 40477 9873 40511
rect 9907 40477 9919 40511
rect 9861 40471 9919 40477
rect 4856 40412 9720 40440
rect 4856 40400 4862 40412
rect 6472 40384 6500 40412
rect 3234 40332 3240 40384
rect 3292 40372 3298 40384
rect 3329 40375 3387 40381
rect 3329 40372 3341 40375
rect 3292 40344 3341 40372
rect 3292 40332 3298 40344
rect 3329 40341 3341 40344
rect 3375 40341 3387 40375
rect 3329 40335 3387 40341
rect 5350 40332 5356 40384
rect 5408 40332 5414 40384
rect 6454 40332 6460 40384
rect 6512 40332 6518 40384
rect 6730 40332 6736 40384
rect 6788 40332 6794 40384
rect 8478 40332 8484 40384
rect 8536 40332 8542 40384
rect 9876 40372 9904 40471
rect 10870 40468 10876 40520
rect 10928 40517 10934 40520
rect 10928 40511 10956 40517
rect 10944 40477 10956 40511
rect 10928 40471 10956 40477
rect 19337 40511 19395 40517
rect 19337 40477 19349 40511
rect 19383 40508 19395 40511
rect 19426 40508 19432 40520
rect 19383 40480 19432 40508
rect 19383 40477 19395 40480
rect 19337 40471 19395 40477
rect 10928 40468 10934 40471
rect 19426 40468 19432 40480
rect 19484 40468 19490 40520
rect 19797 40511 19855 40517
rect 19797 40477 19809 40511
rect 19843 40477 19855 40511
rect 19797 40471 19855 40477
rect 19812 40440 19840 40471
rect 11532 40412 19840 40440
rect 19904 40440 19932 40548
rect 20530 40536 20536 40588
rect 20588 40536 20594 40588
rect 21652 40576 21680 40616
rect 22002 40604 22008 40656
rect 22060 40644 22066 40656
rect 23934 40644 23940 40656
rect 22060 40616 23940 40644
rect 22060 40604 22066 40616
rect 23934 40604 23940 40616
rect 23992 40604 23998 40656
rect 24118 40604 24124 40656
rect 24176 40604 24182 40656
rect 24136 40576 24164 40604
rect 21100 40548 21588 40576
rect 21652 40548 24164 40576
rect 20070 40468 20076 40520
rect 20128 40468 20134 40520
rect 20349 40511 20407 40517
rect 20349 40477 20361 40511
rect 20395 40508 20407 40511
rect 20548 40508 20576 40536
rect 20395 40480 20576 40508
rect 20625 40511 20683 40517
rect 20395 40477 20407 40480
rect 20349 40471 20407 40477
rect 20625 40477 20637 40511
rect 20671 40508 20683 40511
rect 20806 40508 20812 40520
rect 20671 40480 20812 40508
rect 20671 40477 20683 40480
rect 20625 40471 20683 40477
rect 20806 40468 20812 40480
rect 20864 40468 20870 40520
rect 20898 40468 20904 40520
rect 20956 40468 20962 40520
rect 20714 40440 20720 40452
rect 19904 40412 20720 40440
rect 11146 40372 11152 40384
rect 9876 40344 11152 40372
rect 11146 40332 11152 40344
rect 11204 40332 11210 40384
rect 11330 40332 11336 40384
rect 11388 40372 11394 40384
rect 11532 40372 11560 40412
rect 20714 40400 20720 40412
rect 20772 40400 20778 40452
rect 11388 40344 11560 40372
rect 11701 40375 11759 40381
rect 11388 40332 11394 40344
rect 11701 40341 11713 40375
rect 11747 40372 11759 40375
rect 12434 40372 12440 40384
rect 11747 40344 12440 40372
rect 11747 40341 11759 40344
rect 11701 40335 11759 40341
rect 12434 40332 12440 40344
rect 12492 40332 12498 40384
rect 19426 40332 19432 40384
rect 19484 40332 19490 40384
rect 19886 40332 19892 40384
rect 19944 40332 19950 40384
rect 20165 40375 20223 40381
rect 20165 40341 20177 40375
rect 20211 40372 20223 40375
rect 21100 40372 21128 40548
rect 21177 40511 21235 40517
rect 21177 40477 21189 40511
rect 21223 40508 21235 40511
rect 21358 40508 21364 40520
rect 21223 40480 21364 40508
rect 21223 40477 21235 40480
rect 21177 40471 21235 40477
rect 21358 40468 21364 40480
rect 21416 40468 21422 40520
rect 21450 40468 21456 40520
rect 21508 40468 21514 40520
rect 21560 40484 21588 40548
rect 21560 40456 21680 40484
rect 21726 40468 21732 40520
rect 21784 40468 21790 40520
rect 22005 40511 22063 40517
rect 22005 40508 22017 40511
rect 21836 40480 22017 40508
rect 21652 40440 21680 40456
rect 21836 40440 21864 40480
rect 22005 40477 22017 40480
rect 22051 40477 22063 40511
rect 22005 40471 22063 40477
rect 22278 40468 22284 40520
rect 22336 40468 22342 40520
rect 22741 40511 22799 40517
rect 22741 40477 22753 40511
rect 22787 40477 22799 40511
rect 22741 40471 22799 40477
rect 21652 40412 21864 40440
rect 21910 40400 21916 40452
rect 21968 40400 21974 40452
rect 22756 40440 22784 40471
rect 22922 40468 22928 40520
rect 22980 40508 22986 40520
rect 23109 40511 23167 40517
rect 23109 40508 23121 40511
rect 22980 40480 23121 40508
rect 22980 40468 22986 40480
rect 23109 40477 23121 40480
rect 23155 40477 23167 40511
rect 23109 40471 23167 40477
rect 23014 40440 23020 40452
rect 22756 40412 23020 40440
rect 23014 40400 23020 40412
rect 23072 40400 23078 40452
rect 23198 40400 23204 40452
rect 23256 40440 23262 40452
rect 23293 40443 23351 40449
rect 23293 40440 23305 40443
rect 23256 40412 23305 40440
rect 23256 40400 23262 40412
rect 23293 40409 23305 40412
rect 23339 40409 23351 40443
rect 23293 40403 23351 40409
rect 23842 40400 23848 40452
rect 23900 40400 23906 40452
rect 24210 40400 24216 40452
rect 24268 40400 24274 40452
rect 20211 40344 21128 40372
rect 21821 40375 21879 40381
rect 20211 40341 20223 40344
rect 20165 40335 20223 40341
rect 21821 40341 21833 40375
rect 21867 40372 21879 40375
rect 21928 40372 21956 40400
rect 21867 40344 21956 40372
rect 21867 40341 21879 40344
rect 21821 40335 21879 40341
rect 1104 40282 25000 40304
rect 1104 40230 6884 40282
rect 6936 40230 6948 40282
rect 7000 40230 7012 40282
rect 7064 40230 7076 40282
rect 7128 40230 7140 40282
rect 7192 40230 12818 40282
rect 12870 40230 12882 40282
rect 12934 40230 12946 40282
rect 12998 40230 13010 40282
rect 13062 40230 13074 40282
rect 13126 40230 18752 40282
rect 18804 40230 18816 40282
rect 18868 40230 18880 40282
rect 18932 40230 18944 40282
rect 18996 40230 19008 40282
rect 19060 40230 24686 40282
rect 24738 40230 24750 40282
rect 24802 40230 24814 40282
rect 24866 40230 24878 40282
rect 24930 40230 24942 40282
rect 24994 40230 25000 40282
rect 1104 40208 25000 40230
rect 2777 40171 2835 40177
rect 2777 40137 2789 40171
rect 2823 40168 2835 40171
rect 2866 40168 2872 40180
rect 2823 40140 2872 40168
rect 2823 40137 2835 40140
rect 2777 40131 2835 40137
rect 2866 40128 2872 40140
rect 2924 40128 2930 40180
rect 2958 40128 2964 40180
rect 3016 40168 3022 40180
rect 3142 40168 3148 40180
rect 3016 40140 3148 40168
rect 3016 40128 3022 40140
rect 3142 40128 3148 40140
rect 3200 40128 3206 40180
rect 3786 40128 3792 40180
rect 3844 40128 3850 40180
rect 3878 40128 3884 40180
rect 3936 40128 3942 40180
rect 4154 40128 4160 40180
rect 4212 40168 4218 40180
rect 4341 40171 4399 40177
rect 4341 40168 4353 40171
rect 4212 40140 4353 40168
rect 4212 40128 4218 40140
rect 4341 40137 4353 40140
rect 4387 40137 4399 40171
rect 4341 40131 4399 40137
rect 5258 40128 5264 40180
rect 5316 40168 5322 40180
rect 8386 40168 8392 40180
rect 5316 40140 8392 40168
rect 5316 40128 5322 40140
rect 8386 40128 8392 40140
rect 8444 40128 8450 40180
rect 10870 40168 10876 40180
rect 8680 40140 10876 40168
rect 3237 40103 3295 40109
rect 3237 40069 3249 40103
rect 3283 40100 3295 40103
rect 3418 40100 3424 40112
rect 3283 40072 3424 40100
rect 3283 40069 3295 40072
rect 3237 40063 3295 40069
rect 3418 40060 3424 40072
rect 3476 40060 3482 40112
rect 3605 40103 3663 40109
rect 3605 40069 3617 40103
rect 3651 40100 3663 40103
rect 3804 40100 3832 40128
rect 3651 40072 3832 40100
rect 3896 40100 3924 40128
rect 3896 40072 4106 40100
rect 3651 40069 3663 40072
rect 3605 40063 3663 40069
rect 1671 40035 1729 40041
rect 1671 40001 1683 40035
rect 1717 40032 1729 40035
rect 2498 40032 2504 40044
rect 1717 40004 2504 40032
rect 1717 40001 1729 40004
rect 1671 39995 1729 40001
rect 2498 39992 2504 40004
rect 2556 39992 2562 40044
rect 2958 39992 2964 40044
rect 3016 39992 3022 40044
rect 3326 39992 3332 40044
rect 3384 40032 3390 40044
rect 3513 40035 3571 40041
rect 3513 40032 3525 40035
rect 3384 40004 3525 40032
rect 3384 39992 3390 40004
rect 3513 40001 3525 40004
rect 3559 40001 3571 40035
rect 3513 39995 3571 40001
rect 3786 39992 3792 40044
rect 3844 40032 3850 40044
rect 3973 40035 4031 40041
rect 3973 40032 3985 40035
rect 3844 40004 3985 40032
rect 3844 39992 3850 40004
rect 3973 40001 3985 40004
rect 4019 40001 4031 40035
rect 4078 40032 4106 40072
rect 4522 40060 4528 40112
rect 4580 40100 4586 40112
rect 4982 40100 4988 40112
rect 4580 40072 4988 40100
rect 4580 40060 4586 40072
rect 4982 40060 4988 40072
rect 5040 40060 5046 40112
rect 6656 40072 8248 40100
rect 5135 40035 5193 40041
rect 5135 40032 5147 40035
rect 4078 40004 5147 40032
rect 3973 39995 4031 40001
rect 5135 40001 5147 40004
rect 5181 40032 5193 40035
rect 6656 40032 6684 40072
rect 6822 40032 6828 40044
rect 5181 40004 6684 40032
rect 6783 40004 6828 40032
rect 5181 40001 5193 40004
rect 5135 39995 5193 40001
rect 6822 39992 6828 40004
rect 6880 39992 6886 40044
rect 8220 40032 8248 40072
rect 8294 40060 8300 40112
rect 8352 40100 8358 40112
rect 8680 40109 8708 40140
rect 10870 40128 10876 40140
rect 10928 40128 10934 40180
rect 19981 40171 20039 40177
rect 19981 40137 19993 40171
rect 20027 40137 20039 40171
rect 19981 40131 20039 40137
rect 8665 40103 8723 40109
rect 8665 40100 8677 40103
rect 8352 40072 8677 40100
rect 8352 40060 8358 40072
rect 8665 40069 8677 40072
rect 8711 40069 8723 40103
rect 8665 40063 8723 40069
rect 9030 40060 9036 40112
rect 9088 40060 9094 40112
rect 9306 40060 9312 40112
rect 9364 40100 9370 40112
rect 11330 40100 11336 40112
rect 9364 40072 11336 40100
rect 9364 40060 9370 40072
rect 11330 40060 11336 40072
rect 11388 40060 11394 40112
rect 15194 40060 15200 40112
rect 15252 40100 15258 40112
rect 16850 40100 16856 40112
rect 15252 40072 16856 40100
rect 15252 40060 15258 40072
rect 16850 40060 16856 40072
rect 16908 40060 16914 40112
rect 19996 40100 20024 40131
rect 20254 40128 20260 40180
rect 20312 40128 20318 40180
rect 20533 40171 20591 40177
rect 20533 40137 20545 40171
rect 20579 40168 20591 40171
rect 20898 40168 20904 40180
rect 20579 40140 20904 40168
rect 20579 40137 20591 40140
rect 20533 40131 20591 40137
rect 20898 40128 20904 40140
rect 20956 40128 20962 40180
rect 21453 40171 21511 40177
rect 21453 40137 21465 40171
rect 21499 40168 21511 40171
rect 22002 40168 22008 40180
rect 21499 40140 22008 40168
rect 21499 40137 21511 40140
rect 21453 40131 21511 40137
rect 22002 40128 22008 40140
rect 22060 40128 22066 40180
rect 22097 40171 22155 40177
rect 22097 40137 22109 40171
rect 22143 40137 22155 40171
rect 22097 40131 22155 40137
rect 20622 40100 20628 40112
rect 19996 40072 20628 40100
rect 20622 40060 20628 40072
rect 20680 40060 20686 40112
rect 20806 40060 20812 40112
rect 20864 40060 20870 40112
rect 21726 40060 21732 40112
rect 21784 40100 21790 40112
rect 22112 40100 22140 40131
rect 22186 40128 22192 40180
rect 22244 40168 22250 40180
rect 22373 40171 22431 40177
rect 22373 40168 22385 40171
rect 22244 40140 22385 40168
rect 22244 40128 22250 40140
rect 22373 40137 22385 40140
rect 22419 40137 22431 40171
rect 22373 40131 22431 40137
rect 22833 40171 22891 40177
rect 22833 40137 22845 40171
rect 22879 40168 22891 40171
rect 23106 40168 23112 40180
rect 22879 40140 23112 40168
rect 22879 40137 22891 40140
rect 22833 40131 22891 40137
rect 23106 40128 23112 40140
rect 23164 40128 23170 40180
rect 23385 40171 23443 40177
rect 23385 40137 23397 40171
rect 23431 40168 23443 40171
rect 23658 40168 23664 40180
rect 23431 40140 23664 40168
rect 23431 40137 23443 40140
rect 23385 40131 23443 40137
rect 23658 40128 23664 40140
rect 23716 40128 23722 40180
rect 23750 40128 23756 40180
rect 23808 40128 23814 40180
rect 21784 40072 22048 40100
rect 22112 40072 23060 40100
rect 21784 40060 21790 40072
rect 8570 40042 8576 40044
rect 8404 40032 8576 40042
rect 8220 40014 8576 40032
rect 8220 40004 8432 40014
rect 8570 39992 8576 40014
rect 8628 39992 8634 40044
rect 8754 39992 8760 40044
rect 8812 40032 8818 40044
rect 8938 40032 8944 40044
rect 8812 40004 8944 40032
rect 8812 39992 8818 40004
rect 8938 39992 8944 40004
rect 8996 39992 9002 40044
rect 9214 39992 9220 40044
rect 9272 40032 9278 40044
rect 9401 40035 9459 40041
rect 9401 40032 9413 40035
rect 9272 40004 9413 40032
rect 9272 39992 9278 40004
rect 9401 40001 9413 40004
rect 9447 40001 9459 40035
rect 9401 39995 9459 40001
rect 9766 39992 9772 40044
rect 9824 40041 9830 40044
rect 9824 40035 9841 40041
rect 9829 40001 9841 40035
rect 9824 39995 9841 40001
rect 9824 39992 9830 39995
rect 20162 39992 20168 40044
rect 20220 39992 20226 40044
rect 20438 39992 20444 40044
rect 20496 39992 20502 40044
rect 20714 39992 20720 40044
rect 20772 39992 20778 40044
rect 3240 39976 3292 39982
rect 8484 39976 8536 39982
rect 1397 39967 1455 39973
rect 1397 39933 1409 39967
rect 1443 39933 1455 39967
rect 1397 39927 1455 39933
rect 1412 39828 1440 39927
rect 4798 39924 4804 39976
rect 4856 39964 4862 39976
rect 4893 39967 4951 39973
rect 4893 39964 4905 39967
rect 4856 39936 4905 39964
rect 4856 39924 4862 39936
rect 4893 39933 4905 39936
rect 4939 39933 4951 39967
rect 4893 39927 4951 39933
rect 6454 39924 6460 39976
rect 6512 39964 6518 39976
rect 6549 39967 6607 39973
rect 6549 39964 6561 39967
rect 6512 39936 6561 39964
rect 6512 39924 6518 39936
rect 6549 39933 6561 39936
rect 6595 39933 6607 39967
rect 6549 39927 6607 39933
rect 20824 39964 20852 40060
rect 21376 40044 21588 40056
rect 21082 39992 21088 40044
rect 21140 39992 21146 40044
rect 21376 40041 21548 40044
rect 21361 40035 21548 40041
rect 21361 40001 21373 40035
rect 21407 40028 21548 40035
rect 21407 40001 21419 40028
rect 21361 39995 21419 40001
rect 21542 39992 21548 40028
rect 21600 39992 21606 40044
rect 22020 40041 22048 40072
rect 21637 40035 21695 40041
rect 21637 40001 21649 40035
rect 21683 40032 21695 40035
rect 22005 40035 22063 40041
rect 21683 40004 21956 40032
rect 21683 40001 21695 40004
rect 21637 39995 21695 40001
rect 21928 39964 21956 40004
rect 22005 40001 22017 40035
rect 22051 40001 22063 40035
rect 22005 39995 22063 40001
rect 22094 39992 22100 40044
rect 22152 40032 22158 40044
rect 22281 40035 22339 40041
rect 22281 40032 22293 40035
rect 22152 40004 22293 40032
rect 22152 39992 22158 40004
rect 22281 40001 22293 40004
rect 22327 40001 22339 40035
rect 22281 39995 22339 40001
rect 22554 39992 22560 40044
rect 22612 39992 22618 40044
rect 23032 40041 23060 40072
rect 23474 40060 23480 40112
rect 23532 40100 23538 40112
rect 23532 40072 23612 40100
rect 23532 40060 23538 40072
rect 23017 40035 23075 40041
rect 23017 40001 23029 40035
rect 23063 40001 23075 40035
rect 23017 39995 23075 40001
rect 23290 39992 23296 40044
rect 23348 39992 23354 40044
rect 23584 40041 23612 40072
rect 23569 40035 23627 40041
rect 23569 40001 23581 40035
rect 23615 40001 23627 40035
rect 23569 39995 23627 40001
rect 23658 39992 23664 40044
rect 23716 40032 23722 40044
rect 23937 40035 23995 40041
rect 23937 40032 23949 40035
rect 23716 40004 23949 40032
rect 23716 39992 23722 40004
rect 23937 40001 23949 40004
rect 23983 40001 23995 40035
rect 23937 39995 23995 40001
rect 24026 39992 24032 40044
rect 24084 40032 24090 40044
rect 24121 40035 24179 40041
rect 24121 40032 24133 40035
rect 24084 40004 24133 40032
rect 24084 39992 24090 40004
rect 24121 40001 24133 40004
rect 24167 40001 24179 40035
rect 24121 39995 24179 40001
rect 22462 39964 22468 39976
rect 20824 39936 21680 39964
rect 21928 39936 22468 39964
rect 3240 39918 3292 39924
rect 8484 39918 8536 39924
rect 20898 39856 20904 39908
rect 20956 39856 20962 39908
rect 21177 39899 21235 39905
rect 21177 39865 21189 39899
rect 21223 39896 21235 39899
rect 21266 39896 21272 39908
rect 21223 39868 21272 39896
rect 21223 39865 21235 39868
rect 21177 39859 21235 39865
rect 21266 39856 21272 39868
rect 21324 39856 21330 39908
rect 1854 39828 1860 39840
rect 1412 39800 1860 39828
rect 1854 39788 1860 39800
rect 1912 39788 1918 39840
rect 2409 39831 2467 39837
rect 2409 39797 2421 39831
rect 2455 39828 2467 39831
rect 2590 39828 2596 39840
rect 2455 39800 2596 39828
rect 2455 39797 2467 39800
rect 2409 39791 2467 39797
rect 2590 39788 2596 39800
rect 2648 39788 2654 39840
rect 4525 39831 4583 39837
rect 4525 39797 4537 39831
rect 4571 39828 4583 39831
rect 5166 39828 5172 39840
rect 4571 39800 5172 39828
rect 4571 39797 4583 39800
rect 4525 39791 4583 39797
rect 5166 39788 5172 39800
rect 5224 39788 5230 39840
rect 5902 39788 5908 39840
rect 5960 39788 5966 39840
rect 7466 39788 7472 39840
rect 7524 39828 7530 39840
rect 7561 39831 7619 39837
rect 7561 39828 7573 39831
rect 7524 39800 7573 39828
rect 7524 39788 7530 39800
rect 7561 39797 7573 39800
rect 7607 39797 7619 39831
rect 7561 39791 7619 39797
rect 9953 39831 10011 39837
rect 9953 39797 9965 39831
rect 9999 39828 10011 39831
rect 10226 39828 10232 39840
rect 9999 39800 10232 39828
rect 9999 39797 10011 39800
rect 9953 39791 10011 39797
rect 10226 39788 10232 39800
rect 10284 39828 10290 39840
rect 10410 39828 10416 39840
rect 10284 39800 10416 39828
rect 10284 39788 10290 39800
rect 10410 39788 10416 39800
rect 10468 39788 10474 39840
rect 12526 39788 12532 39840
rect 12584 39828 12590 39840
rect 16942 39828 16948 39840
rect 12584 39800 16948 39828
rect 12584 39788 12590 39800
rect 16942 39788 16948 39800
rect 17000 39828 17006 39840
rect 21358 39828 21364 39840
rect 17000 39800 21364 39828
rect 17000 39788 17006 39800
rect 21358 39788 21364 39800
rect 21416 39788 21422 39840
rect 21652 39828 21680 39936
rect 22462 39924 22468 39936
rect 22520 39924 22526 39976
rect 23109 39899 23167 39905
rect 23109 39865 23121 39899
rect 23155 39896 23167 39899
rect 23382 39896 23388 39908
rect 23155 39868 23388 39896
rect 23155 39865 23167 39868
rect 23109 39859 23167 39865
rect 23382 39856 23388 39868
rect 23440 39856 23446 39908
rect 21821 39831 21879 39837
rect 21821 39828 21833 39831
rect 21652 39800 21833 39828
rect 21821 39797 21833 39800
rect 21867 39797 21879 39831
rect 21821 39791 21879 39797
rect 24394 39788 24400 39840
rect 24452 39788 24458 39840
rect 1104 39738 24840 39760
rect 1104 39686 3917 39738
rect 3969 39686 3981 39738
rect 4033 39686 4045 39738
rect 4097 39686 4109 39738
rect 4161 39686 4173 39738
rect 4225 39686 9851 39738
rect 9903 39686 9915 39738
rect 9967 39686 9979 39738
rect 10031 39686 10043 39738
rect 10095 39686 10107 39738
rect 10159 39686 15785 39738
rect 15837 39686 15849 39738
rect 15901 39686 15913 39738
rect 15965 39686 15977 39738
rect 16029 39686 16041 39738
rect 16093 39686 21719 39738
rect 21771 39686 21783 39738
rect 21835 39686 21847 39738
rect 21899 39686 21911 39738
rect 21963 39686 21975 39738
rect 22027 39686 24840 39738
rect 1104 39664 24840 39686
rect 566 39584 572 39636
rect 624 39624 630 39636
rect 3789 39627 3847 39633
rect 624 39596 2728 39624
rect 624 39584 630 39596
rect 1854 39516 1860 39568
rect 1912 39556 1918 39568
rect 1912 39528 2084 39556
rect 1912 39516 1918 39528
rect 2056 39497 2084 39528
rect 2041 39491 2099 39497
rect 2041 39457 2053 39491
rect 2087 39457 2099 39491
rect 2700 39488 2728 39596
rect 3789 39593 3801 39627
rect 3835 39624 3847 39627
rect 4338 39624 4344 39636
rect 3835 39596 4344 39624
rect 3835 39593 3847 39596
rect 3789 39587 3847 39593
rect 4338 39584 4344 39596
rect 4396 39584 4402 39636
rect 5350 39624 5356 39636
rect 4816 39596 5356 39624
rect 3050 39516 3056 39568
rect 3108 39556 3114 39568
rect 3421 39559 3479 39565
rect 3421 39556 3433 39559
rect 3108 39528 3433 39556
rect 3108 39516 3114 39528
rect 3421 39525 3433 39528
rect 3467 39525 3479 39559
rect 3421 39519 3479 39525
rect 4430 39516 4436 39568
rect 4488 39556 4494 39568
rect 4816 39565 4844 39596
rect 5350 39584 5356 39596
rect 5408 39584 5414 39636
rect 5902 39584 5908 39636
rect 5960 39584 5966 39636
rect 5994 39584 6000 39636
rect 6052 39624 6058 39636
rect 7929 39627 7987 39633
rect 7929 39624 7941 39627
rect 6052 39596 7941 39624
rect 6052 39584 6058 39596
rect 7929 39593 7941 39596
rect 7975 39593 7987 39627
rect 7929 39587 7987 39593
rect 8386 39584 8392 39636
rect 8444 39624 8450 39636
rect 12158 39624 12164 39636
rect 8444 39596 12164 39624
rect 8444 39584 8450 39596
rect 12158 39584 12164 39596
rect 12216 39584 12222 39636
rect 12526 39624 12532 39636
rect 12268 39596 12532 39624
rect 4801 39559 4859 39565
rect 4488 39528 4752 39556
rect 4488 39516 4494 39528
rect 4157 39491 4215 39497
rect 2700 39460 4016 39488
rect 2041 39451 2099 39457
rect 1397 39423 1455 39429
rect 1397 39389 1409 39423
rect 1443 39420 1455 39423
rect 1578 39420 1584 39432
rect 1443 39392 1584 39420
rect 1443 39389 1455 39392
rect 1397 39383 1455 39389
rect 1578 39380 1584 39392
rect 1636 39380 1642 39432
rect 1946 39380 1952 39432
rect 2004 39420 2010 39432
rect 3988 39429 4016 39460
rect 4157 39457 4169 39491
rect 4203 39488 4215 39491
rect 4522 39488 4528 39500
rect 4203 39460 4528 39488
rect 4203 39457 4215 39460
rect 4157 39451 4215 39457
rect 4522 39448 4528 39460
rect 4580 39448 4586 39500
rect 4724 39488 4752 39528
rect 4801 39525 4813 39559
rect 4847 39525 4859 39559
rect 4801 39519 4859 39525
rect 5077 39491 5135 39497
rect 5077 39488 5089 39491
rect 4724 39460 5089 39488
rect 5077 39457 5089 39460
rect 5123 39457 5135 39491
rect 5077 39451 5135 39457
rect 5353 39491 5411 39497
rect 5353 39457 5365 39491
rect 5399 39488 5411 39491
rect 5920 39488 5948 39584
rect 6730 39516 6736 39568
rect 6788 39516 6794 39568
rect 9122 39516 9128 39568
rect 9180 39556 9186 39568
rect 9180 39528 9260 39556
rect 9180 39516 9186 39528
rect 5399 39460 5948 39488
rect 6089 39491 6147 39497
rect 5399 39457 5411 39460
rect 5353 39451 5411 39457
rect 6089 39457 6101 39491
rect 6135 39488 6147 39491
rect 6638 39488 6644 39500
rect 6135 39460 6644 39488
rect 6135 39457 6147 39460
rect 6089 39451 6147 39457
rect 6638 39448 6644 39460
rect 6696 39448 6702 39500
rect 7285 39491 7343 39497
rect 7285 39457 7297 39491
rect 7331 39488 7343 39491
rect 7466 39488 7472 39500
rect 7331 39460 7472 39488
rect 7331 39457 7343 39460
rect 7285 39451 7343 39457
rect 7466 39448 7472 39460
rect 7524 39448 7530 39500
rect 8202 39448 8208 39500
rect 8260 39488 8266 39500
rect 9232 39497 9260 39528
rect 12268 39497 12296 39596
rect 12526 39584 12532 39596
rect 12584 39584 12590 39636
rect 21085 39627 21143 39633
rect 21085 39593 21097 39627
rect 21131 39624 21143 39627
rect 21450 39624 21456 39636
rect 21131 39596 21456 39624
rect 21131 39593 21143 39596
rect 21085 39587 21143 39593
rect 21450 39584 21456 39596
rect 21508 39584 21514 39636
rect 21634 39584 21640 39636
rect 21692 39584 21698 39636
rect 21913 39627 21971 39633
rect 21913 39593 21925 39627
rect 21959 39624 21971 39627
rect 21959 39596 22048 39624
rect 21959 39593 21971 39596
rect 21913 39587 21971 39593
rect 20806 39516 20812 39568
rect 20864 39516 20870 39568
rect 21361 39559 21419 39565
rect 21361 39525 21373 39559
rect 21407 39525 21419 39559
rect 21361 39519 21419 39525
rect 9217 39491 9275 39497
rect 9217 39488 9229 39491
rect 8260 39460 9229 39488
rect 8260 39448 8266 39460
rect 9217 39457 9229 39460
rect 9263 39457 9275 39491
rect 9217 39451 9275 39457
rect 12253 39491 12311 39497
rect 12253 39457 12265 39491
rect 12299 39457 12311 39491
rect 21376 39488 21404 39519
rect 21910 39488 21916 39500
rect 21376 39460 21916 39488
rect 12253 39451 12311 39457
rect 21910 39448 21916 39460
rect 21968 39448 21974 39500
rect 2283 39423 2341 39429
rect 2283 39420 2295 39423
rect 2004 39392 2295 39420
rect 2004 39380 2010 39392
rect 2283 39389 2295 39392
rect 2329 39389 2341 39423
rect 3605 39423 3663 39429
rect 3605 39420 3617 39423
rect 2283 39383 2341 39389
rect 2746 39392 3617 39420
rect 1673 39355 1731 39361
rect 1673 39321 1685 39355
rect 1719 39352 1731 39355
rect 2038 39352 2044 39364
rect 1719 39324 2044 39352
rect 1719 39321 1731 39324
rect 1673 39315 1731 39321
rect 2038 39312 2044 39324
rect 2096 39312 2102 39364
rect 934 39244 940 39296
rect 992 39284 998 39296
rect 2746 39284 2774 39392
rect 3605 39389 3617 39392
rect 3651 39389 3663 39423
rect 3605 39383 3663 39389
rect 3973 39423 4031 39429
rect 3973 39389 3985 39423
rect 4019 39389 4031 39423
rect 3973 39383 4031 39389
rect 4246 39380 4252 39432
rect 4304 39420 4310 39432
rect 4341 39423 4399 39429
rect 4341 39420 4353 39423
rect 4304 39392 4353 39420
rect 4304 39380 4310 39392
rect 4341 39389 4353 39392
rect 4387 39389 4399 39423
rect 4341 39383 4399 39389
rect 5166 39380 5172 39432
rect 5224 39429 5230 39432
rect 5224 39423 5252 39429
rect 5240 39389 5252 39423
rect 5224 39383 5252 39389
rect 6273 39423 6331 39429
rect 6273 39389 6285 39423
rect 6319 39389 6331 39423
rect 6273 39383 6331 39389
rect 5224 39380 5230 39383
rect 3142 39312 3148 39364
rect 3200 39312 3206 39364
rect 992 39256 2774 39284
rect 992 39244 998 39256
rect 3050 39244 3056 39296
rect 3108 39244 3114 39296
rect 3160 39284 3188 39312
rect 5997 39287 6055 39293
rect 5997 39284 6009 39287
rect 3160 39256 6009 39284
rect 5997 39253 6009 39256
rect 6043 39253 6055 39287
rect 5997 39247 6055 39253
rect 6086 39244 6092 39296
rect 6144 39284 6150 39296
rect 6288 39284 6316 39383
rect 7006 39380 7012 39432
rect 7064 39380 7070 39432
rect 7190 39429 7196 39432
rect 7147 39423 7196 39429
rect 7147 39389 7159 39423
rect 7193 39389 7196 39423
rect 7147 39383 7196 39389
rect 7190 39380 7196 39383
rect 7248 39380 7254 39432
rect 9490 39420 9496 39432
rect 9451 39392 9496 39420
rect 9490 39380 9496 39392
rect 9548 39380 9554 39432
rect 10873 39423 10931 39429
rect 10873 39389 10885 39423
rect 10919 39420 10931 39423
rect 11147 39423 11205 39429
rect 10919 39392 11100 39420
rect 10919 39389 10931 39392
rect 10873 39383 10931 39389
rect 7926 39312 7932 39364
rect 7984 39352 7990 39364
rect 11072 39352 11100 39392
rect 11147 39389 11159 39423
rect 11193 39420 11205 39423
rect 11606 39420 11612 39432
rect 11193 39392 11612 39420
rect 11193 39389 11205 39392
rect 11147 39383 11205 39389
rect 11606 39380 11612 39392
rect 11664 39380 11670 39432
rect 12495 39423 12553 39429
rect 12495 39420 12507 39423
rect 11716 39392 12507 39420
rect 11330 39352 11336 39364
rect 7984 39324 10824 39352
rect 11072 39324 11336 39352
rect 7984 39312 7990 39324
rect 6144 39256 6316 39284
rect 6144 39244 6150 39256
rect 7190 39244 7196 39296
rect 7248 39284 7254 39296
rect 10134 39284 10140 39296
rect 7248 39256 10140 39284
rect 7248 39244 7254 39256
rect 10134 39244 10140 39256
rect 10192 39244 10198 39296
rect 10226 39244 10232 39296
rect 10284 39244 10290 39296
rect 10796 39284 10824 39324
rect 11330 39312 11336 39324
rect 11388 39312 11394 39364
rect 11716 39284 11744 39392
rect 12495 39389 12507 39392
rect 12541 39389 12553 39423
rect 12495 39383 12553 39389
rect 20162 39380 20168 39432
rect 20220 39420 20226 39432
rect 20993 39423 21051 39429
rect 20993 39420 21005 39423
rect 20220 39392 21005 39420
rect 20220 39380 20226 39392
rect 20993 39389 21005 39392
rect 21039 39389 21051 39423
rect 20993 39383 21051 39389
rect 21266 39380 21272 39432
rect 21324 39380 21330 39432
rect 21545 39423 21603 39429
rect 21545 39389 21557 39423
rect 21591 39389 21603 39423
rect 21545 39383 21603 39389
rect 21821 39423 21879 39429
rect 21821 39389 21833 39423
rect 21867 39420 21879 39423
rect 22020 39420 22048 39596
rect 22462 39584 22468 39636
rect 22520 39584 22526 39636
rect 22554 39584 22560 39636
rect 22612 39584 22618 39636
rect 22741 39627 22799 39633
rect 22741 39593 22753 39627
rect 22787 39624 22799 39627
rect 23566 39624 23572 39636
rect 22787 39596 23572 39624
rect 22787 39593 22799 39596
rect 22741 39587 22799 39593
rect 23566 39584 23572 39596
rect 23624 39584 23630 39636
rect 22189 39559 22247 39565
rect 22189 39525 22201 39559
rect 22235 39556 22247 39559
rect 22572 39556 22600 39584
rect 22235 39528 22600 39556
rect 23477 39559 23535 39565
rect 22235 39525 22247 39528
rect 22189 39519 22247 39525
rect 23477 39525 23489 39559
rect 23523 39525 23535 39559
rect 23477 39519 23535 39525
rect 22554 39448 22560 39500
rect 22612 39488 22618 39500
rect 23492 39488 23520 39519
rect 22612 39460 23336 39488
rect 23492 39460 23980 39488
rect 22612 39448 22618 39460
rect 21867 39392 22048 39420
rect 22097 39423 22155 39429
rect 21867 39389 21879 39392
rect 21821 39383 21879 39389
rect 22097 39389 22109 39423
rect 22143 39389 22155 39423
rect 22373 39423 22431 39429
rect 22373 39420 22385 39423
rect 22097 39383 22155 39389
rect 22204 39392 22385 39420
rect 19334 39312 19340 39364
rect 19392 39352 19398 39364
rect 21560 39352 21588 39383
rect 19392 39324 21588 39352
rect 19392 39312 19398 39324
rect 22002 39312 22008 39364
rect 22060 39352 22066 39364
rect 22112 39352 22140 39383
rect 22060 39324 22140 39352
rect 22060 39312 22066 39324
rect 10796 39256 11744 39284
rect 11885 39287 11943 39293
rect 11885 39253 11897 39287
rect 11931 39284 11943 39287
rect 12710 39284 12716 39296
rect 11931 39256 12716 39284
rect 11931 39253 11943 39256
rect 11885 39247 11943 39253
rect 12710 39244 12716 39256
rect 12768 39244 12774 39296
rect 13262 39244 13268 39296
rect 13320 39244 13326 39296
rect 17954 39244 17960 39296
rect 18012 39284 18018 39296
rect 21634 39284 21640 39296
rect 18012 39256 21640 39284
rect 18012 39244 18018 39256
rect 21634 39244 21640 39256
rect 21692 39244 21698 39296
rect 22094 39244 22100 39296
rect 22152 39284 22158 39296
rect 22204 39284 22232 39392
rect 22373 39389 22385 39392
rect 22419 39389 22431 39423
rect 22373 39383 22431 39389
rect 22462 39380 22468 39432
rect 22520 39420 22526 39432
rect 22649 39423 22707 39429
rect 22649 39420 22661 39423
rect 22520 39392 22661 39420
rect 22520 39380 22526 39392
rect 22649 39389 22661 39392
rect 22695 39389 22707 39423
rect 22649 39383 22707 39389
rect 22738 39380 22744 39432
rect 22796 39420 22802 39432
rect 22925 39423 22983 39429
rect 22925 39420 22937 39423
rect 22796 39392 22937 39420
rect 22796 39380 22802 39392
rect 22925 39389 22937 39392
rect 22971 39389 22983 39423
rect 22925 39383 22983 39389
rect 23201 39423 23259 39429
rect 23201 39389 23213 39423
rect 23247 39389 23259 39423
rect 23308 39420 23336 39460
rect 23952 39429 23980 39460
rect 23661 39423 23719 39429
rect 23661 39420 23673 39423
rect 23308 39392 23673 39420
rect 23201 39383 23259 39389
rect 23661 39389 23673 39392
rect 23707 39389 23719 39423
rect 23661 39383 23719 39389
rect 23937 39423 23995 39429
rect 23937 39389 23949 39423
rect 23983 39389 23995 39423
rect 23937 39383 23995 39389
rect 22278 39312 22284 39364
rect 22336 39352 22342 39364
rect 23216 39352 23244 39383
rect 22336 39324 23244 39352
rect 22336 39312 22342 39324
rect 22152 39256 22232 39284
rect 22152 39244 22158 39256
rect 23014 39244 23020 39296
rect 23072 39244 23078 39296
rect 24118 39244 24124 39296
rect 24176 39244 24182 39296
rect 1104 39194 25000 39216
rect 1104 39142 6884 39194
rect 6936 39142 6948 39194
rect 7000 39142 7012 39194
rect 7064 39142 7076 39194
rect 7128 39142 7140 39194
rect 7192 39142 12818 39194
rect 12870 39142 12882 39194
rect 12934 39142 12946 39194
rect 12998 39142 13010 39194
rect 13062 39142 13074 39194
rect 13126 39142 18752 39194
rect 18804 39142 18816 39194
rect 18868 39142 18880 39194
rect 18932 39142 18944 39194
rect 18996 39142 19008 39194
rect 19060 39142 24686 39194
rect 24738 39142 24750 39194
rect 24802 39142 24814 39194
rect 24866 39142 24878 39194
rect 24930 39142 24942 39194
rect 24994 39142 25000 39194
rect 1104 39120 25000 39142
rect 1854 39040 1860 39092
rect 1912 39080 1918 39092
rect 1912 39052 2774 39080
rect 1912 39040 1918 39052
rect 2746 39012 2774 39052
rect 3142 39040 3148 39092
rect 3200 39080 3206 39092
rect 3418 39080 3424 39092
rect 3200 39052 3424 39080
rect 3200 39040 3206 39052
rect 3418 39040 3424 39052
rect 3476 39040 3482 39092
rect 3786 39040 3792 39092
rect 3844 39080 3850 39092
rect 6086 39080 6092 39092
rect 3844 39052 6092 39080
rect 3844 39040 3850 39052
rect 6086 39040 6092 39052
rect 6144 39040 6150 39092
rect 6270 39040 6276 39092
rect 6328 39080 6334 39092
rect 6454 39080 6460 39092
rect 6328 39052 6460 39080
rect 6328 39040 6334 39052
rect 6454 39040 6460 39052
rect 6512 39040 6518 39092
rect 6638 39040 6644 39092
rect 6696 39080 6702 39092
rect 8386 39080 8392 39092
rect 6696 39052 8392 39080
rect 6696 39040 6702 39052
rect 8386 39040 8392 39052
rect 8444 39040 8450 39092
rect 10226 39080 10232 39092
rect 9140 39052 10232 39080
rect 3513 39015 3571 39021
rect 2746 38984 3280 39012
rect 3252 38956 3280 38984
rect 3513 38981 3525 39015
rect 3559 39012 3571 39015
rect 4249 39015 4307 39021
rect 3559 38984 4200 39012
rect 3559 38981 3571 38984
rect 3513 38975 3571 38981
rect 1394 38904 1400 38956
rect 1452 38904 1458 38956
rect 1854 38904 1860 38956
rect 1912 38944 1918 38956
rect 2038 38944 2044 38956
rect 1912 38916 2044 38944
rect 1912 38904 1918 38916
rect 2038 38904 2044 38916
rect 2096 38904 2102 38956
rect 2409 38947 2467 38953
rect 2409 38913 2421 38947
rect 2455 38944 2467 38947
rect 2774 38944 2780 38956
rect 2455 38916 2780 38944
rect 2455 38913 2467 38916
rect 2409 38907 2467 38913
rect 2774 38904 2780 38916
rect 2832 38904 2838 38956
rect 3234 38904 3240 38956
rect 3292 38904 3298 38956
rect 3418 38904 3424 38956
rect 3476 38904 3482 38956
rect 3786 38904 3792 38956
rect 3844 38944 3850 38956
rect 3881 38947 3939 38953
rect 3881 38944 3893 38947
rect 3844 38916 3893 38944
rect 3844 38904 3850 38916
rect 3881 38913 3893 38916
rect 3927 38913 3939 38947
rect 4172 38944 4200 38984
rect 4249 38981 4261 39015
rect 4295 39012 4307 39015
rect 4338 39012 4344 39024
rect 4295 38984 4344 39012
rect 4295 38981 4307 38984
rect 4249 38975 4307 38981
rect 4338 38972 4344 38984
rect 4396 38972 4402 39024
rect 4522 38972 4528 39024
rect 4580 39012 4586 39024
rect 4580 38984 8064 39012
rect 4580 38972 4586 38984
rect 4798 38944 4804 38956
rect 4172 38916 4804 38944
rect 3881 38907 3939 38913
rect 4798 38904 4804 38916
rect 4856 38904 4862 38956
rect 5350 38904 5356 38956
rect 5408 38944 5414 38956
rect 7009 38947 7067 38953
rect 7009 38944 7021 38947
rect 5408 38916 7021 38944
rect 5408 38904 5414 38916
rect 7009 38913 7021 38916
rect 7055 38944 7067 38947
rect 7190 38944 7196 38956
rect 7055 38916 7196 38944
rect 7055 38913 7067 38916
rect 7009 38907 7067 38913
rect 7190 38904 7196 38916
rect 7248 38904 7254 38956
rect 7283 38947 7341 38953
rect 7283 38913 7295 38947
rect 7329 38944 7341 38947
rect 7926 38944 7932 38956
rect 7329 38916 7932 38944
rect 7329 38913 7341 38916
rect 7283 38907 7341 38913
rect 7926 38904 7932 38916
rect 7984 38904 7990 38956
rect 8036 38944 8064 38984
rect 8294 38972 8300 39024
rect 8352 39012 8358 39024
rect 8573 39015 8631 39021
rect 8573 39012 8585 39015
rect 8352 38984 8585 39012
rect 8352 38972 8358 38984
rect 8573 38981 8585 38984
rect 8619 38981 8631 39015
rect 8573 38975 8631 38981
rect 8662 38944 8668 38956
rect 8036 38916 8668 38944
rect 8662 38904 8668 38916
rect 8720 38944 8726 38956
rect 8849 38947 8907 38953
rect 8849 38944 8861 38947
rect 8720 38916 8861 38944
rect 8720 38904 8726 38916
rect 8849 38913 8861 38916
rect 8895 38913 8907 38947
rect 8849 38907 8907 38913
rect 8941 38947 8999 38953
rect 8941 38913 8953 38947
rect 8987 38944 8999 38947
rect 9140 38944 9168 39052
rect 10226 39040 10232 39052
rect 10284 39040 10290 39092
rect 12250 39040 12256 39092
rect 12308 39080 12314 39092
rect 13357 39083 13415 39089
rect 13357 39080 13369 39083
rect 12308 39052 13369 39080
rect 12308 39040 12314 39052
rect 13357 39049 13369 39052
rect 13403 39049 13415 39083
rect 13357 39043 13415 39049
rect 20162 39040 20168 39092
rect 20220 39040 20226 39092
rect 20441 39083 20499 39089
rect 20441 39049 20453 39083
rect 20487 39080 20499 39083
rect 20714 39080 20720 39092
rect 20487 39052 20720 39080
rect 20487 39049 20499 39052
rect 20441 39043 20499 39049
rect 20714 39040 20720 39052
rect 20772 39040 20778 39092
rect 21085 39083 21143 39089
rect 21085 39049 21097 39083
rect 21131 39049 21143 39083
rect 21085 39043 21143 39049
rect 22281 39083 22339 39089
rect 22281 39049 22293 39083
rect 22327 39080 22339 39083
rect 22327 39052 22792 39080
rect 22327 39049 22339 39052
rect 22281 39043 22339 39049
rect 9398 38972 9404 39024
rect 9456 39012 9462 39024
rect 9456 38984 9812 39012
rect 9456 38972 9462 38984
rect 8987 38916 9168 38944
rect 8987 38913 8999 38916
rect 8941 38907 8999 38913
rect 9214 38904 9220 38956
rect 9272 38944 9278 38956
rect 9309 38947 9367 38953
rect 9309 38944 9321 38947
rect 9272 38916 9321 38944
rect 9272 38904 9278 38916
rect 9309 38913 9321 38916
rect 9355 38913 9367 38947
rect 9309 38907 9367 38913
rect 9674 38904 9680 38956
rect 9732 38953 9738 38956
rect 9732 38947 9749 38953
rect 9737 38913 9749 38947
rect 9732 38907 9749 38913
rect 9732 38904 9738 38907
rect 2222 38836 2228 38888
rect 2280 38836 2286 38888
rect 2593 38879 2651 38885
rect 2593 38845 2605 38879
rect 2639 38845 2651 38879
rect 2593 38839 2651 38845
rect 2038 38768 2044 38820
rect 2096 38808 2102 38820
rect 2608 38808 2636 38839
rect 3050 38836 3056 38888
rect 3108 38836 3114 38888
rect 4246 38836 4252 38888
rect 4304 38876 4310 38888
rect 4304 38848 4660 38876
rect 4304 38836 4310 38848
rect 2096 38780 2636 38808
rect 2096 38768 2102 38780
rect 4433 38743 4491 38749
rect 4433 38709 4445 38743
rect 4479 38740 4491 38743
rect 4522 38740 4528 38752
rect 4479 38712 4528 38740
rect 4479 38709 4491 38712
rect 4433 38703 4491 38709
rect 4522 38700 4528 38712
rect 4580 38700 4586 38752
rect 4632 38740 4660 38848
rect 8036 38848 8418 38876
rect 8036 38817 8064 38848
rect 8021 38811 8079 38817
rect 8021 38777 8033 38811
rect 8067 38777 8079 38811
rect 9784 38808 9812 38984
rect 10060 38984 11376 39012
rect 10060 38953 10088 38984
rect 11348 38956 11376 38984
rect 18322 38972 18328 39024
rect 18380 39012 18386 39024
rect 21100 39012 21128 39043
rect 22646 39012 22652 39024
rect 18380 38984 21036 39012
rect 21100 38984 21864 39012
rect 18380 38972 18386 38984
rect 10045 38947 10103 38953
rect 10045 38913 10057 38947
rect 10091 38913 10103 38947
rect 10045 38907 10103 38913
rect 10226 38904 10232 38956
rect 10284 38944 10290 38956
rect 10319 38947 10377 38953
rect 10319 38944 10331 38947
rect 10284 38916 10331 38944
rect 10284 38904 10290 38916
rect 10319 38913 10331 38916
rect 10365 38913 10377 38947
rect 10319 38907 10377 38913
rect 11330 38904 11336 38956
rect 11388 38904 11394 38956
rect 12434 38904 12440 38956
rect 12492 38904 12498 38956
rect 12710 38904 12716 38956
rect 12768 38904 12774 38956
rect 19426 38904 19432 38956
rect 19484 38904 19490 38956
rect 20346 38904 20352 38956
rect 20404 38904 20410 38956
rect 20625 38947 20683 38953
rect 20625 38913 20637 38947
rect 20671 38913 20683 38947
rect 20625 38907 20683 38913
rect 11514 38836 11520 38888
rect 11572 38836 11578 38888
rect 11698 38836 11704 38888
rect 11756 38836 11762 38888
rect 12554 38879 12612 38885
rect 12554 38876 12566 38879
rect 12268 38848 12566 38876
rect 9861 38811 9919 38817
rect 9861 38808 9873 38811
rect 9784 38780 9873 38808
rect 8021 38771 8079 38777
rect 9861 38777 9873 38780
rect 9907 38777 9919 38811
rect 9861 38771 9919 38777
rect 11057 38811 11115 38817
rect 11057 38777 11069 38811
rect 11103 38808 11115 38811
rect 12161 38811 12219 38817
rect 12161 38808 12173 38811
rect 11103 38780 12173 38808
rect 11103 38777 11115 38780
rect 11057 38771 11115 38777
rect 12161 38777 12173 38780
rect 12207 38777 12219 38811
rect 12161 38771 12219 38777
rect 8386 38740 8392 38752
rect 4632 38712 8392 38740
rect 8386 38700 8392 38712
rect 8444 38700 8450 38752
rect 9876 38740 9904 38771
rect 11790 38740 11796 38752
rect 9876 38712 11796 38740
rect 11790 38700 11796 38712
rect 11848 38740 11854 38752
rect 12268 38740 12296 38848
rect 12554 38845 12566 38848
rect 12600 38845 12612 38879
rect 20640 38876 20668 38907
rect 12554 38839 12612 38845
rect 15212 38848 20668 38876
rect 15212 38808 15240 38848
rect 13096 38780 15240 38808
rect 19245 38811 19303 38817
rect 11848 38712 12296 38740
rect 11848 38700 11854 38712
rect 12618 38700 12624 38752
rect 12676 38740 12682 38752
rect 13096 38740 13124 38780
rect 19245 38777 19257 38811
rect 19291 38808 19303 38811
rect 21008 38808 21036 38984
rect 21836 38953 21864 38984
rect 21928 38984 22652 39012
rect 21269 38947 21327 38953
rect 21269 38913 21281 38947
rect 21315 38913 21327 38947
rect 21269 38907 21327 38913
rect 21821 38947 21879 38953
rect 21821 38913 21833 38947
rect 21867 38913 21879 38947
rect 21821 38907 21879 38913
rect 21284 38876 21312 38907
rect 21358 38876 21364 38888
rect 21284 38848 21364 38876
rect 21358 38836 21364 38848
rect 21416 38836 21422 38888
rect 21928 38876 21956 38984
rect 22646 38972 22652 38984
rect 22704 38972 22710 39024
rect 22764 38959 22792 39052
rect 22922 39040 22928 39092
rect 22980 39040 22986 39092
rect 23014 39040 23020 39092
rect 23072 39040 23078 39092
rect 23106 39040 23112 39092
rect 23164 39080 23170 39092
rect 23201 39083 23259 39089
rect 23201 39080 23213 39083
rect 23164 39052 23213 39080
rect 23164 39040 23170 39052
rect 23201 39049 23213 39052
rect 23247 39049 23259 39083
rect 23201 39043 23259 39049
rect 23290 39040 23296 39092
rect 23348 39080 23354 39092
rect 23753 39083 23811 39089
rect 23753 39080 23765 39083
rect 23348 39052 23765 39080
rect 23348 39040 23354 39052
rect 23753 39049 23765 39052
rect 23799 39049 23811 39083
rect 23753 39043 23811 39049
rect 22462 38904 22468 38956
rect 22520 38904 22526 38956
rect 22749 38953 22807 38959
rect 22557 38947 22615 38953
rect 22557 38913 22569 38947
rect 22603 38944 22615 38947
rect 22603 38916 22692 38944
rect 22603 38913 22615 38916
rect 22557 38907 22615 38913
rect 21468 38848 21956 38876
rect 22664 38876 22692 38916
rect 22749 38919 22761 38953
rect 22795 38919 22807 38953
rect 22749 38913 22807 38919
rect 23032 38944 23060 39040
rect 25222 39012 25228 39024
rect 23676 38984 25228 39012
rect 23109 38947 23167 38953
rect 23109 38944 23121 38947
rect 23032 38916 23121 38944
rect 23109 38913 23121 38916
rect 23155 38913 23167 38947
rect 23109 38907 23167 38913
rect 23382 38904 23388 38956
rect 23440 38904 23446 38956
rect 23676 38953 23704 38984
rect 25222 38972 25228 38984
rect 25280 38972 25286 39024
rect 23661 38947 23719 38953
rect 23661 38913 23673 38947
rect 23707 38913 23719 38947
rect 23661 38907 23719 38913
rect 23937 38947 23995 38953
rect 23937 38913 23949 38947
rect 23983 38913 23995 38947
rect 23937 38907 23995 38913
rect 22922 38876 22928 38888
rect 22664 38848 22928 38876
rect 21468 38808 21496 38848
rect 22922 38836 22928 38848
rect 22980 38836 22986 38888
rect 23566 38836 23572 38888
rect 23624 38876 23630 38888
rect 23952 38876 23980 38907
rect 24026 38904 24032 38956
rect 24084 38944 24090 38956
rect 24121 38947 24179 38953
rect 24121 38944 24133 38947
rect 24084 38916 24133 38944
rect 24084 38904 24090 38916
rect 24121 38913 24133 38916
rect 24167 38913 24179 38947
rect 24121 38907 24179 38913
rect 23624 38848 23980 38876
rect 23624 38836 23630 38848
rect 19291 38780 20944 38808
rect 21008 38780 21496 38808
rect 21560 38780 22784 38808
rect 19291 38777 19303 38780
rect 19245 38771 19303 38777
rect 12676 38712 13124 38740
rect 12676 38700 12682 38712
rect 13630 38700 13636 38752
rect 13688 38700 13694 38752
rect 14274 38700 14280 38752
rect 14332 38740 14338 38752
rect 16114 38740 16120 38752
rect 14332 38712 16120 38740
rect 14332 38700 14338 38712
rect 16114 38700 16120 38712
rect 16172 38700 16178 38752
rect 20916 38740 20944 38780
rect 21560 38740 21588 38780
rect 20916 38712 21588 38740
rect 21913 38743 21971 38749
rect 21913 38709 21925 38743
rect 21959 38740 21971 38743
rect 22370 38740 22376 38752
rect 21959 38712 22376 38740
rect 21959 38709 21971 38712
rect 21913 38703 21971 38709
rect 22370 38700 22376 38712
rect 22428 38700 22434 38752
rect 22646 38700 22652 38752
rect 22704 38700 22710 38752
rect 22756 38740 22784 38780
rect 23474 38768 23480 38820
rect 23532 38768 23538 38820
rect 23934 38768 23940 38820
rect 23992 38768 23998 38820
rect 23952 38740 23980 38768
rect 22756 38712 23980 38740
rect 24394 38700 24400 38752
rect 24452 38700 24458 38752
rect 1104 38650 24840 38672
rect 1104 38598 3917 38650
rect 3969 38598 3981 38650
rect 4033 38598 4045 38650
rect 4097 38598 4109 38650
rect 4161 38598 4173 38650
rect 4225 38598 9851 38650
rect 9903 38598 9915 38650
rect 9967 38598 9979 38650
rect 10031 38598 10043 38650
rect 10095 38598 10107 38650
rect 10159 38598 15785 38650
rect 15837 38598 15849 38650
rect 15901 38598 15913 38650
rect 15965 38598 15977 38650
rect 16029 38598 16041 38650
rect 16093 38598 21719 38650
rect 21771 38598 21783 38650
rect 21835 38598 21847 38650
rect 21899 38598 21911 38650
rect 21963 38598 21975 38650
rect 22027 38598 24840 38650
rect 1104 38576 24840 38598
rect 3804 38508 4752 38536
rect 2225 38403 2283 38409
rect 2225 38369 2237 38403
rect 2271 38400 2283 38403
rect 2498 38400 2504 38412
rect 2271 38372 2504 38400
rect 2271 38369 2283 38372
rect 2225 38363 2283 38369
rect 2498 38360 2504 38372
rect 2556 38360 2562 38412
rect 3050 38400 3056 38412
rect 2884 38372 3056 38400
rect 1394 38292 1400 38344
rect 1452 38292 1458 38344
rect 2409 38335 2467 38341
rect 2409 38301 2421 38335
rect 2455 38332 2467 38335
rect 2884 38332 2912 38372
rect 3050 38360 3056 38372
rect 3108 38360 3114 38412
rect 3145 38403 3203 38409
rect 3145 38369 3157 38403
rect 3191 38400 3203 38403
rect 3191 38372 3280 38400
rect 3191 38369 3203 38372
rect 3145 38363 3203 38369
rect 3252 38344 3280 38372
rect 2455 38304 2912 38332
rect 2961 38335 3019 38341
rect 2455 38301 2467 38304
rect 2409 38295 2467 38301
rect 2961 38301 2973 38335
rect 3007 38301 3019 38335
rect 2961 38295 3019 38301
rect 2682 38224 2688 38276
rect 2740 38224 2746 38276
rect 1210 38156 1216 38208
rect 1268 38196 1274 38208
rect 2976 38196 3004 38295
rect 3234 38292 3240 38344
rect 3292 38292 3298 38344
rect 3510 38292 3516 38344
rect 3568 38332 3574 38344
rect 3804 38341 3832 38508
rect 4724 38468 4752 38508
rect 4798 38496 4804 38548
rect 4856 38496 4862 38548
rect 6730 38496 6736 38548
rect 6788 38536 6794 38548
rect 6788 38508 8156 38536
rect 6788 38496 6794 38508
rect 5350 38468 5356 38480
rect 4724 38440 5356 38468
rect 5350 38428 5356 38440
rect 5408 38428 5414 38480
rect 8128 38468 8156 38508
rect 8386 38496 8392 38548
rect 8444 38536 8450 38548
rect 9214 38536 9220 38548
rect 8444 38508 9220 38536
rect 8444 38496 8450 38508
rect 9214 38496 9220 38508
rect 9272 38496 9278 38548
rect 12618 38536 12624 38548
rect 10244 38508 12624 38536
rect 8938 38468 8944 38480
rect 8128 38440 8944 38468
rect 8938 38428 8944 38440
rect 8996 38468 9002 38480
rect 9306 38468 9312 38480
rect 8996 38440 9312 38468
rect 8996 38428 9002 38440
rect 9306 38428 9312 38440
rect 9364 38428 9370 38480
rect 3789 38335 3847 38341
rect 3789 38332 3801 38335
rect 3568 38304 3801 38332
rect 3568 38292 3574 38304
rect 3789 38301 3801 38304
rect 3835 38301 3847 38335
rect 4062 38332 4068 38344
rect 4023 38304 4068 38332
rect 3789 38295 3847 38301
rect 4062 38292 4068 38304
rect 4120 38292 4126 38344
rect 7282 38292 7288 38344
rect 7340 38332 7346 38344
rect 7469 38335 7527 38341
rect 7469 38332 7481 38335
rect 7340 38304 7481 38332
rect 7340 38292 7346 38304
rect 7469 38301 7481 38304
rect 7515 38301 7527 38335
rect 10134 38332 10140 38344
rect 7742 38311 10140 38332
rect 7469 38295 7527 38301
rect 7727 38305 10140 38311
rect 7727 38271 7739 38305
rect 7773 38304 10140 38305
rect 7773 38271 7785 38304
rect 10134 38292 10140 38304
rect 10192 38292 10198 38344
rect 10244 38341 10272 38508
rect 12618 38496 12624 38508
rect 12676 38496 12682 38548
rect 13262 38536 13268 38548
rect 12728 38508 13268 38536
rect 12728 38477 12756 38508
rect 13262 38496 13268 38508
rect 13320 38496 13326 38548
rect 18693 38539 18751 38545
rect 18693 38505 18705 38539
rect 18739 38536 18751 38539
rect 19426 38536 19432 38548
rect 18739 38508 19432 38536
rect 18739 38505 18751 38508
rect 18693 38499 18751 38505
rect 19426 38496 19432 38508
rect 19484 38496 19490 38548
rect 22005 38539 22063 38545
rect 22005 38505 22017 38539
rect 22051 38536 22063 38539
rect 22462 38536 22468 38548
rect 22051 38508 22468 38536
rect 22051 38505 22063 38508
rect 22005 38499 22063 38505
rect 22462 38496 22468 38508
rect 22520 38496 22526 38548
rect 23477 38539 23535 38545
rect 23477 38505 23489 38539
rect 23523 38536 23535 38539
rect 24026 38536 24032 38548
rect 23523 38508 24032 38536
rect 23523 38505 23535 38508
rect 23477 38499 23535 38505
rect 24026 38496 24032 38508
rect 24084 38496 24090 38548
rect 12713 38471 12771 38477
rect 12713 38437 12725 38471
rect 12759 38437 12771 38471
rect 12713 38431 12771 38437
rect 11698 38360 11704 38412
rect 11756 38400 11762 38412
rect 12253 38403 12311 38409
rect 12253 38400 12265 38403
rect 11756 38372 12265 38400
rect 11756 38360 11762 38372
rect 12253 38369 12265 38372
rect 12299 38400 12311 38403
rect 12342 38400 12348 38412
rect 12299 38372 12348 38400
rect 12299 38369 12311 38372
rect 12253 38363 12311 38369
rect 12342 38360 12348 38372
rect 12400 38360 12406 38412
rect 12989 38403 13047 38409
rect 12989 38369 13001 38403
rect 13035 38400 13047 38403
rect 13630 38400 13636 38412
rect 13035 38372 13636 38400
rect 13035 38369 13047 38372
rect 12989 38363 13047 38369
rect 13630 38360 13636 38372
rect 13688 38360 13694 38412
rect 19242 38360 19248 38412
rect 19300 38400 19306 38412
rect 19702 38400 19708 38412
rect 19300 38372 19708 38400
rect 19300 38360 19306 38372
rect 19702 38360 19708 38372
rect 19760 38400 19766 38412
rect 20625 38403 20683 38409
rect 20625 38400 20637 38403
rect 19760 38372 20637 38400
rect 19760 38360 19766 38372
rect 20625 38369 20637 38372
rect 20671 38369 20683 38403
rect 20625 38363 20683 38369
rect 10229 38335 10287 38341
rect 10229 38301 10241 38335
rect 10275 38301 10287 38335
rect 10229 38295 10287 38301
rect 10487 38305 10545 38311
rect 7727 38265 7785 38271
rect 1268 38168 3004 38196
rect 1268 38156 1274 38168
rect 5994 38156 6000 38208
rect 6052 38196 6058 38208
rect 7742 38196 7770 38265
rect 8202 38224 8208 38276
rect 8260 38264 8266 38276
rect 8260 38236 9812 38264
rect 8260 38224 8266 38236
rect 9784 38208 9812 38236
rect 6052 38168 7770 38196
rect 6052 38156 6058 38168
rect 8478 38156 8484 38208
rect 8536 38156 8542 38208
rect 9766 38156 9772 38208
rect 9824 38156 9830 38208
rect 10244 38196 10272 38295
rect 10487 38271 10499 38305
rect 10533 38302 10545 38305
rect 10533 38271 10546 38302
rect 11146 38292 11152 38344
rect 11204 38332 11210 38344
rect 12069 38335 12127 38341
rect 12069 38332 12081 38335
rect 11204 38304 12081 38332
rect 11204 38292 11210 38304
rect 12069 38301 12081 38304
rect 12115 38301 12127 38335
rect 12069 38295 12127 38301
rect 13078 38292 13084 38344
rect 13136 38341 13142 38344
rect 13136 38335 13164 38341
rect 13152 38301 13164 38335
rect 13136 38295 13164 38301
rect 13136 38292 13142 38295
rect 13262 38292 13268 38344
rect 13320 38292 13326 38344
rect 18138 38292 18144 38344
rect 18196 38332 18202 38344
rect 18877 38335 18935 38341
rect 18877 38332 18889 38335
rect 18196 38304 18889 38332
rect 18196 38292 18202 38304
rect 18877 38301 18889 38304
rect 18923 38301 18935 38335
rect 18877 38295 18935 38301
rect 19610 38292 19616 38344
rect 19668 38292 19674 38344
rect 22094 38292 22100 38344
rect 22152 38292 22158 38344
rect 22370 38341 22376 38344
rect 22339 38335 22376 38341
rect 22339 38301 22351 38335
rect 22339 38295 22376 38301
rect 22370 38292 22376 38295
rect 22428 38292 22434 38344
rect 22462 38292 22468 38344
rect 22520 38332 22526 38344
rect 23661 38335 23719 38341
rect 23661 38332 23673 38335
rect 22520 38304 23673 38332
rect 22520 38292 22526 38304
rect 23661 38301 23673 38304
rect 23707 38301 23719 38335
rect 23661 38295 23719 38301
rect 23937 38335 23995 38341
rect 23937 38301 23949 38335
rect 23983 38301 23995 38335
rect 23937 38295 23995 38301
rect 10487 38265 10546 38271
rect 10518 38264 10546 38265
rect 10594 38264 10600 38276
rect 10518 38236 10600 38264
rect 10594 38224 10600 38236
rect 10652 38264 10658 38276
rect 13909 38267 13967 38273
rect 10652 38236 11376 38264
rect 10652 38224 10658 38236
rect 10318 38196 10324 38208
rect 10244 38168 10324 38196
rect 10318 38156 10324 38168
rect 10376 38156 10382 38208
rect 11238 38156 11244 38208
rect 11296 38156 11302 38208
rect 11348 38196 11376 38236
rect 13909 38233 13921 38267
rect 13955 38264 13967 38267
rect 20870 38267 20928 38273
rect 20870 38264 20882 38267
rect 13955 38236 20882 38264
rect 13955 38233 13967 38236
rect 13909 38227 13967 38233
rect 20870 38233 20882 38236
rect 20916 38264 20928 38267
rect 21358 38264 21364 38276
rect 20916 38236 21364 38264
rect 20916 38233 20928 38236
rect 20870 38227 20928 38233
rect 21358 38224 21364 38236
rect 21416 38224 21422 38276
rect 23952 38264 23980 38295
rect 22066 38236 23980 38264
rect 12434 38196 12440 38208
rect 11348 38168 12440 38196
rect 12434 38156 12440 38168
rect 12492 38156 12498 38208
rect 12526 38156 12532 38208
rect 12584 38196 12590 38208
rect 13078 38196 13084 38208
rect 12584 38168 13084 38196
rect 12584 38156 12590 38168
rect 13078 38156 13084 38168
rect 13136 38156 13142 38208
rect 19429 38199 19487 38205
rect 19429 38165 19441 38199
rect 19475 38196 19487 38199
rect 20346 38196 20352 38208
rect 19475 38168 20352 38196
rect 19475 38165 19487 38168
rect 19429 38159 19487 38165
rect 20346 38156 20352 38168
rect 20404 38156 20410 38208
rect 21450 38156 21456 38208
rect 21508 38196 21514 38208
rect 22066 38196 22094 38236
rect 21508 38168 22094 38196
rect 21508 38156 21514 38168
rect 22278 38156 22284 38208
rect 22336 38196 22342 38208
rect 22922 38196 22928 38208
rect 22336 38168 22928 38196
rect 22336 38156 22342 38168
rect 22922 38156 22928 38168
rect 22980 38196 22986 38208
rect 23109 38199 23167 38205
rect 23109 38196 23121 38199
rect 22980 38168 23121 38196
rect 22980 38156 22986 38168
rect 23109 38165 23121 38168
rect 23155 38165 23167 38199
rect 23109 38159 23167 38165
rect 24118 38156 24124 38208
rect 24176 38156 24182 38208
rect 1104 38106 25000 38128
rect 1104 38054 6884 38106
rect 6936 38054 6948 38106
rect 7000 38054 7012 38106
rect 7064 38054 7076 38106
rect 7128 38054 7140 38106
rect 7192 38054 12818 38106
rect 12870 38054 12882 38106
rect 12934 38054 12946 38106
rect 12998 38054 13010 38106
rect 13062 38054 13074 38106
rect 13126 38054 18752 38106
rect 18804 38054 18816 38106
rect 18868 38054 18880 38106
rect 18932 38054 18944 38106
rect 18996 38054 19008 38106
rect 19060 38054 24686 38106
rect 24738 38054 24750 38106
rect 24802 38054 24814 38106
rect 24866 38054 24878 38106
rect 24930 38054 24942 38106
rect 24994 38054 25000 38106
rect 1104 38032 25000 38054
rect 1302 37952 1308 38004
rect 1360 37992 1366 38004
rect 1360 37964 3924 37992
rect 1360 37952 1366 37964
rect 2590 37816 2596 37868
rect 2648 37816 2654 37868
rect 3326 37816 3332 37868
rect 3384 37816 3390 37868
rect 3896 37865 3924 37964
rect 6730 37952 6736 38004
rect 6788 37992 6794 38004
rect 9490 37992 9496 38004
rect 6788 37964 9496 37992
rect 6788 37952 6794 37964
rect 9490 37952 9496 37964
rect 9548 37992 9554 38004
rect 10594 37992 10600 38004
rect 9548 37964 10600 37992
rect 9548 37952 9554 37964
rect 10594 37952 10600 37964
rect 10652 37952 10658 38004
rect 13262 37952 13268 38004
rect 13320 37992 13326 38004
rect 13725 37995 13783 38001
rect 13725 37992 13737 37995
rect 13320 37964 13737 37992
rect 13320 37952 13326 37964
rect 13725 37961 13737 37964
rect 13771 37961 13783 37995
rect 13725 37955 13783 37961
rect 18138 37952 18144 38004
rect 18196 37952 18202 38004
rect 20901 37995 20959 38001
rect 20901 37961 20913 37995
rect 20947 37992 20959 37995
rect 21450 37992 21456 38004
rect 20947 37964 21456 37992
rect 20947 37961 20959 37964
rect 20901 37955 20959 37961
rect 21450 37952 21456 37964
rect 21508 37952 21514 38004
rect 21913 37995 21971 38001
rect 21913 37961 21925 37995
rect 21959 37992 21971 37995
rect 23014 37992 23020 38004
rect 21959 37964 23020 37992
rect 21959 37961 21971 37964
rect 21913 37955 21971 37961
rect 23014 37952 23020 37964
rect 23072 37952 23078 38004
rect 23382 37952 23388 38004
rect 23440 37952 23446 38004
rect 8294 37884 8300 37936
rect 8352 37924 8358 37936
rect 8481 37927 8539 37933
rect 8481 37924 8493 37927
rect 8352 37896 8493 37924
rect 8352 37884 8358 37896
rect 8481 37893 8493 37896
rect 8527 37893 8539 37927
rect 8481 37887 8539 37893
rect 8662 37884 8668 37936
rect 8720 37924 8726 37936
rect 8757 37927 8815 37933
rect 8757 37924 8769 37927
rect 8720 37896 8769 37924
rect 8720 37884 8726 37896
rect 8757 37893 8769 37896
rect 8803 37893 8815 37927
rect 8757 37887 8815 37893
rect 8849 37927 8907 37933
rect 8849 37893 8861 37927
rect 8895 37924 8907 37927
rect 8895 37896 9536 37924
rect 8895 37893 8907 37896
rect 8849 37887 8907 37893
rect 3881 37859 3939 37865
rect 3881 37825 3893 37859
rect 3927 37825 3939 37859
rect 3881 37819 3939 37825
rect 4062 37816 4068 37868
rect 4120 37856 4126 37868
rect 4859 37859 4917 37865
rect 4859 37856 4871 37859
rect 4120 37828 4871 37856
rect 4120 37816 4126 37828
rect 4859 37825 4871 37828
rect 4905 37825 4917 37859
rect 4859 37819 4917 37825
rect 7377 37859 7435 37865
rect 7377 37825 7389 37859
rect 7423 37825 7435 37859
rect 7377 37819 7435 37825
rect 1397 37791 1455 37797
rect 1397 37757 1409 37791
rect 1443 37757 1455 37791
rect 1397 37751 1455 37757
rect 1581 37791 1639 37797
rect 1581 37757 1593 37791
rect 1627 37788 1639 37791
rect 1762 37788 1768 37800
rect 1627 37760 1768 37788
rect 1627 37757 1639 37760
rect 1581 37751 1639 37757
rect 1412 37720 1440 37751
rect 1762 37748 1768 37760
rect 1820 37748 1826 37800
rect 2314 37748 2320 37800
rect 2372 37748 2378 37800
rect 2455 37791 2513 37797
rect 2455 37757 2467 37791
rect 2501 37788 2513 37791
rect 3142 37788 3148 37800
rect 2501 37760 3148 37788
rect 2501 37757 2513 37760
rect 2455 37751 2513 37757
rect 3142 37748 3148 37760
rect 3200 37788 3206 37800
rect 3418 37788 3424 37800
rect 3200 37760 3424 37788
rect 3200 37748 3206 37760
rect 3418 37748 3424 37760
rect 3476 37748 3482 37800
rect 3513 37791 3571 37797
rect 3513 37757 3525 37791
rect 3559 37757 3571 37791
rect 3513 37751 3571 37757
rect 1854 37720 1860 37732
rect 1412 37692 1860 37720
rect 1854 37680 1860 37692
rect 1912 37680 1918 37732
rect 2041 37723 2099 37729
rect 2041 37689 2053 37723
rect 2087 37720 2099 37723
rect 2130 37720 2136 37732
rect 2087 37692 2136 37720
rect 2087 37689 2099 37692
rect 2041 37683 2099 37689
rect 2130 37680 2136 37692
rect 2188 37680 2194 37732
rect 3528 37720 3556 37751
rect 4154 37748 4160 37800
rect 4212 37748 4218 37800
rect 4522 37748 4528 37800
rect 4580 37788 4586 37800
rect 4617 37791 4675 37797
rect 4617 37788 4629 37791
rect 4580 37760 4629 37788
rect 4580 37748 4586 37760
rect 4617 37757 4629 37760
rect 4663 37757 4675 37791
rect 7392 37788 7420 37819
rect 7558 37816 7564 37868
rect 7616 37816 7622 37868
rect 9214 37816 9220 37868
rect 9272 37816 9278 37868
rect 9508 37856 9536 37896
rect 9582 37884 9588 37936
rect 9640 37884 9646 37936
rect 9766 37884 9772 37936
rect 9824 37924 9830 37936
rect 15194 37924 15200 37936
rect 9824 37896 15200 37924
rect 9824 37884 9830 37896
rect 15194 37884 15200 37896
rect 15252 37924 15258 37936
rect 15252 37896 18368 37924
rect 15252 37884 15258 37896
rect 9674 37856 9680 37868
rect 9508 37828 9680 37856
rect 9674 37816 9680 37828
rect 9732 37816 9738 37868
rect 12434 37816 12440 37868
rect 12492 37856 12498 37868
rect 18340 37865 18368 37896
rect 22646 37884 22652 37936
rect 22704 37924 22710 37936
rect 22833 37927 22891 37933
rect 22833 37924 22845 37927
rect 22704 37896 22845 37924
rect 22704 37884 22710 37896
rect 22833 37893 22845 37896
rect 22879 37893 22891 37927
rect 22833 37887 22891 37893
rect 12955 37859 13013 37865
rect 12955 37856 12967 37859
rect 12492 37828 12967 37856
rect 12492 37816 12498 37828
rect 8484 37800 8536 37806
rect 7650 37788 7656 37800
rect 7392 37760 7656 37788
rect 4617 37751 4675 37757
rect 2976 37692 3556 37720
rect 2498 37612 2504 37664
rect 2556 37652 2562 37664
rect 2976 37652 3004 37692
rect 2556 37624 3004 37652
rect 2556 37612 2562 37624
rect 3142 37612 3148 37664
rect 3200 37652 3206 37664
rect 3237 37655 3295 37661
rect 3237 37652 3249 37655
rect 3200 37624 3249 37652
rect 3200 37612 3206 37624
rect 3237 37621 3249 37624
rect 3283 37621 3295 37655
rect 3528 37652 3556 37692
rect 4430 37652 4436 37664
rect 3528 37624 4436 37652
rect 3237 37615 3295 37621
rect 4430 37612 4436 37624
rect 4488 37612 4494 37664
rect 4632 37652 4660 37751
rect 7650 37748 7656 37760
rect 7708 37748 7714 37800
rect 8484 37742 8536 37748
rect 5810 37720 5816 37732
rect 5552 37692 5816 37720
rect 5552 37652 5580 37692
rect 5810 37680 5816 37692
rect 5868 37720 5874 37732
rect 6454 37720 6460 37732
rect 5868 37692 6460 37720
rect 5868 37680 5874 37692
rect 6454 37680 6460 37692
rect 6512 37680 6518 37732
rect 6638 37680 6644 37732
rect 6696 37720 6702 37732
rect 7926 37720 7932 37732
rect 6696 37692 7932 37720
rect 6696 37680 6702 37692
rect 7926 37680 7932 37692
rect 7984 37680 7990 37732
rect 12636 37720 12664 37828
rect 12955 37825 12967 37828
rect 13001 37825 13013 37859
rect 12955 37819 13013 37825
rect 18325 37859 18383 37865
rect 18325 37825 18337 37859
rect 18371 37825 18383 37859
rect 18325 37819 18383 37825
rect 21082 37816 21088 37868
rect 21140 37816 21146 37868
rect 22097 37859 22155 37865
rect 22097 37825 22109 37859
rect 22143 37825 22155 37859
rect 22097 37819 22155 37825
rect 12710 37748 12716 37800
rect 12768 37748 12774 37800
rect 15654 37748 15660 37800
rect 15712 37788 15718 37800
rect 20254 37788 20260 37800
rect 15712 37760 20260 37788
rect 15712 37748 15718 37760
rect 20254 37748 20260 37760
rect 20312 37748 20318 37800
rect 20530 37748 20536 37800
rect 20588 37788 20594 37800
rect 22112 37788 22140 37819
rect 22186 37816 22192 37868
rect 22244 37856 22250 37868
rect 22465 37859 22523 37865
rect 22465 37856 22477 37859
rect 22244 37828 22477 37856
rect 22244 37816 22250 37828
rect 22465 37825 22477 37828
rect 22511 37825 22523 37859
rect 22465 37819 22523 37825
rect 23014 37816 23020 37868
rect 23072 37856 23078 37868
rect 23109 37859 23167 37865
rect 23109 37856 23121 37859
rect 23072 37828 23121 37856
rect 23072 37816 23078 37828
rect 23109 37825 23121 37828
rect 23155 37825 23167 37859
rect 23109 37819 23167 37825
rect 23290 37816 23296 37868
rect 23348 37856 23354 37868
rect 23569 37859 23627 37865
rect 23569 37856 23581 37859
rect 23348 37828 23581 37856
rect 23348 37816 23354 37828
rect 23569 37825 23581 37828
rect 23615 37825 23627 37859
rect 23569 37819 23627 37825
rect 23842 37816 23848 37868
rect 23900 37816 23906 37868
rect 24121 37859 24179 37865
rect 24121 37825 24133 37859
rect 24167 37825 24179 37859
rect 24121 37819 24179 37825
rect 20588 37760 22140 37788
rect 20588 37748 20594 37760
rect 22278 37748 22284 37800
rect 22336 37748 22342 37800
rect 24136 37788 24164 37819
rect 22480 37760 24164 37788
rect 12636 37692 12756 37720
rect 12728 37664 12756 37692
rect 20898 37680 20904 37732
rect 20956 37720 20962 37732
rect 22480 37720 22508 37760
rect 20956 37692 22508 37720
rect 20956 37680 20962 37692
rect 22554 37680 22560 37732
rect 22612 37720 22618 37732
rect 22925 37723 22983 37729
rect 22925 37720 22937 37723
rect 22612 37692 22937 37720
rect 22612 37680 22618 37692
rect 22925 37689 22937 37692
rect 22971 37689 22983 37723
rect 22925 37683 22983 37689
rect 4632 37624 5580 37652
rect 5626 37612 5632 37664
rect 5684 37612 5690 37664
rect 7469 37655 7527 37661
rect 7469 37621 7481 37655
rect 7515 37652 7527 37655
rect 8202 37652 8208 37664
rect 7515 37624 8208 37652
rect 7515 37621 7527 37624
rect 7469 37615 7527 37621
rect 8202 37612 8208 37624
rect 8260 37612 8266 37664
rect 9769 37655 9827 37661
rect 9769 37621 9781 37655
rect 9815 37652 9827 37655
rect 11054 37652 11060 37664
rect 9815 37624 11060 37652
rect 9815 37621 9827 37624
rect 9769 37615 9827 37621
rect 11054 37612 11060 37624
rect 11112 37612 11118 37664
rect 12710 37612 12716 37664
rect 12768 37612 12774 37664
rect 22741 37655 22799 37661
rect 22741 37621 22753 37655
rect 22787 37652 22799 37655
rect 23382 37652 23388 37664
rect 22787 37624 23388 37652
rect 22787 37621 22799 37624
rect 22741 37615 22799 37621
rect 23382 37612 23388 37624
rect 23440 37612 23446 37664
rect 23661 37655 23719 37661
rect 23661 37621 23673 37655
rect 23707 37652 23719 37655
rect 24026 37652 24032 37664
rect 23707 37624 24032 37652
rect 23707 37621 23719 37624
rect 23661 37615 23719 37621
rect 24026 37612 24032 37624
rect 24084 37612 24090 37664
rect 24394 37612 24400 37664
rect 24452 37612 24458 37664
rect 1104 37562 24840 37584
rect 1104 37510 3917 37562
rect 3969 37510 3981 37562
rect 4033 37510 4045 37562
rect 4097 37510 4109 37562
rect 4161 37510 4173 37562
rect 4225 37510 9851 37562
rect 9903 37510 9915 37562
rect 9967 37510 9979 37562
rect 10031 37510 10043 37562
rect 10095 37510 10107 37562
rect 10159 37510 15785 37562
rect 15837 37510 15849 37562
rect 15901 37510 15913 37562
rect 15965 37510 15977 37562
rect 16029 37510 16041 37562
rect 16093 37510 21719 37562
rect 21771 37510 21783 37562
rect 21835 37510 21847 37562
rect 21899 37510 21911 37562
rect 21963 37510 21975 37562
rect 22027 37510 24840 37562
rect 1104 37488 24840 37510
rect 1762 37408 1768 37460
rect 1820 37448 1826 37460
rect 1820 37420 2084 37448
rect 1820 37408 1826 37420
rect 2056 37380 2084 37420
rect 2130 37408 2136 37460
rect 2188 37448 2194 37460
rect 2409 37451 2467 37457
rect 2409 37448 2421 37451
rect 2188 37420 2421 37448
rect 2188 37408 2194 37420
rect 2409 37417 2421 37420
rect 2455 37417 2467 37451
rect 7561 37451 7619 37457
rect 2409 37411 2467 37417
rect 5000 37420 7512 37448
rect 5000 37392 5028 37420
rect 7484 37392 7512 37420
rect 7561 37417 7573 37451
rect 7607 37448 7619 37451
rect 7650 37448 7656 37460
rect 7607 37420 7656 37448
rect 7607 37417 7619 37420
rect 7561 37411 7619 37417
rect 7650 37408 7656 37420
rect 7708 37408 7714 37460
rect 8128 37420 9628 37448
rect 4338 37380 4344 37392
rect 2056 37352 4344 37380
rect 4338 37340 4344 37352
rect 4396 37340 4402 37392
rect 4982 37340 4988 37392
rect 5040 37340 5046 37392
rect 7466 37340 7472 37392
rect 7524 37380 7530 37392
rect 8128 37380 8156 37420
rect 7524 37352 8156 37380
rect 9600 37380 9628 37420
rect 9674 37408 9680 37460
rect 9732 37448 9738 37460
rect 9953 37451 10011 37457
rect 9953 37448 9965 37451
rect 9732 37420 9965 37448
rect 9732 37408 9738 37420
rect 9953 37417 9965 37420
rect 9999 37417 10011 37451
rect 19610 37448 19616 37460
rect 9953 37411 10011 37417
rect 12406 37420 19616 37448
rect 12406 37380 12434 37420
rect 19610 37408 19616 37420
rect 19668 37408 19674 37460
rect 22462 37408 22468 37460
rect 22520 37408 22526 37460
rect 23109 37451 23167 37457
rect 23109 37417 23121 37451
rect 23155 37448 23167 37451
rect 23290 37448 23296 37460
rect 23155 37420 23296 37448
rect 23155 37417 23167 37420
rect 23109 37411 23167 37417
rect 23290 37408 23296 37420
rect 23348 37408 23354 37460
rect 23661 37451 23719 37457
rect 23661 37417 23673 37451
rect 23707 37448 23719 37451
rect 23842 37448 23848 37460
rect 23707 37420 23848 37448
rect 23707 37417 23719 37420
rect 23661 37411 23719 37417
rect 23842 37408 23848 37420
rect 23900 37408 23906 37460
rect 9600 37352 12434 37380
rect 7524 37340 7530 37352
rect 19150 37340 19156 37392
rect 19208 37380 19214 37392
rect 23750 37380 23756 37392
rect 19208 37352 23756 37380
rect 19208 37340 19214 37352
rect 23750 37340 23756 37352
rect 23808 37340 23814 37392
rect 3510 37312 3516 37324
rect 2884 37284 3516 37312
rect 1397 37247 1455 37253
rect 1397 37213 1409 37247
rect 1443 37213 1455 37247
rect 1397 37207 1455 37213
rect 1671 37247 1729 37253
rect 1671 37213 1683 37247
rect 1717 37244 1729 37247
rect 2130 37244 2136 37256
rect 1717 37216 2136 37244
rect 1717 37213 1729 37216
rect 1671 37207 1729 37213
rect 1412 37176 1440 37207
rect 2130 37204 2136 37216
rect 2188 37204 2194 37256
rect 2774 37204 2780 37256
rect 2832 37204 2838 37256
rect 2884 37176 2912 37284
rect 3510 37272 3516 37284
rect 3568 37272 3574 37324
rect 4522 37272 4528 37324
rect 4580 37312 4586 37324
rect 5077 37315 5135 37321
rect 5077 37312 5089 37315
rect 4580 37284 5089 37312
rect 4580 37272 4586 37284
rect 5077 37281 5089 37284
rect 5123 37281 5135 37315
rect 5077 37275 5135 37281
rect 6454 37272 6460 37324
rect 6512 37312 6518 37324
rect 6512 37284 6592 37312
rect 6512 37272 6518 37284
rect 3789 37247 3847 37253
rect 3789 37244 3801 37247
rect 1412 37148 2912 37176
rect 2976 37216 3801 37244
rect 1302 37068 1308 37120
rect 1360 37108 1366 37120
rect 2976 37108 3004 37216
rect 3789 37213 3801 37216
rect 3835 37213 3847 37247
rect 3789 37207 3847 37213
rect 3878 37204 3884 37256
rect 3936 37244 3942 37256
rect 6564 37253 6592 37284
rect 8202 37272 8208 37324
rect 8260 37272 8266 37324
rect 13814 37272 13820 37324
rect 13872 37312 13878 37324
rect 19334 37312 19340 37324
rect 13872 37284 19340 37312
rect 13872 37272 13878 37284
rect 19334 37272 19340 37284
rect 19392 37272 19398 37324
rect 23290 37312 23296 37324
rect 21836 37284 23296 37312
rect 4341 37247 4399 37253
rect 4341 37244 4353 37247
rect 3936 37216 4353 37244
rect 3936 37204 3942 37216
rect 4341 37213 4353 37216
rect 4387 37213 4399 37247
rect 4341 37207 4399 37213
rect 5351 37247 5409 37253
rect 5351 37213 5363 37247
rect 5397 37244 5409 37247
rect 6549 37247 6607 37253
rect 5397 37216 6500 37244
rect 5397 37213 5409 37216
rect 5351 37207 5409 37213
rect 3053 37179 3111 37185
rect 3053 37145 3065 37179
rect 3099 37145 3111 37179
rect 3053 37139 3111 37145
rect 4065 37179 4123 37185
rect 4065 37145 4077 37179
rect 4111 37176 4123 37179
rect 4522 37176 4528 37188
rect 4111 37148 4528 37176
rect 4111 37145 4123 37148
rect 4065 37139 4123 37145
rect 1360 37080 3004 37108
rect 3068 37108 3096 37139
rect 4522 37136 4528 37148
rect 4580 37136 4586 37188
rect 4617 37179 4675 37185
rect 4617 37145 4629 37179
rect 4663 37176 4675 37179
rect 5166 37176 5172 37188
rect 4663 37148 5172 37176
rect 4663 37145 4675 37148
rect 4617 37139 4675 37145
rect 5166 37136 5172 37148
rect 5224 37136 5230 37188
rect 6472 37176 6500 37216
rect 6549 37213 6561 37247
rect 6595 37213 6607 37247
rect 6549 37207 6607 37213
rect 6823 37237 6881 37243
rect 6823 37203 6835 37237
rect 6869 37203 6881 37237
rect 7650 37204 7656 37256
rect 7708 37244 7714 37256
rect 7929 37247 7987 37253
rect 7929 37244 7941 37247
rect 7708 37216 7941 37244
rect 7708 37204 7714 37216
rect 7929 37213 7941 37216
rect 7975 37213 7987 37247
rect 7929 37207 7987 37213
rect 8018 37204 8024 37256
rect 8076 37204 8082 37256
rect 8110 37204 8116 37256
rect 8168 37204 8174 37256
rect 8941 37247 8999 37253
rect 8941 37213 8953 37247
rect 8987 37244 8999 37247
rect 9122 37244 9128 37256
rect 8987 37216 9128 37244
rect 8987 37213 8999 37216
rect 8941 37207 8999 37213
rect 6823 37197 6881 37203
rect 6638 37176 6644 37188
rect 6472 37148 6644 37176
rect 6638 37136 6644 37148
rect 6696 37136 6702 37188
rect 5258 37108 5264 37120
rect 3068 37080 5264 37108
rect 1360 37068 1366 37080
rect 5258 37068 5264 37080
rect 5316 37068 5322 37120
rect 6089 37111 6147 37117
rect 6089 37077 6101 37111
rect 6135 37108 6147 37111
rect 6178 37108 6184 37120
rect 6135 37080 6184 37108
rect 6135 37077 6147 37080
rect 6089 37071 6147 37077
rect 6178 37068 6184 37080
rect 6236 37068 6242 37120
rect 6730 37068 6736 37120
rect 6788 37108 6794 37120
rect 6840 37108 6868 37197
rect 8128 37176 8156 37204
rect 8205 37179 8263 37185
rect 8205 37176 8217 37179
rect 8128 37148 8217 37176
rect 8205 37145 8217 37148
rect 8251 37145 8263 37179
rect 8956 37176 8984 37207
rect 9122 37204 9128 37216
rect 9180 37204 9186 37256
rect 9215 37237 9273 37243
rect 9215 37203 9227 37237
rect 9261 37234 9273 37237
rect 9306 37234 9312 37256
rect 9261 37206 9312 37234
rect 9261 37203 9273 37206
rect 9306 37204 9312 37206
rect 9364 37204 9370 37256
rect 12618 37244 12624 37256
rect 9416 37216 12624 37244
rect 9215 37197 9273 37203
rect 9416 37188 9444 37216
rect 12618 37204 12624 37216
rect 12676 37244 12682 37256
rect 16482 37244 16488 37256
rect 12676 37216 16488 37244
rect 12676 37204 12682 37216
rect 16482 37204 16488 37216
rect 16540 37204 16546 37256
rect 19426 37204 19432 37256
rect 19484 37204 19490 37256
rect 19981 37247 20039 37253
rect 19981 37213 19993 37247
rect 20027 37213 20039 37247
rect 19981 37207 20039 37213
rect 8205 37139 8263 37145
rect 8312 37148 8984 37176
rect 6788 37080 6868 37108
rect 6788 37068 6794 37080
rect 7282 37068 7288 37120
rect 7340 37108 7346 37120
rect 7742 37108 7748 37120
rect 7340 37080 7748 37108
rect 7340 37068 7346 37080
rect 7742 37068 7748 37080
rect 7800 37108 7806 37120
rect 8312 37108 8340 37148
rect 9398 37136 9404 37188
rect 9456 37136 9462 37188
rect 19996 37176 20024 37207
rect 20346 37204 20352 37256
rect 20404 37204 20410 37256
rect 20898 37204 20904 37256
rect 20956 37204 20962 37256
rect 21082 37204 21088 37256
rect 21140 37204 21146 37256
rect 21450 37204 21456 37256
rect 21508 37244 21514 37256
rect 21836 37244 21864 37284
rect 23290 37272 23296 37284
rect 23348 37272 23354 37324
rect 21508 37216 21864 37244
rect 21913 37247 21971 37253
rect 21508 37204 21514 37216
rect 21913 37213 21925 37247
rect 21959 37213 21971 37247
rect 22649 37247 22707 37253
rect 22649 37244 22661 37247
rect 21913 37207 21971 37213
rect 22066 37216 22661 37244
rect 20916 37176 20944 37204
rect 9646 37148 11652 37176
rect 7800 37080 8340 37108
rect 7800 37068 7806 37080
rect 8386 37068 8392 37120
rect 8444 37108 8450 37120
rect 9306 37108 9312 37120
rect 8444 37080 9312 37108
rect 8444 37068 8450 37080
rect 9306 37068 9312 37080
rect 9364 37108 9370 37120
rect 9646 37108 9674 37148
rect 11624 37120 11652 37148
rect 19260 37148 20024 37176
rect 20088 37148 20944 37176
rect 9364 37080 9674 37108
rect 9364 37068 9370 37080
rect 11606 37068 11612 37120
rect 11664 37108 11670 37120
rect 13630 37108 13636 37120
rect 11664 37080 13636 37108
rect 11664 37068 11670 37080
rect 13630 37068 13636 37080
rect 13688 37068 13694 37120
rect 19260 37117 19288 37148
rect 19245 37111 19303 37117
rect 19245 37077 19257 37111
rect 19291 37077 19303 37111
rect 19245 37071 19303 37077
rect 19797 37111 19855 37117
rect 19797 37077 19809 37111
rect 19843 37108 19855 37111
rect 20088 37108 20116 37148
rect 19843 37080 20116 37108
rect 20165 37111 20223 37117
rect 19843 37077 19855 37080
rect 19797 37071 19855 37077
rect 20165 37077 20177 37111
rect 20211 37108 20223 37111
rect 21100 37108 21128 37204
rect 21928 37176 21956 37207
rect 21284 37148 21956 37176
rect 21284 37120 21312 37148
rect 20211 37080 21128 37108
rect 20211 37077 20223 37080
rect 20165 37071 20223 37077
rect 21266 37068 21272 37120
rect 21324 37068 21330 37120
rect 21729 37111 21787 37117
rect 21729 37077 21741 37111
rect 21775 37108 21787 37111
rect 22066 37108 22094 37216
rect 22649 37213 22661 37216
rect 22695 37213 22707 37247
rect 22649 37207 22707 37213
rect 23385 37247 23443 37253
rect 23385 37213 23397 37247
rect 23431 37244 23443 37247
rect 23474 37244 23480 37256
rect 23431 37216 23480 37244
rect 23431 37213 23443 37216
rect 23385 37207 23443 37213
rect 23474 37204 23480 37216
rect 23532 37204 23538 37256
rect 23658 37204 23664 37256
rect 23716 37204 23722 37256
rect 23842 37204 23848 37256
rect 23900 37204 23906 37256
rect 23934 37204 23940 37256
rect 23992 37204 23998 37256
rect 21775 37080 22094 37108
rect 23201 37111 23259 37117
rect 21775 37077 21787 37080
rect 21729 37071 21787 37077
rect 23201 37077 23213 37111
rect 23247 37108 23259 37111
rect 23676 37108 23704 37204
rect 23247 37080 23704 37108
rect 23247 37077 23259 37080
rect 23201 37071 23259 37077
rect 24118 37068 24124 37120
rect 24176 37068 24182 37120
rect 1104 37018 25000 37040
rect 1104 36966 6884 37018
rect 6936 36966 6948 37018
rect 7000 36966 7012 37018
rect 7064 36966 7076 37018
rect 7128 36966 7140 37018
rect 7192 36966 12818 37018
rect 12870 36966 12882 37018
rect 12934 36966 12946 37018
rect 12998 36966 13010 37018
rect 13062 36966 13074 37018
rect 13126 36966 18752 37018
rect 18804 36966 18816 37018
rect 18868 36966 18880 37018
rect 18932 36966 18944 37018
rect 18996 36966 19008 37018
rect 19060 36966 24686 37018
rect 24738 36966 24750 37018
rect 24802 36966 24814 37018
rect 24866 36966 24878 37018
rect 24930 36966 24942 37018
rect 24994 36966 25000 37018
rect 1104 36944 25000 36966
rect 3145 36907 3203 36913
rect 3145 36873 3157 36907
rect 3191 36904 3203 36907
rect 3418 36904 3424 36916
rect 3191 36876 3424 36904
rect 3191 36873 3203 36876
rect 3145 36867 3203 36873
rect 3418 36864 3424 36876
rect 3476 36864 3482 36916
rect 5629 36907 5687 36913
rect 5629 36904 5641 36907
rect 3528 36876 5641 36904
rect 3528 36845 3556 36876
rect 5629 36873 5641 36876
rect 5675 36873 5687 36907
rect 5629 36867 5687 36873
rect 5718 36864 5724 36916
rect 5776 36904 5782 36916
rect 7190 36904 7196 36916
rect 5776 36876 7196 36904
rect 5776 36864 5782 36876
rect 7190 36864 7196 36876
rect 7248 36864 7254 36916
rect 7469 36907 7527 36913
rect 7469 36873 7481 36907
rect 7515 36904 7527 36907
rect 7558 36904 7564 36916
rect 7515 36876 7564 36904
rect 7515 36873 7527 36876
rect 7469 36867 7527 36873
rect 7558 36864 7564 36876
rect 7616 36864 7622 36916
rect 8018 36864 8024 36916
rect 8076 36864 8082 36916
rect 9122 36864 9128 36916
rect 9180 36904 9186 36916
rect 9398 36904 9404 36916
rect 9180 36876 9404 36904
rect 9180 36864 9186 36876
rect 9398 36864 9404 36876
rect 9456 36864 9462 36916
rect 10134 36904 10140 36916
rect 9646 36876 10140 36904
rect 3513 36839 3571 36845
rect 3513 36805 3525 36839
rect 3559 36805 3571 36839
rect 3513 36799 3571 36805
rect 3602 36796 3608 36848
rect 3660 36836 3666 36848
rect 4154 36836 4160 36848
rect 3660 36808 4160 36836
rect 3660 36796 3666 36808
rect 4154 36796 4160 36808
rect 4212 36796 4218 36848
rect 4249 36839 4307 36845
rect 4249 36805 4261 36839
rect 4295 36836 4307 36839
rect 4338 36836 4344 36848
rect 4295 36808 4344 36836
rect 4295 36805 4307 36808
rect 4249 36799 4307 36805
rect 4338 36796 4344 36808
rect 4396 36836 4402 36848
rect 4982 36836 4988 36848
rect 4396 36808 4988 36836
rect 4396 36796 4402 36808
rect 4982 36796 4988 36808
rect 5040 36796 5046 36848
rect 5166 36796 5172 36848
rect 5224 36836 5230 36848
rect 5442 36836 5448 36848
rect 5224 36808 5448 36836
rect 5224 36796 5230 36808
rect 5442 36796 5448 36808
rect 5500 36836 5506 36848
rect 7285 36839 7343 36845
rect 5500 36808 5948 36836
rect 5500 36796 5506 36808
rect 1210 36728 1216 36780
rect 1268 36768 1274 36780
rect 1397 36771 1455 36777
rect 1397 36768 1409 36771
rect 1268 36740 1409 36768
rect 1268 36728 1274 36740
rect 1397 36737 1409 36740
rect 1443 36737 1455 36771
rect 1397 36731 1455 36737
rect 1949 36771 2007 36777
rect 1949 36737 1961 36771
rect 1995 36768 2007 36771
rect 2866 36768 2872 36780
rect 1995 36740 2872 36768
rect 1995 36737 2007 36740
rect 1949 36731 2007 36737
rect 2866 36728 2872 36740
rect 2924 36728 2930 36780
rect 3421 36771 3479 36777
rect 3421 36737 3433 36771
rect 3467 36768 3479 36771
rect 3620 36768 3648 36796
rect 3467 36740 3648 36768
rect 3467 36737 3479 36740
rect 3421 36731 3479 36737
rect 3786 36728 3792 36780
rect 3844 36768 3850 36780
rect 3881 36771 3939 36777
rect 3881 36768 3893 36771
rect 3844 36740 3893 36768
rect 3844 36728 3850 36740
rect 3881 36737 3893 36740
rect 3927 36737 3939 36771
rect 3881 36731 3939 36737
rect 4430 36728 4436 36780
rect 4488 36768 4494 36780
rect 4891 36771 4949 36777
rect 4891 36768 4903 36771
rect 4488 36740 4903 36768
rect 4488 36728 4494 36740
rect 4891 36737 4903 36740
rect 4937 36768 4949 36771
rect 4937 36740 5854 36768
rect 4937 36737 4949 36740
rect 4891 36731 4949 36737
rect 14 36660 20 36712
rect 72 36660 78 36712
rect 1673 36703 1731 36709
rect 1673 36669 1685 36703
rect 1719 36700 1731 36703
rect 1762 36700 1768 36712
rect 1719 36672 1768 36700
rect 1719 36669 1731 36672
rect 1673 36663 1731 36669
rect 1762 36660 1768 36672
rect 1820 36660 1826 36712
rect 2133 36703 2191 36709
rect 2133 36669 2145 36703
rect 2179 36669 2191 36703
rect 2133 36663 2191 36669
rect 32 36632 60 36660
rect 2148 36632 2176 36663
rect 2314 36660 2320 36712
rect 2372 36660 2378 36712
rect 3326 36660 3332 36712
rect 3384 36660 3390 36712
rect 4617 36703 4675 36709
rect 4617 36669 4629 36703
rect 4663 36669 4675 36703
rect 5718 36700 5724 36712
rect 4617 36663 4675 36669
rect 5276 36672 5724 36700
rect 32 36604 2176 36632
rect 2332 36632 2360 36660
rect 2685 36635 2743 36641
rect 2685 36632 2697 36635
rect 2332 36604 2697 36632
rect 2685 36601 2697 36604
rect 2731 36601 2743 36635
rect 2685 36595 2743 36601
rect 4338 36592 4344 36644
rect 4396 36632 4402 36644
rect 4632 36632 4660 36663
rect 4396 36604 4660 36632
rect 4396 36592 4402 36604
rect 4430 36524 4436 36576
rect 4488 36524 4494 36576
rect 4632 36564 4660 36604
rect 5276 36564 5304 36672
rect 5718 36660 5724 36672
rect 5776 36660 5782 36712
rect 4632 36536 5304 36564
rect 5826 36564 5854 36740
rect 5920 36700 5948 36808
rect 7285 36805 7297 36839
rect 7331 36836 7343 36839
rect 8036 36836 8064 36864
rect 9646 36836 9674 36876
rect 10134 36864 10140 36876
rect 10192 36904 10198 36916
rect 18601 36907 18659 36913
rect 10192 36876 10916 36904
rect 10192 36864 10198 36876
rect 10888 36836 10916 36876
rect 18601 36873 18613 36907
rect 18647 36904 18659 36907
rect 19426 36904 19432 36916
rect 18647 36876 19432 36904
rect 18647 36873 18659 36876
rect 18601 36867 18659 36873
rect 19426 36864 19432 36876
rect 19484 36864 19490 36916
rect 19521 36907 19579 36913
rect 19521 36873 19533 36907
rect 19567 36904 19579 36907
rect 20346 36904 20352 36916
rect 19567 36876 20352 36904
rect 19567 36873 19579 36876
rect 19521 36867 19579 36873
rect 20346 36864 20352 36876
rect 20404 36864 20410 36916
rect 22373 36907 22431 36913
rect 22373 36873 22385 36907
rect 22419 36873 22431 36907
rect 22373 36867 22431 36873
rect 23385 36907 23443 36913
rect 23385 36873 23397 36907
rect 23431 36904 23443 36907
rect 23566 36904 23572 36916
rect 23431 36876 23572 36904
rect 23431 36873 23443 36876
rect 23385 36867 23443 36873
rect 22388 36836 22416 36867
rect 23566 36864 23572 36876
rect 23624 36864 23630 36916
rect 23661 36907 23719 36913
rect 23661 36873 23673 36907
rect 23707 36904 23719 36907
rect 23934 36904 23940 36916
rect 23707 36876 23940 36904
rect 23707 36873 23719 36876
rect 23661 36867 23719 36873
rect 23934 36864 23940 36876
rect 23992 36864 23998 36916
rect 7331 36808 8064 36836
rect 8128 36808 9674 36836
rect 9876 36808 10824 36836
rect 10888 36808 19748 36836
rect 22388 36808 23888 36836
rect 7331 36805 7343 36808
rect 7285 36799 7343 36805
rect 7190 36728 7196 36780
rect 7248 36728 7254 36780
rect 7650 36728 7656 36780
rect 7708 36728 7714 36780
rect 7558 36700 7564 36712
rect 5920 36672 7564 36700
rect 7558 36660 7564 36672
rect 7616 36700 7622 36712
rect 8128 36700 8156 36808
rect 9876 36777 9904 36808
rect 9861 36771 9919 36777
rect 9861 36737 9873 36771
rect 9907 36737 9919 36771
rect 10134 36768 10140 36780
rect 10095 36740 10140 36768
rect 9861 36731 9919 36737
rect 10134 36728 10140 36740
rect 10192 36728 10198 36780
rect 10796 36712 10824 36808
rect 19720 36777 19748 36808
rect 18785 36771 18843 36777
rect 18785 36768 18797 36771
rect 18156 36740 18797 36768
rect 7616 36672 8156 36700
rect 7616 36660 7622 36672
rect 10778 36660 10784 36712
rect 10836 36660 10842 36712
rect 18156 36644 18184 36740
rect 18785 36737 18797 36740
rect 18831 36737 18843 36771
rect 18785 36731 18843 36737
rect 19705 36771 19763 36777
rect 19705 36737 19717 36771
rect 19751 36737 19763 36771
rect 19705 36731 19763 36737
rect 22278 36728 22284 36780
rect 22336 36768 22342 36780
rect 23860 36777 23888 36808
rect 24026 36796 24032 36848
rect 24084 36836 24090 36848
rect 24121 36839 24179 36845
rect 24121 36836 24133 36839
rect 24084 36808 24133 36836
rect 24084 36796 24090 36808
rect 24121 36805 24133 36808
rect 24167 36805 24179 36839
rect 24121 36799 24179 36805
rect 22557 36771 22615 36777
rect 22557 36768 22569 36771
rect 22336 36740 22569 36768
rect 22336 36728 22342 36740
rect 22557 36737 22569 36740
rect 22603 36737 22615 36771
rect 23569 36771 23627 36777
rect 23569 36768 23581 36771
rect 22557 36731 22615 36737
rect 23032 36740 23581 36768
rect 10796 36604 13492 36632
rect 10796 36564 10824 36604
rect 13464 36576 13492 36604
rect 16758 36592 16764 36644
rect 16816 36632 16822 36644
rect 17770 36632 17776 36644
rect 16816 36604 17776 36632
rect 16816 36592 16822 36604
rect 17770 36592 17776 36604
rect 17828 36592 17834 36644
rect 18138 36592 18144 36644
rect 18196 36592 18202 36644
rect 23032 36576 23060 36740
rect 23569 36737 23581 36740
rect 23615 36737 23627 36771
rect 23569 36731 23627 36737
rect 23845 36771 23903 36777
rect 23845 36737 23857 36771
rect 23891 36737 23903 36771
rect 23845 36731 23903 36737
rect 5826 36536 10824 36564
rect 10870 36524 10876 36576
rect 10928 36524 10934 36576
rect 12066 36524 12072 36576
rect 12124 36564 12130 36576
rect 12526 36564 12532 36576
rect 12124 36536 12532 36564
rect 12124 36524 12130 36536
rect 12526 36524 12532 36536
rect 12584 36524 12590 36576
rect 13446 36524 13452 36576
rect 13504 36524 13510 36576
rect 13722 36524 13728 36576
rect 13780 36564 13786 36576
rect 22922 36564 22928 36576
rect 13780 36536 22928 36564
rect 13780 36524 13786 36536
rect 22922 36524 22928 36536
rect 22980 36524 22986 36576
rect 23014 36524 23020 36576
rect 23072 36524 23078 36576
rect 24394 36524 24400 36576
rect 24452 36524 24458 36576
rect 1104 36474 24840 36496
rect 1104 36422 3917 36474
rect 3969 36422 3981 36474
rect 4033 36422 4045 36474
rect 4097 36422 4109 36474
rect 4161 36422 4173 36474
rect 4225 36422 9851 36474
rect 9903 36422 9915 36474
rect 9967 36422 9979 36474
rect 10031 36422 10043 36474
rect 10095 36422 10107 36474
rect 10159 36422 15785 36474
rect 15837 36422 15849 36474
rect 15901 36422 15913 36474
rect 15965 36422 15977 36474
rect 16029 36422 16041 36474
rect 16093 36422 21719 36474
rect 21771 36422 21783 36474
rect 21835 36422 21847 36474
rect 21899 36422 21911 36474
rect 21963 36422 21975 36474
rect 22027 36422 24840 36474
rect 1104 36400 24840 36422
rect 2424 36332 3096 36360
rect 2424 36292 2452 36332
rect 2332 36264 2452 36292
rect 2332 36233 2360 36264
rect 2317 36227 2375 36233
rect 2317 36193 2329 36227
rect 2363 36193 2375 36227
rect 2317 36187 2375 36193
rect 3068 36224 3096 36332
rect 3326 36320 3332 36372
rect 3384 36320 3390 36372
rect 4338 36320 4344 36372
rect 4396 36320 4402 36372
rect 6917 36363 6975 36369
rect 6917 36329 6929 36363
rect 6963 36360 6975 36363
rect 7190 36360 7196 36372
rect 6963 36332 7196 36360
rect 6963 36329 6975 36332
rect 6917 36323 6975 36329
rect 7190 36320 7196 36332
rect 7248 36320 7254 36372
rect 7650 36320 7656 36372
rect 7708 36320 7714 36372
rect 8110 36320 8116 36372
rect 8168 36360 8174 36372
rect 8168 36332 10180 36360
rect 8168 36320 8174 36332
rect 4356 36224 4384 36320
rect 4430 36252 4436 36304
rect 4488 36252 4494 36304
rect 4614 36252 4620 36304
rect 4672 36292 4678 36304
rect 4672 36264 5304 36292
rect 4672 36252 4678 36264
rect 3068 36196 4384 36224
rect 4448 36224 4476 36252
rect 5169 36227 5227 36233
rect 5169 36224 5181 36227
rect 4448 36196 5181 36224
rect 3068 36168 3096 36196
rect 5169 36193 5181 36196
rect 5215 36193 5227 36227
rect 5276 36224 5304 36264
rect 5626 36252 5632 36304
rect 5684 36252 5690 36304
rect 6825 36295 6883 36301
rect 6825 36261 6837 36295
rect 6871 36292 6883 36295
rect 7668 36292 7696 36320
rect 6871 36264 7696 36292
rect 6871 36261 6883 36264
rect 6825 36255 6883 36261
rect 5718 36224 5724 36236
rect 5276 36196 5724 36224
rect 5169 36187 5227 36193
rect 5718 36184 5724 36196
rect 5776 36224 5782 36236
rect 6022 36227 6080 36233
rect 6022 36224 6034 36227
rect 5776 36196 6034 36224
rect 5776 36184 5782 36196
rect 6022 36193 6034 36196
rect 6068 36193 6080 36227
rect 6022 36187 6080 36193
rect 6178 36184 6184 36236
rect 6236 36184 6242 36236
rect 1394 36116 1400 36168
rect 1452 36116 1458 36168
rect 2559 36159 2617 36165
rect 2559 36156 2571 36159
rect 1596 36128 2571 36156
rect 1118 35980 1124 36032
rect 1176 36020 1182 36032
rect 1596 36020 1624 36128
rect 2559 36125 2571 36128
rect 2605 36156 2617 36159
rect 2682 36156 2688 36168
rect 2605 36128 2688 36156
rect 2605 36125 2617 36128
rect 2559 36119 2617 36125
rect 2682 36116 2688 36128
rect 2740 36116 2746 36168
rect 3050 36116 3056 36168
rect 3108 36116 3114 36168
rect 3786 36116 3792 36168
rect 3844 36116 3850 36168
rect 4338 36116 4344 36168
rect 4396 36116 4402 36168
rect 4430 36116 4436 36168
rect 4488 36156 4494 36168
rect 4985 36159 5043 36165
rect 4985 36156 4997 36159
rect 4488 36128 4997 36156
rect 4488 36116 4494 36128
rect 4985 36125 4997 36128
rect 5031 36156 5043 36159
rect 5074 36156 5080 36168
rect 5031 36128 5080 36156
rect 5031 36125 5043 36128
rect 4985 36119 5043 36125
rect 5074 36116 5080 36128
rect 5132 36116 5138 36168
rect 5902 36116 5908 36168
rect 5960 36116 5966 36168
rect 7101 36159 7159 36165
rect 7101 36125 7113 36159
rect 7147 36156 7159 36159
rect 7282 36156 7288 36168
rect 7147 36128 7288 36156
rect 7147 36125 7159 36128
rect 7101 36119 7159 36125
rect 7282 36116 7288 36128
rect 7340 36116 7346 36168
rect 9401 36159 9459 36165
rect 9401 36125 9413 36159
rect 9447 36125 9459 36159
rect 9401 36119 9459 36125
rect 9675 36159 9733 36165
rect 9675 36125 9687 36159
rect 9721 36156 9733 36159
rect 10042 36156 10048 36168
rect 9721 36128 10048 36156
rect 9721 36125 9733 36128
rect 9675 36119 9733 36125
rect 1673 36091 1731 36097
rect 1673 36057 1685 36091
rect 1719 36088 1731 36091
rect 1719 36060 2728 36088
rect 1719 36057 1731 36060
rect 1673 36051 1731 36057
rect 2700 36032 2728 36060
rect 4062 36048 4068 36100
rect 4120 36048 4126 36100
rect 4617 36091 4675 36097
rect 4617 36057 4629 36091
rect 4663 36088 4675 36091
rect 5166 36088 5172 36100
rect 4663 36060 5172 36088
rect 4663 36057 4675 36060
rect 4617 36051 4675 36057
rect 5166 36048 5172 36060
rect 5224 36048 5230 36100
rect 9416 36088 9444 36119
rect 10042 36116 10048 36128
rect 10100 36116 10106 36168
rect 10152 36156 10180 36332
rect 10778 36320 10784 36372
rect 10836 36360 10842 36372
rect 14550 36360 14556 36372
rect 10836 36332 14556 36360
rect 10836 36320 10842 36332
rect 14550 36320 14556 36332
rect 14608 36360 14614 36372
rect 16574 36360 16580 36372
rect 14608 36332 16580 36360
rect 14608 36320 14614 36332
rect 16574 36320 16580 36332
rect 16632 36320 16638 36372
rect 21545 36363 21603 36369
rect 21545 36329 21557 36363
rect 21591 36360 21603 36363
rect 22278 36360 22284 36372
rect 21591 36332 22284 36360
rect 21591 36329 21603 36332
rect 21545 36323 21603 36329
rect 22278 36320 22284 36332
rect 22336 36320 22342 36372
rect 22480 36332 22692 36360
rect 10796 36233 10824 36320
rect 15102 36252 15108 36304
rect 15160 36292 15166 36304
rect 18322 36292 18328 36304
rect 15160 36264 18328 36292
rect 15160 36252 15166 36264
rect 18322 36252 18328 36264
rect 18380 36252 18386 36304
rect 19978 36252 19984 36304
rect 20036 36292 20042 36304
rect 22480 36292 22508 36332
rect 20036 36264 22508 36292
rect 22557 36295 22615 36301
rect 20036 36252 20042 36264
rect 22557 36261 22569 36295
rect 22603 36261 22615 36295
rect 22664 36292 22692 36332
rect 22830 36320 22836 36372
rect 22888 36320 22894 36372
rect 23201 36295 23259 36301
rect 23201 36292 23213 36295
rect 22664 36264 23213 36292
rect 22557 36255 22615 36261
rect 23201 36261 23213 36264
rect 23247 36261 23259 36295
rect 23201 36255 23259 36261
rect 10781 36227 10839 36233
rect 10781 36193 10793 36227
rect 10827 36193 10839 36227
rect 20346 36224 20352 36236
rect 10781 36187 10839 36193
rect 11992 36196 12204 36224
rect 11023 36159 11081 36165
rect 11023 36156 11035 36159
rect 10152 36128 11035 36156
rect 11023 36125 11035 36128
rect 11069 36156 11081 36159
rect 11992 36156 12020 36196
rect 11069 36128 12020 36156
rect 11069 36125 11081 36128
rect 11023 36119 11081 36125
rect 10318 36088 10324 36100
rect 9416 36060 10324 36088
rect 10318 36048 10324 36060
rect 10376 36088 10382 36100
rect 11882 36088 11888 36100
rect 10376 36060 11888 36088
rect 10376 36048 10382 36060
rect 11882 36048 11888 36060
rect 11940 36048 11946 36100
rect 12176 36088 12204 36196
rect 17880 36196 20352 36224
rect 12250 36116 12256 36168
rect 12308 36116 12314 36168
rect 12434 36116 12440 36168
rect 12492 36156 12498 36168
rect 12527 36159 12585 36165
rect 12527 36156 12539 36159
rect 12492 36128 12539 36156
rect 12492 36116 12498 36128
rect 12527 36125 12539 36128
rect 12573 36156 12585 36159
rect 13722 36156 13728 36168
rect 12573 36128 13728 36156
rect 12573 36125 12585 36128
rect 12527 36119 12585 36125
rect 13722 36116 13728 36128
rect 13780 36116 13786 36168
rect 17880 36088 17908 36196
rect 20346 36184 20352 36196
rect 20404 36224 20410 36236
rect 21266 36224 21272 36236
rect 20404 36196 21272 36224
rect 20404 36184 20410 36196
rect 21266 36184 21272 36196
rect 21324 36184 21330 36236
rect 22572 36224 22600 36255
rect 23474 36252 23480 36304
rect 23532 36292 23538 36304
rect 24302 36292 24308 36304
rect 23532 36264 24308 36292
rect 23532 36252 23538 36264
rect 24302 36252 24308 36264
rect 24360 36252 24366 36304
rect 22572 36196 23060 36224
rect 18325 36159 18383 36165
rect 18325 36156 18337 36159
rect 12176 36060 17908 36088
rect 17972 36128 18337 36156
rect 17972 36032 18000 36128
rect 18325 36125 18337 36128
rect 18371 36125 18383 36159
rect 18325 36119 18383 36125
rect 18693 36159 18751 36165
rect 18693 36125 18705 36159
rect 18739 36125 18751 36159
rect 18693 36119 18751 36125
rect 18785 36159 18843 36165
rect 18785 36125 18797 36159
rect 18831 36156 18843 36159
rect 19242 36156 19248 36168
rect 18831 36128 19248 36156
rect 18831 36125 18843 36128
rect 18785 36119 18843 36125
rect 18708 36088 18736 36119
rect 19242 36116 19248 36128
rect 19300 36116 19306 36168
rect 19426 36116 19432 36168
rect 19484 36116 19490 36168
rect 20257 36159 20315 36165
rect 20257 36156 20269 36159
rect 19904 36128 20269 36156
rect 18156 36060 18736 36088
rect 1176 35992 1624 36020
rect 1176 35980 1182 35992
rect 2682 35980 2688 36032
rect 2740 35980 2746 36032
rect 4154 35980 4160 36032
rect 4212 36020 4218 36032
rect 8386 36020 8392 36032
rect 4212 35992 8392 36020
rect 4212 35980 4218 35992
rect 8386 35980 8392 35992
rect 8444 35980 8450 36032
rect 9950 35980 9956 36032
rect 10008 36020 10014 36032
rect 10413 36023 10471 36029
rect 10413 36020 10425 36023
rect 10008 35992 10425 36020
rect 10008 35980 10014 35992
rect 10413 35989 10425 35992
rect 10459 35989 10471 36023
rect 10413 35983 10471 35989
rect 11330 35980 11336 36032
rect 11388 36020 11394 36032
rect 11793 36023 11851 36029
rect 11793 36020 11805 36023
rect 11388 35992 11805 36020
rect 11388 35980 11394 35992
rect 11793 35989 11805 35992
rect 11839 35989 11851 36023
rect 11793 35983 11851 35989
rect 12158 35980 12164 36032
rect 12216 36020 12222 36032
rect 13265 36023 13323 36029
rect 13265 36020 13277 36023
rect 12216 35992 13277 36020
rect 12216 35980 12222 35992
rect 13265 35989 13277 35992
rect 13311 35989 13323 36023
rect 13265 35983 13323 35989
rect 17954 35980 17960 36032
rect 18012 35980 18018 36032
rect 18156 36029 18184 36060
rect 19904 36032 19932 36128
rect 20257 36125 20269 36128
rect 20303 36125 20315 36159
rect 20257 36119 20315 36125
rect 20622 36116 20628 36168
rect 20680 36156 20686 36168
rect 21729 36159 21787 36165
rect 21729 36156 21741 36159
rect 20680 36128 21741 36156
rect 20680 36116 20686 36128
rect 21729 36125 21741 36128
rect 21775 36125 21787 36159
rect 21729 36119 21787 36125
rect 22738 36116 22744 36168
rect 22796 36116 22802 36168
rect 23032 36165 23060 36196
rect 23290 36184 23296 36236
rect 23348 36224 23354 36236
rect 23348 36196 23888 36224
rect 23348 36184 23354 36196
rect 23860 36165 23888 36196
rect 23017 36159 23075 36165
rect 23017 36125 23029 36159
rect 23063 36125 23075 36159
rect 23017 36119 23075 36125
rect 23385 36159 23443 36165
rect 23385 36125 23397 36159
rect 23431 36156 23443 36159
rect 23661 36159 23719 36165
rect 23431 36128 23520 36156
rect 23431 36125 23443 36128
rect 23385 36119 23443 36125
rect 18141 36023 18199 36029
rect 18141 35989 18153 36023
rect 18187 35989 18199 36023
rect 18141 35983 18199 35989
rect 19245 36023 19303 36029
rect 19245 35989 19257 36023
rect 19291 36020 19303 36023
rect 19334 36020 19340 36032
rect 19291 35992 19340 36020
rect 19291 35989 19303 35992
rect 19245 35983 19303 35989
rect 19334 35980 19340 35992
rect 19392 35980 19398 36032
rect 19886 35980 19892 36032
rect 19944 35980 19950 36032
rect 20073 36023 20131 36029
rect 20073 35989 20085 36023
rect 20119 36020 20131 36023
rect 21542 36020 21548 36032
rect 20119 35992 21548 36020
rect 20119 35989 20131 35992
rect 20073 35983 20131 35989
rect 21542 35980 21548 35992
rect 21600 35980 21606 36032
rect 23492 36029 23520 36128
rect 23661 36125 23673 36159
rect 23707 36125 23719 36159
rect 23661 36119 23719 36125
rect 23845 36159 23903 36165
rect 23845 36125 23857 36159
rect 23891 36125 23903 36159
rect 23845 36119 23903 36125
rect 23676 36088 23704 36119
rect 25406 36088 25412 36100
rect 23676 36060 25412 36088
rect 25406 36048 25412 36060
rect 25464 36048 25470 36100
rect 23477 36023 23535 36029
rect 23477 35989 23489 36023
rect 23523 35989 23535 36023
rect 23477 35983 23535 35989
rect 24118 35980 24124 36032
rect 24176 35980 24182 36032
rect 1104 35930 25000 35952
rect 1104 35878 6884 35930
rect 6936 35878 6948 35930
rect 7000 35878 7012 35930
rect 7064 35878 7076 35930
rect 7128 35878 7140 35930
rect 7192 35878 12818 35930
rect 12870 35878 12882 35930
rect 12934 35878 12946 35930
rect 12998 35878 13010 35930
rect 13062 35878 13074 35930
rect 13126 35878 18752 35930
rect 18804 35878 18816 35930
rect 18868 35878 18880 35930
rect 18932 35878 18944 35930
rect 18996 35878 19008 35930
rect 19060 35878 24686 35930
rect 24738 35878 24750 35930
rect 24802 35878 24814 35930
rect 24866 35878 24878 35930
rect 24930 35878 24942 35930
rect 24994 35878 25000 35930
rect 1104 35856 25000 35878
rect 3510 35776 3516 35828
rect 3568 35816 3574 35828
rect 4706 35816 4712 35828
rect 3568 35788 4712 35816
rect 3568 35776 3574 35788
rect 4706 35776 4712 35788
rect 4764 35776 4770 35828
rect 6181 35819 6239 35825
rect 6181 35785 6193 35819
rect 6227 35816 6239 35819
rect 7282 35816 7288 35828
rect 6227 35788 7288 35816
rect 6227 35785 6239 35788
rect 6181 35779 6239 35785
rect 7282 35776 7288 35788
rect 7340 35776 7346 35828
rect 9398 35776 9404 35828
rect 9456 35816 9462 35828
rect 9456 35788 9720 35816
rect 9456 35776 9462 35788
rect 1302 35708 1308 35760
rect 1360 35748 1366 35760
rect 1360 35720 3832 35748
rect 1360 35708 1366 35720
rect 1397 35683 1455 35689
rect 1397 35649 1409 35683
rect 1443 35680 1455 35683
rect 1486 35680 1492 35692
rect 1443 35652 1492 35680
rect 1443 35649 1455 35652
rect 1397 35643 1455 35649
rect 1486 35640 1492 35652
rect 1544 35640 1550 35692
rect 2682 35680 2688 35692
rect 2643 35652 2688 35680
rect 2682 35640 2688 35652
rect 2740 35640 2746 35692
rect 3050 35640 3056 35692
rect 3108 35640 3114 35692
rect 3804 35689 3832 35720
rect 6454 35708 6460 35760
rect 6512 35748 6518 35760
rect 7374 35748 7380 35760
rect 6512 35720 7380 35748
rect 6512 35708 6518 35720
rect 7374 35708 7380 35720
rect 7432 35708 7438 35760
rect 8021 35751 8079 35757
rect 8021 35717 8033 35751
rect 8067 35748 8079 35751
rect 8202 35748 8208 35760
rect 8067 35720 8208 35748
rect 8067 35717 8079 35720
rect 8021 35711 8079 35717
rect 8202 35708 8208 35720
rect 8260 35708 8266 35760
rect 8297 35751 8355 35757
rect 8297 35717 8309 35751
rect 8343 35748 8355 35751
rect 9125 35751 9183 35757
rect 9125 35748 9137 35751
rect 8343 35720 8524 35748
rect 8343 35717 8355 35720
rect 8297 35711 8355 35717
rect 8496 35692 8524 35720
rect 8680 35720 9137 35748
rect 8680 35692 8708 35720
rect 9125 35717 9137 35720
rect 9171 35748 9183 35751
rect 9582 35748 9588 35760
rect 9171 35720 9588 35748
rect 9171 35717 9183 35720
rect 9125 35711 9183 35717
rect 9582 35708 9588 35720
rect 9640 35708 9646 35760
rect 3789 35683 3847 35689
rect 3789 35649 3801 35683
rect 3835 35649 3847 35683
rect 3789 35643 3847 35649
rect 6178 35640 6184 35692
rect 6236 35640 6242 35692
rect 8386 35640 8392 35692
rect 8444 35640 8450 35692
rect 8478 35640 8484 35692
rect 8536 35640 8542 35692
rect 8662 35640 8668 35692
rect 8720 35640 8726 35692
rect 8754 35640 8760 35692
rect 8812 35680 8818 35692
rect 9214 35680 9220 35692
rect 8812 35652 9220 35680
rect 8812 35640 8818 35652
rect 9214 35640 9220 35652
rect 9272 35640 9278 35692
rect 9692 35689 9720 35788
rect 10226 35776 10232 35828
rect 10284 35816 10290 35828
rect 10284 35788 11192 35816
rect 10284 35776 10290 35788
rect 11164 35748 11192 35788
rect 11790 35776 11796 35828
rect 11848 35776 11854 35828
rect 11900 35788 12572 35816
rect 11900 35748 11928 35788
rect 12544 35757 12572 35788
rect 13446 35776 13452 35828
rect 13504 35816 13510 35828
rect 18138 35816 18144 35828
rect 13504 35788 18144 35816
rect 13504 35776 13510 35788
rect 11164 35720 11928 35748
rect 12529 35751 12587 35757
rect 12529 35717 12541 35751
rect 12575 35717 12587 35751
rect 12529 35711 12587 35717
rect 12894 35708 12900 35760
rect 12952 35708 12958 35760
rect 14382 35719 14410 35788
rect 18138 35776 18144 35788
rect 18196 35776 18202 35828
rect 19061 35819 19119 35825
rect 19061 35785 19073 35819
rect 19107 35816 19119 35819
rect 19426 35816 19432 35828
rect 19107 35788 19432 35816
rect 19107 35785 19119 35788
rect 19061 35779 19119 35785
rect 19426 35776 19432 35788
rect 19484 35776 19490 35828
rect 19702 35816 19708 35828
rect 19628 35788 19708 35816
rect 19628 35748 19656 35788
rect 19702 35776 19708 35788
rect 19760 35776 19766 35828
rect 20993 35819 21051 35825
rect 20993 35785 21005 35819
rect 21039 35816 21051 35819
rect 22649 35819 22707 35825
rect 21039 35788 21956 35816
rect 21039 35785 21051 35788
rect 20993 35779 21051 35785
rect 19886 35757 19892 35760
rect 19858 35751 19892 35757
rect 19858 35748 19870 35751
rect 14351 35713 14410 35719
rect 9677 35683 9735 35689
rect 9677 35649 9689 35683
rect 9723 35649 9735 35683
rect 9677 35643 9735 35649
rect 10410 35640 10416 35692
rect 10468 35640 10474 35692
rect 10530 35683 10588 35689
rect 10530 35680 10542 35683
rect 10518 35649 10542 35680
rect 10576 35649 10588 35683
rect 10518 35643 10588 35649
rect 11333 35683 11391 35689
rect 11333 35649 11345 35683
rect 11379 35680 11391 35683
rect 11974 35680 11980 35692
rect 11379 35652 11980 35680
rect 11379 35649 11391 35652
rect 11333 35643 11391 35649
rect 1670 35572 1676 35624
rect 1728 35572 1734 35624
rect 2409 35615 2467 35621
rect 2409 35581 2421 35615
rect 2455 35581 2467 35615
rect 2409 35575 2467 35581
rect 2424 35476 2452 35575
rect 3068 35476 3096 35640
rect 3326 35572 3332 35624
rect 3384 35612 3390 35624
rect 3973 35615 4031 35621
rect 3973 35612 3985 35615
rect 3384 35584 3985 35612
rect 3384 35572 3390 35584
rect 3973 35581 3985 35584
rect 4019 35612 4031 35615
rect 4154 35612 4160 35624
rect 4019 35584 4160 35612
rect 4019 35581 4031 35584
rect 3973 35575 4031 35581
rect 4154 35572 4160 35584
rect 4212 35572 4218 35624
rect 4341 35615 4399 35621
rect 4341 35581 4353 35615
rect 4387 35581 4399 35615
rect 4341 35575 4399 35581
rect 4356 35544 4384 35575
rect 4522 35572 4528 35624
rect 4580 35572 4586 35624
rect 5258 35572 5264 35624
rect 5316 35572 5322 35624
rect 5350 35572 5356 35624
rect 5408 35621 5414 35624
rect 5408 35615 5436 35621
rect 5424 35581 5436 35615
rect 5408 35575 5436 35581
rect 5537 35615 5595 35621
rect 5537 35581 5549 35615
rect 5583 35612 5595 35615
rect 6196 35612 6224 35640
rect 5583 35584 6224 35612
rect 5583 35581 5595 35584
rect 5537 35575 5595 35581
rect 5408 35572 5414 35575
rect 8202 35572 8208 35624
rect 8260 35572 8266 35624
rect 9493 35615 9551 35621
rect 9493 35581 9505 35615
rect 9539 35581 9551 35615
rect 9493 35575 9551 35581
rect 4614 35544 4620 35556
rect 4356 35516 4620 35544
rect 4614 35504 4620 35516
rect 4672 35504 4678 35556
rect 4985 35547 5043 35553
rect 4985 35513 4997 35547
rect 5031 35513 5043 35547
rect 4985 35507 5043 35513
rect 2424 35448 3096 35476
rect 3418 35436 3424 35488
rect 3476 35436 3482 35488
rect 5000 35476 5028 35507
rect 9508 35488 9536 35575
rect 10226 35572 10232 35624
rect 10284 35612 10290 35624
rect 10518 35612 10546 35643
rect 11974 35640 11980 35652
rect 12032 35640 12038 35692
rect 12066 35640 12072 35692
rect 12124 35640 12130 35692
rect 12158 35640 12164 35692
rect 12216 35640 12222 35692
rect 12250 35640 12256 35692
rect 12308 35680 12314 35692
rect 12308 35652 14136 35680
rect 14351 35679 14363 35713
rect 14397 35682 14410 35713
rect 17696 35720 19656 35748
rect 14397 35679 14409 35682
rect 14351 35673 14409 35679
rect 12308 35640 12314 35652
rect 10284 35584 10546 35612
rect 10699 35615 10757 35621
rect 10284 35572 10290 35584
rect 10699 35581 10711 35615
rect 10745 35612 10757 35615
rect 11238 35612 11244 35624
rect 10745 35584 11244 35612
rect 10745 35581 10757 35584
rect 10699 35575 10757 35581
rect 11238 35572 11244 35584
rect 11296 35572 11302 35624
rect 13078 35612 13084 35624
rect 12834 35584 13084 35612
rect 13078 35572 13084 35584
rect 13136 35572 13142 35624
rect 14108 35621 14136 35652
rect 17696 35624 17724 35720
rect 17954 35689 17960 35692
rect 17948 35680 17960 35689
rect 17915 35652 17960 35680
rect 17948 35643 17960 35652
rect 17954 35640 17960 35643
rect 18012 35640 18018 35692
rect 19150 35640 19156 35692
rect 19208 35640 19214 35692
rect 19242 35640 19248 35692
rect 19300 35640 19306 35692
rect 19628 35689 19656 35720
rect 19720 35720 19870 35748
rect 19613 35683 19671 35689
rect 19613 35649 19625 35683
rect 19659 35649 19671 35683
rect 19613 35643 19671 35649
rect 14093 35615 14151 35621
rect 14093 35581 14105 35615
rect 14139 35581 14151 35615
rect 14093 35575 14151 35581
rect 9950 35504 9956 35556
rect 10008 35544 10014 35556
rect 10137 35547 10195 35553
rect 10137 35544 10149 35547
rect 10008 35516 10149 35544
rect 10008 35504 10014 35516
rect 10137 35513 10149 35516
rect 10183 35513 10195 35547
rect 14108 35544 14136 35575
rect 17678 35572 17684 35624
rect 17736 35572 17742 35624
rect 19426 35572 19432 35624
rect 19484 35572 19490 35624
rect 19720 35612 19748 35720
rect 19858 35717 19870 35720
rect 19858 35711 19892 35717
rect 19886 35708 19892 35711
rect 19944 35708 19950 35760
rect 21361 35751 21419 35757
rect 21361 35717 21373 35751
rect 21407 35748 21419 35751
rect 21726 35748 21732 35760
rect 21407 35720 21732 35748
rect 21407 35717 21419 35720
rect 21361 35711 21419 35717
rect 21726 35708 21732 35720
rect 21784 35708 21790 35760
rect 21085 35683 21143 35689
rect 21085 35649 21097 35683
rect 21131 35680 21143 35683
rect 21266 35680 21272 35692
rect 21131 35652 21272 35680
rect 21131 35649 21143 35652
rect 21085 35643 21143 35649
rect 21266 35640 21272 35652
rect 21324 35640 21330 35692
rect 21453 35683 21511 35689
rect 21453 35649 21465 35683
rect 21499 35678 21511 35683
rect 21542 35678 21548 35692
rect 21499 35650 21548 35678
rect 21499 35649 21511 35650
rect 21453 35643 21511 35649
rect 21542 35640 21548 35650
rect 21600 35640 21606 35692
rect 21928 35684 21956 35788
rect 22649 35785 22661 35819
rect 22695 35816 22707 35819
rect 22738 35816 22744 35828
rect 22695 35788 22744 35816
rect 22695 35785 22707 35788
rect 22649 35779 22707 35785
rect 22738 35776 22744 35788
rect 22796 35776 22802 35828
rect 22925 35819 22983 35825
rect 22925 35785 22937 35819
rect 22971 35785 22983 35819
rect 22925 35779 22983 35785
rect 22186 35708 22192 35760
rect 22244 35748 22250 35760
rect 22940 35748 22968 35779
rect 23290 35776 23296 35828
rect 23348 35776 23354 35828
rect 23569 35819 23627 35825
rect 23569 35785 23581 35819
rect 23615 35816 23627 35819
rect 23842 35816 23848 35828
rect 23615 35788 23848 35816
rect 23615 35785 23627 35788
rect 23569 35779 23627 35785
rect 23842 35776 23848 35788
rect 23900 35776 23906 35828
rect 22244 35720 22876 35748
rect 22940 35720 23520 35748
rect 22244 35708 22250 35720
rect 21997 35687 22055 35693
rect 21997 35684 22009 35687
rect 21928 35656 22009 35684
rect 21997 35653 22009 35656
rect 22043 35653 22055 35687
rect 21997 35647 22055 35653
rect 22094 35640 22100 35692
rect 22152 35640 22158 35692
rect 22281 35683 22339 35689
rect 22281 35649 22293 35683
rect 22327 35649 22339 35683
rect 22281 35643 22339 35649
rect 19628 35584 19748 35612
rect 21361 35615 21419 35621
rect 14108 35516 14228 35544
rect 10137 35507 10195 35513
rect 14200 35488 14228 35516
rect 15286 35504 15292 35556
rect 15344 35504 15350 35556
rect 19628 35544 19656 35584
rect 21361 35581 21373 35615
rect 21407 35612 21419 35615
rect 22189 35615 22247 35621
rect 22189 35612 22201 35615
rect 21407 35584 22201 35612
rect 21407 35581 21419 35584
rect 21361 35575 21419 35581
rect 22189 35581 22201 35584
rect 22235 35581 22247 35615
rect 22189 35575 22247 35581
rect 18616 35516 19656 35544
rect 21177 35547 21235 35553
rect 5626 35476 5632 35488
rect 5000 35448 5632 35476
rect 5626 35436 5632 35448
rect 5684 35436 5690 35488
rect 9306 35436 9312 35488
rect 9364 35436 9370 35488
rect 9490 35436 9496 35488
rect 9548 35436 9554 35488
rect 13081 35479 13139 35485
rect 13081 35445 13093 35479
rect 13127 35476 13139 35479
rect 13906 35476 13912 35488
rect 13127 35448 13912 35476
rect 13127 35445 13139 35448
rect 13081 35439 13139 35445
rect 13906 35436 13912 35448
rect 13964 35436 13970 35488
rect 14182 35436 14188 35488
rect 14240 35436 14246 35488
rect 14458 35436 14464 35488
rect 14516 35476 14522 35488
rect 15105 35479 15163 35485
rect 15105 35476 15117 35479
rect 14516 35448 15117 35476
rect 14516 35436 14522 35448
rect 15105 35445 15117 35448
rect 15151 35445 15163 35479
rect 15304 35476 15332 35504
rect 18616 35476 18644 35516
rect 21177 35513 21189 35547
rect 21223 35544 21235 35547
rect 21545 35547 21603 35553
rect 21545 35544 21557 35547
rect 21223 35516 21312 35544
rect 21223 35513 21235 35516
rect 21177 35507 21235 35513
rect 15304 35448 18644 35476
rect 19337 35479 19395 35485
rect 15105 35439 15163 35445
rect 19337 35445 19349 35479
rect 19383 35476 19395 35479
rect 20714 35476 20720 35488
rect 19383 35448 20720 35476
rect 19383 35445 19395 35448
rect 19337 35439 19395 35445
rect 20714 35436 20720 35448
rect 20772 35436 20778 35488
rect 21284 35476 21312 35516
rect 21468 35516 21557 35544
rect 21468 35476 21496 35516
rect 21545 35513 21557 35516
rect 21591 35513 21603 35547
rect 21545 35507 21603 35513
rect 21821 35547 21879 35553
rect 21821 35513 21833 35547
rect 21867 35544 21879 35547
rect 22296 35544 22324 35643
rect 22554 35640 22560 35692
rect 22612 35640 22618 35692
rect 22848 35689 22876 35720
rect 23492 35689 23520 35720
rect 22833 35683 22891 35689
rect 22833 35649 22845 35683
rect 22879 35649 22891 35683
rect 22833 35643 22891 35649
rect 23109 35683 23167 35689
rect 23109 35649 23121 35683
rect 23155 35649 23167 35683
rect 23109 35643 23167 35649
rect 23477 35683 23535 35689
rect 23477 35649 23489 35683
rect 23523 35649 23535 35683
rect 23477 35643 23535 35649
rect 23753 35683 23811 35689
rect 23753 35649 23765 35683
rect 23799 35649 23811 35683
rect 23753 35643 23811 35649
rect 23124 35612 23152 35643
rect 22388 35584 23152 35612
rect 22388 35553 22416 35584
rect 21867 35516 22324 35544
rect 22373 35547 22431 35553
rect 21867 35513 21879 35516
rect 21821 35507 21879 35513
rect 22373 35513 22385 35547
rect 22419 35513 22431 35547
rect 22373 35507 22431 35513
rect 22922 35504 22928 35556
rect 22980 35544 22986 35556
rect 23768 35544 23796 35643
rect 24118 35640 24124 35692
rect 24176 35640 24182 35692
rect 25682 35544 25688 35556
rect 22980 35516 23796 35544
rect 24320 35516 25688 35544
rect 22980 35504 22986 35516
rect 21284 35448 21496 35476
rect 21726 35436 21732 35488
rect 21784 35476 21790 35488
rect 24320 35476 24348 35516
rect 25682 35504 25688 35516
rect 25740 35504 25746 35556
rect 21784 35448 24348 35476
rect 21784 35436 21790 35448
rect 24394 35436 24400 35488
rect 24452 35436 24458 35488
rect 1104 35386 24840 35408
rect 1104 35334 3917 35386
rect 3969 35334 3981 35386
rect 4033 35334 4045 35386
rect 4097 35334 4109 35386
rect 4161 35334 4173 35386
rect 4225 35334 9851 35386
rect 9903 35334 9915 35386
rect 9967 35334 9979 35386
rect 10031 35334 10043 35386
rect 10095 35334 10107 35386
rect 10159 35334 15785 35386
rect 15837 35334 15849 35386
rect 15901 35334 15913 35386
rect 15965 35334 15977 35386
rect 16029 35334 16041 35386
rect 16093 35334 21719 35386
rect 21771 35334 21783 35386
rect 21835 35334 21847 35386
rect 21899 35334 21911 35386
rect 21963 35334 21975 35386
rect 22027 35334 24840 35386
rect 1104 35312 24840 35334
rect 3142 35272 3148 35284
rect 2332 35244 3148 35272
rect 1581 35139 1639 35145
rect 1581 35105 1593 35139
rect 1627 35136 1639 35139
rect 1670 35136 1676 35148
rect 1627 35108 1676 35136
rect 1627 35105 1639 35108
rect 1581 35099 1639 35105
rect 1670 35096 1676 35108
rect 1728 35096 1734 35148
rect 2222 35096 2228 35148
rect 2280 35096 2286 35148
rect 2332 35136 2360 35244
rect 3142 35232 3148 35244
rect 3200 35232 3206 35284
rect 3421 35275 3479 35281
rect 3421 35241 3433 35275
rect 3467 35272 3479 35275
rect 3694 35272 3700 35284
rect 3467 35244 3700 35272
rect 3467 35241 3479 35244
rect 3421 35235 3479 35241
rect 3694 35232 3700 35244
rect 3752 35232 3758 35284
rect 5810 35232 5816 35284
rect 5868 35272 5874 35284
rect 6178 35272 6184 35284
rect 5868 35244 6184 35272
rect 5868 35232 5874 35244
rect 6178 35232 6184 35244
rect 6236 35232 6242 35284
rect 7742 35272 7748 35284
rect 7300 35244 7748 35272
rect 5828 35204 5856 35232
rect 5736 35176 5856 35204
rect 2501 35139 2559 35145
rect 2501 35136 2513 35139
rect 2332 35108 2513 35136
rect 2501 35105 2513 35108
rect 2547 35105 2559 35139
rect 2501 35099 2559 35105
rect 2639 35139 2697 35145
rect 2639 35105 2651 35139
rect 2685 35136 2697 35139
rect 2685 35108 3372 35136
rect 2685 35105 2697 35108
rect 2639 35099 2697 35105
rect 1765 35071 1823 35077
rect 1765 35037 1777 35071
rect 1811 35037 1823 35071
rect 1765 35031 1823 35037
rect 1780 34932 1808 35031
rect 2774 35028 2780 35080
rect 2832 35028 2838 35080
rect 3344 35068 3372 35108
rect 3418 35096 3424 35148
rect 3476 35136 3482 35148
rect 5736 35145 5764 35176
rect 7300 35145 7328 35244
rect 7742 35232 7748 35244
rect 7800 35232 7806 35284
rect 8202 35232 8208 35284
rect 8260 35272 8266 35284
rect 8297 35275 8355 35281
rect 8297 35272 8309 35275
rect 8260 35244 8309 35272
rect 8260 35232 8266 35244
rect 8297 35241 8309 35244
rect 8343 35241 8355 35275
rect 8297 35235 8355 35241
rect 8662 35232 8668 35284
rect 8720 35272 8726 35284
rect 10318 35272 10324 35284
rect 8720 35244 10324 35272
rect 8720 35232 8726 35244
rect 10318 35232 10324 35244
rect 10376 35232 10382 35284
rect 13078 35232 13084 35284
rect 13136 35232 13142 35284
rect 13722 35232 13728 35284
rect 13780 35272 13786 35284
rect 19337 35275 19395 35281
rect 13780 35244 19288 35272
rect 13780 35232 13786 35244
rect 9398 35204 9404 35216
rect 7944 35176 9404 35204
rect 5721 35139 5779 35145
rect 3476 35108 3818 35136
rect 3476 35096 3482 35108
rect 5721 35105 5733 35139
rect 5767 35105 5779 35139
rect 5721 35099 5779 35105
rect 7285 35139 7343 35145
rect 7285 35105 7297 35139
rect 7331 35105 7343 35139
rect 7285 35099 7343 35105
rect 7944 35080 7972 35176
rect 9398 35164 9404 35176
rect 9456 35204 9462 35216
rect 10781 35207 10839 35213
rect 9456 35176 9812 35204
rect 9456 35164 9462 35176
rect 9784 35136 9812 35176
rect 10781 35173 10793 35207
rect 10827 35204 10839 35207
rect 10870 35204 10876 35216
rect 10827 35176 10876 35204
rect 10827 35173 10839 35176
rect 10781 35167 10839 35173
rect 10870 35164 10876 35176
rect 10928 35164 10934 35216
rect 18785 35207 18843 35213
rect 18785 35173 18797 35207
rect 18831 35204 18843 35207
rect 19150 35204 19156 35216
rect 18831 35176 19156 35204
rect 18831 35173 18843 35176
rect 18785 35167 18843 35173
rect 19150 35164 19156 35176
rect 19208 35164 19214 35216
rect 19260 35204 19288 35244
rect 19337 35241 19349 35275
rect 19383 35272 19395 35275
rect 19426 35272 19432 35284
rect 19383 35244 19432 35272
rect 19383 35241 19395 35244
rect 19337 35235 19395 35241
rect 19426 35232 19432 35244
rect 19484 35232 19490 35284
rect 20364 35244 21220 35272
rect 20364 35204 20392 35244
rect 21192 35216 21220 35244
rect 21266 35232 21272 35284
rect 21324 35272 21330 35284
rect 21910 35272 21916 35284
rect 21324 35244 21916 35272
rect 21324 35232 21330 35244
rect 21910 35232 21916 35244
rect 21968 35232 21974 35284
rect 22554 35272 22560 35284
rect 22020 35244 22560 35272
rect 19260 35176 20392 35204
rect 21174 35164 21180 35216
rect 21232 35164 21238 35216
rect 10321 35139 10379 35145
rect 10321 35136 10333 35139
rect 8036 35108 9674 35136
rect 9784 35108 10333 35136
rect 8036 35080 8064 35108
rect 4062 35068 4068 35080
rect 3344 35040 4068 35068
rect 4062 35028 4068 35040
rect 4120 35028 4126 35080
rect 4246 35028 4252 35080
rect 4304 35028 4310 35080
rect 5166 35028 5172 35080
rect 5224 35068 5230 35080
rect 5995 35071 6053 35077
rect 5995 35068 6007 35071
rect 5224 35040 6007 35068
rect 5224 35028 5230 35040
rect 5995 35037 6007 35040
rect 6041 35068 6053 35071
rect 7558 35068 7564 35080
rect 6041 35040 7144 35068
rect 7519 35040 7564 35068
rect 6041 35037 6053 35040
rect 5995 35031 6053 35037
rect 3252 34972 4106 35000
rect 3252 34932 3280 34972
rect 1780 34904 3280 34932
rect 3418 34892 3424 34944
rect 3476 34932 3482 34944
rect 3973 34935 4031 34941
rect 3973 34932 3985 34935
rect 3476 34904 3985 34932
rect 3476 34892 3482 34904
rect 3973 34901 3985 34904
rect 4019 34901 4031 34935
rect 4078 34932 4106 34972
rect 4154 34960 4160 35012
rect 4212 35000 4218 35012
rect 4341 35003 4399 35009
rect 4341 35000 4353 35003
rect 4212 34972 4353 35000
rect 4212 34960 4218 34972
rect 4341 34969 4353 34972
rect 4387 34969 4399 35003
rect 4341 34963 4399 34969
rect 4709 35003 4767 35009
rect 4709 34969 4721 35003
rect 4755 35000 4767 35003
rect 4798 35000 4804 35012
rect 4755 34972 4804 35000
rect 4755 34969 4767 34972
rect 4709 34963 4767 34969
rect 4798 34960 4804 34972
rect 4856 34960 4862 35012
rect 7116 35000 7144 35040
rect 7558 35028 7564 35040
rect 7616 35028 7622 35080
rect 7926 35028 7932 35080
rect 7984 35028 7990 35080
rect 8018 35028 8024 35080
rect 8076 35028 8082 35080
rect 8294 35028 8300 35080
rect 8352 35068 8358 35080
rect 8478 35068 8484 35080
rect 8352 35040 8484 35068
rect 8352 35028 8358 35040
rect 8478 35028 8484 35040
rect 8536 35028 8542 35080
rect 9646 35068 9674 35108
rect 10321 35105 10333 35108
rect 10367 35105 10379 35139
rect 10321 35099 10379 35105
rect 12066 35096 12072 35148
rect 12124 35096 12130 35148
rect 19334 35096 19340 35148
rect 19392 35096 19398 35148
rect 22020 35136 22048 35244
rect 22554 35232 22560 35244
rect 22612 35232 22618 35284
rect 23198 35232 23204 35284
rect 23256 35232 23262 35284
rect 24118 35232 24124 35284
rect 24176 35232 24182 35284
rect 22189 35207 22247 35213
rect 22189 35173 22201 35207
rect 22235 35204 22247 35207
rect 24136 35204 24164 35232
rect 22235 35176 24164 35204
rect 22235 35173 22247 35176
rect 22189 35167 22247 35173
rect 21284 35108 22048 35136
rect 10042 35068 10048 35080
rect 9646 35040 10048 35068
rect 10042 35028 10048 35040
rect 10100 35028 10106 35080
rect 10137 35071 10195 35077
rect 10137 35037 10149 35071
rect 10183 35037 10195 35071
rect 10137 35031 10195 35037
rect 9858 35000 9864 35012
rect 7116 34972 9864 35000
rect 9858 34960 9864 34972
rect 9916 34960 9922 35012
rect 10152 35000 10180 35031
rect 11054 35028 11060 35080
rect 11112 35028 11118 35080
rect 11146 35028 11152 35080
rect 11204 35077 11210 35080
rect 11204 35071 11232 35077
rect 11220 35037 11232 35071
rect 11204 35031 11232 35037
rect 11204 35028 11210 35031
rect 11330 35028 11336 35080
rect 11388 35028 11394 35080
rect 12250 35068 12256 35080
rect 11900 35040 12256 35068
rect 9968 34972 10180 35000
rect 4522 34932 4528 34944
rect 4078 34904 4528 34932
rect 3973 34895 4031 34901
rect 4522 34892 4528 34904
rect 4580 34932 4586 34944
rect 4982 34932 4988 34944
rect 4580 34904 4988 34932
rect 4580 34892 4586 34904
rect 4982 34892 4988 34904
rect 5040 34892 5046 34944
rect 5074 34892 5080 34944
rect 5132 34892 5138 34944
rect 5166 34892 5172 34944
rect 5224 34932 5230 34944
rect 5261 34935 5319 34941
rect 5261 34932 5273 34935
rect 5224 34904 5273 34932
rect 5224 34892 5230 34904
rect 5261 34901 5273 34904
rect 5307 34901 5319 34935
rect 5261 34895 5319 34901
rect 5718 34892 5724 34944
rect 5776 34932 5782 34944
rect 6733 34935 6791 34941
rect 6733 34932 6745 34935
rect 5776 34904 6745 34932
rect 5776 34892 5782 34904
rect 6733 34901 6745 34904
rect 6779 34901 6791 34935
rect 6733 34895 6791 34901
rect 7558 34892 7564 34944
rect 7616 34932 7622 34944
rect 9490 34932 9496 34944
rect 7616 34904 9496 34932
rect 7616 34892 7622 34904
rect 9490 34892 9496 34904
rect 9548 34932 9554 34944
rect 9968 34932 9996 34972
rect 9548 34904 9996 34932
rect 9548 34892 9554 34904
rect 10042 34892 10048 34944
rect 10100 34932 10106 34944
rect 11900 34932 11928 35040
rect 12250 35028 12256 35040
rect 12308 35068 12314 35080
rect 12343 35071 12401 35077
rect 12343 35068 12355 35071
rect 12308 35040 12355 35068
rect 12308 35028 12314 35040
rect 12343 35037 12355 35040
rect 12389 35068 12401 35071
rect 17773 35071 17831 35077
rect 12389 35040 13492 35068
rect 12389 35037 12401 35040
rect 12343 35031 12401 35037
rect 13464 35012 13492 35040
rect 17773 35037 17785 35071
rect 17819 35037 17831 35071
rect 18046 35068 18052 35080
rect 18007 35040 18052 35068
rect 17773 35031 17831 35037
rect 12618 34960 12624 35012
rect 12676 35000 12682 35012
rect 12894 35000 12900 35012
rect 12676 34972 12900 35000
rect 12676 34960 12682 34972
rect 12894 34960 12900 34972
rect 12952 34960 12958 35012
rect 13446 34960 13452 35012
rect 13504 34960 13510 35012
rect 14182 34960 14188 35012
rect 14240 35000 14246 35012
rect 15470 35000 15476 35012
rect 14240 34972 15476 35000
rect 14240 34960 14246 34972
rect 15470 34960 15476 34972
rect 15528 34960 15534 35012
rect 17788 35000 17816 35031
rect 18046 35028 18052 35040
rect 18104 35028 18110 35080
rect 19150 35028 19156 35080
rect 19208 35068 19214 35080
rect 19245 35071 19303 35077
rect 19245 35068 19257 35071
rect 19208 35040 19257 35068
rect 19208 35028 19214 35040
rect 19245 35037 19257 35040
rect 19291 35037 19303 35071
rect 19352 35068 19380 35096
rect 19429 35071 19487 35077
rect 19429 35068 19441 35071
rect 19352 35040 19441 35068
rect 19245 35031 19303 35037
rect 19429 35037 19441 35040
rect 19475 35037 19487 35071
rect 19429 35031 19487 35037
rect 20257 35071 20315 35077
rect 20257 35037 20269 35071
rect 20303 35068 20315 35071
rect 20438 35068 20444 35080
rect 20303 35040 20444 35068
rect 20303 35037 20315 35040
rect 20257 35031 20315 35037
rect 20438 35028 20444 35040
rect 20496 35028 20502 35080
rect 20531 35071 20589 35077
rect 20531 35037 20543 35071
rect 20577 35068 20589 35071
rect 20622 35068 20628 35080
rect 20577 35040 20628 35068
rect 20577 35037 20589 35040
rect 20531 35031 20589 35037
rect 20622 35028 20628 35040
rect 20680 35028 20686 35080
rect 21284 35068 21312 35108
rect 22738 35096 22744 35148
rect 22796 35136 22802 35148
rect 22796 35108 23704 35136
rect 22796 35096 22802 35108
rect 20916 35040 21312 35068
rect 17788 34972 18000 35000
rect 10100 34904 11928 34932
rect 11977 34935 12035 34941
rect 10100 34892 10106 34904
rect 11977 34901 11989 34935
rect 12023 34932 12035 34935
rect 17862 34932 17868 34944
rect 12023 34904 17868 34932
rect 12023 34901 12035 34904
rect 11977 34895 12035 34901
rect 17862 34892 17868 34904
rect 17920 34892 17926 34944
rect 17972 34932 18000 34972
rect 18230 34960 18236 35012
rect 18288 35000 18294 35012
rect 20916 35000 20944 35040
rect 21450 35028 21456 35080
rect 21508 35068 21514 35080
rect 23676 35077 23704 35108
rect 22373 35071 22431 35077
rect 22373 35068 22385 35071
rect 21508 35040 22385 35068
rect 21508 35028 21514 35040
rect 22373 35037 22385 35040
rect 22419 35037 22431 35071
rect 22373 35031 22431 35037
rect 23385 35071 23443 35077
rect 23385 35037 23397 35071
rect 23431 35068 23443 35071
rect 23661 35071 23719 35077
rect 23431 35040 23520 35068
rect 23431 35037 23443 35040
rect 23385 35031 23443 35037
rect 18288 34972 20944 35000
rect 18288 34960 18294 34972
rect 21174 34960 21180 35012
rect 21232 35000 21238 35012
rect 21232 34972 23244 35000
rect 21232 34960 21238 34972
rect 23216 34944 23244 34972
rect 19702 34932 19708 34944
rect 17972 34904 19708 34932
rect 19702 34892 19708 34904
rect 19760 34932 19766 34944
rect 20438 34932 20444 34944
rect 19760 34904 20444 34932
rect 19760 34892 19766 34904
rect 20438 34892 20444 34904
rect 20496 34932 20502 34944
rect 22094 34932 22100 34944
rect 20496 34904 22100 34932
rect 20496 34892 20502 34904
rect 22094 34892 22100 34904
rect 22152 34892 22158 34944
rect 23198 34892 23204 34944
rect 23256 34892 23262 34944
rect 23492 34941 23520 35040
rect 23661 35037 23673 35071
rect 23707 35037 23719 35071
rect 23661 35031 23719 35037
rect 23566 34960 23572 35012
rect 23624 35000 23630 35012
rect 23845 35003 23903 35009
rect 23845 35000 23857 35003
rect 23624 34972 23857 35000
rect 23624 34960 23630 34972
rect 23845 34969 23857 34972
rect 23891 34969 23903 35003
rect 23845 34963 23903 34969
rect 24210 34960 24216 35012
rect 24268 34960 24274 35012
rect 23477 34935 23535 34941
rect 23477 34901 23489 34935
rect 23523 34901 23535 34935
rect 23477 34895 23535 34901
rect 1104 34842 25000 34864
rect 1104 34790 6884 34842
rect 6936 34790 6948 34842
rect 7000 34790 7012 34842
rect 7064 34790 7076 34842
rect 7128 34790 7140 34842
rect 7192 34790 12818 34842
rect 12870 34790 12882 34842
rect 12934 34790 12946 34842
rect 12998 34790 13010 34842
rect 13062 34790 13074 34842
rect 13126 34790 18752 34842
rect 18804 34790 18816 34842
rect 18868 34790 18880 34842
rect 18932 34790 18944 34842
rect 18996 34790 19008 34842
rect 19060 34790 24686 34842
rect 24738 34790 24750 34842
rect 24802 34790 24814 34842
rect 24866 34790 24878 34842
rect 24930 34790 24942 34842
rect 24994 34790 25000 34842
rect 1104 34768 25000 34790
rect 1762 34688 1768 34740
rect 1820 34688 1826 34740
rect 2501 34731 2559 34737
rect 2501 34697 2513 34731
rect 2547 34728 2559 34731
rect 2774 34728 2780 34740
rect 2547 34700 2780 34728
rect 2547 34697 2559 34700
rect 2501 34691 2559 34697
rect 2774 34688 2780 34700
rect 2832 34688 2838 34740
rect 3142 34688 3148 34740
rect 3200 34728 3206 34740
rect 3418 34728 3424 34740
rect 3200 34700 3424 34728
rect 3200 34688 3206 34700
rect 3418 34688 3424 34700
rect 3476 34688 3482 34740
rect 4154 34688 4160 34740
rect 4212 34728 4218 34740
rect 4249 34731 4307 34737
rect 4249 34728 4261 34731
rect 4212 34700 4261 34728
rect 4212 34688 4218 34700
rect 4249 34697 4261 34700
rect 4295 34697 4307 34731
rect 4249 34691 4307 34697
rect 4614 34688 4620 34740
rect 4672 34728 4678 34740
rect 4672 34700 5120 34728
rect 4672 34688 4678 34700
rect 1780 34601 1808 34688
rect 4062 34620 4068 34672
rect 4120 34660 4126 34672
rect 4798 34660 4804 34672
rect 4120 34632 4804 34660
rect 4120 34620 4126 34632
rect 4798 34620 4804 34632
rect 4856 34620 4862 34672
rect 5092 34669 5120 34700
rect 5718 34688 5724 34740
rect 5776 34688 5782 34740
rect 7377 34731 7435 34737
rect 7377 34728 7389 34731
rect 5828 34700 7389 34728
rect 5077 34663 5135 34669
rect 5077 34629 5089 34663
rect 5123 34629 5135 34663
rect 5077 34623 5135 34629
rect 5169 34663 5227 34669
rect 5169 34629 5181 34663
rect 5215 34660 5227 34663
rect 5736 34660 5764 34688
rect 5215 34632 5764 34660
rect 5215 34629 5227 34632
rect 5169 34623 5227 34629
rect 1763 34595 1821 34601
rect 1763 34561 1775 34595
rect 1809 34592 1821 34595
rect 3511 34595 3569 34601
rect 3511 34592 3523 34595
rect 1809 34564 3523 34592
rect 1809 34561 1821 34564
rect 1763 34555 1821 34561
rect 3511 34561 3523 34564
rect 3557 34592 3569 34595
rect 4338 34592 4344 34604
rect 3557 34564 4344 34592
rect 3557 34561 3569 34564
rect 3511 34555 3569 34561
rect 4338 34552 4344 34564
rect 4396 34552 4402 34604
rect 4522 34552 4528 34604
rect 4580 34592 4586 34604
rect 5350 34592 5356 34604
rect 4580 34564 5356 34592
rect 4580 34552 4586 34564
rect 5350 34552 5356 34564
rect 5408 34592 5414 34604
rect 5537 34595 5595 34601
rect 5537 34592 5549 34595
rect 5408 34564 5549 34592
rect 5408 34552 5414 34564
rect 5537 34561 5549 34564
rect 5583 34561 5595 34595
rect 5537 34555 5595 34561
rect 1486 34484 1492 34536
rect 1544 34484 1550 34536
rect 2866 34484 2872 34536
rect 2924 34524 2930 34536
rect 3050 34524 3056 34536
rect 2924 34496 3056 34524
rect 2924 34484 2930 34496
rect 3050 34484 3056 34496
rect 3108 34524 3114 34536
rect 3237 34527 3295 34533
rect 3237 34524 3249 34527
rect 3108 34496 3249 34524
rect 3108 34484 3114 34496
rect 3237 34493 3249 34496
rect 3283 34493 3295 34527
rect 5828 34510 5856 34700
rect 7377 34697 7389 34700
rect 7423 34697 7435 34731
rect 7377 34691 7435 34697
rect 8294 34688 8300 34740
rect 8352 34688 8358 34740
rect 8386 34688 8392 34740
rect 8444 34728 8450 34740
rect 9033 34731 9091 34737
rect 9033 34728 9045 34731
rect 8444 34700 9045 34728
rect 8444 34688 8450 34700
rect 9033 34697 9045 34700
rect 9079 34697 9091 34731
rect 9033 34691 9091 34697
rect 9858 34688 9864 34740
rect 9916 34728 9922 34740
rect 9916 34700 14410 34728
rect 9916 34688 9922 34700
rect 5905 34663 5963 34669
rect 5905 34629 5917 34663
rect 5951 34629 5963 34663
rect 6638 34631 6644 34672
rect 5905 34623 5963 34629
rect 6623 34625 6644 34631
rect 3237 34487 3295 34493
rect 5920 34456 5948 34623
rect 6178 34552 6184 34604
rect 6236 34592 6242 34604
rect 6365 34595 6423 34601
rect 6365 34592 6377 34595
rect 6236 34564 6377 34592
rect 6236 34552 6242 34564
rect 6365 34561 6377 34564
rect 6411 34561 6423 34595
rect 6623 34591 6635 34625
rect 6696 34620 6702 34672
rect 8018 34620 8024 34672
rect 8076 34620 8082 34672
rect 8312 34660 8340 34688
rect 11146 34660 11152 34672
rect 8312 34632 11152 34660
rect 11146 34620 11152 34632
rect 11204 34620 11210 34672
rect 14382 34660 14410 34700
rect 15470 34688 15476 34740
rect 15528 34728 15534 34740
rect 16666 34728 16672 34740
rect 15528 34700 16672 34728
rect 15528 34688 15534 34700
rect 16666 34688 16672 34700
rect 16724 34688 16730 34740
rect 17402 34728 17408 34740
rect 16868 34700 17408 34728
rect 16114 34660 16120 34672
rect 14382 34632 16120 34660
rect 14382 34631 14410 34632
rect 14351 34625 14410 34631
rect 6669 34594 6682 34620
rect 6669 34591 6681 34594
rect 6623 34585 6681 34591
rect 6365 34555 6423 34561
rect 5920 34428 6224 34456
rect 6196 34400 6224 34428
rect 1762 34348 1768 34400
rect 1820 34388 1826 34400
rect 2406 34388 2412 34400
rect 1820 34360 2412 34388
rect 1820 34348 1826 34360
rect 2406 34348 2412 34360
rect 2464 34348 2470 34400
rect 6086 34348 6092 34400
rect 6144 34348 6150 34400
rect 6178 34348 6184 34400
rect 6236 34348 6242 34400
rect 6380 34388 6408 34555
rect 7742 34552 7748 34604
rect 7800 34552 7806 34604
rect 8036 34592 8064 34620
rect 8263 34595 8321 34601
rect 8263 34592 8275 34595
rect 8036 34564 8275 34592
rect 8263 34561 8275 34564
rect 8309 34561 8321 34595
rect 8263 34555 8321 34561
rect 10594 34552 10600 34604
rect 10652 34592 10658 34604
rect 11054 34592 11060 34604
rect 10652 34564 11060 34592
rect 10652 34552 10658 34564
rect 11054 34552 11060 34564
rect 11112 34552 11118 34604
rect 14351 34591 14363 34625
rect 14397 34594 14410 34625
rect 16114 34620 16120 34632
rect 16172 34620 16178 34672
rect 16868 34660 16896 34700
rect 17402 34688 17408 34700
rect 17460 34728 17466 34740
rect 17681 34731 17739 34737
rect 17681 34728 17693 34731
rect 17460 34700 17693 34728
rect 17460 34688 17466 34700
rect 17681 34697 17693 34700
rect 17727 34697 17739 34731
rect 17681 34691 17739 34697
rect 20625 34731 20683 34737
rect 20625 34697 20637 34731
rect 20671 34697 20683 34731
rect 20625 34691 20683 34697
rect 16224 34632 16896 34660
rect 16224 34601 16252 34632
rect 17218 34620 17224 34672
rect 17276 34660 17282 34672
rect 19334 34660 19340 34672
rect 17276 34632 19340 34660
rect 17276 34620 17282 34632
rect 19334 34620 19340 34632
rect 19392 34620 19398 34672
rect 20640 34660 20668 34691
rect 21450 34688 21456 34740
rect 21508 34688 21514 34740
rect 21821 34731 21879 34737
rect 21821 34697 21833 34731
rect 21867 34728 21879 34731
rect 22741 34731 22799 34737
rect 21867 34700 22692 34728
rect 21867 34697 21879 34700
rect 21821 34691 21879 34697
rect 20640 34632 21680 34660
rect 16943 34605 17001 34611
rect 16209 34595 16267 34601
rect 14397 34591 14409 34594
rect 14351 34585 14409 34591
rect 16209 34561 16221 34595
rect 16255 34561 16267 34595
rect 16209 34555 16267 34561
rect 16666 34552 16672 34604
rect 16724 34552 16730 34604
rect 16943 34571 16955 34605
rect 16989 34598 17001 34605
rect 16989 34592 17172 34598
rect 17236 34592 17264 34620
rect 16989 34571 17264 34592
rect 16943 34570 17264 34571
rect 16943 34565 17001 34570
rect 17144 34564 17264 34570
rect 17862 34552 17868 34604
rect 17920 34592 17926 34604
rect 20162 34592 20168 34604
rect 17920 34564 20168 34592
rect 17920 34552 17926 34564
rect 20162 34552 20168 34564
rect 20220 34592 20226 34604
rect 21652 34601 21680 34632
rect 22664 34601 22692 34700
rect 22741 34697 22753 34731
rect 22787 34697 22799 34731
rect 22741 34691 22799 34697
rect 23293 34731 23351 34737
rect 23293 34697 23305 34731
rect 23339 34728 23351 34731
rect 23566 34728 23572 34740
rect 23339 34700 23572 34728
rect 23339 34697 23351 34700
rect 23293 34691 23351 34697
rect 22756 34660 22784 34691
rect 23566 34688 23572 34700
rect 23624 34688 23630 34740
rect 23661 34731 23719 34737
rect 23661 34697 23673 34731
rect 23707 34697 23719 34731
rect 23661 34691 23719 34697
rect 23676 34660 23704 34691
rect 24121 34663 24179 34669
rect 24121 34660 24133 34663
rect 22756 34632 23612 34660
rect 23676 34632 24133 34660
rect 20809 34595 20867 34601
rect 20809 34592 20821 34595
rect 20220 34564 20821 34592
rect 20220 34552 20226 34564
rect 20809 34561 20821 34564
rect 20855 34561 20867 34595
rect 20809 34555 20867 34561
rect 21637 34595 21695 34601
rect 21637 34561 21649 34595
rect 21683 34561 21695 34595
rect 21637 34555 21695 34561
rect 22005 34595 22063 34601
rect 22005 34561 22017 34595
rect 22051 34561 22063 34595
rect 22005 34555 22063 34561
rect 22649 34595 22707 34601
rect 22649 34561 22661 34595
rect 22695 34561 22707 34595
rect 22649 34555 22707 34561
rect 22925 34595 22983 34601
rect 22925 34561 22937 34595
rect 22971 34592 22983 34595
rect 23014 34592 23020 34604
rect 22971 34564 23020 34592
rect 22971 34561 22983 34564
rect 22925 34555 22983 34561
rect 7760 34524 7788 34552
rect 8021 34527 8079 34533
rect 8021 34524 8033 34527
rect 7760 34496 8033 34524
rect 8021 34493 8033 34496
rect 8067 34493 8079 34527
rect 8021 34487 8079 34493
rect 8938 34484 8944 34536
rect 8996 34524 9002 34536
rect 10410 34524 10416 34536
rect 8996 34496 10416 34524
rect 8996 34484 9002 34496
rect 10410 34484 10416 34496
rect 10468 34484 10474 34536
rect 14090 34484 14096 34536
rect 14148 34484 14154 34536
rect 16390 34484 16396 34536
rect 16448 34484 16454 34536
rect 16485 34527 16543 34533
rect 16485 34493 16497 34527
rect 16531 34524 16543 34527
rect 16531 34496 16620 34524
rect 16531 34493 16543 34496
rect 16485 34487 16543 34493
rect 9122 34416 9128 34468
rect 9180 34456 9186 34468
rect 9582 34456 9588 34468
rect 9180 34428 9588 34456
rect 9180 34416 9186 34428
rect 9582 34416 9588 34428
rect 9640 34416 9646 34468
rect 6822 34388 6828 34400
rect 6380 34360 6828 34388
rect 6822 34348 6828 34360
rect 6880 34348 6886 34400
rect 15102 34348 15108 34400
rect 15160 34348 15166 34400
rect 16298 34348 16304 34400
rect 16356 34348 16362 34400
rect 16408 34397 16436 34484
rect 16393 34391 16451 34397
rect 16393 34357 16405 34391
rect 16439 34357 16451 34391
rect 16592 34388 16620 34496
rect 19426 34484 19432 34536
rect 19484 34524 19490 34536
rect 22020 34524 22048 34555
rect 23014 34552 23020 34564
rect 23072 34552 23078 34604
rect 23198 34552 23204 34604
rect 23256 34552 23262 34604
rect 23477 34595 23535 34601
rect 23477 34561 23489 34595
rect 23523 34561 23535 34595
rect 23584 34592 23612 34632
rect 24121 34629 24133 34632
rect 24167 34629 24179 34663
rect 24121 34623 24179 34629
rect 23845 34595 23903 34601
rect 23845 34592 23857 34595
rect 23584 34564 23857 34592
rect 23477 34555 23535 34561
rect 23845 34561 23857 34564
rect 23891 34561 23903 34595
rect 23845 34555 23903 34561
rect 23492 34524 23520 34555
rect 19484 34496 20116 34524
rect 19484 34484 19490 34496
rect 20088 34456 20116 34496
rect 20916 34496 22048 34524
rect 22480 34496 23520 34524
rect 20916 34456 20944 34496
rect 22480 34465 22508 34496
rect 24394 34484 24400 34536
rect 24452 34484 24458 34536
rect 20088 34428 20944 34456
rect 22465 34459 22523 34465
rect 22465 34425 22477 34459
rect 22511 34425 22523 34459
rect 22465 34419 22523 34425
rect 23014 34416 23020 34468
rect 23072 34416 23078 34468
rect 23382 34416 23388 34468
rect 23440 34456 23446 34468
rect 25590 34456 25596 34468
rect 23440 34428 25596 34456
rect 23440 34416 23446 34428
rect 25590 34416 25596 34428
rect 25648 34416 25654 34468
rect 17494 34388 17500 34400
rect 16592 34360 17500 34388
rect 16393 34351 16451 34357
rect 17494 34348 17500 34360
rect 17552 34348 17558 34400
rect 20254 34348 20260 34400
rect 20312 34388 20318 34400
rect 25498 34388 25504 34400
rect 20312 34360 25504 34388
rect 20312 34348 20318 34360
rect 25498 34348 25504 34360
rect 25556 34348 25562 34400
rect 1104 34298 24840 34320
rect 1104 34246 3917 34298
rect 3969 34246 3981 34298
rect 4033 34246 4045 34298
rect 4097 34246 4109 34298
rect 4161 34246 4173 34298
rect 4225 34246 9851 34298
rect 9903 34246 9915 34298
rect 9967 34246 9979 34298
rect 10031 34246 10043 34298
rect 10095 34246 10107 34298
rect 10159 34246 15785 34298
rect 15837 34246 15849 34298
rect 15901 34246 15913 34298
rect 15965 34246 15977 34298
rect 16029 34246 16041 34298
rect 16093 34246 21719 34298
rect 21771 34246 21783 34298
rect 21835 34246 21847 34298
rect 21899 34246 21911 34298
rect 21963 34246 21975 34298
rect 22027 34246 24840 34298
rect 1104 34224 24840 34246
rect 2222 34144 2228 34196
rect 2280 34184 2286 34196
rect 2409 34187 2467 34193
rect 2409 34184 2421 34187
rect 2280 34156 2421 34184
rect 2280 34144 2286 34156
rect 2409 34153 2421 34156
rect 2455 34153 2467 34187
rect 2409 34147 2467 34153
rect 2682 34144 2688 34196
rect 2740 34184 2746 34196
rect 4614 34184 4620 34196
rect 2740 34156 4620 34184
rect 2740 34144 2746 34156
rect 4614 34144 4620 34156
rect 4672 34144 4678 34196
rect 9214 34184 9220 34196
rect 5644 34156 9220 34184
rect 1397 33983 1455 33989
rect 1397 33949 1409 33983
rect 1443 33980 1455 33983
rect 1671 33983 1729 33989
rect 1443 33952 1532 33980
rect 1443 33949 1455 33952
rect 1397 33943 1455 33949
rect 1504 33856 1532 33952
rect 1671 33949 1683 33983
rect 1717 33980 1729 33983
rect 2700 33980 2728 34144
rect 3602 34076 3608 34128
rect 3660 34116 3666 34128
rect 5644 34116 5672 34156
rect 9214 34144 9220 34156
rect 9272 34144 9278 34196
rect 9582 34144 9588 34196
rect 9640 34184 9646 34196
rect 10321 34187 10379 34193
rect 10321 34184 10333 34187
rect 9640 34156 10333 34184
rect 9640 34144 9646 34156
rect 10321 34153 10333 34156
rect 10367 34153 10379 34187
rect 10321 34147 10379 34153
rect 10502 34144 10508 34196
rect 10560 34144 10566 34196
rect 14090 34144 14096 34196
rect 14148 34184 14154 34196
rect 14148 34156 16160 34184
rect 14148 34144 14154 34156
rect 3660 34088 4568 34116
rect 3660 34076 3666 34088
rect 3053 34051 3111 34057
rect 3053 34017 3065 34051
rect 3099 34048 3111 34051
rect 3099 34020 4476 34048
rect 3099 34017 3111 34020
rect 3053 34011 3111 34017
rect 1717 33952 2728 33980
rect 1717 33949 1729 33952
rect 1671 33943 1729 33949
rect 2774 33940 2780 33992
rect 2832 33940 2838 33992
rect 3786 33940 3792 33992
rect 3844 33940 3850 33992
rect 3878 33940 3884 33992
rect 3936 33980 3942 33992
rect 4341 33983 4399 33989
rect 4341 33980 4353 33983
rect 3936 33952 4353 33980
rect 3936 33940 3942 33952
rect 4341 33949 4353 33952
rect 4387 33949 4399 33983
rect 4341 33943 4399 33949
rect 2314 33872 2320 33924
rect 2372 33912 2378 33924
rect 2498 33912 2504 33924
rect 2372 33884 2504 33912
rect 2372 33872 2378 33884
rect 2498 33872 2504 33884
rect 2556 33872 2562 33924
rect 4065 33915 4123 33921
rect 4065 33881 4077 33915
rect 4111 33912 4123 33915
rect 4246 33912 4252 33924
rect 4111 33884 4252 33912
rect 4111 33881 4123 33884
rect 4065 33875 4123 33881
rect 4246 33872 4252 33884
rect 4304 33872 4310 33924
rect 4448 33912 4476 34020
rect 4540 33980 4568 34088
rect 4632 34088 5672 34116
rect 4632 34057 4660 34088
rect 9122 34076 9128 34128
rect 9180 34076 9186 34128
rect 9401 34119 9459 34125
rect 9401 34085 9413 34119
rect 9447 34116 9459 34119
rect 10520 34116 10548 34144
rect 9447 34088 10548 34116
rect 9447 34085 9459 34088
rect 9401 34079 9459 34085
rect 4617 34051 4675 34057
rect 4617 34017 4629 34051
rect 4663 34017 4675 34051
rect 4617 34011 4675 34017
rect 6822 34008 6828 34060
rect 6880 34048 6886 34060
rect 7009 34051 7067 34057
rect 7009 34048 7021 34051
rect 6880 34020 7021 34048
rect 6880 34008 6886 34020
rect 7009 34017 7021 34020
rect 7055 34017 7067 34051
rect 9140 34048 9168 34076
rect 9309 34051 9367 34057
rect 9309 34048 9321 34051
rect 9140 34020 9321 34048
rect 7009 34011 7067 34017
rect 9309 34017 9321 34020
rect 9355 34017 9367 34051
rect 9309 34011 9367 34017
rect 9493 34051 9551 34057
rect 9493 34017 9505 34051
rect 9539 34048 9551 34051
rect 10045 34051 10103 34057
rect 10045 34048 10057 34051
rect 9539 34020 10057 34048
rect 9539 34017 9551 34020
rect 9493 34011 9551 34017
rect 10045 34017 10057 34020
rect 10091 34017 10103 34051
rect 10045 34011 10103 34017
rect 11882 34008 11888 34060
rect 11940 34048 11946 34060
rect 14108 34057 14136 34144
rect 16132 34116 16160 34156
rect 16298 34144 16304 34196
rect 16356 34184 16362 34196
rect 17221 34187 17279 34193
rect 17221 34184 17233 34187
rect 16356 34156 17233 34184
rect 16356 34144 16362 34156
rect 17221 34153 17233 34156
rect 17267 34153 17279 34187
rect 17221 34147 17279 34153
rect 17494 34144 17500 34196
rect 17552 34144 17558 34196
rect 22094 34184 22100 34196
rect 17604 34156 22100 34184
rect 17604 34116 17632 34156
rect 22094 34144 22100 34156
rect 22152 34144 22158 34196
rect 23845 34187 23903 34193
rect 23845 34153 23857 34187
rect 23891 34184 23903 34187
rect 24486 34184 24492 34196
rect 23891 34156 24492 34184
rect 23891 34153 23903 34156
rect 23845 34147 23903 34153
rect 24486 34144 24492 34156
rect 24544 34144 24550 34196
rect 16132 34088 17632 34116
rect 21453 34119 21511 34125
rect 21453 34085 21465 34119
rect 21499 34085 21511 34119
rect 21453 34079 21511 34085
rect 22465 34119 22523 34125
rect 22465 34085 22477 34119
rect 22511 34116 22523 34119
rect 22511 34088 23244 34116
rect 22511 34085 22523 34088
rect 22465 34079 22523 34085
rect 12161 34051 12219 34057
rect 12161 34048 12173 34051
rect 11940 34020 12173 34048
rect 11940 34008 11946 34020
rect 12161 34017 12173 34020
rect 12207 34017 12219 34051
rect 12161 34011 12219 34017
rect 14093 34051 14151 34057
rect 14093 34017 14105 34051
rect 14139 34017 14151 34051
rect 14093 34011 14151 34017
rect 15470 34008 15476 34060
rect 15528 34008 15534 34060
rect 21468 34048 21496 34079
rect 21468 34020 22692 34048
rect 5258 33980 5264 33992
rect 4540 33952 5264 33980
rect 5258 33940 5264 33952
rect 5316 33980 5322 33992
rect 5537 33983 5595 33989
rect 5537 33980 5549 33983
rect 5316 33952 5549 33980
rect 5316 33940 5322 33952
rect 5537 33949 5549 33952
rect 5583 33949 5595 33983
rect 5537 33943 5595 33949
rect 5718 33940 5724 33992
rect 5776 33980 5782 33992
rect 5811 33983 5869 33989
rect 5811 33980 5823 33983
rect 5776 33952 5823 33980
rect 5776 33940 5782 33952
rect 5811 33949 5823 33952
rect 5857 33980 5869 33983
rect 5902 33980 5908 33992
rect 5857 33952 5908 33980
rect 5857 33949 5869 33952
rect 5811 33943 5869 33949
rect 5902 33940 5908 33952
rect 5960 33940 5966 33992
rect 6012 33979 7326 33980
rect 6012 33973 7341 33979
rect 6012 33952 7295 33973
rect 6012 33912 6040 33952
rect 7283 33939 7295 33952
rect 7329 33939 7341 33973
rect 9122 33940 9128 33992
rect 9180 33980 9186 33992
rect 9217 33983 9275 33989
rect 9217 33980 9229 33983
rect 9180 33952 9229 33980
rect 9180 33940 9186 33952
rect 9217 33949 9229 33952
rect 9263 33949 9275 33983
rect 9217 33943 9275 33949
rect 9769 33983 9827 33989
rect 9769 33949 9781 33983
rect 9815 33949 9827 33983
rect 9769 33943 9827 33949
rect 9953 33983 10011 33989
rect 9953 33949 9965 33983
rect 9999 33949 10011 33983
rect 9953 33943 10011 33949
rect 7283 33933 7341 33939
rect 4448 33884 6040 33912
rect 6086 33872 6092 33924
rect 6144 33872 6150 33924
rect 1486 33804 1492 33856
rect 1544 33804 1550 33856
rect 1946 33804 1952 33856
rect 2004 33844 2010 33856
rect 2222 33844 2228 33856
rect 2004 33816 2228 33844
rect 2004 33804 2010 33816
rect 2222 33804 2228 33816
rect 2280 33804 2286 33856
rect 2682 33804 2688 33856
rect 2740 33844 2746 33856
rect 6104 33844 6132 33872
rect 2740 33816 6132 33844
rect 2740 33804 2746 33816
rect 6546 33804 6552 33856
rect 6604 33804 6610 33856
rect 7298 33844 7326 33933
rect 7374 33844 7380 33856
rect 7298 33816 7380 33844
rect 7374 33804 7380 33816
rect 7432 33804 7438 33856
rect 8021 33847 8079 33853
rect 8021 33813 8033 33847
rect 8067 33844 8079 33847
rect 8110 33844 8116 33856
rect 8067 33816 8116 33844
rect 8067 33813 8079 33816
rect 8021 33807 8079 33813
rect 8110 33804 8116 33816
rect 8168 33804 8174 33856
rect 9398 33804 9404 33856
rect 9456 33844 9462 33856
rect 9585 33847 9643 33853
rect 9585 33844 9597 33847
rect 9456 33816 9597 33844
rect 9456 33804 9462 33816
rect 9585 33813 9597 33816
rect 9631 33813 9643 33847
rect 9585 33807 9643 33813
rect 9674 33804 9680 33856
rect 9732 33844 9738 33856
rect 9784 33844 9812 33943
rect 9732 33816 9812 33844
rect 9974 33844 10002 33943
rect 10134 33940 10140 33992
rect 10192 33940 10198 33992
rect 10229 33983 10287 33989
rect 10229 33949 10241 33983
rect 10275 33949 10287 33983
rect 10229 33943 10287 33949
rect 12435 33983 12493 33989
rect 12435 33949 12447 33983
rect 12481 33980 12493 33983
rect 13722 33980 13728 33992
rect 12481 33952 13728 33980
rect 12481 33949 12493 33952
rect 12435 33943 12493 33949
rect 10042 33872 10048 33924
rect 10100 33912 10106 33924
rect 10244 33912 10272 33943
rect 13722 33940 13728 33952
rect 13780 33940 13786 33992
rect 14367 33983 14425 33989
rect 14367 33980 14379 33983
rect 13832 33952 14379 33980
rect 10100 33884 10272 33912
rect 10100 33872 10106 33884
rect 11330 33872 11336 33924
rect 11388 33912 11394 33924
rect 13832 33912 13860 33952
rect 14367 33949 14379 33952
rect 14413 33980 14425 33983
rect 15378 33980 15384 33992
rect 14413 33952 15384 33980
rect 14413 33949 14425 33952
rect 14367 33943 14425 33949
rect 15378 33940 15384 33952
rect 15436 33940 15442 33992
rect 15715 33983 15773 33989
rect 15715 33980 15727 33983
rect 15470 33952 15727 33980
rect 11388 33884 13860 33912
rect 11388 33872 11394 33884
rect 14918 33872 14924 33924
rect 14976 33912 14982 33924
rect 15470 33912 15498 33952
rect 15715 33949 15727 33952
rect 15761 33980 15773 33983
rect 15761 33949 15774 33980
rect 15715 33943 15774 33949
rect 14976 33884 15498 33912
rect 15746 33912 15774 33943
rect 17126 33940 17132 33992
rect 17184 33940 17190 33992
rect 17402 33989 17408 33992
rect 17395 33983 17408 33989
rect 17395 33980 17407 33983
rect 17363 33952 17407 33980
rect 17395 33949 17407 33952
rect 17395 33943 17408 33949
rect 17402 33940 17408 33943
rect 17460 33940 17466 33992
rect 17586 33940 17592 33992
rect 17644 33940 17650 33992
rect 19334 33940 19340 33992
rect 19392 33980 19398 33992
rect 20254 33980 20260 33992
rect 19392 33952 20260 33980
rect 19392 33940 19398 33952
rect 20254 33940 20260 33952
rect 20312 33980 20318 33992
rect 20312 33952 21312 33980
rect 20312 33940 20318 33952
rect 21174 33912 21180 33924
rect 15746 33884 21180 33912
rect 14976 33872 14982 33884
rect 21174 33872 21180 33884
rect 21232 33872 21238 33924
rect 21284 33912 21312 33952
rect 21358 33940 21364 33992
rect 21416 33980 21422 33992
rect 22664 33989 22692 34020
rect 23216 33989 23244 34088
rect 21637 33983 21695 33989
rect 21637 33980 21649 33983
rect 21416 33952 21649 33980
rect 21416 33940 21422 33952
rect 21637 33949 21649 33952
rect 21683 33949 21695 33983
rect 22373 33983 22431 33989
rect 22373 33980 22385 33983
rect 21637 33943 21695 33949
rect 22066 33952 22385 33980
rect 22066 33912 22094 33952
rect 22373 33949 22385 33952
rect 22419 33949 22431 33983
rect 22373 33943 22431 33949
rect 22649 33983 22707 33989
rect 22649 33949 22661 33983
rect 22695 33949 22707 33983
rect 22649 33943 22707 33949
rect 23201 33983 23259 33989
rect 23201 33949 23213 33983
rect 23247 33949 23259 33983
rect 23201 33943 23259 33949
rect 23290 33940 23296 33992
rect 23348 33980 23354 33992
rect 23569 33983 23627 33989
rect 23569 33980 23581 33983
rect 23348 33952 23581 33980
rect 23348 33940 23354 33952
rect 23569 33949 23581 33952
rect 23615 33949 23627 33983
rect 23569 33943 23627 33949
rect 23658 33940 23664 33992
rect 23716 33940 23722 33992
rect 23937 33983 23995 33989
rect 23937 33949 23949 33983
rect 23983 33949 23995 33983
rect 23937 33943 23995 33949
rect 23952 33912 23980 33943
rect 21284 33884 22094 33912
rect 23032 33884 23980 33912
rect 10502 33844 10508 33856
rect 9974 33816 10508 33844
rect 9732 33804 9738 33816
rect 10502 33804 10508 33816
rect 10560 33804 10566 33856
rect 13170 33804 13176 33856
rect 13228 33804 13234 33856
rect 14642 33804 14648 33856
rect 14700 33844 14706 33856
rect 15105 33847 15163 33853
rect 15105 33844 15117 33847
rect 14700 33816 15117 33844
rect 14700 33804 14706 33816
rect 15105 33813 15117 33816
rect 15151 33813 15163 33847
rect 15105 33807 15163 33813
rect 16482 33804 16488 33856
rect 16540 33804 16546 33856
rect 22186 33804 22192 33856
rect 22244 33804 22250 33856
rect 23032 33853 23060 33884
rect 23017 33847 23075 33853
rect 23017 33813 23029 33847
rect 23063 33813 23075 33847
rect 23017 33807 23075 33813
rect 23382 33804 23388 33856
rect 23440 33804 23446 33856
rect 24118 33804 24124 33856
rect 24176 33804 24182 33856
rect 1104 33754 25000 33776
rect 14 33668 20 33720
rect 72 33668 78 33720
rect 1104 33702 6884 33754
rect 6936 33702 6948 33754
rect 7000 33702 7012 33754
rect 7064 33702 7076 33754
rect 7128 33702 7140 33754
rect 7192 33702 12818 33754
rect 12870 33702 12882 33754
rect 12934 33702 12946 33754
rect 12998 33702 13010 33754
rect 13062 33702 13074 33754
rect 13126 33702 18752 33754
rect 18804 33702 18816 33754
rect 18868 33702 18880 33754
rect 18932 33702 18944 33754
rect 18996 33702 19008 33754
rect 19060 33702 24686 33754
rect 24738 33702 24750 33754
rect 24802 33702 24814 33754
rect 24866 33702 24878 33754
rect 24930 33702 24942 33754
rect 24994 33702 25000 33754
rect 1104 33680 25000 33702
rect 32 33640 60 33668
rect 5718 33640 5724 33652
rect 32 33612 5724 33640
rect 5718 33600 5724 33612
rect 5776 33640 5782 33652
rect 7650 33640 7656 33652
rect 5776 33612 7656 33640
rect 5776 33600 5782 33612
rect 7650 33600 7656 33612
rect 7708 33600 7714 33652
rect 9401 33643 9459 33649
rect 7760 33612 9352 33640
rect 106 33532 112 33584
rect 164 33572 170 33584
rect 2682 33572 2688 33584
rect 164 33544 2688 33572
rect 164 33532 170 33544
rect 2682 33532 2688 33544
rect 2740 33532 2746 33584
rect 2777 33575 2835 33581
rect 2777 33541 2789 33575
rect 2823 33572 2835 33575
rect 6730 33572 6736 33584
rect 2823 33544 6736 33572
rect 2823 33541 2835 33544
rect 2777 33535 2835 33541
rect 842 33464 848 33516
rect 900 33504 906 33516
rect 1118 33504 1124 33516
rect 900 33476 1124 33504
rect 900 33464 906 33476
rect 1118 33464 1124 33476
rect 1176 33464 1182 33516
rect 1394 33464 1400 33516
rect 1452 33464 1458 33516
rect 1670 33464 1676 33516
rect 1728 33464 1734 33516
rect 1946 33464 1952 33516
rect 2004 33464 2010 33516
rect 2498 33464 2504 33516
rect 2556 33464 2562 33516
rect 3387 33507 3445 33513
rect 3387 33504 3399 33507
rect 3068 33476 3399 33504
rect 1688 33368 1716 33464
rect 2225 33439 2283 33445
rect 2225 33405 2237 33439
rect 2271 33436 2283 33439
rect 2590 33436 2596 33448
rect 2271 33408 2596 33436
rect 2271 33405 2283 33408
rect 2225 33399 2283 33405
rect 2590 33396 2596 33408
rect 2648 33396 2654 33448
rect 3068 33380 3096 33476
rect 3387 33473 3399 33476
rect 3433 33473 3445 33507
rect 3387 33467 3445 33473
rect 4338 33464 4344 33516
rect 4396 33504 4402 33516
rect 5350 33504 5356 33516
rect 4396 33476 5356 33504
rect 4396 33464 4402 33476
rect 5350 33464 5356 33476
rect 5408 33464 5414 33516
rect 6288 33448 6316 33544
rect 6730 33532 6736 33544
rect 6788 33532 6794 33584
rect 7760 33572 7788 33612
rect 6840 33544 7788 33572
rect 6840 33516 6868 33544
rect 6822 33464 6828 33516
rect 6880 33464 6886 33516
rect 8662 33513 8668 33516
rect 7561 33507 7619 33513
rect 7561 33473 7573 33507
rect 7607 33504 7619 33507
rect 8619 33507 8668 33513
rect 7607 33476 7972 33504
rect 7607 33473 7619 33476
rect 7561 33467 7619 33473
rect 7944 33448 7972 33476
rect 8619 33473 8631 33507
rect 8665 33473 8668 33507
rect 8619 33467 8668 33473
rect 8662 33464 8668 33467
rect 8720 33464 8726 33516
rect 8754 33464 8760 33516
rect 8812 33464 8818 33516
rect 3145 33439 3203 33445
rect 3145 33405 3157 33439
rect 3191 33405 3203 33439
rect 3145 33399 3203 33405
rect 3050 33368 3056 33380
rect 1688 33340 3056 33368
rect 3050 33328 3056 33340
rect 3108 33328 3114 33380
rect 2866 33260 2872 33312
rect 2924 33300 2930 33312
rect 3160 33300 3188 33399
rect 4982 33396 4988 33448
rect 5040 33436 5046 33448
rect 6178 33436 6184 33448
rect 5040 33408 6184 33436
rect 5040 33396 5046 33408
rect 6178 33396 6184 33408
rect 6236 33396 6242 33448
rect 6270 33396 6276 33448
rect 6328 33396 6334 33448
rect 7745 33439 7803 33445
rect 7745 33405 7757 33439
rect 7791 33405 7803 33439
rect 7745 33399 7803 33405
rect 4798 33328 4804 33380
rect 4856 33368 4862 33380
rect 5626 33368 5632 33380
rect 4856 33340 5632 33368
rect 4856 33328 4862 33340
rect 5626 33328 5632 33340
rect 5684 33328 5690 33380
rect 7760 33368 7788 33399
rect 7926 33396 7932 33448
rect 7984 33396 7990 33448
rect 8110 33396 8116 33448
rect 8168 33436 8174 33448
rect 8205 33439 8263 33445
rect 8205 33436 8217 33439
rect 8168 33408 8217 33436
rect 8168 33396 8174 33408
rect 8205 33405 8217 33408
rect 8251 33405 8263 33439
rect 8481 33439 8539 33445
rect 8481 33436 8493 33439
rect 8205 33399 8263 33405
rect 8312 33408 8493 33436
rect 7760 33340 8248 33368
rect 8220 33312 8248 33340
rect 2924 33272 3188 33300
rect 2924 33260 2930 33272
rect 3878 33260 3884 33312
rect 3936 33300 3942 33312
rect 4157 33303 4215 33309
rect 4157 33300 4169 33303
rect 3936 33272 4169 33300
rect 3936 33260 3942 33272
rect 4157 33269 4169 33272
rect 4203 33269 4215 33303
rect 4157 33263 4215 33269
rect 4246 33260 4252 33312
rect 4304 33300 4310 33312
rect 4709 33303 4767 33309
rect 4709 33300 4721 33303
rect 4304 33272 4721 33300
rect 4304 33260 4310 33272
rect 4709 33269 4721 33272
rect 4755 33269 4767 33303
rect 4709 33263 4767 33269
rect 5810 33260 5816 33312
rect 5868 33300 5874 33312
rect 6086 33300 6092 33312
rect 5868 33272 6092 33300
rect 5868 33260 5874 33272
rect 6086 33260 6092 33272
rect 6144 33260 6150 33312
rect 8202 33260 8208 33312
rect 8260 33260 8266 33312
rect 8312 33300 8340 33408
rect 8481 33405 8493 33408
rect 8527 33405 8539 33439
rect 9324 33436 9352 33612
rect 9401 33609 9413 33643
rect 9447 33640 9459 33643
rect 9582 33640 9588 33652
rect 9447 33612 9588 33640
rect 9447 33609 9459 33612
rect 9401 33603 9459 33609
rect 9582 33600 9588 33612
rect 9640 33600 9646 33652
rect 10134 33640 10140 33652
rect 9690 33612 10140 33640
rect 9398 33464 9404 33516
rect 9456 33504 9462 33516
rect 9690 33504 9718 33612
rect 10134 33600 10140 33612
rect 10192 33600 10198 33652
rect 10502 33600 10508 33652
rect 10560 33600 10566 33652
rect 12342 33640 12348 33652
rect 11808 33612 12348 33640
rect 10318 33572 10324 33584
rect 10158 33544 10324 33572
rect 9456 33476 9718 33504
rect 9751 33507 9809 33513
rect 9456 33464 9462 33476
rect 9751 33473 9763 33507
rect 9797 33502 9809 33507
rect 10158 33504 10186 33544
rect 10318 33532 10324 33544
rect 10376 33572 10382 33584
rect 10962 33572 10968 33584
rect 10376 33544 10968 33572
rect 10376 33532 10382 33544
rect 10962 33532 10968 33544
rect 11020 33532 11026 33584
rect 11808 33513 11836 33612
rect 12342 33600 12348 33612
rect 12400 33600 12406 33652
rect 12710 33600 12716 33652
rect 12768 33640 12774 33652
rect 13722 33640 13728 33652
rect 12768 33612 13728 33640
rect 12768 33600 12774 33612
rect 13722 33600 13728 33612
rect 13780 33600 13786 33652
rect 14826 33600 14832 33652
rect 14884 33640 14890 33652
rect 15749 33643 15807 33649
rect 15749 33640 15761 33643
rect 14884 33612 15761 33640
rect 14884 33600 14890 33612
rect 15749 33609 15761 33612
rect 15795 33609 15807 33643
rect 15749 33603 15807 33609
rect 17129 33643 17187 33649
rect 17129 33609 17141 33643
rect 17175 33640 17187 33643
rect 17586 33640 17592 33652
rect 17175 33612 17592 33640
rect 17175 33609 17187 33612
rect 17129 33603 17187 33609
rect 17586 33600 17592 33612
rect 17644 33600 17650 33652
rect 19705 33643 19763 33649
rect 19705 33609 19717 33643
rect 19751 33640 19763 33643
rect 19751 33612 20208 33640
rect 19751 33609 19763 33612
rect 19705 33603 19763 33609
rect 16850 33532 16856 33584
rect 16908 33572 16914 33584
rect 17402 33572 17408 33584
rect 16908 33544 17408 33572
rect 16908 33532 16914 33544
rect 17402 33532 17408 33544
rect 17460 33532 17466 33584
rect 19518 33572 19524 33584
rect 17604 33544 19524 33572
rect 11793 33507 11851 33513
rect 11793 33504 11805 33507
rect 9864 33502 10186 33504
rect 9797 33476 10186 33502
rect 10244 33476 11805 33504
rect 9797 33474 9892 33476
rect 9797 33473 9809 33474
rect 9751 33467 9809 33473
rect 9490 33436 9496 33448
rect 9324 33408 9496 33436
rect 8481 33399 8539 33405
rect 9490 33396 9496 33408
rect 9548 33396 9554 33448
rect 9858 33300 9864 33312
rect 8312 33272 9864 33300
rect 9858 33260 9864 33272
rect 9916 33260 9922 33312
rect 9950 33260 9956 33312
rect 10008 33300 10014 33312
rect 10244 33300 10272 33476
rect 11793 33473 11805 33476
rect 11839 33473 11851 33507
rect 11793 33467 11851 33473
rect 15102 33464 15108 33516
rect 15160 33464 15166 33516
rect 17310 33464 17316 33516
rect 17368 33464 17374 33516
rect 10318 33396 10324 33448
rect 10376 33436 10382 33448
rect 11609 33439 11667 33445
rect 11609 33436 11621 33439
rect 10376 33408 11621 33436
rect 10376 33396 10382 33408
rect 11609 33405 11621 33408
rect 11655 33405 11667 33439
rect 12529 33439 12587 33445
rect 12529 33436 12541 33439
rect 11609 33399 11667 33405
rect 11716 33408 12541 33436
rect 11238 33328 11244 33380
rect 11296 33368 11302 33380
rect 11716 33368 11744 33408
rect 12529 33405 12541 33408
rect 12575 33405 12587 33439
rect 12529 33399 12587 33405
rect 12618 33396 12624 33448
rect 12676 33445 12682 33448
rect 12676 33439 12704 33445
rect 12692 33405 12704 33439
rect 12676 33399 12704 33405
rect 12805 33439 12863 33445
rect 12805 33405 12817 33439
rect 12851 33436 12863 33439
rect 13170 33436 13176 33448
rect 12851 33408 13176 33436
rect 12851 33405 12863 33408
rect 12805 33399 12863 33405
rect 12676 33396 12682 33399
rect 13170 33396 13176 33408
rect 13228 33396 13234 33448
rect 13909 33439 13967 33445
rect 13909 33405 13921 33439
rect 13955 33405 13967 33439
rect 13909 33399 13967 33405
rect 14093 33439 14151 33445
rect 14093 33405 14105 33439
rect 14139 33436 14151 33439
rect 14553 33439 14611 33445
rect 14139 33408 14412 33436
rect 14139 33405 14151 33408
rect 14093 33399 14151 33405
rect 11790 33368 11796 33380
rect 11296 33340 11796 33368
rect 11296 33328 11302 33340
rect 11790 33328 11796 33340
rect 11848 33328 11854 33380
rect 12250 33328 12256 33380
rect 12308 33328 12314 33380
rect 13924 33368 13952 33399
rect 14384 33380 14412 33408
rect 14553 33405 14565 33439
rect 14599 33436 14611 33439
rect 14642 33436 14648 33448
rect 14599 33408 14648 33436
rect 14599 33405 14611 33408
rect 14553 33399 14611 33405
rect 14642 33396 14648 33408
rect 14700 33396 14706 33448
rect 14826 33396 14832 33448
rect 14884 33396 14890 33448
rect 14918 33396 14924 33448
rect 14976 33445 14982 33448
rect 14976 33439 15004 33445
rect 14992 33405 15004 33439
rect 14976 33399 15004 33405
rect 14976 33396 14982 33399
rect 14182 33368 14188 33380
rect 13924 33340 14188 33368
rect 14182 33328 14188 33340
rect 14240 33328 14246 33380
rect 14366 33328 14372 33380
rect 14424 33328 14430 33380
rect 10008 33272 10272 33300
rect 10008 33260 10014 33272
rect 10410 33260 10416 33312
rect 10468 33300 10474 33312
rect 12618 33300 12624 33312
rect 10468 33272 12624 33300
rect 10468 33260 10474 33272
rect 12618 33260 12624 33272
rect 12676 33260 12682 33312
rect 13449 33303 13507 33309
rect 13449 33269 13461 33303
rect 13495 33300 13507 33303
rect 17604 33300 17632 33544
rect 19518 33532 19524 33544
rect 19576 33572 19582 33584
rect 19576 33544 19748 33572
rect 19576 33532 19582 33544
rect 17954 33464 17960 33516
rect 18012 33504 18018 33516
rect 18325 33507 18383 33513
rect 18325 33504 18337 33507
rect 18012 33476 18337 33504
rect 18012 33464 18018 33476
rect 18325 33473 18337 33476
rect 18371 33473 18383 33507
rect 18325 33467 18383 33473
rect 18693 33507 18751 33513
rect 18693 33473 18705 33507
rect 18739 33473 18751 33507
rect 18693 33467 18751 33473
rect 19061 33507 19119 33513
rect 19061 33473 19073 33507
rect 19107 33504 19119 33507
rect 19429 33507 19487 33513
rect 19429 33504 19441 33507
rect 19107 33476 19441 33504
rect 19107 33473 19119 33476
rect 19061 33467 19119 33473
rect 18708 33436 18736 33467
rect 19168 33448 19196 33476
rect 19429 33473 19441 33476
rect 19475 33473 19487 33507
rect 19429 33467 19487 33473
rect 19610 33464 19616 33516
rect 19668 33464 19674 33516
rect 19720 33504 19748 33544
rect 20180 33513 20208 33612
rect 22186 33600 22192 33652
rect 22244 33600 22250 33652
rect 22738 33600 22744 33652
rect 22796 33600 22802 33652
rect 23017 33643 23075 33649
rect 23017 33609 23029 33643
rect 23063 33640 23075 33643
rect 23290 33640 23296 33652
rect 23063 33612 23296 33640
rect 23063 33609 23075 33612
rect 23017 33603 23075 33609
rect 23290 33600 23296 33612
rect 23348 33600 23354 33652
rect 23382 33600 23388 33652
rect 23440 33600 23446 33652
rect 23658 33600 23664 33652
rect 23716 33640 23722 33652
rect 23753 33643 23811 33649
rect 23753 33640 23765 33643
rect 23716 33612 23765 33640
rect 23716 33600 23722 33612
rect 23753 33609 23765 33612
rect 23799 33609 23811 33643
rect 23753 33603 23811 33609
rect 22204 33572 22232 33600
rect 23400 33572 23428 33600
rect 24121 33575 24179 33581
rect 24121 33572 24133 33575
rect 22204 33544 23244 33572
rect 23400 33544 24133 33572
rect 19889 33507 19947 33513
rect 19889 33504 19901 33507
rect 19720 33476 19901 33504
rect 19889 33473 19901 33476
rect 19935 33473 19947 33507
rect 19889 33467 19947 33473
rect 20165 33507 20223 33513
rect 20165 33473 20177 33507
rect 20211 33473 20223 33507
rect 22281 33507 22339 33513
rect 22281 33504 22293 33507
rect 20165 33467 20223 33473
rect 22066 33476 22293 33504
rect 18156 33408 18736 33436
rect 18156 33377 18184 33408
rect 19150 33396 19156 33448
rect 19208 33396 19214 33448
rect 19337 33439 19395 33445
rect 19337 33405 19349 33439
rect 19383 33436 19395 33439
rect 19521 33439 19579 33445
rect 19521 33436 19533 33439
rect 19383 33408 19533 33436
rect 19383 33405 19395 33408
rect 19337 33399 19395 33405
rect 19521 33405 19533 33408
rect 19567 33405 19579 33439
rect 19521 33399 19579 33405
rect 18141 33371 18199 33377
rect 18141 33337 18153 33371
rect 18187 33337 18199 33371
rect 18141 33331 18199 33337
rect 18598 33328 18604 33380
rect 18656 33368 18662 33380
rect 22066 33368 22094 33476
rect 22281 33473 22293 33476
rect 22327 33473 22339 33507
rect 22281 33467 22339 33473
rect 22646 33464 22652 33516
rect 22704 33504 22710 33516
rect 23216 33513 23244 33544
rect 24121 33541 24133 33544
rect 24167 33541 24179 33575
rect 24121 33535 24179 33541
rect 22925 33507 22983 33513
rect 22925 33504 22937 33507
rect 22704 33476 22937 33504
rect 22704 33464 22710 33476
rect 22925 33473 22937 33476
rect 22971 33473 22983 33507
rect 22925 33467 22983 33473
rect 23201 33507 23259 33513
rect 23201 33473 23213 33507
rect 23247 33473 23259 33507
rect 23201 33467 23259 33473
rect 23290 33464 23296 33516
rect 23348 33504 23354 33516
rect 23569 33507 23627 33513
rect 23569 33504 23581 33507
rect 23348 33476 23581 33504
rect 23348 33464 23354 33476
rect 23569 33473 23581 33476
rect 23615 33473 23627 33507
rect 23569 33467 23627 33473
rect 23934 33464 23940 33516
rect 23992 33464 23998 33516
rect 18656 33340 19288 33368
rect 18656 33328 18662 33340
rect 19260 33309 19288 33340
rect 19352 33340 22094 33368
rect 19352 33312 19380 33340
rect 13495 33272 17632 33300
rect 18785 33303 18843 33309
rect 13495 33269 13507 33272
rect 13449 33263 13507 33269
rect 18785 33269 18797 33303
rect 18831 33300 18843 33303
rect 19153 33303 19211 33309
rect 19153 33300 19165 33303
rect 18831 33272 19165 33300
rect 18831 33269 18843 33272
rect 18785 33263 18843 33269
rect 19153 33269 19165 33272
rect 19199 33269 19211 33303
rect 19153 33263 19211 33269
rect 19245 33303 19303 33309
rect 19245 33269 19257 33303
rect 19291 33269 19303 33303
rect 19245 33263 19303 33269
rect 19334 33260 19340 33312
rect 19392 33260 19398 33312
rect 20257 33303 20315 33309
rect 20257 33269 20269 33303
rect 20303 33300 20315 33303
rect 20806 33300 20812 33312
rect 20303 33272 20812 33300
rect 20303 33269 20315 33272
rect 20257 33263 20315 33269
rect 20806 33260 20812 33272
rect 20864 33260 20870 33312
rect 22094 33260 22100 33312
rect 22152 33260 22158 33312
rect 23385 33303 23443 33309
rect 23385 33269 23397 33303
rect 23431 33300 23443 33303
rect 23842 33300 23848 33312
rect 23431 33272 23848 33300
rect 23431 33269 23443 33272
rect 23385 33263 23443 33269
rect 23842 33260 23848 33272
rect 23900 33260 23906 33312
rect 24394 33260 24400 33312
rect 24452 33260 24458 33312
rect 1104 33210 24840 33232
rect 1104 33158 3917 33210
rect 3969 33158 3981 33210
rect 4033 33158 4045 33210
rect 4097 33158 4109 33210
rect 4161 33158 4173 33210
rect 4225 33158 9851 33210
rect 9903 33158 9915 33210
rect 9967 33158 9979 33210
rect 10031 33158 10043 33210
rect 10095 33158 10107 33210
rect 10159 33158 15785 33210
rect 15837 33158 15849 33210
rect 15901 33158 15913 33210
rect 15965 33158 15977 33210
rect 16029 33158 16041 33210
rect 16093 33158 21719 33210
rect 21771 33158 21783 33210
rect 21835 33158 21847 33210
rect 21899 33158 21911 33210
rect 21963 33158 21975 33210
rect 22027 33158 24840 33210
rect 1104 33136 24840 33158
rect 1854 33056 1860 33108
rect 1912 33096 1918 33108
rect 1912 33068 2544 33096
rect 1912 33056 1918 33068
rect 2516 33028 2544 33068
rect 5258 33056 5264 33108
rect 5316 33056 5322 33108
rect 7466 33056 7472 33108
rect 7524 33056 7530 33108
rect 8018 33056 8024 33108
rect 8076 33096 8082 33108
rect 8662 33096 8668 33108
rect 8076 33068 8668 33096
rect 8076 33056 8082 33068
rect 8662 33056 8668 33068
rect 8720 33056 8726 33108
rect 9309 33099 9367 33105
rect 9309 33065 9321 33099
rect 9355 33096 9367 33099
rect 9398 33096 9404 33108
rect 9355 33068 9404 33096
rect 9355 33065 9367 33068
rect 9309 33059 9367 33065
rect 9398 33056 9404 33068
rect 9456 33056 9462 33108
rect 11974 33096 11980 33108
rect 9646 33068 11192 33096
rect 2516 33000 3740 33028
rect 3050 32920 3056 32972
rect 3108 32960 3114 32972
rect 3510 32960 3516 32972
rect 3108 32932 3516 32960
rect 3108 32920 3114 32932
rect 3510 32920 3516 32932
rect 3568 32920 3574 32972
rect 1397 32895 1455 32901
rect 1397 32861 1409 32895
rect 1443 32892 1455 32895
rect 1578 32892 1584 32904
rect 1443 32864 1584 32892
rect 1443 32861 1455 32864
rect 1397 32855 1455 32861
rect 1578 32852 1584 32864
rect 1636 32852 1642 32904
rect 1670 32852 1676 32904
rect 1728 32892 1734 32904
rect 2777 32895 2835 32901
rect 1728 32864 1771 32892
rect 1728 32852 1734 32864
rect 2777 32861 2789 32895
rect 2823 32861 2835 32895
rect 2777 32855 2835 32861
rect 1302 32784 1308 32836
rect 1360 32824 1366 32836
rect 2792 32824 2820 32855
rect 3602 32852 3608 32904
rect 3660 32852 3666 32904
rect 3712 32882 3740 33000
rect 3792 32972 3844 32978
rect 5074 32920 5080 32972
rect 5132 32960 5138 32972
rect 5276 32960 5304 33056
rect 5132 32932 5304 32960
rect 5132 32920 5138 32932
rect 6546 32920 6552 32972
rect 6604 32920 6610 32972
rect 7282 32920 7288 32972
rect 7340 32960 7346 32972
rect 7484 32960 7512 33056
rect 7650 32988 7656 33040
rect 7708 33028 7714 33040
rect 9646 33028 9674 33068
rect 7708 33000 9674 33028
rect 7708 32988 7714 33000
rect 7340 32932 7512 32960
rect 9416 32932 9628 32960
rect 7340 32920 7346 32932
rect 3792 32914 3844 32920
rect 3878 32882 3884 32904
rect 3712 32854 3884 32882
rect 3878 32852 3884 32854
rect 3936 32892 3942 32904
rect 3936 32864 4200 32892
rect 3936 32852 3942 32864
rect 1360 32796 2820 32824
rect 1360 32784 1366 32796
rect 3050 32784 3056 32836
rect 3108 32784 3114 32836
rect 4172 32824 4200 32864
rect 4246 32852 4252 32904
rect 4304 32852 4310 32904
rect 4338 32852 4344 32904
rect 4396 32852 4402 32904
rect 9416 32892 9444 32932
rect 4816 32864 9444 32892
rect 4709 32827 4767 32833
rect 4709 32824 4721 32827
rect 3344 32796 4108 32824
rect 4172 32796 4721 32824
rect 1486 32716 1492 32768
rect 1544 32756 1550 32768
rect 2409 32759 2467 32765
rect 2409 32756 2421 32759
rect 1544 32728 2421 32756
rect 1544 32716 1550 32728
rect 2409 32725 2421 32728
rect 2455 32725 2467 32759
rect 2409 32719 2467 32725
rect 2590 32716 2596 32768
rect 2648 32756 2654 32768
rect 3344 32756 3372 32796
rect 2648 32728 3372 32756
rect 3421 32759 3479 32765
rect 2648 32716 2654 32728
rect 3421 32725 3433 32759
rect 3467 32756 3479 32759
rect 3602 32756 3608 32768
rect 3467 32728 3608 32756
rect 3467 32725 3479 32728
rect 3421 32719 3479 32725
rect 3602 32716 3608 32728
rect 3660 32716 3666 32768
rect 3694 32716 3700 32768
rect 3752 32756 3758 32768
rect 3973 32759 4031 32765
rect 3973 32756 3985 32759
rect 3752 32728 3985 32756
rect 3752 32716 3758 32728
rect 3973 32725 3985 32728
rect 4019 32725 4031 32759
rect 4080 32756 4108 32796
rect 4709 32793 4721 32796
rect 4755 32793 4767 32827
rect 4709 32787 4767 32793
rect 4816 32756 4844 32864
rect 9490 32852 9496 32904
rect 9548 32852 9554 32904
rect 9600 32892 9628 32932
rect 9674 32920 9680 32972
rect 9732 32960 9738 32972
rect 9769 32963 9827 32969
rect 9769 32960 9781 32963
rect 9732 32932 9781 32960
rect 9732 32920 9738 32932
rect 9769 32929 9781 32932
rect 9815 32929 9827 32963
rect 9769 32923 9827 32929
rect 9600 32864 9996 32892
rect 5718 32784 5724 32836
rect 5776 32784 5782 32836
rect 6454 32784 6460 32836
rect 6512 32784 6518 32836
rect 6546 32784 6552 32836
rect 6604 32784 6610 32836
rect 6914 32784 6920 32836
rect 6972 32784 6978 32836
rect 7098 32784 7104 32836
rect 7156 32824 7162 32836
rect 7285 32827 7343 32833
rect 7285 32824 7297 32827
rect 7156 32796 7297 32824
rect 7156 32784 7162 32796
rect 7285 32793 7297 32796
rect 7331 32793 7343 32827
rect 9858 32824 9864 32836
rect 7285 32787 7343 32793
rect 7392 32796 9864 32824
rect 4080 32728 4844 32756
rect 3973 32719 4031 32725
rect 4982 32716 4988 32768
rect 5040 32756 5046 32768
rect 5077 32759 5135 32765
rect 5077 32756 5089 32759
rect 5040 32728 5089 32756
rect 5040 32716 5046 32728
rect 5077 32725 5089 32728
rect 5123 32725 5135 32759
rect 5077 32719 5135 32725
rect 5258 32716 5264 32768
rect 5316 32716 5322 32768
rect 6181 32759 6239 32765
rect 6181 32725 6193 32759
rect 6227 32756 6239 32759
rect 7392 32756 7420 32796
rect 9858 32784 9864 32796
rect 9916 32784 9922 32836
rect 9968 32824 9996 32864
rect 10042 32852 10048 32904
rect 10100 32852 10106 32904
rect 11164 32892 11192 33068
rect 11256 33068 11980 33096
rect 11256 32969 11284 33068
rect 11974 33056 11980 33068
rect 12032 33056 12038 33108
rect 12250 33056 12256 33108
rect 12308 33056 12314 33108
rect 14090 33096 14096 33108
rect 12636 33068 14096 33096
rect 11241 32963 11299 32969
rect 11241 32929 11253 32963
rect 11287 32929 11299 32963
rect 11241 32923 11299 32929
rect 12526 32920 12532 32972
rect 12584 32960 12590 32972
rect 12636 32969 12664 33068
rect 14090 33056 14096 33068
rect 14148 33056 14154 33108
rect 14826 33096 14832 33108
rect 14292 33068 14832 33096
rect 12621 32963 12679 32969
rect 12621 32960 12633 32963
rect 12584 32932 12633 32960
rect 12584 32920 12590 32932
rect 12621 32929 12633 32932
rect 12667 32929 12679 32963
rect 12621 32923 12679 32929
rect 11515 32895 11573 32901
rect 11515 32892 11527 32895
rect 11164 32864 11527 32892
rect 11515 32861 11527 32864
rect 11561 32892 11573 32895
rect 12895 32895 12953 32901
rect 11561 32864 11652 32892
rect 11561 32861 11573 32864
rect 11515 32855 11573 32861
rect 11624 32824 11652 32864
rect 12895 32861 12907 32895
rect 12941 32892 12953 32895
rect 13998 32892 14004 32904
rect 12941 32864 14004 32892
rect 12941 32861 12953 32864
rect 12895 32855 12953 32861
rect 11974 32824 11980 32836
rect 9968 32796 10916 32824
rect 11624 32796 11980 32824
rect 6227 32728 7420 32756
rect 6227 32725 6239 32728
rect 6181 32719 6239 32725
rect 7466 32716 7472 32768
rect 7524 32756 7530 32768
rect 8202 32756 8208 32768
rect 7524 32728 8208 32756
rect 7524 32716 7530 32728
rect 8202 32716 8208 32728
rect 8260 32716 8266 32768
rect 10778 32716 10784 32768
rect 10836 32716 10842 32768
rect 10888 32756 10916 32796
rect 11974 32784 11980 32796
rect 12032 32824 12038 32836
rect 13078 32824 13084 32836
rect 12032 32796 13084 32824
rect 12032 32784 12038 32796
rect 13078 32784 13084 32796
rect 13136 32784 13142 32836
rect 13188 32756 13216 32864
rect 13998 32852 14004 32864
rect 14056 32852 14062 32904
rect 14292 32824 14320 33068
rect 14826 33056 14832 33068
rect 14884 33056 14890 33108
rect 16482 33096 16488 33108
rect 16040 33068 16488 33096
rect 14366 32988 14372 33040
rect 14424 33028 14430 33040
rect 15562 33028 15568 33040
rect 14424 33000 15568 33028
rect 14424 32988 14430 33000
rect 15562 32988 15568 33000
rect 15620 32988 15626 33040
rect 16040 33037 16068 33068
rect 16482 33056 16488 33068
rect 16540 33056 16546 33108
rect 17126 33056 17132 33108
rect 17184 33096 17190 33108
rect 17313 33099 17371 33105
rect 17313 33096 17325 33099
rect 17184 33068 17325 33096
rect 17184 33056 17190 33068
rect 17313 33065 17325 33068
rect 17359 33065 17371 33099
rect 17313 33059 17371 33065
rect 18046 33056 18052 33108
rect 18104 33096 18110 33108
rect 19242 33096 19248 33108
rect 18104 33068 19248 33096
rect 18104 33056 18110 33068
rect 19242 33056 19248 33068
rect 19300 33056 19306 33108
rect 20806 33056 20812 33108
rect 20864 33056 20870 33108
rect 21284 33068 21496 33096
rect 16025 33031 16083 33037
rect 16025 32997 16037 33031
rect 16071 32997 16083 33031
rect 16025 32991 16083 32997
rect 20625 33031 20683 33037
rect 20625 32997 20637 33031
rect 20671 33028 20683 33031
rect 21284 33028 21312 33068
rect 20671 33000 21312 33028
rect 21361 33031 21419 33037
rect 20671 32997 20683 33000
rect 20625 32991 20683 32997
rect 21361 32997 21373 33031
rect 21407 32997 21419 33031
rect 21361 32991 21419 32997
rect 16418 32963 16476 32969
rect 16418 32960 16430 32963
rect 14844 32932 16430 32960
rect 14844 32904 14872 32932
rect 16418 32929 16430 32932
rect 16464 32929 16476 32963
rect 16418 32923 16476 32929
rect 16577 32963 16635 32969
rect 16577 32929 16589 32963
rect 16623 32960 16635 32963
rect 16758 32960 16764 32972
rect 16623 32932 16764 32960
rect 16623 32929 16635 32932
rect 16577 32923 16635 32929
rect 16758 32920 16764 32932
rect 16816 32920 16822 32972
rect 20993 32963 21051 32969
rect 20993 32929 21005 32963
rect 21039 32960 21051 32963
rect 21177 32963 21235 32969
rect 21177 32960 21189 32963
rect 21039 32932 21189 32960
rect 21039 32929 21051 32932
rect 20993 32923 21051 32929
rect 21177 32929 21189 32932
rect 21223 32929 21235 32963
rect 21177 32923 21235 32929
rect 14826 32852 14832 32904
rect 14884 32852 14890 32904
rect 15378 32852 15384 32904
rect 15436 32852 15442 32904
rect 15562 32852 15568 32904
rect 15620 32852 15626 32904
rect 16298 32852 16304 32904
rect 16356 32852 16362 32904
rect 17221 32895 17279 32901
rect 17221 32861 17233 32895
rect 17267 32892 17279 32895
rect 17497 32895 17555 32901
rect 17497 32892 17509 32895
rect 17267 32864 17509 32892
rect 17267 32861 17279 32864
rect 17221 32855 17279 32861
rect 17497 32861 17509 32864
rect 17543 32861 17555 32895
rect 17497 32855 17555 32861
rect 17586 32852 17592 32904
rect 17644 32892 17650 32904
rect 17681 32895 17739 32901
rect 17681 32892 17693 32895
rect 17644 32864 17693 32892
rect 17644 32852 17650 32864
rect 17681 32861 17693 32864
rect 17727 32892 17739 32895
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 17727 32864 19257 32892
rect 17727 32861 17739 32864
rect 17681 32855 17739 32861
rect 19245 32861 19257 32864
rect 19291 32892 19303 32895
rect 20622 32892 20628 32904
rect 19291 32864 20628 32892
rect 19291 32861 19303 32864
rect 19245 32855 19303 32861
rect 20622 32852 20628 32864
rect 20680 32852 20686 32904
rect 20717 32895 20775 32901
rect 20717 32861 20729 32895
rect 20763 32892 20775 32895
rect 21085 32895 21143 32901
rect 21085 32892 21097 32895
rect 20763 32864 21097 32892
rect 20763 32861 20775 32864
rect 20717 32855 20775 32861
rect 21085 32861 21097 32864
rect 21131 32861 21143 32895
rect 21085 32855 21143 32861
rect 21269 32895 21327 32901
rect 21269 32861 21281 32895
rect 21315 32892 21327 32895
rect 21376 32892 21404 32991
rect 21315 32864 21404 32892
rect 21468 32892 21496 33068
rect 22094 33056 22100 33108
rect 22152 33056 22158 33108
rect 23017 33099 23075 33105
rect 23017 33065 23029 33099
rect 23063 33096 23075 33099
rect 23290 33096 23296 33108
rect 23063 33068 23296 33096
rect 23063 33065 23075 33068
rect 23017 33059 23075 33065
rect 23290 33056 23296 33068
rect 23348 33056 23354 33108
rect 22112 32960 22140 33056
rect 22649 33031 22707 33037
rect 22649 32997 22661 33031
rect 22695 33028 22707 33031
rect 22695 33000 23612 33028
rect 22695 32997 22707 33000
rect 22649 32991 22707 32997
rect 22112 32932 23244 32960
rect 23216 32901 23244 32932
rect 21545 32895 21603 32901
rect 21545 32892 21557 32895
rect 21468 32864 21557 32892
rect 21315 32861 21327 32864
rect 21269 32855 21327 32861
rect 21545 32861 21557 32864
rect 21591 32861 21603 32895
rect 22005 32895 22063 32901
rect 22005 32892 22017 32895
rect 21545 32855 21603 32861
rect 21652 32864 22017 32892
rect 14366 32824 14372 32836
rect 14292 32796 14372 32824
rect 14366 32784 14372 32796
rect 14424 32784 14430 32836
rect 17954 32833 17960 32836
rect 17926 32827 17960 32833
rect 17926 32824 17938 32827
rect 17696 32796 17938 32824
rect 10888 32728 13216 32756
rect 13630 32716 13636 32768
rect 13688 32716 13694 32768
rect 13998 32716 14004 32768
rect 14056 32756 14062 32768
rect 17696 32756 17724 32796
rect 17926 32793 17938 32796
rect 17926 32787 17960 32793
rect 17954 32784 17960 32787
rect 18012 32784 18018 32836
rect 19518 32833 19524 32836
rect 19512 32824 19524 32833
rect 19479 32796 19524 32824
rect 19512 32787 19524 32796
rect 19518 32784 19524 32787
rect 19576 32784 19582 32836
rect 20732 32768 20760 32855
rect 21652 32836 21680 32864
rect 22005 32861 22017 32864
rect 22051 32861 22063 32895
rect 22005 32855 22063 32861
rect 22833 32895 22891 32901
rect 22833 32861 22845 32895
rect 22879 32861 22891 32895
rect 22833 32855 22891 32861
rect 23201 32895 23259 32901
rect 23201 32861 23213 32895
rect 23247 32861 23259 32895
rect 23201 32855 23259 32861
rect 21174 32784 21180 32836
rect 21232 32824 21238 32836
rect 21634 32824 21640 32836
rect 21232 32796 21640 32824
rect 21232 32784 21238 32796
rect 21634 32784 21640 32796
rect 21692 32784 21698 32836
rect 22848 32824 22876 32855
rect 23474 32852 23480 32904
rect 23532 32852 23538 32904
rect 23584 32892 23612 33000
rect 23753 32895 23811 32901
rect 23753 32892 23765 32895
rect 23584 32864 23765 32892
rect 23753 32861 23765 32864
rect 23799 32861 23811 32895
rect 23753 32855 23811 32861
rect 23842 32852 23848 32904
rect 23900 32892 23906 32904
rect 23937 32895 23995 32901
rect 23937 32892 23949 32895
rect 23900 32864 23949 32892
rect 23900 32852 23906 32864
rect 23937 32861 23949 32864
rect 23983 32861 23995 32895
rect 23937 32855 23995 32861
rect 22066 32796 22876 32824
rect 14056 32728 17724 32756
rect 19061 32759 19119 32765
rect 14056 32716 14062 32728
rect 19061 32725 19073 32759
rect 19107 32756 19119 32759
rect 19334 32756 19340 32768
rect 19107 32728 19340 32756
rect 19107 32725 19119 32728
rect 19061 32719 19119 32725
rect 19334 32716 19340 32728
rect 19392 32716 19398 32768
rect 20714 32716 20720 32768
rect 20772 32716 20778 32768
rect 20990 32716 20996 32768
rect 21048 32716 21054 32768
rect 21821 32759 21879 32765
rect 21821 32725 21833 32759
rect 21867 32756 21879 32759
rect 22066 32756 22094 32796
rect 21867 32728 22094 32756
rect 21867 32725 21879 32728
rect 21821 32719 21879 32725
rect 23290 32716 23296 32768
rect 23348 32716 23354 32768
rect 23566 32716 23572 32768
rect 23624 32716 23630 32768
rect 24118 32716 24124 32768
rect 24176 32716 24182 32768
rect 1104 32666 25000 32688
rect 1104 32614 6884 32666
rect 6936 32614 6948 32666
rect 7000 32614 7012 32666
rect 7064 32614 7076 32666
rect 7128 32614 7140 32666
rect 7192 32614 12818 32666
rect 12870 32614 12882 32666
rect 12934 32614 12946 32666
rect 12998 32614 13010 32666
rect 13062 32614 13074 32666
rect 13126 32614 18752 32666
rect 18804 32614 18816 32666
rect 18868 32614 18880 32666
rect 18932 32614 18944 32666
rect 18996 32614 19008 32666
rect 19060 32614 24686 32666
rect 24738 32614 24750 32666
rect 24802 32614 24814 32666
rect 24866 32614 24878 32666
rect 24930 32614 24942 32666
rect 24994 32614 25000 32666
rect 1104 32592 25000 32614
rect 1210 32512 1216 32564
rect 1268 32552 1274 32564
rect 2590 32552 2596 32564
rect 1268 32524 2596 32552
rect 1268 32512 1274 32524
rect 2590 32512 2596 32524
rect 2648 32512 2654 32564
rect 2866 32512 2872 32564
rect 2924 32552 2930 32564
rect 2924 32524 3188 32552
rect 2924 32512 2930 32524
rect 2317 32419 2375 32425
rect 1504 32388 1808 32416
rect 1504 32360 1532 32388
rect 1397 32351 1455 32357
rect 1397 32317 1409 32351
rect 1443 32317 1455 32351
rect 1397 32311 1455 32317
rect 1412 32280 1440 32311
rect 1486 32308 1492 32360
rect 1544 32308 1550 32360
rect 1581 32351 1639 32357
rect 1581 32317 1593 32351
rect 1627 32348 1639 32351
rect 1670 32348 1676 32360
rect 1627 32320 1676 32348
rect 1627 32317 1639 32320
rect 1581 32311 1639 32317
rect 1670 32308 1676 32320
rect 1728 32308 1734 32360
rect 1780 32348 1808 32388
rect 2317 32385 2329 32419
rect 2363 32385 2375 32419
rect 3160 32416 3188 32524
rect 3234 32512 3240 32564
rect 3292 32512 3298 32564
rect 3602 32512 3608 32564
rect 3660 32552 3666 32564
rect 3660 32524 4200 32552
rect 3660 32512 3666 32524
rect 3789 32419 3847 32425
rect 3789 32416 3801 32419
rect 3160 32388 3801 32416
rect 2317 32379 2375 32385
rect 3789 32385 3801 32388
rect 3835 32385 3847 32419
rect 3789 32379 3847 32385
rect 2041 32351 2099 32357
rect 2041 32348 2053 32351
rect 1780 32320 2053 32348
rect 2041 32317 2053 32320
rect 2087 32317 2099 32351
rect 2041 32311 2099 32317
rect 2130 32308 2136 32360
rect 2188 32348 2194 32360
rect 2332 32348 2360 32379
rect 3970 32376 3976 32428
rect 4028 32416 4034 32428
rect 4063 32419 4121 32425
rect 4063 32416 4075 32419
rect 4028 32388 4075 32416
rect 4028 32376 4034 32388
rect 4063 32385 4075 32388
rect 4109 32385 4121 32419
rect 4172 32416 4200 32524
rect 4338 32512 4344 32564
rect 4396 32552 4402 32564
rect 4801 32555 4859 32561
rect 4801 32552 4813 32555
rect 4396 32524 4813 32552
rect 4396 32512 4402 32524
rect 4801 32521 4813 32524
rect 4847 32521 4859 32555
rect 4801 32515 4859 32521
rect 5258 32512 5264 32564
rect 5316 32552 5322 32564
rect 9401 32555 9459 32561
rect 5316 32524 9352 32552
rect 5316 32512 5322 32524
rect 4246 32444 4252 32496
rect 4304 32484 4310 32496
rect 5442 32484 5448 32496
rect 4304 32456 5448 32484
rect 4304 32444 4310 32456
rect 5442 32444 5448 32456
rect 5500 32444 5506 32496
rect 5534 32444 5540 32496
rect 5592 32444 5598 32496
rect 6730 32444 6736 32496
rect 6788 32484 6794 32496
rect 7466 32484 7472 32496
rect 6788 32456 7472 32484
rect 6788 32444 6794 32456
rect 7466 32444 7472 32456
rect 7524 32444 7530 32496
rect 7742 32484 7748 32496
rect 7576 32456 7748 32484
rect 5552 32416 5580 32444
rect 4172 32388 5580 32416
rect 4063 32379 4121 32385
rect 2188 32320 2360 32348
rect 2188 32308 2194 32320
rect 2406 32308 2412 32360
rect 2464 32357 2470 32360
rect 2464 32351 2492 32357
rect 2480 32317 2492 32351
rect 2464 32311 2492 32317
rect 2464 32308 2470 32311
rect 2590 32308 2596 32360
rect 2648 32308 2654 32360
rect 1854 32280 1860 32292
rect 1412 32252 1860 32280
rect 1854 32240 1860 32252
rect 1912 32240 1918 32292
rect 7484 32280 7512 32444
rect 7576 32357 7604 32456
rect 7742 32444 7748 32456
rect 7800 32444 7806 32496
rect 9324 32484 9352 32524
rect 9401 32521 9413 32555
rect 9447 32552 9459 32555
rect 9490 32552 9496 32564
rect 9447 32524 9496 32552
rect 9447 32521 9459 32524
rect 9401 32515 9459 32521
rect 9490 32512 9496 32524
rect 9548 32512 9554 32564
rect 19061 32555 19119 32561
rect 9600 32524 19012 32552
rect 9600 32484 9628 32524
rect 9324 32456 9628 32484
rect 9858 32444 9864 32496
rect 9916 32484 9922 32496
rect 11701 32487 11759 32493
rect 11701 32484 11713 32487
rect 9916 32456 11713 32484
rect 9916 32444 9922 32456
rect 11701 32453 11713 32456
rect 11747 32484 11759 32487
rect 13262 32484 13268 32496
rect 11747 32456 13268 32484
rect 11747 32453 11759 32456
rect 11701 32447 11759 32453
rect 13262 32444 13268 32456
rect 13320 32444 13326 32496
rect 14090 32444 14096 32496
rect 14148 32444 14154 32496
rect 14458 32444 14464 32496
rect 14516 32444 14522 32496
rect 14826 32444 14832 32496
rect 14884 32444 14890 32496
rect 15197 32487 15255 32493
rect 15197 32453 15209 32487
rect 15243 32484 15255 32487
rect 15562 32484 15568 32496
rect 15243 32456 15568 32484
rect 15243 32453 15255 32456
rect 15197 32447 15255 32453
rect 15562 32444 15568 32456
rect 15620 32484 15626 32496
rect 15620 32456 16160 32484
rect 15620 32444 15626 32456
rect 16132 32428 16160 32456
rect 16758 32444 16764 32496
rect 16816 32484 16822 32496
rect 18046 32484 18052 32496
rect 16816 32456 18052 32484
rect 16816 32444 16822 32456
rect 18046 32444 18052 32456
rect 18104 32444 18110 32496
rect 18984 32484 19012 32524
rect 19061 32521 19073 32555
rect 19107 32552 19119 32555
rect 19150 32552 19156 32564
rect 19107 32524 19156 32552
rect 19107 32521 19119 32524
rect 19061 32515 19119 32521
rect 19150 32512 19156 32524
rect 19208 32512 19214 32564
rect 19429 32555 19487 32561
rect 19429 32521 19441 32555
rect 19475 32552 19487 32555
rect 19610 32552 19616 32564
rect 19475 32524 19616 32552
rect 19475 32521 19487 32524
rect 19429 32515 19487 32521
rect 19610 32512 19616 32524
rect 19668 32512 19674 32564
rect 20714 32512 20720 32564
rect 20772 32512 20778 32564
rect 20806 32512 20812 32564
rect 20864 32552 20870 32564
rect 23201 32555 23259 32561
rect 20864 32524 23152 32552
rect 20864 32512 20870 32524
rect 22066 32487 22124 32493
rect 22066 32484 22078 32487
rect 18984 32456 22078 32484
rect 18307 32449 18365 32455
rect 7668 32388 7880 32416
rect 7561 32351 7619 32357
rect 7561 32317 7573 32351
rect 7607 32317 7619 32351
rect 7561 32311 7619 32317
rect 7668 32280 7696 32388
rect 7745 32351 7803 32357
rect 7745 32317 7757 32351
rect 7791 32317 7803 32351
rect 7852 32348 7880 32388
rect 8754 32376 8760 32428
rect 8812 32376 8818 32428
rect 9674 32376 9680 32428
rect 9732 32416 9738 32428
rect 10045 32419 10103 32425
rect 10045 32416 10057 32419
rect 9732 32388 10057 32416
rect 9732 32376 9738 32388
rect 10045 32385 10057 32388
rect 10091 32385 10103 32419
rect 10045 32379 10103 32385
rect 10226 32376 10232 32428
rect 10284 32416 10290 32428
rect 10319 32419 10377 32425
rect 10319 32416 10331 32419
rect 10284 32388 10331 32416
rect 10284 32376 10290 32388
rect 10319 32385 10331 32388
rect 10365 32385 10377 32419
rect 10319 32379 10377 32385
rect 10686 32376 10692 32428
rect 10744 32416 10750 32428
rect 10744 32388 11560 32416
rect 10744 32376 10750 32388
rect 11532 32360 11560 32388
rect 14366 32376 14372 32428
rect 14424 32376 14430 32428
rect 16114 32376 16120 32428
rect 16172 32376 16178 32428
rect 16666 32376 16672 32428
rect 16724 32376 16730 32428
rect 16776 32416 16804 32444
rect 16911 32419 16969 32425
rect 16911 32416 16923 32419
rect 16776 32388 16923 32416
rect 16911 32385 16923 32388
rect 16957 32385 16969 32419
rect 16911 32379 16969 32385
rect 17034 32376 17040 32428
rect 17092 32416 17098 32428
rect 18307 32416 18319 32449
rect 17092 32415 18319 32416
rect 18353 32446 18365 32449
rect 18353 32416 18368 32446
rect 18353 32415 18736 32416
rect 17092 32388 18736 32415
rect 17092 32376 17098 32388
rect 8481 32351 8539 32357
rect 8481 32348 8493 32351
rect 7852 32320 8493 32348
rect 7745 32311 7803 32317
rect 8481 32317 8493 32320
rect 8527 32317 8539 32351
rect 8481 32311 8539 32317
rect 8619 32351 8677 32357
rect 8619 32317 8631 32351
rect 8665 32348 8677 32351
rect 9490 32348 9496 32360
rect 8665 32320 9496 32348
rect 8665 32317 8677 32320
rect 8619 32311 8677 32317
rect 7484 32252 7696 32280
rect 7760 32280 7788 32311
rect 9490 32308 9496 32320
rect 9548 32308 9554 32360
rect 11514 32308 11520 32360
rect 11572 32308 11578 32360
rect 13630 32308 13636 32360
rect 13688 32348 13694 32360
rect 13688 32320 13938 32348
rect 13688 32308 13694 32320
rect 17862 32308 17868 32360
rect 17920 32348 17926 32360
rect 18049 32351 18107 32357
rect 18049 32348 18061 32351
rect 17920 32320 18061 32348
rect 17920 32308 17926 32320
rect 18049 32317 18061 32320
rect 18095 32317 18107 32351
rect 18708 32348 18736 32388
rect 19334 32376 19340 32428
rect 19392 32416 19398 32428
rect 19613 32419 19671 32425
rect 19613 32416 19625 32419
rect 19392 32388 19625 32416
rect 19392 32376 19398 32388
rect 19613 32385 19625 32388
rect 19659 32385 19671 32419
rect 19613 32379 19671 32385
rect 19702 32376 19708 32428
rect 19760 32376 19766 32428
rect 19979 32419 20037 32425
rect 19979 32385 19991 32419
rect 20025 32416 20037 32419
rect 20070 32416 20076 32428
rect 20025 32388 20076 32416
rect 20025 32385 20037 32388
rect 19979 32379 20037 32385
rect 20070 32376 20076 32388
rect 20128 32416 20134 32428
rect 20530 32416 20536 32428
rect 20128 32388 20536 32416
rect 20128 32376 20134 32388
rect 20530 32376 20536 32388
rect 20588 32376 20594 32428
rect 20622 32376 20628 32428
rect 20680 32376 20686 32428
rect 21652 32425 21680 32456
rect 22066 32453 22078 32456
rect 22112 32453 22124 32487
rect 23124 32484 23152 32524
rect 23201 32521 23213 32555
rect 23247 32552 23259 32555
rect 23474 32552 23480 32564
rect 23247 32524 23480 32552
rect 23247 32521 23259 32524
rect 23201 32515 23259 32521
rect 23474 32512 23480 32524
rect 23532 32512 23538 32564
rect 23566 32512 23572 32564
rect 23624 32552 23630 32564
rect 23624 32524 24164 32552
rect 23624 32512 23630 32524
rect 23750 32484 23756 32496
rect 23124 32456 23756 32484
rect 22066 32447 22124 32453
rect 23750 32444 23756 32456
rect 23808 32444 23814 32496
rect 24136 32493 24164 32524
rect 24121 32487 24179 32493
rect 24121 32453 24133 32487
rect 24167 32453 24179 32487
rect 24121 32447 24179 32453
rect 21637 32419 21695 32425
rect 21637 32385 21649 32419
rect 21683 32385 21695 32419
rect 21637 32379 21695 32385
rect 23382 32376 23388 32428
rect 23440 32416 23446 32428
rect 23661 32419 23719 32425
rect 23661 32416 23673 32419
rect 23440 32388 23673 32416
rect 23440 32376 23446 32388
rect 23661 32385 23673 32388
rect 23707 32385 23719 32419
rect 23661 32379 23719 32385
rect 23937 32419 23995 32425
rect 23937 32385 23949 32419
rect 23983 32385 23995 32419
rect 23937 32379 23995 32385
rect 19426 32348 19432 32360
rect 18708 32320 19432 32348
rect 18049 32311 18107 32317
rect 7760 32252 7878 32280
rect 1210 32172 1216 32224
rect 1268 32212 1274 32224
rect 1670 32212 1676 32224
rect 1268 32184 1676 32212
rect 1268 32172 1274 32184
rect 1670 32172 1676 32184
rect 1728 32172 1734 32224
rect 7850 32212 7878 32252
rect 8110 32240 8116 32292
rect 8168 32280 8174 32292
rect 8205 32283 8263 32289
rect 8205 32280 8217 32283
rect 8168 32252 8217 32280
rect 8168 32240 8174 32252
rect 8205 32249 8217 32252
rect 8251 32249 8263 32283
rect 8205 32243 8263 32249
rect 11882 32240 11888 32292
rect 11940 32240 11946 32292
rect 9306 32212 9312 32224
rect 7850 32184 9312 32212
rect 9306 32172 9312 32184
rect 9364 32212 9370 32224
rect 10502 32212 10508 32224
rect 9364 32184 10508 32212
rect 9364 32172 9370 32184
rect 10502 32172 10508 32184
rect 10560 32172 10566 32224
rect 11054 32172 11060 32224
rect 11112 32172 11118 32224
rect 15381 32215 15439 32221
rect 15381 32181 15393 32215
rect 15427 32212 15439 32215
rect 15562 32212 15568 32224
rect 15427 32184 15568 32212
rect 15427 32181 15439 32184
rect 15381 32175 15439 32181
rect 15562 32172 15568 32184
rect 15620 32172 15626 32224
rect 16942 32172 16948 32224
rect 17000 32212 17006 32224
rect 17681 32215 17739 32221
rect 17681 32212 17693 32215
rect 17000 32184 17693 32212
rect 17000 32172 17006 32184
rect 17681 32181 17693 32184
rect 17727 32181 17739 32215
rect 18064 32212 18092 32311
rect 19426 32308 19432 32320
rect 19484 32308 19490 32360
rect 19720 32212 19748 32376
rect 20640 32348 20668 32376
rect 21821 32351 21879 32357
rect 21821 32348 21833 32351
rect 20640 32320 21833 32348
rect 21821 32317 21833 32320
rect 21867 32317 21879 32351
rect 21821 32311 21879 32317
rect 23566 32308 23572 32360
rect 23624 32348 23630 32360
rect 23952 32348 23980 32379
rect 23624 32320 23980 32348
rect 23624 32308 23630 32320
rect 23106 32240 23112 32292
rect 23164 32280 23170 32292
rect 23164 32252 23796 32280
rect 23164 32240 23170 32252
rect 18064 32184 19748 32212
rect 17681 32175 17739 32181
rect 21450 32172 21456 32224
rect 21508 32172 21514 32224
rect 23474 32172 23480 32224
rect 23532 32172 23538 32224
rect 23768 32221 23796 32252
rect 23753 32215 23811 32221
rect 23753 32181 23765 32215
rect 23799 32181 23811 32215
rect 23753 32175 23811 32181
rect 24394 32172 24400 32224
rect 24452 32172 24458 32224
rect 1104 32122 24840 32144
rect 1104 32070 3917 32122
rect 3969 32070 3981 32122
rect 4033 32070 4045 32122
rect 4097 32070 4109 32122
rect 4161 32070 4173 32122
rect 4225 32070 9851 32122
rect 9903 32070 9915 32122
rect 9967 32070 9979 32122
rect 10031 32070 10043 32122
rect 10095 32070 10107 32122
rect 10159 32070 15785 32122
rect 15837 32070 15849 32122
rect 15901 32070 15913 32122
rect 15965 32070 15977 32122
rect 16029 32070 16041 32122
rect 16093 32070 21719 32122
rect 21771 32070 21783 32122
rect 21835 32070 21847 32122
rect 21899 32070 21911 32122
rect 21963 32070 21975 32122
rect 22027 32070 24840 32122
rect 1104 32048 24840 32070
rect 2409 32011 2467 32017
rect 2409 31977 2421 32011
rect 2455 32008 2467 32011
rect 2590 32008 2596 32020
rect 2455 31980 2596 32008
rect 2455 31977 2467 31980
rect 2409 31971 2467 31977
rect 2590 31968 2596 31980
rect 2648 31968 2654 32020
rect 6454 32008 6460 32020
rect 2976 31980 6460 32008
rect 2976 31881 3004 31980
rect 6454 31968 6460 31980
rect 6512 31968 6518 32020
rect 6546 31968 6552 32020
rect 6604 32008 6610 32020
rect 7101 32011 7159 32017
rect 7101 32008 7113 32011
rect 6604 31980 7113 32008
rect 6604 31968 6610 31980
rect 7101 31977 7113 31980
rect 7147 31977 7159 32011
rect 8481 32011 8539 32017
rect 7101 31971 7159 31977
rect 7576 31980 8432 32008
rect 7576 31940 7604 31980
rect 6840 31912 7604 31940
rect 8404 31940 8432 31980
rect 8481 31977 8493 32011
rect 8527 32008 8539 32011
rect 8754 32008 8760 32020
rect 8527 31980 8760 32008
rect 8527 31977 8539 31980
rect 8481 31971 8539 31977
rect 8754 31968 8760 31980
rect 8812 31968 8818 32020
rect 10226 31968 10232 32020
rect 10284 31968 10290 32020
rect 10778 32008 10784 32020
rect 10336 31980 10784 32008
rect 10244 31940 10272 31968
rect 10336 31949 10364 31980
rect 10778 31968 10784 31980
rect 10836 31968 10842 32020
rect 11517 32011 11575 32017
rect 11517 31977 11529 32011
rect 11563 32008 11575 32011
rect 13998 32008 14004 32020
rect 11563 31980 14004 32008
rect 11563 31977 11575 31980
rect 11517 31971 11575 31977
rect 13998 31968 14004 31980
rect 14056 31968 14062 32020
rect 14090 31968 14096 32020
rect 14148 32008 14154 32020
rect 14918 32008 14924 32020
rect 14148 31980 14924 32008
rect 14148 31968 14154 31980
rect 14918 31968 14924 31980
rect 14976 32008 14982 32020
rect 16666 32008 16672 32020
rect 14976 31980 16672 32008
rect 14976 31968 14982 31980
rect 16666 31968 16672 31980
rect 16724 31968 16730 32020
rect 17310 31968 17316 32020
rect 17368 32008 17374 32020
rect 17497 32011 17555 32017
rect 17497 32008 17509 32011
rect 17368 31980 17509 32008
rect 17368 31968 17374 31980
rect 17497 31977 17509 31980
rect 17543 31977 17555 32011
rect 17497 31971 17555 31977
rect 18414 31968 18420 32020
rect 18472 32008 18478 32020
rect 19150 32008 19156 32020
rect 18472 31980 19156 32008
rect 18472 31968 18478 31980
rect 19150 31968 19156 31980
rect 19208 31968 19214 32020
rect 21450 31968 21456 32020
rect 21508 32008 21514 32020
rect 21508 31980 22094 32008
rect 21508 31968 21514 31980
rect 8404 31912 10272 31940
rect 10321 31943 10379 31949
rect 2961 31875 3019 31881
rect 2961 31841 2973 31875
rect 3007 31841 3019 31875
rect 2961 31835 3019 31841
rect 5074 31832 5080 31884
rect 5132 31872 5138 31884
rect 5350 31872 5356 31884
rect 5132 31844 5356 31872
rect 5132 31832 5138 31844
rect 5350 31832 5356 31844
rect 5408 31872 5414 31884
rect 6089 31875 6147 31881
rect 6089 31872 6101 31875
rect 5408 31844 6101 31872
rect 5408 31832 5414 31844
rect 6089 31841 6101 31844
rect 6135 31841 6147 31875
rect 6089 31835 6147 31841
rect 1397 31807 1455 31813
rect 1397 31773 1409 31807
rect 1443 31773 1455 31807
rect 1397 31767 1455 31773
rect 1655 31777 1713 31783
rect 474 31628 480 31680
rect 532 31668 538 31680
rect 658 31668 664 31680
rect 532 31640 664 31668
rect 532 31628 538 31640
rect 658 31628 664 31640
rect 716 31628 722 31680
rect 1412 31668 1440 31767
rect 1655 31743 1667 31777
rect 1701 31774 1713 31777
rect 1701 31743 1714 31774
rect 1762 31764 1768 31816
rect 1820 31804 1826 31816
rect 1820 31776 2084 31804
rect 1820 31764 1826 31776
rect 1655 31737 1714 31743
rect 1686 31736 1714 31737
rect 2056 31736 2084 31776
rect 2774 31764 2780 31816
rect 2832 31764 2838 31816
rect 4157 31807 4215 31813
rect 4157 31773 4169 31807
rect 4203 31804 4215 31807
rect 4431 31807 4489 31813
rect 4431 31804 4443 31807
rect 4203 31776 4292 31804
rect 4203 31773 4215 31776
rect 4157 31767 4215 31773
rect 1686 31708 1900 31736
rect 2056 31708 3280 31736
rect 1578 31668 1584 31680
rect 1412 31640 1584 31668
rect 1578 31628 1584 31640
rect 1636 31668 1642 31680
rect 1762 31668 1768 31680
rect 1636 31640 1768 31668
rect 1636 31628 1642 31640
rect 1762 31628 1768 31640
rect 1820 31628 1826 31680
rect 1872 31668 1900 31708
rect 3252 31680 3280 31708
rect 2222 31668 2228 31680
rect 1872 31640 2228 31668
rect 2222 31628 2228 31640
rect 2280 31628 2286 31680
rect 3234 31628 3240 31680
rect 3292 31628 3298 31680
rect 4264 31668 4292 31776
rect 4430 31774 4443 31804
rect 4356 31773 4443 31774
rect 4477 31804 4489 31807
rect 4477 31776 4660 31804
rect 4477 31773 4489 31776
rect 4356 31767 4489 31773
rect 4356 31748 4458 31767
rect 4632 31748 4660 31776
rect 4338 31696 4344 31748
rect 4396 31746 4458 31748
rect 4396 31696 4402 31746
rect 4614 31696 4620 31748
rect 4672 31696 4678 31748
rect 4798 31736 4804 31748
rect 4724 31708 4804 31736
rect 4724 31668 4752 31708
rect 4798 31696 4804 31708
rect 4856 31736 4862 31748
rect 5092 31736 5120 31832
rect 6840 31816 6868 31912
rect 6914 31832 6920 31884
rect 6972 31872 6978 31884
rect 7466 31872 7472 31884
rect 6972 31844 7472 31872
rect 6972 31832 6978 31844
rect 7466 31832 7472 31844
rect 7524 31832 7530 31884
rect 9864 31881 9892 31912
rect 10321 31909 10333 31943
rect 10367 31909 10379 31943
rect 10321 31903 10379 31909
rect 16301 31943 16359 31949
rect 16301 31909 16313 31943
rect 16347 31940 16359 31943
rect 16390 31940 16396 31952
rect 16347 31912 16396 31940
rect 16347 31909 16359 31912
rect 16301 31903 16359 31909
rect 16390 31900 16396 31912
rect 16448 31900 16454 31952
rect 18138 31900 18144 31952
rect 18196 31940 18202 31952
rect 21358 31940 21364 31952
rect 18196 31912 21364 31940
rect 18196 31900 18202 31912
rect 21358 31900 21364 31912
rect 21416 31900 21422 31952
rect 9677 31875 9735 31881
rect 9677 31841 9689 31875
rect 9723 31872 9735 31875
rect 9861 31875 9919 31881
rect 9723 31844 9757 31872
rect 9723 31841 9735 31844
rect 9677 31835 9735 31841
rect 9861 31841 9873 31875
rect 9907 31841 9919 31875
rect 10410 31872 10416 31884
rect 9861 31835 9919 31841
rect 10060 31844 10416 31872
rect 6331 31807 6389 31813
rect 6331 31773 6343 31807
rect 6377 31773 6389 31807
rect 6331 31767 6389 31773
rect 4856 31708 5120 31736
rect 4856 31696 4862 31708
rect 6178 31696 6184 31748
rect 6236 31736 6242 31748
rect 6346 31736 6374 31767
rect 6454 31764 6460 31816
rect 6512 31804 6518 31816
rect 6512 31776 6776 31804
rect 6512 31764 6518 31776
rect 6236 31708 6374 31736
rect 6748 31736 6776 31776
rect 6822 31764 6828 31816
rect 6880 31764 6886 31816
rect 7650 31804 7656 31816
rect 7024 31776 7656 31804
rect 7024 31736 7052 31776
rect 7650 31764 7656 31776
rect 7708 31764 7714 31816
rect 7743 31807 7801 31813
rect 7743 31773 7755 31807
rect 7789 31773 7801 31807
rect 9692 31804 9720 31835
rect 10060 31804 10088 31844
rect 10410 31832 10416 31844
rect 10468 31832 10474 31884
rect 10686 31832 10692 31884
rect 10744 31881 10750 31884
rect 10744 31875 10772 31881
rect 10760 31841 10772 31875
rect 10744 31835 10772 31841
rect 10873 31875 10931 31881
rect 10873 31841 10885 31875
rect 10919 31872 10931 31875
rect 11054 31872 11060 31884
rect 10919 31844 11060 31872
rect 10919 31841 10931 31844
rect 10873 31835 10931 31841
rect 10744 31832 10750 31835
rect 11054 31832 11060 31844
rect 11112 31832 11118 31884
rect 11238 31832 11244 31884
rect 11296 31872 11302 31884
rect 11885 31875 11943 31881
rect 11885 31872 11897 31875
rect 11296 31844 11897 31872
rect 11296 31832 11302 31844
rect 11885 31841 11897 31844
rect 11931 31841 11943 31875
rect 12161 31875 12219 31881
rect 12161 31872 12173 31875
rect 11885 31835 11943 31841
rect 12084 31844 12173 31872
rect 7743 31767 7801 31773
rect 9416 31776 10088 31804
rect 6748 31708 7052 31736
rect 6236 31696 6242 31708
rect 7558 31696 7564 31748
rect 7616 31736 7622 31748
rect 7758 31736 7786 31767
rect 7616 31708 7786 31736
rect 7616 31696 7622 31708
rect 9416 31680 9444 31776
rect 10594 31764 10600 31816
rect 10652 31764 10658 31816
rect 11900 31736 11928 31835
rect 12084 31816 12112 31844
rect 12161 31841 12173 31844
rect 12207 31841 12219 31875
rect 12161 31835 12219 31841
rect 13170 31832 13176 31884
rect 13228 31872 13234 31884
rect 16577 31875 16635 31881
rect 16577 31872 16589 31875
rect 13228 31844 16589 31872
rect 13228 31832 13234 31844
rect 16577 31841 16589 31844
rect 16623 31841 16635 31875
rect 16577 31835 16635 31841
rect 16850 31832 16856 31884
rect 16908 31832 16914 31884
rect 12066 31764 12072 31816
rect 12124 31764 12130 31816
rect 12403 31797 12461 31803
rect 12403 31794 12415 31797
rect 12268 31766 12415 31794
rect 12268 31736 12296 31766
rect 12403 31763 12415 31766
rect 12449 31763 12461 31797
rect 12526 31764 12532 31816
rect 12584 31764 12590 31816
rect 15562 31764 15568 31816
rect 15620 31804 15626 31816
rect 15657 31807 15715 31813
rect 15657 31804 15669 31807
rect 15620 31776 15669 31804
rect 15620 31764 15626 31776
rect 15657 31773 15669 31776
rect 15703 31773 15715 31807
rect 15657 31767 15715 31773
rect 15841 31807 15899 31813
rect 15841 31773 15853 31807
rect 15887 31773 15899 31807
rect 15841 31767 15899 31773
rect 12403 31757 12461 31763
rect 11900 31708 12296 31736
rect 4264 31640 4752 31668
rect 5074 31628 5080 31680
rect 5132 31668 5138 31680
rect 5169 31671 5227 31677
rect 5169 31668 5181 31671
rect 5132 31640 5181 31668
rect 5132 31628 5138 31640
rect 5169 31637 5181 31640
rect 5215 31637 5227 31671
rect 5169 31631 5227 31637
rect 5902 31628 5908 31680
rect 5960 31668 5966 31680
rect 8846 31668 8852 31680
rect 5960 31640 8852 31668
rect 5960 31628 5966 31640
rect 8846 31628 8852 31640
rect 8904 31628 8910 31680
rect 9398 31628 9404 31680
rect 9456 31628 9462 31680
rect 9582 31628 9588 31680
rect 9640 31668 9646 31680
rect 11790 31668 11796 31680
rect 9640 31640 11796 31668
rect 9640 31628 9646 31640
rect 11790 31628 11796 31640
rect 11848 31628 11854 31680
rect 12066 31628 12072 31680
rect 12124 31668 12130 31680
rect 12544 31668 12572 31764
rect 12710 31696 12716 31748
rect 12768 31736 12774 31748
rect 14826 31736 14832 31748
rect 12768 31708 14832 31736
rect 12768 31696 12774 31708
rect 14826 31696 14832 31708
rect 14884 31696 14890 31748
rect 12124 31640 12572 31668
rect 13173 31671 13231 31677
rect 12124 31628 12130 31640
rect 13173 31637 13185 31671
rect 13219 31668 13231 31671
rect 13262 31668 13268 31680
rect 13219 31640 13268 31668
rect 13219 31637 13231 31640
rect 13173 31631 13231 31637
rect 13262 31628 13268 31640
rect 13320 31628 13326 31680
rect 14182 31628 14188 31680
rect 14240 31668 14246 31680
rect 15102 31668 15108 31680
rect 14240 31640 15108 31668
rect 14240 31628 14246 31640
rect 15102 31628 15108 31640
rect 15160 31628 15166 31680
rect 15856 31668 15884 31767
rect 16666 31764 16672 31816
rect 16724 31813 16730 31816
rect 16724 31807 16752 31813
rect 16740 31773 16752 31807
rect 16724 31767 16752 31773
rect 16724 31764 16730 31767
rect 17494 31764 17500 31816
rect 17552 31804 17558 31816
rect 17770 31804 17776 31816
rect 17552 31776 17776 31804
rect 17552 31764 17558 31776
rect 17770 31764 17776 31776
rect 17828 31764 17834 31816
rect 22066 31804 22094 31980
rect 23017 31943 23075 31949
rect 23017 31909 23029 31943
rect 23063 31940 23075 31943
rect 24486 31940 24492 31952
rect 23063 31912 24492 31940
rect 23063 31909 23075 31912
rect 23017 31903 23075 31909
rect 24486 31900 24492 31912
rect 24544 31900 24550 31952
rect 22373 31875 22431 31881
rect 22373 31841 22385 31875
rect 22419 31872 22431 31875
rect 23293 31875 23351 31881
rect 23293 31872 23305 31875
rect 22419 31844 22784 31872
rect 22419 31841 22431 31844
rect 22373 31835 22431 31841
rect 22756 31813 22784 31844
rect 23124 31844 23305 31872
rect 23124 31813 23152 31844
rect 23293 31841 23305 31844
rect 23339 31841 23351 31875
rect 23293 31835 23351 31841
rect 23474 31832 23480 31884
rect 23532 31872 23538 31884
rect 23532 31844 23888 31872
rect 23532 31832 23538 31844
rect 22281 31807 22339 31813
rect 22281 31804 22293 31807
rect 22066 31776 22293 31804
rect 22281 31773 22293 31776
rect 22327 31773 22339 31807
rect 22281 31767 22339 31773
rect 22741 31807 22799 31813
rect 22741 31773 22753 31807
rect 22787 31773 22799 31807
rect 22741 31767 22799 31773
rect 22925 31807 22983 31813
rect 22925 31773 22937 31807
rect 22971 31773 22983 31807
rect 22925 31767 22983 31773
rect 23109 31807 23167 31813
rect 23109 31773 23121 31807
rect 23155 31773 23167 31807
rect 23109 31767 23167 31773
rect 23201 31807 23259 31813
rect 23201 31773 23213 31807
rect 23247 31773 23259 31807
rect 23385 31807 23443 31813
rect 23385 31804 23397 31807
rect 23201 31767 23259 31773
rect 23308 31776 23397 31804
rect 22940 31736 22968 31767
rect 23216 31736 23244 31767
rect 23308 31748 23336 31776
rect 23385 31773 23397 31776
rect 23431 31773 23443 31807
rect 23566 31804 23572 31816
rect 23385 31767 23443 31773
rect 23492 31776 23572 31804
rect 22940 31708 23244 31736
rect 16758 31668 16764 31680
rect 15856 31640 16764 31668
rect 16758 31628 16764 31640
rect 16816 31628 16822 31680
rect 22830 31628 22836 31680
rect 22888 31668 22894 31680
rect 22940 31668 22968 31708
rect 23290 31696 23296 31748
rect 23348 31696 23354 31748
rect 23492 31677 23520 31776
rect 23566 31764 23572 31776
rect 23624 31764 23630 31816
rect 23658 31764 23664 31816
rect 23716 31764 23722 31816
rect 23860 31813 23888 31844
rect 23845 31807 23903 31813
rect 23845 31773 23857 31807
rect 23891 31773 23903 31807
rect 23845 31767 23903 31773
rect 24210 31764 24216 31816
rect 24268 31764 24274 31816
rect 22888 31640 22968 31668
rect 23477 31671 23535 31677
rect 22888 31628 22894 31640
rect 23477 31637 23489 31671
rect 23523 31637 23535 31671
rect 23477 31631 23535 31637
rect 1104 31578 25000 31600
rect 1104 31526 6884 31578
rect 6936 31526 6948 31578
rect 7000 31526 7012 31578
rect 7064 31526 7076 31578
rect 7128 31526 7140 31578
rect 7192 31526 12818 31578
rect 12870 31526 12882 31578
rect 12934 31526 12946 31578
rect 12998 31526 13010 31578
rect 13062 31526 13074 31578
rect 13126 31526 18752 31578
rect 18804 31526 18816 31578
rect 18868 31526 18880 31578
rect 18932 31526 18944 31578
rect 18996 31526 19008 31578
rect 19060 31526 24686 31578
rect 24738 31526 24750 31578
rect 24802 31526 24814 31578
rect 24866 31526 24878 31578
rect 24930 31526 24942 31578
rect 24994 31526 25000 31578
rect 1104 31504 25000 31526
rect 3878 31464 3884 31476
rect 3804 31436 3884 31464
rect 1118 31356 1124 31408
rect 1176 31396 1182 31408
rect 1176 31368 3556 31396
rect 1176 31356 1182 31368
rect 1489 31331 1547 31337
rect 1489 31297 1501 31331
rect 1535 31328 1547 31331
rect 1578 31328 1584 31340
rect 1535 31300 1584 31328
rect 1535 31297 1547 31300
rect 1489 31291 1547 31297
rect 1578 31288 1584 31300
rect 1636 31288 1642 31340
rect 2038 31288 2044 31340
rect 2096 31328 2102 31340
rect 2131 31331 2189 31337
rect 2131 31328 2143 31331
rect 2096 31300 2143 31328
rect 2096 31288 2102 31300
rect 2131 31297 2143 31300
rect 2177 31328 2189 31331
rect 2590 31328 2596 31340
rect 2177 31300 2596 31328
rect 2177 31297 2189 31300
rect 2131 31291 2189 31297
rect 2590 31288 2596 31300
rect 2648 31288 2654 31340
rect 3528 31337 3556 31368
rect 3804 31337 3832 31436
rect 3878 31424 3884 31436
rect 3936 31424 3942 31476
rect 3973 31467 4031 31473
rect 3973 31433 3985 31467
rect 4019 31464 4031 31467
rect 4614 31464 4620 31476
rect 4019 31436 4620 31464
rect 4019 31433 4031 31436
rect 3973 31427 4031 31433
rect 4614 31424 4620 31436
rect 4672 31424 4678 31476
rect 4724 31436 5488 31464
rect 3237 31331 3295 31337
rect 3237 31297 3249 31331
rect 3283 31297 3295 31331
rect 3237 31291 3295 31297
rect 3513 31331 3571 31337
rect 3513 31297 3525 31331
rect 3559 31297 3571 31331
rect 3513 31291 3571 31297
rect 3789 31331 3847 31337
rect 3789 31297 3801 31331
rect 3835 31297 3847 31331
rect 3789 31291 3847 31297
rect 1762 31220 1768 31272
rect 1820 31260 1826 31272
rect 1857 31263 1915 31269
rect 1857 31260 1869 31263
rect 1820 31232 1869 31260
rect 1820 31220 1826 31232
rect 1857 31229 1869 31232
rect 1903 31229 1915 31263
rect 1857 31223 1915 31229
rect 2774 31220 2780 31272
rect 2832 31260 2838 31272
rect 3252 31260 3280 31291
rect 4724 31260 4752 31436
rect 5460 31396 5488 31436
rect 5534 31424 5540 31476
rect 5592 31464 5598 31476
rect 12710 31464 12716 31476
rect 5592 31436 12716 31464
rect 5592 31424 5598 31436
rect 12710 31424 12716 31436
rect 12768 31464 12774 31476
rect 12805 31467 12863 31473
rect 12805 31464 12817 31467
rect 12768 31436 12817 31464
rect 12768 31424 12774 31436
rect 12805 31433 12817 31436
rect 12851 31433 12863 31467
rect 12805 31427 12863 31433
rect 12894 31424 12900 31476
rect 12952 31464 12958 31476
rect 12952 31436 13492 31464
rect 12952 31424 12958 31436
rect 7558 31396 7564 31408
rect 5460 31368 7564 31396
rect 7558 31356 7564 31368
rect 7616 31396 7622 31408
rect 11882 31396 11888 31408
rect 7616 31368 11888 31396
rect 7616 31356 7622 31368
rect 11882 31356 11888 31368
rect 11940 31356 11946 31408
rect 13464 31396 13492 31436
rect 14366 31424 14372 31476
rect 14424 31464 14430 31476
rect 18046 31464 18052 31476
rect 14424 31436 18052 31464
rect 14424 31424 14430 31436
rect 18046 31424 18052 31436
rect 18104 31424 18110 31476
rect 18598 31424 18604 31476
rect 18656 31464 18662 31476
rect 18656 31436 22094 31464
rect 18656 31424 18662 31436
rect 13464 31368 13584 31396
rect 4798 31288 4804 31340
rect 4856 31328 4862 31340
rect 4893 31331 4951 31337
rect 4893 31328 4905 31331
rect 4856 31300 4905 31328
rect 4856 31288 4862 31300
rect 4893 31297 4905 31300
rect 4939 31297 4951 31331
rect 4893 31291 4951 31297
rect 5167 31331 5225 31337
rect 5167 31297 5179 31331
rect 5213 31328 5225 31331
rect 5258 31328 5264 31340
rect 5213 31300 5264 31328
rect 5213 31297 5225 31300
rect 5167 31291 5225 31297
rect 5258 31288 5264 31300
rect 5316 31288 5322 31340
rect 5534 31288 5540 31340
rect 5592 31328 5598 31340
rect 5718 31328 5724 31340
rect 5592 31300 5724 31328
rect 5592 31288 5598 31300
rect 5718 31288 5724 31300
rect 5776 31288 5782 31340
rect 7466 31288 7472 31340
rect 7524 31328 7530 31340
rect 8113 31331 8171 31337
rect 8113 31328 8125 31331
rect 7524 31300 8125 31328
rect 7524 31288 7530 31300
rect 8113 31297 8125 31300
rect 8159 31297 8171 31331
rect 8113 31291 8171 31297
rect 8387 31331 8445 31337
rect 8387 31297 8399 31331
rect 8433 31328 8445 31331
rect 8433 31300 8800 31328
rect 8433 31297 8445 31300
rect 8387 31291 8445 31297
rect 2832 31232 3280 31260
rect 3620 31232 4752 31260
rect 8772 31260 8800 31300
rect 8938 31288 8944 31340
rect 8996 31328 9002 31340
rect 12894 31328 12900 31340
rect 8996 31300 12900 31328
rect 8996 31288 9002 31300
rect 12894 31288 12900 31300
rect 12952 31288 12958 31340
rect 13078 31288 13084 31340
rect 13136 31288 13142 31340
rect 13173 31331 13231 31337
rect 13173 31297 13185 31331
rect 13219 31328 13231 31331
rect 13446 31328 13452 31340
rect 13219 31300 13452 31328
rect 13219 31297 13231 31300
rect 13173 31291 13231 31297
rect 13446 31288 13452 31300
rect 13504 31288 13510 31340
rect 13556 31337 13584 31368
rect 13906 31356 13912 31408
rect 13964 31356 13970 31408
rect 22066 31396 22094 31436
rect 22830 31424 22836 31476
rect 22888 31424 22894 31476
rect 23474 31464 23480 31476
rect 22940 31436 23480 31464
rect 22940 31396 22968 31436
rect 23474 31424 23480 31436
rect 23532 31424 23538 31476
rect 23661 31467 23719 31473
rect 23661 31433 23673 31467
rect 23707 31464 23719 31467
rect 23934 31464 23940 31476
rect 23707 31436 23940 31464
rect 23707 31433 23719 31436
rect 23661 31427 23719 31433
rect 23934 31424 23940 31436
rect 23992 31424 23998 31476
rect 22066 31368 22968 31396
rect 15455 31361 15513 31367
rect 13541 31331 13599 31337
rect 13541 31297 13553 31331
rect 13587 31297 13599 31331
rect 15455 31327 15467 31361
rect 15501 31358 15513 31361
rect 15501 31328 15516 31358
rect 23014 31356 23020 31408
rect 23072 31396 23078 31408
rect 24121 31399 24179 31405
rect 24121 31396 24133 31399
rect 23072 31368 24133 31396
rect 23072 31356 23078 31368
rect 24121 31365 24133 31368
rect 24167 31365 24179 31399
rect 24121 31359 24179 31365
rect 16022 31328 16028 31340
rect 15501 31327 16028 31328
rect 15455 31321 16028 31327
rect 15488 31300 16028 31321
rect 13541 31291 13599 31297
rect 16022 31288 16028 31300
rect 16080 31288 16086 31340
rect 18138 31288 18144 31340
rect 18196 31288 18202 31340
rect 22063 31331 22121 31337
rect 22063 31297 22075 31331
rect 22109 31328 22121 31331
rect 22186 31328 22192 31340
rect 22109 31300 22192 31328
rect 22109 31297 22121 31300
rect 22063 31291 22121 31297
rect 22186 31288 22192 31300
rect 22244 31288 22250 31340
rect 23385 31331 23443 31337
rect 23385 31297 23397 31331
rect 23431 31297 23443 31331
rect 23385 31291 23443 31297
rect 23845 31331 23903 31337
rect 23845 31297 23857 31331
rect 23891 31328 23903 31331
rect 25038 31328 25044 31340
rect 23891 31300 25044 31328
rect 23891 31297 23903 31300
rect 23845 31291 23903 31297
rect 9030 31260 9036 31272
rect 8772 31232 9036 31260
rect 2832 31220 2838 31232
rect 1673 31195 1731 31201
rect 1673 31161 1685 31195
rect 1719 31161 1731 31195
rect 3620 31192 3648 31232
rect 9030 31220 9036 31232
rect 9088 31260 9094 31272
rect 12434 31260 12440 31272
rect 9088 31232 12440 31260
rect 9088 31220 9094 31232
rect 12434 31220 12440 31232
rect 12492 31220 12498 31272
rect 13262 31220 13268 31272
rect 13320 31220 13326 31272
rect 14182 31220 14188 31272
rect 14240 31260 14246 31272
rect 15197 31263 15255 31269
rect 15197 31260 15209 31263
rect 14240 31232 15209 31260
rect 14240 31220 14246 31232
rect 15197 31229 15209 31232
rect 15243 31229 15255 31263
rect 15197 31223 15255 31229
rect 19702 31220 19708 31272
rect 19760 31260 19766 31272
rect 21818 31260 21824 31272
rect 19760 31232 21824 31260
rect 19760 31220 19766 31232
rect 21818 31220 21824 31232
rect 21876 31220 21882 31272
rect 1673 31155 1731 31161
rect 2792 31164 3648 31192
rect 3697 31195 3755 31201
rect 1688 31124 1716 31155
rect 2792 31124 2820 31164
rect 3697 31161 3709 31195
rect 3743 31192 3755 31195
rect 4614 31192 4620 31204
rect 3743 31164 4620 31192
rect 3743 31161 3755 31164
rect 3697 31155 3755 31161
rect 4614 31152 4620 31164
rect 4672 31152 4678 31204
rect 6362 31192 6368 31204
rect 5552 31164 6368 31192
rect 1688 31096 2820 31124
rect 2869 31127 2927 31133
rect 2869 31093 2881 31127
rect 2915 31124 2927 31127
rect 3050 31124 3056 31136
rect 2915 31096 3056 31124
rect 2915 31093 2927 31096
rect 2869 31087 2927 31093
rect 3050 31084 3056 31096
rect 3108 31084 3114 31136
rect 3421 31127 3479 31133
rect 3421 31093 3433 31127
rect 3467 31124 3479 31127
rect 4522 31124 4528 31136
rect 3467 31096 4528 31124
rect 3467 31093 3479 31096
rect 3421 31087 3479 31093
rect 4522 31084 4528 31096
rect 4580 31084 4586 31136
rect 4798 31084 4804 31136
rect 4856 31124 4862 31136
rect 5552 31124 5580 31164
rect 6362 31152 6368 31164
rect 6420 31152 6426 31204
rect 12250 31192 12256 31204
rect 9232 31164 12256 31192
rect 9232 31136 9260 31164
rect 12250 31152 12256 31164
rect 12308 31152 12314 31204
rect 18690 31192 18696 31204
rect 16132 31164 18696 31192
rect 4856 31096 5580 31124
rect 4856 31084 4862 31096
rect 5902 31084 5908 31136
rect 5960 31084 5966 31136
rect 8570 31084 8576 31136
rect 8628 31124 8634 31136
rect 9125 31127 9183 31133
rect 9125 31124 9137 31127
rect 8628 31096 9137 31124
rect 8628 31084 8634 31096
rect 9125 31093 9137 31096
rect 9171 31093 9183 31127
rect 9125 31087 9183 31093
rect 9214 31084 9220 31136
rect 9272 31084 9278 31136
rect 9674 31084 9680 31136
rect 9732 31124 9738 31136
rect 10686 31124 10692 31136
rect 9732 31096 10692 31124
rect 9732 31084 9738 31096
rect 10686 31084 10692 31096
rect 10744 31084 10750 31136
rect 10962 31084 10968 31136
rect 11020 31124 11026 31136
rect 12618 31124 12624 31136
rect 11020 31096 12624 31124
rect 11020 31084 11026 31096
rect 12618 31084 12624 31096
rect 12676 31084 12682 31136
rect 14093 31127 14151 31133
rect 14093 31093 14105 31127
rect 14139 31124 14151 31127
rect 16132 31124 16160 31164
rect 18690 31152 18696 31164
rect 18748 31152 18754 31204
rect 23400 31192 23428 31291
rect 25038 31288 25044 31300
rect 25096 31288 25102 31340
rect 22756 31164 23428 31192
rect 14139 31096 16160 31124
rect 16209 31127 16267 31133
rect 14139 31093 14151 31096
rect 14093 31087 14151 31093
rect 16209 31093 16221 31127
rect 16255 31124 16267 31127
rect 16482 31124 16488 31136
rect 16255 31096 16488 31124
rect 16255 31093 16267 31096
rect 16209 31087 16267 31093
rect 16482 31084 16488 31096
rect 16540 31084 16546 31136
rect 17957 31127 18015 31133
rect 17957 31093 17969 31127
rect 18003 31124 18015 31127
rect 18598 31124 18604 31136
rect 18003 31096 18604 31124
rect 18003 31093 18015 31096
rect 17957 31087 18015 31093
rect 18598 31084 18604 31096
rect 18656 31084 18662 31136
rect 20530 31084 20536 31136
rect 20588 31124 20594 31136
rect 22756 31124 22784 31164
rect 20588 31096 22784 31124
rect 20588 31084 20594 31096
rect 23198 31084 23204 31136
rect 23256 31084 23262 31136
rect 24394 31084 24400 31136
rect 24452 31084 24458 31136
rect 1104 31034 24840 31056
rect 1104 30982 3917 31034
rect 3969 30982 3981 31034
rect 4033 30982 4045 31034
rect 4097 30982 4109 31034
rect 4161 30982 4173 31034
rect 4225 30982 9851 31034
rect 9903 30982 9915 31034
rect 9967 30982 9979 31034
rect 10031 30982 10043 31034
rect 10095 30982 10107 31034
rect 10159 30982 15785 31034
rect 15837 30982 15849 31034
rect 15901 30982 15913 31034
rect 15965 30982 15977 31034
rect 16029 30982 16041 31034
rect 16093 30982 21719 31034
rect 21771 30982 21783 31034
rect 21835 30982 21847 31034
rect 21899 30982 21911 31034
rect 21963 30982 21975 31034
rect 22027 30982 24840 31034
rect 1104 30960 24840 30982
rect 3602 30920 3608 30932
rect 492 30892 3608 30920
rect 492 30864 520 30892
rect 3602 30880 3608 30892
rect 3660 30880 3666 30932
rect 3973 30923 4031 30929
rect 3973 30889 3985 30923
rect 4019 30920 4031 30923
rect 4798 30920 4804 30932
rect 4019 30892 4804 30920
rect 4019 30889 4031 30892
rect 3973 30883 4031 30889
rect 4798 30880 4804 30892
rect 4856 30880 4862 30932
rect 6086 30880 6092 30932
rect 6144 30920 6150 30932
rect 6454 30920 6460 30932
rect 6144 30892 6460 30920
rect 6144 30880 6150 30892
rect 6454 30880 6460 30892
rect 6512 30880 6518 30932
rect 7374 30880 7380 30932
rect 7432 30920 7438 30932
rect 9674 30920 9680 30932
rect 7432 30892 9680 30920
rect 7432 30880 7438 30892
rect 9674 30880 9680 30892
rect 9732 30880 9738 30932
rect 10502 30920 10508 30932
rect 9766 30892 10508 30920
rect 474 30812 480 30864
rect 532 30812 538 30864
rect 3620 30784 3648 30880
rect 9766 30852 9794 30892
rect 10502 30880 10508 30892
rect 10560 30880 10566 30932
rect 12250 30880 12256 30932
rect 12308 30880 12314 30932
rect 12434 30880 12440 30932
rect 12492 30920 12498 30932
rect 12492 30892 13308 30920
rect 12492 30880 12498 30892
rect 8128 30824 9794 30852
rect 3620 30756 3832 30784
rect 1394 30676 1400 30728
rect 1452 30676 1458 30728
rect 1673 30719 1731 30725
rect 1673 30685 1685 30719
rect 1719 30685 1731 30719
rect 1673 30679 1731 30685
rect 1688 30648 1716 30679
rect 1762 30676 1768 30728
rect 1820 30716 1826 30728
rect 1946 30716 1952 30728
rect 1820 30688 1952 30716
rect 1820 30676 1826 30688
rect 1946 30676 1952 30688
rect 2004 30716 2010 30728
rect 2317 30719 2375 30725
rect 2317 30716 2329 30719
rect 2004 30688 2329 30716
rect 2004 30676 2010 30688
rect 2317 30685 2329 30688
rect 2363 30685 2375 30719
rect 2317 30679 2375 30685
rect 2498 30676 2504 30728
rect 2556 30716 2562 30728
rect 2591 30719 2649 30725
rect 2591 30716 2603 30719
rect 2556 30688 2603 30716
rect 2556 30676 2562 30688
rect 2591 30685 2603 30688
rect 2637 30716 2649 30719
rect 2682 30716 2688 30728
rect 2637 30688 2688 30716
rect 2637 30685 2649 30688
rect 2591 30679 2649 30685
rect 2682 30676 2688 30688
rect 2740 30676 2746 30728
rect 3804 30725 3832 30756
rect 5074 30744 5080 30796
rect 5132 30744 5138 30796
rect 5902 30744 5908 30796
rect 5960 30744 5966 30796
rect 7466 30744 7472 30796
rect 7524 30744 7530 30796
rect 3789 30719 3847 30725
rect 3789 30685 3801 30719
rect 3835 30685 3847 30719
rect 3789 30679 3847 30685
rect 3970 30676 3976 30728
rect 4028 30716 4034 30728
rect 4890 30716 4896 30728
rect 4028 30688 4896 30716
rect 4028 30676 4034 30688
rect 4890 30676 4896 30688
rect 4948 30676 4954 30728
rect 5169 30719 5227 30725
rect 5169 30685 5181 30719
rect 5215 30712 5227 30719
rect 5920 30716 5948 30744
rect 5276 30712 5948 30716
rect 5215 30688 5948 30712
rect 5215 30685 5304 30688
rect 5169 30684 5304 30685
rect 5169 30679 5227 30684
rect 7282 30676 7288 30728
rect 7340 30716 7346 30728
rect 7711 30719 7769 30725
rect 7711 30716 7723 30719
rect 7340 30688 7723 30716
rect 7340 30676 7346 30688
rect 7711 30685 7723 30688
rect 7757 30685 7769 30719
rect 8128 30716 8156 30824
rect 9950 30744 9956 30796
rect 10008 30784 10014 30796
rect 10045 30787 10103 30793
rect 10045 30784 10057 30787
rect 10008 30756 10057 30784
rect 10008 30744 10014 30756
rect 10045 30753 10057 30756
rect 10091 30753 10103 30787
rect 10045 30747 10103 30753
rect 7711 30679 7769 30685
rect 7852 30688 8156 30716
rect 1688 30620 5028 30648
rect 3326 30540 3332 30592
rect 3384 30540 3390 30592
rect 3510 30540 3516 30592
rect 3568 30580 3574 30592
rect 4062 30580 4068 30592
rect 3568 30552 4068 30580
rect 3568 30540 3574 30552
rect 4062 30540 4068 30552
rect 4120 30540 4126 30592
rect 4798 30540 4804 30592
rect 4856 30540 4862 30592
rect 5000 30580 5028 30620
rect 5074 30608 5080 30660
rect 5132 30608 5138 30660
rect 5537 30651 5595 30657
rect 5537 30617 5549 30651
rect 5583 30648 5595 30651
rect 5718 30648 5724 30660
rect 5583 30620 5724 30648
rect 5583 30617 5595 30620
rect 5537 30611 5595 30617
rect 5718 30608 5724 30620
rect 5776 30608 5782 30660
rect 7852 30648 7880 30688
rect 8662 30676 8668 30728
rect 8720 30716 8726 30728
rect 10319 30719 10377 30725
rect 10319 30716 10331 30719
rect 8720 30688 10331 30716
rect 8720 30676 8726 30688
rect 10319 30685 10331 30688
rect 10365 30716 10377 30719
rect 11698 30716 11704 30728
rect 10365 30688 11704 30716
rect 10365 30685 10377 30688
rect 10319 30679 10377 30685
rect 11698 30676 11704 30688
rect 11756 30676 11762 30728
rect 12268 30716 12296 30880
rect 13280 30852 13308 30892
rect 13446 30880 13452 30932
rect 13504 30920 13510 30932
rect 13633 30923 13691 30929
rect 13633 30920 13645 30923
rect 13504 30892 13645 30920
rect 13504 30880 13510 30892
rect 13633 30889 13645 30892
rect 13679 30889 13691 30923
rect 13633 30883 13691 30889
rect 14826 30880 14832 30932
rect 14884 30920 14890 30932
rect 16298 30920 16304 30932
rect 14884 30892 16304 30920
rect 14884 30880 14890 30892
rect 16298 30880 16304 30892
rect 16356 30880 16362 30932
rect 18598 30880 18604 30932
rect 18656 30880 18662 30932
rect 23014 30880 23020 30932
rect 23072 30880 23078 30932
rect 23198 30880 23204 30932
rect 23256 30880 23262 30932
rect 23293 30923 23351 30929
rect 23293 30889 23305 30923
rect 23339 30920 23351 30923
rect 23382 30920 23388 30932
rect 23339 30892 23388 30920
rect 23339 30889 23351 30892
rect 23293 30883 23351 30889
rect 23382 30880 23388 30892
rect 23440 30880 23446 30932
rect 13280 30824 13492 30852
rect 13464 30796 13492 30824
rect 15580 30824 16068 30852
rect 15580 30796 15608 30824
rect 12526 30744 12532 30796
rect 12584 30784 12590 30796
rect 12621 30787 12679 30793
rect 12621 30784 12633 30787
rect 12584 30756 12633 30784
rect 12584 30744 12590 30756
rect 12621 30753 12633 30756
rect 12667 30753 12679 30787
rect 12621 30747 12679 30753
rect 13446 30744 13452 30796
rect 13504 30784 13510 30796
rect 13814 30784 13820 30796
rect 13504 30756 13820 30784
rect 13504 30744 13510 30756
rect 13814 30744 13820 30756
rect 13872 30744 13878 30796
rect 14458 30744 14464 30796
rect 14516 30784 14522 30796
rect 15010 30784 15016 30796
rect 14516 30756 15016 30784
rect 14516 30744 14522 30756
rect 15010 30744 15016 30756
rect 15068 30744 15074 30796
rect 15562 30744 15568 30796
rect 15620 30744 15626 30796
rect 15930 30744 15936 30796
rect 15988 30744 15994 30796
rect 16040 30784 16068 30824
rect 16209 30787 16267 30793
rect 16209 30784 16221 30787
rect 16040 30756 16221 30784
rect 16209 30753 16221 30756
rect 16255 30753 16267 30787
rect 16209 30747 16267 30753
rect 16298 30744 16304 30796
rect 16356 30793 16362 30796
rect 16356 30787 16384 30793
rect 16372 30753 16384 30787
rect 16356 30747 16384 30753
rect 16356 30744 16362 30747
rect 16482 30744 16488 30796
rect 16540 30744 16546 30796
rect 17494 30744 17500 30796
rect 17552 30744 17558 30796
rect 12863 30719 12921 30725
rect 12863 30716 12875 30719
rect 12268 30688 12875 30716
rect 12863 30685 12875 30688
rect 12909 30685 12921 30719
rect 12863 30679 12921 30685
rect 14734 30676 14740 30728
rect 14792 30676 14798 30728
rect 15286 30676 15292 30728
rect 15344 30676 15350 30728
rect 15470 30676 15476 30728
rect 15528 30716 15534 30728
rect 15654 30716 15660 30728
rect 15528 30688 15660 30716
rect 15528 30676 15534 30688
rect 15654 30676 15660 30688
rect 15712 30676 15718 30728
rect 17129 30719 17187 30725
rect 17129 30685 17141 30719
rect 17175 30716 17187 30719
rect 17764 30719 17822 30725
rect 17764 30716 17776 30719
rect 17175 30688 17776 30716
rect 17175 30685 17187 30688
rect 17129 30679 17187 30685
rect 17764 30685 17776 30688
rect 17810 30716 17822 30719
rect 18138 30716 18144 30728
rect 17810 30688 18144 30716
rect 17810 30685 17822 30688
rect 17764 30679 17822 30685
rect 18138 30676 18144 30688
rect 18196 30676 18202 30728
rect 18616 30716 18644 30880
rect 18877 30855 18935 30861
rect 18877 30821 18889 30855
rect 18923 30821 18935 30855
rect 18877 30815 18935 30821
rect 18892 30784 18920 30815
rect 18966 30812 18972 30864
rect 19024 30852 19030 30864
rect 20070 30852 20076 30864
rect 19024 30824 20076 30852
rect 19024 30812 19030 30824
rect 20070 30812 20076 30824
rect 20128 30812 20134 30864
rect 23216 30784 23244 30880
rect 18892 30756 20024 30784
rect 23216 30756 23520 30784
rect 19996 30725 20024 30756
rect 19245 30719 19303 30725
rect 19245 30716 19257 30719
rect 18616 30688 19257 30716
rect 19245 30685 19257 30688
rect 19291 30685 19303 30719
rect 19245 30679 19303 30685
rect 19521 30719 19579 30725
rect 19521 30685 19533 30719
rect 19567 30685 19579 30719
rect 19521 30679 19579 30685
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30716 19763 30719
rect 19981 30719 20039 30725
rect 19751 30688 19840 30716
rect 19751 30685 19763 30688
rect 19705 30679 19763 30685
rect 8938 30648 8944 30660
rect 5828 30620 7328 30648
rect 5828 30580 5856 30620
rect 5000 30552 5856 30580
rect 5902 30540 5908 30592
rect 5960 30540 5966 30592
rect 7300 30580 7328 30620
rect 7484 30620 7880 30648
rect 7944 30620 8944 30648
rect 7484 30580 7512 30620
rect 7944 30592 7972 30620
rect 8938 30608 8944 30620
rect 8996 30608 9002 30660
rect 9030 30608 9036 30660
rect 9088 30648 9094 30660
rect 11517 30651 11575 30657
rect 11517 30648 11529 30651
rect 9088 30620 11529 30648
rect 9088 30608 9094 30620
rect 11517 30617 11529 30620
rect 11563 30648 11575 30651
rect 14752 30648 14780 30676
rect 11563 30620 14780 30648
rect 11563 30617 11575 30620
rect 11517 30611 11575 30617
rect 18966 30608 18972 30660
rect 19024 30608 19030 30660
rect 19536 30648 19564 30679
rect 19260 30620 19564 30648
rect 7300 30552 7512 30580
rect 7558 30540 7564 30592
rect 7616 30580 7622 30592
rect 7742 30580 7748 30592
rect 7616 30552 7748 30580
rect 7616 30540 7622 30552
rect 7742 30540 7748 30552
rect 7800 30540 7806 30592
rect 7926 30540 7932 30592
rect 7984 30540 7990 30592
rect 8110 30540 8116 30592
rect 8168 30580 8174 30592
rect 8481 30583 8539 30589
rect 8481 30580 8493 30583
rect 8168 30552 8493 30580
rect 8168 30540 8174 30552
rect 8481 30549 8493 30552
rect 8527 30549 8539 30583
rect 8481 30543 8539 30549
rect 9490 30540 9496 30592
rect 9548 30580 9554 30592
rect 10502 30580 10508 30592
rect 9548 30552 10508 30580
rect 9548 30540 9554 30552
rect 10502 30540 10508 30552
rect 10560 30540 10566 30592
rect 11054 30540 11060 30592
rect 11112 30540 11118 30592
rect 11606 30540 11612 30592
rect 11664 30540 11670 30592
rect 14826 30540 14832 30592
rect 14884 30580 14890 30592
rect 18984 30580 19012 30608
rect 19260 30592 19288 30620
rect 14884 30552 19012 30580
rect 14884 30540 14890 30552
rect 19242 30540 19248 30592
rect 19300 30540 19306 30592
rect 19334 30540 19340 30592
rect 19392 30540 19398 30592
rect 19610 30540 19616 30592
rect 19668 30540 19674 30592
rect 19812 30589 19840 30688
rect 19981 30685 19993 30719
rect 20027 30685 20039 30719
rect 19981 30679 20039 30685
rect 20901 30719 20959 30725
rect 20901 30685 20913 30719
rect 20947 30685 20959 30719
rect 20901 30679 20959 30685
rect 21085 30719 21143 30725
rect 21085 30685 21097 30719
rect 21131 30716 21143 30719
rect 21450 30716 21456 30728
rect 21131 30688 21456 30716
rect 21131 30685 21143 30688
rect 21085 30679 21143 30685
rect 20916 30592 20944 30679
rect 21450 30676 21456 30688
rect 21508 30676 21514 30728
rect 23198 30676 23204 30728
rect 23256 30676 23262 30728
rect 23492 30725 23520 30756
rect 23477 30719 23535 30725
rect 23477 30685 23489 30719
rect 23523 30685 23535 30719
rect 23477 30679 23535 30685
rect 23842 30608 23848 30660
rect 23900 30608 23906 30660
rect 24210 30608 24216 30660
rect 24268 30608 24274 30660
rect 19797 30583 19855 30589
rect 19797 30549 19809 30583
rect 19843 30549 19855 30583
rect 19797 30543 19855 30549
rect 20346 30540 20352 30592
rect 20404 30580 20410 30592
rect 20806 30580 20812 30592
rect 20404 30552 20812 30580
rect 20404 30540 20410 30552
rect 20806 30540 20812 30552
rect 20864 30540 20870 30592
rect 20898 30540 20904 30592
rect 20956 30540 20962 30592
rect 21082 30540 21088 30592
rect 21140 30540 21146 30592
rect 22830 30540 22836 30592
rect 22888 30580 22894 30592
rect 23566 30580 23572 30592
rect 22888 30552 23572 30580
rect 22888 30540 22894 30552
rect 23566 30540 23572 30552
rect 23624 30540 23630 30592
rect 1104 30490 25000 30512
rect 1104 30438 6884 30490
rect 6936 30438 6948 30490
rect 7000 30438 7012 30490
rect 7064 30438 7076 30490
rect 7128 30438 7140 30490
rect 7192 30438 12818 30490
rect 12870 30438 12882 30490
rect 12934 30438 12946 30490
rect 12998 30438 13010 30490
rect 13062 30438 13074 30490
rect 13126 30438 18752 30490
rect 18804 30438 18816 30490
rect 18868 30438 18880 30490
rect 18932 30438 18944 30490
rect 18996 30438 19008 30490
rect 19060 30438 24686 30490
rect 24738 30438 24750 30490
rect 24802 30438 24814 30490
rect 24866 30438 24878 30490
rect 24930 30438 24942 30490
rect 24994 30438 25000 30490
rect 1104 30416 25000 30438
rect 1302 30336 1308 30388
rect 1360 30376 1366 30388
rect 2774 30376 2780 30388
rect 1360 30348 2780 30376
rect 1360 30336 1366 30348
rect 2774 30336 2780 30348
rect 2832 30336 2838 30388
rect 3326 30376 3332 30388
rect 3252 30348 3332 30376
rect 2682 30268 2688 30320
rect 2740 30268 2746 30320
rect 3053 30311 3111 30317
rect 3053 30277 3065 30311
rect 3099 30308 3111 30311
rect 3252 30308 3280 30348
rect 3326 30336 3332 30348
rect 3384 30336 3390 30388
rect 3970 30336 3976 30388
rect 4028 30336 4034 30388
rect 4172 30348 4844 30376
rect 3789 30311 3847 30317
rect 3789 30308 3801 30311
rect 3099 30280 3280 30308
rect 3344 30280 3801 30308
rect 3099 30277 3111 30280
rect 3053 30271 3111 30277
rect 1397 30243 1455 30249
rect 1397 30209 1409 30243
rect 1443 30240 1455 30243
rect 1486 30240 1492 30252
rect 1443 30212 1492 30240
rect 1443 30209 1455 30212
rect 1397 30203 1455 30209
rect 1486 30200 1492 30212
rect 1544 30200 1550 30252
rect 1670 30200 1676 30252
rect 1728 30240 1734 30252
rect 2041 30243 2099 30249
rect 2041 30240 2053 30243
rect 1728 30212 2053 30240
rect 1728 30200 1734 30212
rect 2041 30209 2053 30212
rect 2087 30209 2099 30243
rect 2041 30203 2099 30209
rect 2774 30200 2780 30252
rect 2832 30240 2838 30252
rect 2961 30243 3019 30249
rect 2961 30240 2973 30243
rect 2832 30212 2973 30240
rect 2832 30200 2838 30212
rect 2961 30209 2973 30212
rect 3007 30209 3019 30243
rect 2961 30203 3019 30209
rect 3234 30200 3240 30252
rect 3292 30240 3298 30252
rect 3344 30240 3372 30280
rect 3789 30277 3801 30280
rect 3835 30277 3847 30311
rect 3789 30271 3847 30277
rect 3292 30212 3372 30240
rect 3292 30200 3298 30212
rect 3418 30200 3424 30252
rect 3476 30238 3482 30252
rect 4172 30240 4200 30348
rect 4246 30268 4252 30320
rect 4304 30308 4310 30320
rect 4816 30308 4844 30348
rect 6178 30336 6184 30388
rect 6236 30376 6242 30388
rect 8018 30376 8024 30388
rect 6236 30348 8024 30376
rect 6236 30336 6242 30348
rect 7944 30317 7972 30348
rect 8018 30336 8024 30348
rect 8076 30336 8082 30388
rect 9674 30336 9680 30388
rect 9732 30376 9738 30388
rect 15565 30379 15623 30385
rect 9732 30348 14136 30376
rect 9732 30336 9738 30348
rect 7929 30311 7987 30317
rect 4304 30280 4752 30308
rect 4816 30280 7236 30308
rect 4304 30268 4310 30280
rect 3528 30238 4200 30240
rect 3476 30212 4200 30238
rect 4617 30243 4675 30249
rect 3476 30210 3556 30212
rect 3476 30200 3482 30210
rect 4617 30209 4629 30243
rect 4663 30209 4675 30243
rect 4724 30240 4752 30280
rect 5166 30249 5172 30252
rect 5135 30243 5172 30249
rect 5135 30240 5147 30243
rect 4724 30212 5147 30240
rect 4617 30203 4675 30209
rect 5135 30209 5147 30212
rect 5135 30203 5172 30209
rect 1578 30132 1584 30184
rect 1636 30132 1642 30184
rect 2130 30132 2136 30184
rect 2188 30132 2194 30184
rect 3050 30132 3056 30184
rect 3108 30132 3114 30184
rect 4632 30172 4660 30203
rect 5166 30200 5172 30203
rect 5224 30200 5230 30252
rect 5534 30200 5540 30252
rect 5592 30240 5598 30252
rect 6270 30240 6276 30252
rect 5592 30212 6276 30240
rect 5592 30200 5598 30212
rect 6270 30200 6276 30212
rect 6328 30240 6334 30252
rect 6607 30243 6665 30249
rect 6607 30240 6619 30243
rect 6328 30212 6619 30240
rect 6328 30200 6334 30212
rect 6607 30209 6619 30212
rect 6653 30209 6665 30243
rect 6607 30203 6665 30209
rect 4893 30175 4951 30181
rect 4632 30144 4752 30172
rect 1486 30064 1492 30116
rect 1544 30104 1550 30116
rect 2148 30104 2176 30132
rect 1544 30076 2176 30104
rect 1544 30064 1550 30076
rect 4724 30048 4752 30144
rect 4893 30141 4905 30175
rect 4939 30141 4951 30175
rect 6178 30172 6184 30184
rect 4893 30135 4951 30141
rect 5552 30144 6184 30172
rect 4798 30064 4804 30116
rect 4856 30064 4862 30116
rect 2130 29996 2136 30048
rect 2188 29996 2194 30048
rect 4706 29996 4712 30048
rect 4764 29996 4770 30048
rect 4908 30036 4936 30135
rect 5350 30036 5356 30048
rect 4908 30008 5356 30036
rect 5350 29996 5356 30008
rect 5408 30036 5414 30048
rect 5552 30036 5580 30144
rect 6178 30132 6184 30144
rect 6236 30172 6242 30184
rect 6365 30175 6423 30181
rect 6365 30172 6377 30175
rect 6236 30144 6377 30172
rect 6236 30132 6242 30144
rect 6365 30141 6377 30144
rect 6411 30141 6423 30175
rect 6365 30135 6423 30141
rect 7208 30104 7236 30280
rect 7929 30277 7941 30311
rect 7975 30277 7987 30311
rect 7929 30271 7987 30277
rect 8202 30268 8208 30320
rect 8260 30268 8266 30320
rect 8297 30311 8355 30317
rect 8297 30277 8309 30311
rect 8343 30308 8355 30311
rect 8570 30308 8576 30320
rect 8343 30280 8576 30308
rect 8343 30277 8355 30280
rect 8297 30271 8355 30277
rect 8570 30268 8576 30280
rect 8628 30268 8634 30320
rect 9030 30268 9036 30320
rect 9088 30268 9094 30320
rect 11514 30268 11520 30320
rect 11572 30308 11578 30320
rect 12713 30311 12771 30317
rect 12713 30308 12725 30311
rect 11572 30280 12725 30308
rect 11572 30268 11578 30280
rect 12713 30277 12725 30280
rect 12759 30308 12771 30311
rect 14108 30308 14136 30348
rect 15565 30345 15577 30379
rect 15611 30376 15623 30379
rect 15930 30376 15936 30388
rect 15611 30348 15936 30376
rect 15611 30345 15623 30348
rect 15565 30339 15623 30345
rect 15930 30336 15936 30348
rect 15988 30336 15994 30388
rect 18969 30379 19027 30385
rect 18156 30348 18368 30376
rect 17310 30308 17316 30320
rect 12759 30280 13400 30308
rect 14108 30280 14688 30308
rect 12759 30277 12771 30280
rect 12713 30271 12771 30277
rect 7650 30200 7656 30252
rect 7708 30240 7714 30252
rect 8220 30240 8248 30268
rect 7708 30212 8248 30240
rect 7708 30200 7714 30212
rect 8662 30200 8668 30252
rect 8720 30200 8726 30252
rect 8846 30200 8852 30252
rect 8904 30240 8910 30252
rect 9493 30243 9551 30249
rect 9493 30240 9505 30243
rect 8904 30212 9505 30240
rect 8904 30200 8910 30212
rect 9493 30209 9505 30212
rect 9539 30209 9551 30243
rect 9858 30240 9864 30252
rect 9493 30203 9551 30209
rect 9600 30212 9864 30240
rect 8110 30132 8116 30184
rect 8168 30132 8174 30184
rect 9030 30132 9036 30184
rect 9088 30172 9094 30184
rect 9600 30172 9628 30212
rect 9858 30200 9864 30212
rect 9916 30200 9922 30252
rect 10413 30243 10471 30249
rect 10413 30209 10425 30243
rect 10459 30238 10471 30243
rect 10459 30209 10474 30238
rect 10413 30203 10474 30209
rect 9088 30144 9628 30172
rect 9088 30132 9094 30144
rect 9674 30132 9680 30184
rect 9732 30132 9738 30184
rect 10042 30132 10048 30184
rect 10100 30172 10106 30184
rect 10446 30172 10474 30203
rect 12066 30200 12072 30252
rect 12124 30200 12130 30252
rect 12253 30243 12311 30249
rect 12253 30209 12265 30243
rect 12299 30209 12311 30243
rect 12253 30203 12311 30209
rect 10100 30144 10474 30172
rect 10100 30132 10106 30144
rect 10502 30132 10508 30184
rect 10560 30181 10566 30184
rect 10560 30175 10588 30181
rect 10576 30141 10588 30175
rect 10560 30135 10588 30141
rect 10689 30175 10747 30181
rect 10689 30141 10701 30175
rect 10735 30172 10747 30175
rect 11054 30172 11060 30184
rect 10735 30144 11060 30172
rect 10735 30141 10747 30144
rect 10689 30135 10747 30141
rect 10560 30132 10566 30135
rect 11054 30132 11060 30144
rect 11112 30132 11118 30184
rect 12268 30172 12296 30203
rect 11900 30144 12296 30172
rect 10137 30107 10195 30113
rect 7208 30076 7972 30104
rect 7944 30048 7972 30076
rect 10137 30073 10149 30107
rect 10183 30104 10195 30107
rect 10226 30104 10232 30116
rect 10183 30076 10232 30104
rect 10183 30073 10195 30076
rect 10137 30067 10195 30073
rect 10226 30064 10232 30076
rect 10284 30064 10290 30116
rect 11900 30113 11928 30144
rect 11885 30107 11943 30113
rect 11885 30073 11897 30107
rect 11931 30073 11943 30107
rect 11885 30067 11943 30073
rect 12897 30107 12955 30113
rect 12897 30073 12909 30107
rect 12943 30073 12955 30107
rect 13372 30104 13400 30280
rect 14660 30240 14688 30280
rect 16868 30280 17316 30308
rect 14827 30243 14885 30249
rect 14827 30240 14839 30243
rect 14660 30212 14839 30240
rect 14827 30209 14839 30212
rect 14873 30240 14885 30243
rect 16868 30240 16896 30280
rect 17310 30268 17316 30280
rect 17368 30308 17374 30320
rect 18156 30308 18184 30348
rect 17368 30280 18184 30308
rect 18340 30308 18368 30348
rect 18969 30345 18981 30379
rect 19015 30376 19027 30379
rect 19242 30376 19248 30388
rect 19015 30348 19248 30376
rect 19015 30345 19027 30348
rect 18969 30339 19027 30345
rect 19242 30336 19248 30348
rect 19300 30336 19306 30388
rect 20717 30379 20775 30385
rect 20717 30345 20729 30379
rect 20763 30345 20775 30379
rect 20717 30339 20775 30345
rect 20438 30308 20444 30320
rect 18340 30280 20444 30308
rect 17368 30268 17374 30280
rect 20438 30268 20444 30280
rect 20496 30268 20502 30320
rect 20732 30308 20760 30339
rect 21450 30336 21456 30388
rect 21508 30336 21514 30388
rect 23566 30336 23572 30388
rect 23624 30336 23630 30388
rect 20732 30280 21680 30308
rect 14873 30212 16896 30240
rect 14873 30209 14885 30212
rect 14827 30203 14885 30209
rect 17954 30200 17960 30252
rect 18012 30200 18018 30252
rect 18230 30200 18236 30252
rect 18288 30200 18294 30252
rect 19058 30200 19064 30252
rect 19116 30240 19122 30252
rect 19593 30243 19651 30249
rect 19593 30240 19605 30243
rect 19116 30212 19605 30240
rect 19116 30200 19122 30212
rect 19593 30209 19605 30212
rect 19639 30209 19651 30243
rect 19593 30203 19651 30209
rect 20809 30243 20867 30249
rect 20809 30209 20821 30243
rect 20855 30240 20867 30243
rect 20898 30240 20904 30252
rect 20855 30212 20904 30240
rect 20855 30209 20867 30212
rect 20809 30203 20867 30209
rect 20898 30200 20904 30212
rect 20956 30200 20962 30252
rect 21082 30198 21088 30250
rect 21140 30198 21146 30250
rect 21174 30200 21180 30252
rect 21232 30200 21238 30252
rect 21652 30249 21680 30280
rect 22830 30268 22836 30320
rect 22888 30268 22894 30320
rect 24121 30311 24179 30317
rect 24121 30308 24133 30311
rect 23400 30280 24133 30308
rect 21637 30243 21695 30249
rect 21637 30209 21649 30243
rect 21683 30209 21695 30243
rect 21637 30203 21695 30209
rect 22649 30243 22707 30249
rect 22649 30209 22661 30243
rect 22695 30240 22707 30243
rect 22848 30240 22876 30268
rect 23400 30252 23428 30280
rect 24121 30277 24133 30280
rect 24167 30277 24179 30311
rect 24121 30271 24179 30277
rect 22695 30212 22876 30240
rect 22925 30243 22983 30249
rect 22695 30209 22707 30212
rect 22649 30203 22707 30209
rect 22925 30209 22937 30243
rect 22971 30209 22983 30243
rect 22925 30203 22983 30209
rect 14182 30132 14188 30184
rect 14240 30172 14246 30184
rect 14553 30175 14611 30181
rect 14553 30172 14565 30175
rect 14240 30144 14565 30172
rect 14240 30132 14246 30144
rect 14553 30141 14565 30144
rect 14599 30141 14611 30175
rect 14553 30135 14611 30141
rect 19337 30175 19395 30181
rect 19337 30141 19349 30175
rect 19383 30141 19395 30175
rect 21085 30171 21097 30198
rect 21131 30171 21143 30198
rect 21085 30165 21143 30171
rect 19337 30135 19395 30141
rect 14458 30104 14464 30116
rect 13372 30076 14464 30104
rect 12897 30067 12955 30073
rect 5408 30008 5580 30036
rect 5408 29996 5414 30008
rect 5902 29996 5908 30048
rect 5960 29996 5966 30048
rect 7374 29996 7380 30048
rect 7432 29996 7438 30048
rect 7926 29996 7932 30048
rect 7984 29996 7990 30048
rect 9214 29996 9220 30048
rect 9272 29996 9278 30048
rect 11330 29996 11336 30048
rect 11388 29996 11394 30048
rect 12345 30039 12403 30045
rect 12345 30005 12357 30039
rect 12391 30036 12403 30039
rect 12710 30036 12716 30048
rect 12391 30008 12716 30036
rect 12391 30005 12403 30008
rect 12345 29999 12403 30005
rect 12710 29996 12716 30008
rect 12768 29996 12774 30048
rect 12912 30036 12940 30067
rect 14458 30064 14464 30076
rect 14516 30064 14522 30116
rect 15396 30076 18092 30104
rect 15396 30036 15424 30076
rect 12912 30008 15424 30036
rect 15470 29996 15476 30048
rect 15528 30036 15534 30048
rect 17954 30036 17960 30048
rect 15528 30008 17960 30036
rect 15528 29996 15534 30008
rect 17954 29996 17960 30008
rect 18012 29996 18018 30048
rect 18064 30036 18092 30076
rect 18230 30036 18236 30048
rect 18064 30008 18236 30036
rect 18230 29996 18236 30008
rect 18288 29996 18294 30048
rect 19352 30036 19380 30135
rect 20901 30107 20959 30113
rect 20901 30073 20913 30107
rect 20947 30104 20959 30107
rect 21269 30107 21327 30113
rect 21269 30104 21281 30107
rect 20947 30076 21281 30104
rect 20947 30073 20959 30076
rect 20901 30067 20959 30073
rect 21269 30073 21281 30076
rect 21315 30073 21327 30107
rect 22948 30104 22976 30203
rect 23014 30200 23020 30252
rect 23072 30240 23078 30252
rect 23201 30243 23259 30249
rect 23201 30240 23213 30243
rect 23072 30212 23213 30240
rect 23072 30200 23078 30212
rect 23201 30209 23213 30212
rect 23247 30209 23259 30243
rect 23201 30203 23259 30209
rect 23382 30200 23388 30252
rect 23440 30200 23446 30252
rect 23477 30243 23535 30249
rect 23477 30209 23489 30243
rect 23523 30209 23535 30243
rect 23477 30203 23535 30209
rect 23492 30172 23520 30203
rect 23566 30200 23572 30252
rect 23624 30240 23630 30252
rect 23753 30243 23811 30249
rect 23753 30240 23765 30243
rect 23624 30212 23765 30240
rect 23624 30200 23630 30212
rect 23753 30209 23765 30212
rect 23799 30209 23811 30243
rect 23753 30203 23811 30209
rect 23216 30144 23520 30172
rect 23017 30107 23075 30113
rect 23017 30104 23029 30107
rect 22948 30076 23029 30104
rect 21269 30067 21327 30073
rect 23017 30073 23029 30076
rect 23063 30073 23075 30107
rect 23017 30067 23075 30073
rect 20622 30036 20628 30048
rect 19352 30008 20628 30036
rect 20622 29996 20628 30008
rect 20680 29996 20686 30048
rect 20990 29996 20996 30048
rect 21048 29996 21054 30048
rect 22465 30039 22523 30045
rect 22465 30005 22477 30039
rect 22511 30036 22523 30039
rect 22554 30036 22560 30048
rect 22511 30008 22560 30036
rect 22511 30005 22523 30008
rect 22465 29999 22523 30005
rect 22554 29996 22560 30008
rect 22612 29996 22618 30048
rect 22741 30039 22799 30045
rect 22741 30005 22753 30039
rect 22787 30036 22799 30039
rect 23216 30036 23244 30144
rect 22787 30008 23244 30036
rect 23293 30039 23351 30045
rect 22787 30005 22799 30008
rect 22741 29999 22799 30005
rect 23293 30005 23305 30039
rect 23339 30036 23351 30039
rect 23842 30036 23848 30048
rect 23339 30008 23848 30036
rect 23339 30005 23351 30008
rect 23293 29999 23351 30005
rect 23842 29996 23848 30008
rect 23900 29996 23906 30048
rect 24394 29996 24400 30048
rect 24452 29996 24458 30048
rect 1104 29946 24840 29968
rect 1104 29894 3917 29946
rect 3969 29894 3981 29946
rect 4033 29894 4045 29946
rect 4097 29894 4109 29946
rect 4161 29894 4173 29946
rect 4225 29894 9851 29946
rect 9903 29894 9915 29946
rect 9967 29894 9979 29946
rect 10031 29894 10043 29946
rect 10095 29894 10107 29946
rect 10159 29894 15785 29946
rect 15837 29894 15849 29946
rect 15901 29894 15913 29946
rect 15965 29894 15977 29946
rect 16029 29894 16041 29946
rect 16093 29894 21719 29946
rect 21771 29894 21783 29946
rect 21835 29894 21847 29946
rect 21899 29894 21911 29946
rect 21963 29894 21975 29946
rect 22027 29894 24840 29946
rect 1104 29872 24840 29894
rect 1946 29832 1952 29844
rect 1504 29804 1952 29832
rect 1394 29588 1400 29640
rect 1452 29628 1458 29640
rect 1504 29637 1532 29804
rect 1946 29792 1952 29804
rect 2004 29792 2010 29844
rect 2314 29792 2320 29844
rect 2372 29792 2378 29844
rect 2406 29792 2412 29844
rect 2464 29792 2470 29844
rect 3513 29835 3571 29841
rect 3513 29801 3525 29835
rect 3559 29832 3571 29835
rect 3602 29832 3608 29844
rect 3559 29804 3608 29832
rect 3559 29801 3571 29804
rect 3513 29795 3571 29801
rect 3602 29792 3608 29804
rect 3660 29832 3666 29844
rect 3786 29832 3792 29844
rect 3660 29804 3792 29832
rect 3660 29792 3666 29804
rect 3786 29792 3792 29804
rect 3844 29792 3850 29844
rect 11514 29832 11520 29844
rect 3896 29804 5764 29832
rect 1489 29631 1547 29637
rect 1489 29628 1501 29631
rect 1452 29600 1501 29628
rect 1452 29588 1458 29600
rect 1489 29597 1501 29600
rect 1535 29597 1547 29631
rect 1489 29591 1547 29597
rect 1763 29631 1821 29637
rect 1763 29597 1775 29631
rect 1809 29628 1821 29631
rect 2222 29628 2228 29640
rect 1809 29600 2228 29628
rect 1809 29597 1821 29600
rect 1763 29591 1821 29597
rect 2222 29588 2228 29600
rect 2280 29628 2286 29640
rect 2332 29628 2360 29792
rect 2424 29696 2452 29792
rect 2682 29724 2688 29776
rect 2740 29764 2746 29776
rect 3896 29764 3924 29804
rect 2740 29736 3924 29764
rect 3973 29767 4031 29773
rect 2740 29724 2746 29736
rect 3973 29733 3985 29767
rect 4019 29733 4031 29767
rect 3973 29727 4031 29733
rect 3510 29696 3516 29708
rect 2424 29668 3516 29696
rect 3510 29656 3516 29668
rect 3568 29696 3574 29708
rect 3988 29696 4016 29727
rect 5074 29724 5080 29776
rect 5132 29724 5138 29776
rect 3568 29668 4016 29696
rect 3568 29656 3574 29668
rect 4062 29656 4068 29708
rect 4120 29656 4126 29708
rect 2280 29600 2360 29628
rect 2280 29588 2286 29600
rect 3050 29588 3056 29640
rect 3108 29628 3114 29640
rect 3329 29631 3387 29637
rect 3329 29628 3341 29631
rect 3108 29600 3341 29628
rect 3108 29588 3114 29600
rect 3329 29597 3341 29600
rect 3375 29597 3387 29631
rect 3329 29591 3387 29597
rect 3789 29631 3847 29637
rect 3789 29597 3801 29631
rect 3835 29597 3847 29631
rect 3789 29591 3847 29597
rect 1302 29520 1308 29572
rect 1360 29560 1366 29572
rect 3804 29560 3832 29591
rect 4246 29588 4252 29640
rect 4304 29628 4310 29640
rect 4339 29631 4397 29637
rect 4339 29628 4351 29631
rect 4304 29600 4351 29628
rect 4304 29588 4310 29600
rect 4339 29597 4351 29600
rect 4385 29597 4397 29631
rect 4339 29591 4397 29597
rect 1360 29532 3832 29560
rect 4354 29560 4382 29591
rect 4890 29588 4896 29640
rect 4948 29628 4954 29640
rect 5736 29637 5764 29804
rect 7760 29804 11520 29832
rect 5902 29656 5908 29708
rect 5960 29696 5966 29708
rect 5960 29668 6394 29696
rect 5960 29656 5966 29668
rect 5445 29631 5503 29637
rect 5445 29628 5457 29631
rect 4948 29600 5457 29628
rect 4948 29588 4954 29600
rect 5445 29597 5457 29600
rect 5491 29597 5503 29631
rect 5445 29591 5503 29597
rect 5721 29631 5779 29637
rect 5721 29597 5733 29631
rect 5767 29628 5779 29631
rect 5767 29600 5948 29628
rect 5767 29597 5779 29600
rect 5721 29591 5779 29597
rect 5350 29560 5356 29572
rect 4354 29532 5356 29560
rect 1360 29520 1366 29532
rect 5350 29520 5356 29532
rect 5408 29520 5414 29572
rect 5920 29504 5948 29600
rect 6638 29588 6644 29640
rect 6696 29628 6702 29640
rect 6825 29631 6883 29637
rect 6825 29628 6837 29631
rect 6696 29600 6837 29628
rect 6696 29588 6702 29600
rect 6825 29597 6837 29600
rect 6871 29597 6883 29631
rect 6825 29591 6883 29597
rect 6917 29631 6975 29637
rect 6917 29597 6929 29631
rect 6963 29628 6975 29631
rect 7374 29628 7380 29640
rect 6963 29600 7380 29628
rect 6963 29597 6975 29600
rect 6917 29591 6975 29597
rect 7374 29588 7380 29600
rect 7432 29588 7438 29640
rect 7190 29520 7196 29572
rect 7248 29560 7254 29572
rect 7285 29563 7343 29569
rect 7285 29560 7297 29563
rect 7248 29532 7297 29560
rect 7248 29520 7254 29532
rect 7285 29529 7297 29532
rect 7331 29529 7343 29563
rect 7760 29560 7788 29804
rect 11514 29792 11520 29804
rect 11572 29792 11578 29844
rect 11609 29835 11667 29841
rect 11609 29801 11621 29835
rect 11655 29832 11667 29835
rect 12066 29832 12072 29844
rect 11655 29804 12072 29832
rect 11655 29801 11667 29804
rect 11609 29795 11667 29801
rect 12066 29792 12072 29804
rect 12124 29792 12130 29844
rect 13541 29835 13599 29841
rect 13541 29801 13553 29835
rect 13587 29832 13599 29835
rect 13587 29804 15148 29832
rect 13587 29801 13599 29804
rect 13541 29795 13599 29801
rect 7837 29767 7895 29773
rect 7837 29733 7849 29767
rect 7883 29764 7895 29767
rect 8202 29764 8208 29776
rect 7883 29736 8208 29764
rect 7883 29733 7895 29736
rect 7837 29727 7895 29733
rect 8202 29724 8208 29736
rect 8260 29764 8266 29776
rect 9490 29764 9496 29776
rect 8260 29736 9496 29764
rect 8260 29724 8266 29736
rect 9490 29724 9496 29736
rect 9548 29724 9554 29776
rect 9766 29764 9772 29776
rect 9646 29736 9772 29764
rect 8570 29588 8576 29640
rect 8628 29588 8634 29640
rect 9490 29588 9496 29640
rect 9548 29628 9554 29640
rect 9646 29628 9674 29736
rect 9766 29724 9772 29736
rect 9824 29764 9830 29776
rect 9824 29736 10546 29764
rect 9824 29724 9830 29736
rect 10134 29656 10140 29708
rect 10192 29696 10198 29708
rect 10413 29699 10471 29705
rect 10413 29696 10425 29699
rect 10192 29668 10425 29696
rect 10192 29656 10198 29668
rect 10413 29665 10425 29668
rect 10459 29665 10471 29699
rect 10518 29696 10546 29736
rect 12526 29724 12532 29776
rect 12584 29764 12590 29776
rect 12713 29767 12771 29773
rect 12713 29764 12725 29767
rect 12584 29736 12725 29764
rect 12584 29724 12590 29736
rect 12713 29733 12725 29736
rect 12759 29764 12771 29767
rect 15120 29764 15148 29804
rect 15194 29792 15200 29844
rect 15252 29832 15258 29844
rect 15746 29832 15752 29844
rect 15252 29804 15752 29832
rect 15252 29792 15258 29804
rect 15746 29792 15752 29804
rect 15804 29792 15810 29844
rect 19334 29792 19340 29844
rect 19392 29792 19398 29844
rect 19610 29792 19616 29844
rect 19668 29792 19674 29844
rect 19812 29804 20567 29832
rect 15470 29764 15476 29776
rect 12759 29736 13124 29764
rect 15120 29736 15476 29764
rect 12759 29733 12771 29736
rect 12713 29727 12771 29733
rect 10870 29705 10876 29708
rect 10689 29699 10747 29705
rect 10689 29696 10701 29699
rect 10518 29668 10701 29696
rect 10413 29659 10471 29665
rect 10689 29665 10701 29668
rect 10735 29665 10747 29699
rect 10689 29659 10747 29665
rect 10827 29699 10876 29705
rect 10827 29665 10839 29699
rect 10873 29665 10876 29699
rect 10827 29659 10876 29665
rect 10870 29656 10876 29659
rect 10928 29656 10934 29708
rect 13096 29705 13124 29736
rect 15470 29724 15476 29736
rect 15528 29724 15534 29776
rect 16482 29724 16488 29776
rect 16540 29724 16546 29776
rect 13081 29699 13139 29705
rect 13081 29665 13093 29699
rect 13127 29665 13139 29699
rect 13081 29659 13139 29665
rect 19521 29699 19579 29705
rect 19521 29665 19533 29699
rect 19567 29696 19579 29699
rect 19628 29696 19656 29792
rect 19812 29776 19840 29804
rect 19794 29724 19800 29776
rect 19852 29724 19858 29776
rect 19812 29696 19840 29724
rect 19889 29699 19947 29705
rect 19889 29696 19901 29699
rect 19567 29668 19656 29696
rect 19720 29668 19901 29696
rect 19567 29665 19579 29668
rect 19521 29659 19579 29665
rect 9548 29600 9674 29628
rect 9769 29631 9827 29637
rect 9548 29588 9554 29600
rect 9769 29597 9781 29631
rect 9815 29597 9827 29631
rect 9769 29591 9827 29597
rect 7285 29523 7343 29529
rect 7576 29532 7788 29560
rect 8588 29560 8616 29588
rect 9398 29560 9404 29572
rect 8588 29532 9404 29560
rect 2501 29495 2559 29501
rect 2501 29461 2513 29495
rect 2547 29492 2559 29495
rect 2590 29492 2596 29504
rect 2547 29464 2596 29492
rect 2547 29461 2559 29464
rect 2501 29455 2559 29461
rect 2590 29452 2596 29464
rect 2648 29452 2654 29504
rect 2682 29452 2688 29504
rect 2740 29492 2746 29504
rect 3694 29492 3700 29504
rect 2740 29464 3700 29492
rect 2740 29452 2746 29464
rect 3694 29452 3700 29464
rect 3752 29452 3758 29504
rect 5902 29452 5908 29504
rect 5960 29452 5966 29504
rect 6549 29495 6607 29501
rect 6549 29461 6561 29495
rect 6595 29492 6607 29495
rect 7576 29492 7604 29532
rect 9398 29520 9404 29532
rect 9456 29560 9462 29572
rect 9784 29560 9812 29591
rect 9858 29588 9864 29640
rect 9916 29628 9922 29640
rect 9953 29631 10011 29637
rect 9953 29628 9965 29631
rect 9916 29600 9965 29628
rect 9916 29588 9922 29600
rect 9953 29597 9965 29600
rect 9999 29597 10011 29631
rect 9953 29591 10011 29597
rect 10962 29588 10968 29640
rect 11020 29588 11026 29640
rect 11606 29588 11612 29640
rect 11664 29628 11670 29640
rect 11701 29631 11759 29637
rect 11701 29628 11713 29631
rect 11664 29600 11713 29628
rect 11664 29588 11670 29600
rect 11701 29597 11713 29600
rect 11747 29597 11759 29631
rect 11974 29628 11980 29640
rect 11935 29600 11980 29628
rect 11701 29591 11759 29597
rect 9456 29532 9812 29560
rect 11716 29560 11744 29591
rect 11974 29588 11980 29600
rect 12032 29588 12038 29640
rect 12710 29588 12716 29640
rect 12768 29628 12774 29640
rect 13265 29631 13323 29637
rect 13265 29628 13277 29631
rect 12768 29600 13277 29628
rect 12768 29588 12774 29600
rect 13265 29597 13277 29600
rect 13311 29597 13323 29631
rect 13998 29628 14004 29640
rect 13265 29591 13323 29597
rect 13372 29600 14004 29628
rect 13372 29560 13400 29600
rect 13998 29588 14004 29600
rect 14056 29628 14062 29640
rect 14093 29631 14151 29637
rect 14093 29628 14105 29631
rect 14056 29600 14105 29628
rect 14056 29588 14062 29600
rect 14093 29597 14105 29600
rect 14139 29597 14151 29631
rect 14826 29628 14832 29640
rect 14093 29591 14151 29597
rect 14351 29601 14409 29607
rect 11716 29532 13400 29560
rect 9456 29520 9462 29532
rect 13630 29520 13636 29572
rect 13688 29520 13694 29572
rect 14351 29567 14363 29601
rect 14397 29598 14409 29601
rect 14568 29600 14832 29628
rect 14397 29567 14410 29598
rect 14568 29572 14596 29600
rect 14826 29588 14832 29600
rect 14884 29628 14890 29640
rect 15473 29631 15531 29637
rect 15473 29628 15485 29631
rect 14884 29600 15485 29628
rect 14884 29588 14890 29600
rect 15473 29597 15485 29600
rect 15519 29597 15531 29631
rect 15473 29591 15531 29597
rect 14351 29561 14410 29567
rect 14382 29560 14410 29561
rect 14382 29532 14412 29560
rect 14384 29504 14412 29532
rect 14550 29520 14556 29572
rect 14608 29520 14614 29572
rect 15488 29560 15516 29591
rect 15746 29588 15752 29640
rect 15804 29628 15810 29640
rect 16298 29628 16304 29640
rect 15804 29600 16304 29628
rect 15804 29588 15810 29600
rect 16298 29588 16304 29600
rect 16356 29588 16362 29640
rect 19242 29588 19248 29640
rect 19300 29588 19306 29640
rect 19426 29588 19432 29640
rect 19484 29628 19490 29640
rect 19720 29628 19748 29668
rect 19889 29665 19901 29668
rect 19935 29665 19947 29699
rect 20539 29696 20567 29804
rect 20898 29792 20904 29844
rect 20956 29792 20962 29844
rect 22554 29792 22560 29844
rect 22612 29792 22618 29844
rect 23109 29835 23167 29841
rect 23109 29801 23121 29835
rect 23155 29832 23167 29835
rect 23566 29832 23572 29844
rect 23155 29804 23572 29832
rect 23155 29801 23167 29804
rect 23109 29795 23167 29801
rect 23566 29792 23572 29804
rect 23624 29792 23630 29844
rect 22572 29764 22600 29792
rect 23382 29764 23388 29776
rect 22572 29736 23388 29764
rect 23382 29724 23388 29736
rect 23440 29724 23446 29776
rect 21082 29696 21088 29708
rect 20539 29668 21088 29696
rect 19889 29659 19947 29665
rect 21082 29656 21088 29668
rect 21140 29696 21146 29708
rect 21361 29699 21419 29705
rect 21361 29696 21373 29699
rect 21140 29668 21373 29696
rect 21140 29656 21146 29668
rect 21361 29665 21373 29668
rect 21407 29665 21419 29699
rect 21361 29659 21419 29665
rect 22278 29656 22284 29708
rect 22336 29696 22342 29708
rect 22336 29668 25360 29696
rect 22336 29656 22342 29668
rect 25332 29640 25360 29668
rect 19484 29600 19748 29628
rect 19797 29631 19855 29637
rect 19484 29588 19490 29600
rect 19797 29597 19809 29631
rect 19843 29597 19855 29631
rect 20162 29628 20168 29640
rect 20123 29600 20168 29628
rect 19797 29591 19855 29597
rect 17034 29560 17040 29572
rect 15488 29532 17040 29560
rect 17034 29520 17040 29532
rect 17092 29520 17098 29572
rect 19058 29520 19064 29572
rect 19116 29560 19122 29572
rect 19812 29560 19840 29591
rect 20162 29588 20168 29600
rect 20220 29588 20226 29640
rect 21174 29588 21180 29640
rect 21232 29588 21238 29640
rect 21634 29588 21640 29640
rect 21692 29588 21698 29640
rect 23293 29631 23351 29637
rect 23293 29628 23305 29631
rect 22066 29600 23305 29628
rect 19116 29532 19840 29560
rect 19116 29520 19122 29532
rect 19260 29504 19288 29532
rect 6595 29464 7604 29492
rect 7653 29495 7711 29501
rect 6595 29461 6607 29464
rect 6549 29455 6607 29461
rect 7653 29461 7665 29495
rect 7699 29492 7711 29495
rect 7742 29492 7748 29504
rect 7699 29464 7748 29492
rect 7699 29461 7711 29464
rect 7653 29455 7711 29461
rect 7742 29452 7748 29464
rect 7800 29452 7806 29504
rect 8846 29452 8852 29504
rect 8904 29492 8910 29504
rect 10870 29492 10876 29504
rect 8904 29464 10876 29492
rect 8904 29452 8910 29464
rect 10870 29452 10876 29464
rect 10928 29452 10934 29504
rect 14366 29452 14372 29504
rect 14424 29452 14430 29504
rect 14642 29452 14648 29504
rect 14700 29492 14706 29504
rect 15105 29495 15163 29501
rect 15105 29492 15117 29495
rect 14700 29464 15117 29492
rect 14700 29452 14706 29464
rect 15105 29461 15117 29464
rect 15151 29461 15163 29495
rect 15105 29455 15163 29461
rect 19242 29452 19248 29504
rect 19300 29452 19306 29504
rect 19518 29452 19524 29504
rect 19576 29452 19582 29504
rect 19613 29495 19671 29501
rect 19613 29461 19625 29495
rect 19659 29492 19671 29495
rect 21192 29492 21220 29588
rect 21818 29520 21824 29572
rect 21876 29560 21882 29572
rect 22066 29560 22094 29600
rect 23293 29597 23305 29600
rect 23339 29597 23351 29631
rect 23661 29631 23719 29637
rect 23661 29628 23673 29631
rect 23293 29591 23351 29597
rect 23400 29600 23673 29628
rect 21876 29532 22094 29560
rect 21876 29520 21882 29532
rect 22922 29520 22928 29572
rect 22980 29560 22986 29572
rect 23400 29560 23428 29600
rect 23661 29597 23673 29600
rect 23707 29597 23719 29631
rect 23661 29591 23719 29597
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 23845 29563 23903 29569
rect 23845 29560 23857 29563
rect 22980 29532 23428 29560
rect 23492 29532 23857 29560
rect 22980 29520 22986 29532
rect 19659 29464 21220 29492
rect 19659 29461 19671 29464
rect 19613 29455 19671 29461
rect 22370 29452 22376 29504
rect 22428 29452 22434 29504
rect 23492 29501 23520 29532
rect 23845 29529 23857 29532
rect 23891 29529 23903 29563
rect 23845 29523 23903 29529
rect 24210 29520 24216 29572
rect 24268 29520 24274 29572
rect 23477 29495 23535 29501
rect 23477 29461 23489 29495
rect 23523 29461 23535 29495
rect 23477 29455 23535 29461
rect 1104 29402 25000 29424
rect 1104 29350 6884 29402
rect 6936 29350 6948 29402
rect 7000 29350 7012 29402
rect 7064 29350 7076 29402
rect 7128 29350 7140 29402
rect 7192 29350 12818 29402
rect 12870 29350 12882 29402
rect 12934 29350 12946 29402
rect 12998 29350 13010 29402
rect 13062 29350 13074 29402
rect 13126 29350 18752 29402
rect 18804 29350 18816 29402
rect 18868 29350 18880 29402
rect 18932 29350 18944 29402
rect 18996 29350 19008 29402
rect 19060 29350 24686 29402
rect 24738 29350 24750 29402
rect 24802 29350 24814 29402
rect 24866 29350 24878 29402
rect 24930 29350 24942 29402
rect 24994 29350 25000 29402
rect 1104 29328 25000 29350
rect 1118 29248 1124 29300
rect 1176 29288 1182 29300
rect 1176 29260 3464 29288
rect 1176 29248 1182 29260
rect 2314 29112 2320 29164
rect 2372 29112 2378 29164
rect 2590 29112 2596 29164
rect 2648 29112 2654 29164
rect 3436 29161 3464 29260
rect 4706 29248 4712 29300
rect 4764 29288 4770 29300
rect 7742 29288 7748 29300
rect 4764 29260 7748 29288
rect 4764 29248 4770 29260
rect 7742 29248 7748 29260
rect 7800 29248 7806 29300
rect 9582 29288 9588 29300
rect 9398 29260 9588 29288
rect 3712 29192 6408 29220
rect 3421 29155 3479 29161
rect 3421 29121 3433 29155
rect 3467 29121 3479 29155
rect 3421 29115 3479 29121
rect 1394 29044 1400 29096
rect 1452 29044 1458 29096
rect 3712 29093 3740 29192
rect 3878 29112 3884 29164
rect 3936 29112 3942 29164
rect 4890 29112 4896 29164
rect 4948 29152 4954 29164
rect 4983 29155 5041 29161
rect 4983 29152 4995 29155
rect 4948 29124 4995 29152
rect 4948 29112 4954 29124
rect 4983 29121 4995 29124
rect 5029 29152 5041 29155
rect 6086 29152 6092 29164
rect 5029 29124 6092 29152
rect 5029 29121 5041 29124
rect 4983 29115 5041 29121
rect 6086 29112 6092 29124
rect 6144 29112 6150 29164
rect 6380 29152 6408 29192
rect 9398 29191 9426 29260
rect 9582 29248 9588 29260
rect 9640 29248 9646 29300
rect 10134 29248 10140 29300
rect 10192 29248 10198 29300
rect 10778 29248 10784 29300
rect 10836 29248 10842 29300
rect 11330 29248 11336 29300
rect 11388 29248 11394 29300
rect 11977 29291 12035 29297
rect 11977 29257 11989 29291
rect 12023 29257 12035 29291
rect 11977 29251 12035 29257
rect 12621 29291 12679 29297
rect 12621 29257 12633 29291
rect 12667 29288 12679 29291
rect 13630 29288 13636 29300
rect 12667 29260 13636 29288
rect 12667 29257 12679 29260
rect 12621 29251 12679 29257
rect 9383 29185 9441 29191
rect 8846 29152 8852 29164
rect 6380 29124 8852 29152
rect 8846 29112 8852 29124
rect 8904 29112 8910 29164
rect 9383 29151 9395 29185
rect 9429 29151 9441 29185
rect 9674 29180 9680 29232
rect 9732 29220 9738 29232
rect 10796 29220 10824 29248
rect 9732 29192 10824 29220
rect 9732 29180 9738 29192
rect 9383 29145 9441 29151
rect 9582 29122 9588 29174
rect 9640 29152 9646 29174
rect 11348 29152 11376 29248
rect 11992 29220 12020 29251
rect 13630 29248 13636 29260
rect 13688 29248 13694 29300
rect 14366 29248 14372 29300
rect 14424 29288 14430 29300
rect 14424 29260 23336 29288
rect 14424 29248 14430 29260
rect 11992 29192 12689 29220
rect 12161 29155 12219 29161
rect 12161 29152 12173 29155
rect 9640 29124 10272 29152
rect 11348 29124 12173 29152
rect 9640 29122 9646 29124
rect 1581 29087 1639 29093
rect 1581 29053 1593 29087
rect 1627 29053 1639 29087
rect 1581 29047 1639 29053
rect 2455 29087 2513 29093
rect 2455 29053 2467 29087
rect 2501 29084 2513 29087
rect 3697 29087 3755 29093
rect 3697 29084 3709 29087
rect 2501 29056 3709 29084
rect 2501 29053 2513 29056
rect 2455 29047 2513 29053
rect 3697 29053 3709 29056
rect 3743 29053 3755 29087
rect 3697 29047 3755 29053
rect 1596 29016 1624 29047
rect 1854 29016 1860 29028
rect 1596 28988 1860 29016
rect 1854 28976 1860 28988
rect 1912 28976 1918 29028
rect 2038 28976 2044 29028
rect 2096 28976 2102 29028
rect 3237 29019 3295 29025
rect 3237 28985 3249 29019
rect 3283 29016 3295 29019
rect 3896 29016 3924 29112
rect 4154 29044 4160 29096
rect 4212 29084 4218 29096
rect 4522 29084 4528 29096
rect 4212 29056 4528 29084
rect 4212 29044 4218 29056
rect 4522 29044 4528 29056
rect 4580 29084 4586 29096
rect 4709 29087 4767 29093
rect 4709 29084 4721 29087
rect 4580 29056 4721 29084
rect 4580 29044 4586 29056
rect 4709 29053 4721 29056
rect 4755 29053 4767 29087
rect 6104 29084 6132 29112
rect 6638 29084 6644 29096
rect 6104 29056 6644 29084
rect 4709 29047 4767 29053
rect 6638 29044 6644 29056
rect 6696 29044 6702 29096
rect 7374 29044 7380 29096
rect 7432 29084 7438 29096
rect 9030 29084 9036 29096
rect 7432 29056 9036 29084
rect 7432 29044 7438 29056
rect 9030 29044 9036 29056
rect 9088 29084 9094 29096
rect 9125 29087 9183 29093
rect 9125 29084 9137 29087
rect 9088 29056 9137 29084
rect 9088 29044 9094 29056
rect 9125 29053 9137 29056
rect 9171 29053 9183 29087
rect 9125 29047 9183 29053
rect 10244 29028 10272 29124
rect 12161 29121 12173 29124
rect 12207 29121 12219 29155
rect 12161 29115 12219 29121
rect 12437 29155 12495 29161
rect 12437 29121 12449 29155
rect 12483 29152 12495 29155
rect 12526 29152 12532 29164
rect 12483 29124 12532 29152
rect 12483 29121 12495 29124
rect 12437 29115 12495 29121
rect 12526 29112 12532 29124
rect 12584 29112 12590 29164
rect 12661 29161 12689 29192
rect 13170 29180 13176 29232
rect 13228 29220 13234 29232
rect 22278 29220 22284 29232
rect 13228 29192 22284 29220
rect 13228 29180 13234 29192
rect 22278 29180 22284 29192
rect 22336 29180 22342 29232
rect 12621 29155 12689 29161
rect 12621 29121 12633 29155
rect 12667 29128 12689 29155
rect 12986 29152 12992 29164
rect 12667 29121 12679 29128
rect 12947 29124 12992 29152
rect 12621 29115 12679 29121
rect 12986 29112 12992 29124
rect 13044 29112 13050 29164
rect 13722 29112 13728 29164
rect 13780 29152 13786 29164
rect 14367 29155 14425 29161
rect 14367 29152 14379 29155
rect 13780 29124 14379 29152
rect 13780 29112 13786 29124
rect 14367 29121 14379 29124
rect 14413 29152 14425 29155
rect 14413 29124 15240 29152
rect 14413 29121 14425 29124
rect 14367 29115 14425 29121
rect 12713 29087 12771 29093
rect 12713 29053 12725 29087
rect 12759 29053 12771 29087
rect 12713 29047 12771 29053
rect 3283 28988 3924 29016
rect 4172 28988 4844 29016
rect 3283 28985 3295 28988
rect 3237 28979 3295 28985
rect 1578 28908 1584 28960
rect 1636 28948 1642 28960
rect 3510 28948 3516 28960
rect 1636 28920 3516 28948
rect 1636 28908 1642 28920
rect 3510 28908 3516 28920
rect 3568 28908 3574 28960
rect 3602 28908 3608 28960
rect 3660 28948 3666 28960
rect 4172 28948 4200 28988
rect 3660 28920 4200 28948
rect 4816 28948 4844 28988
rect 5460 28988 5856 29016
rect 5460 28948 5488 28988
rect 4816 28920 5488 28948
rect 3660 28908 3666 28920
rect 5534 28908 5540 28960
rect 5592 28948 5598 28960
rect 5721 28951 5779 28957
rect 5721 28948 5733 28951
rect 5592 28920 5733 28948
rect 5592 28908 5598 28920
rect 5721 28917 5733 28920
rect 5767 28917 5779 28951
rect 5828 28948 5856 28988
rect 7282 28976 7288 29028
rect 7340 29016 7346 29028
rect 7742 29016 7748 29028
rect 7340 28988 7748 29016
rect 7340 28976 7346 28988
rect 7742 28976 7748 28988
rect 7800 28976 7806 29028
rect 8386 29016 8392 29028
rect 8220 28988 8392 29016
rect 8220 28948 8248 28988
rect 8386 28976 8392 28988
rect 8444 28976 8450 29028
rect 10226 28976 10232 29028
rect 10284 28976 10290 29028
rect 12250 28976 12256 29028
rect 12308 29016 12314 29028
rect 12728 29016 12756 29047
rect 13906 29044 13912 29096
rect 13964 29084 13970 29096
rect 14093 29087 14151 29093
rect 14093 29084 14105 29087
rect 13964 29056 14105 29084
rect 13964 29044 13970 29056
rect 14093 29053 14105 29056
rect 14139 29053 14151 29087
rect 14093 29047 14151 29053
rect 13725 29019 13783 29025
rect 12308 28988 12848 29016
rect 12308 28976 12314 28988
rect 5828 28920 8248 28948
rect 5721 28911 5779 28917
rect 8294 28908 8300 28960
rect 8352 28948 8358 28960
rect 8846 28948 8852 28960
rect 8352 28920 8852 28948
rect 8352 28908 8358 28920
rect 8846 28908 8852 28920
rect 8904 28948 8910 28960
rect 9858 28948 9864 28960
rect 8904 28920 9864 28948
rect 8904 28908 8910 28920
rect 9858 28908 9864 28920
rect 9916 28908 9922 28960
rect 12820 28948 12848 28988
rect 13725 28985 13737 29019
rect 13771 29016 13783 29019
rect 13998 29016 14004 29028
rect 13771 28988 14004 29016
rect 13771 28985 13783 28988
rect 13725 28979 13783 28985
rect 13998 28976 14004 28988
rect 14056 28976 14062 29028
rect 15102 28976 15108 29028
rect 15160 28976 15166 29028
rect 15212 29016 15240 29124
rect 16942 29112 16948 29164
rect 17000 29152 17006 29164
rect 17279 29155 17337 29161
rect 17279 29152 17291 29155
rect 17000 29124 17291 29152
rect 17000 29112 17006 29124
rect 17279 29121 17291 29124
rect 17325 29152 17337 29155
rect 17402 29152 17408 29164
rect 17325 29124 17408 29152
rect 17325 29121 17337 29124
rect 17279 29115 17337 29121
rect 17402 29112 17408 29124
rect 17460 29112 17466 29164
rect 17862 29112 17868 29164
rect 17920 29152 17926 29164
rect 20714 29152 20720 29164
rect 17920 29124 20720 29152
rect 17920 29112 17926 29124
rect 20714 29112 20720 29124
rect 20772 29112 20778 29164
rect 21358 29112 21364 29164
rect 21416 29112 21422 29164
rect 21818 29152 21824 29164
rect 21468 29124 21824 29152
rect 17034 29044 17040 29096
rect 17092 29044 17098 29096
rect 21468 29084 21496 29124
rect 21818 29112 21824 29124
rect 21876 29112 21882 29164
rect 22370 29112 22376 29164
rect 22428 29112 22434 29164
rect 22554 29112 22560 29164
rect 22612 29112 22618 29164
rect 23109 29155 23167 29161
rect 23109 29121 23121 29155
rect 23155 29152 23167 29155
rect 23308 29152 23336 29260
rect 23385 29155 23443 29161
rect 23385 29152 23397 29155
rect 23155 29124 23244 29152
rect 23308 29124 23397 29152
rect 23155 29121 23167 29124
rect 23109 29115 23167 29121
rect 17696 29056 21496 29084
rect 15212 28988 17172 29016
rect 14826 28948 14832 28960
rect 12820 28920 14832 28948
rect 14826 28908 14832 28920
rect 14884 28908 14890 28960
rect 17144 28948 17172 28988
rect 17696 28948 17724 29056
rect 21177 29019 21235 29025
rect 21177 28985 21189 29019
rect 21223 29016 21235 29019
rect 22094 29016 22100 29028
rect 21223 28988 22100 29016
rect 21223 28985 21235 28988
rect 21177 28979 21235 28985
rect 22094 28976 22100 28988
rect 22152 28976 22158 29028
rect 22922 28976 22928 29028
rect 22980 28976 22986 29028
rect 23216 29025 23244 29124
rect 23385 29121 23397 29124
rect 23431 29121 23443 29155
rect 23385 29115 23443 29121
rect 23845 29155 23903 29161
rect 23845 29121 23857 29155
rect 23891 29121 23903 29155
rect 23845 29115 23903 29121
rect 23201 29019 23259 29025
rect 23201 28985 23213 29019
rect 23247 28985 23259 29019
rect 23201 28979 23259 28985
rect 23382 28976 23388 29028
rect 23440 29016 23446 29028
rect 23860 29016 23888 29115
rect 24118 29112 24124 29164
rect 24176 29112 24182 29164
rect 23440 28988 23888 29016
rect 23440 28976 23446 28988
rect 24394 28976 24400 29028
rect 24452 28976 24458 29028
rect 17144 28920 17724 28948
rect 18049 28951 18107 28957
rect 18049 28917 18061 28951
rect 18095 28948 18107 28951
rect 18414 28948 18420 28960
rect 18095 28920 18420 28948
rect 18095 28917 18107 28920
rect 18049 28911 18107 28917
rect 18414 28908 18420 28920
rect 18472 28908 18478 28960
rect 18598 28908 18604 28960
rect 18656 28948 18662 28960
rect 21726 28948 21732 28960
rect 18656 28920 21732 28948
rect 18656 28908 18662 28920
rect 21726 28908 21732 28920
rect 21784 28908 21790 28960
rect 22462 28908 22468 28960
rect 22520 28908 22526 28960
rect 23661 28951 23719 28957
rect 23661 28917 23673 28951
rect 23707 28948 23719 28951
rect 23934 28948 23940 28960
rect 23707 28920 23940 28948
rect 23707 28917 23719 28920
rect 23661 28911 23719 28917
rect 23934 28908 23940 28920
rect 23992 28908 23998 28960
rect 1104 28858 24840 28880
rect 1104 28806 3917 28858
rect 3969 28806 3981 28858
rect 4033 28806 4045 28858
rect 4097 28806 4109 28858
rect 4161 28806 4173 28858
rect 4225 28806 9851 28858
rect 9903 28806 9915 28858
rect 9967 28806 9979 28858
rect 10031 28806 10043 28858
rect 10095 28806 10107 28858
rect 10159 28806 15785 28858
rect 15837 28806 15849 28858
rect 15901 28806 15913 28858
rect 15965 28806 15977 28858
rect 16029 28806 16041 28858
rect 16093 28806 21719 28858
rect 21771 28806 21783 28858
rect 21835 28806 21847 28858
rect 21899 28806 21911 28858
rect 21963 28806 21975 28858
rect 22027 28806 24840 28858
rect 1104 28784 24840 28806
rect 1946 28704 1952 28756
rect 2004 28744 2010 28756
rect 3602 28744 3608 28756
rect 2004 28716 3608 28744
rect 2004 28704 2010 28716
rect 3602 28704 3608 28716
rect 3660 28704 3666 28756
rect 5902 28704 5908 28756
rect 5960 28744 5966 28756
rect 8018 28744 8024 28756
rect 5960 28716 8024 28744
rect 5960 28704 5966 28716
rect 8018 28704 8024 28716
rect 8076 28704 8082 28756
rect 10594 28704 10600 28756
rect 10652 28744 10658 28756
rect 18598 28744 18604 28756
rect 10652 28716 18604 28744
rect 10652 28704 10658 28716
rect 18598 28704 18604 28716
rect 18656 28704 18662 28756
rect 19061 28747 19119 28753
rect 19061 28713 19073 28747
rect 19107 28744 19119 28747
rect 19242 28744 19248 28756
rect 19107 28716 19248 28744
rect 19107 28713 19119 28716
rect 19061 28707 19119 28713
rect 19242 28704 19248 28716
rect 19300 28704 19306 28756
rect 19334 28704 19340 28756
rect 19392 28744 19398 28756
rect 20349 28747 20407 28753
rect 19392 28716 20300 28744
rect 19392 28704 19398 28716
rect 3329 28679 3387 28685
rect 3329 28645 3341 28679
rect 3375 28676 3387 28679
rect 5261 28679 5319 28685
rect 3375 28648 3832 28676
rect 3375 28645 3387 28648
rect 3329 28639 3387 28645
rect 3804 28594 3832 28648
rect 5261 28645 5273 28679
rect 5307 28676 5319 28679
rect 8662 28676 8668 28688
rect 5307 28648 6224 28676
rect 5307 28645 5319 28648
rect 5261 28639 5319 28645
rect 1210 28500 1216 28552
rect 1268 28540 1274 28552
rect 1857 28543 1915 28549
rect 1857 28540 1869 28543
rect 1268 28512 1869 28540
rect 1268 28500 1274 28512
rect 1857 28509 1869 28512
rect 1903 28509 1915 28543
rect 1857 28503 1915 28509
rect 2314 28500 2320 28552
rect 2372 28500 2378 28552
rect 2498 28500 2504 28552
rect 2556 28540 2562 28552
rect 2591 28543 2649 28549
rect 2591 28540 2603 28543
rect 2556 28512 2603 28540
rect 2556 28500 2562 28512
rect 2591 28509 2603 28512
rect 2637 28509 2649 28543
rect 2591 28503 2649 28509
rect 2682 28500 2688 28552
rect 2740 28540 2746 28552
rect 4249 28543 4307 28549
rect 2740 28512 4182 28540
rect 2740 28500 2746 28512
rect 750 28432 756 28484
rect 808 28472 814 28484
rect 1489 28475 1547 28481
rect 1489 28472 1501 28475
rect 808 28444 1501 28472
rect 808 28432 814 28444
rect 1489 28441 1501 28444
rect 1535 28441 1547 28475
rect 1489 28435 1547 28441
rect 1673 28475 1731 28481
rect 1673 28441 1685 28475
rect 1719 28472 1731 28475
rect 3878 28472 3884 28484
rect 1719 28444 3884 28472
rect 1719 28441 1731 28444
rect 1673 28435 1731 28441
rect 3878 28432 3884 28444
rect 3936 28432 3942 28484
rect 1946 28364 1952 28416
rect 2004 28364 2010 28416
rect 2590 28364 2596 28416
rect 2648 28404 2654 28416
rect 3786 28404 3792 28416
rect 2648 28376 3792 28404
rect 2648 28364 2654 28376
rect 3786 28364 3792 28376
rect 3844 28404 3850 28416
rect 3973 28407 4031 28413
rect 3973 28404 3985 28407
rect 3844 28376 3985 28404
rect 3844 28364 3850 28376
rect 3973 28373 3985 28376
rect 4019 28373 4031 28407
rect 4154 28404 4182 28512
rect 4249 28509 4261 28543
rect 4295 28540 4307 28543
rect 4295 28512 5304 28540
rect 4295 28509 4307 28512
rect 4249 28503 4307 28509
rect 5276 28484 5304 28512
rect 5534 28500 5540 28552
rect 5592 28540 5598 28552
rect 5902 28540 5908 28552
rect 5592 28512 5908 28540
rect 5592 28500 5598 28512
rect 5902 28500 5908 28512
rect 5960 28500 5966 28552
rect 4338 28432 4344 28484
rect 4396 28432 4402 28484
rect 4709 28475 4767 28481
rect 4709 28441 4721 28475
rect 4755 28472 4767 28475
rect 5166 28472 5172 28484
rect 4755 28444 5172 28472
rect 4755 28441 4767 28444
rect 4709 28435 4767 28441
rect 4724 28404 4752 28435
rect 5166 28432 5172 28444
rect 5224 28432 5230 28484
rect 5258 28432 5264 28484
rect 5316 28432 5322 28484
rect 6196 28472 6224 28648
rect 7484 28648 8668 28676
rect 7484 28620 7512 28648
rect 8662 28636 8668 28648
rect 8720 28636 8726 28688
rect 15470 28636 15476 28688
rect 15528 28676 15534 28688
rect 15528 28648 16068 28676
rect 15528 28636 15534 28648
rect 7466 28568 7472 28620
rect 7524 28568 7530 28620
rect 11606 28608 11612 28620
rect 8128 28580 11612 28608
rect 6270 28500 6276 28552
rect 6328 28500 6334 28552
rect 6546 28549 6552 28552
rect 6515 28543 6552 28549
rect 6515 28509 6527 28543
rect 6515 28503 6552 28509
rect 6546 28500 6552 28503
rect 6604 28500 6610 28552
rect 6638 28500 6644 28552
rect 6696 28540 6702 28552
rect 8128 28540 8156 28580
rect 11606 28568 11612 28580
rect 11664 28568 11670 28620
rect 11882 28568 11888 28620
rect 11940 28608 11946 28620
rect 12158 28608 12164 28620
rect 11940 28580 12164 28608
rect 11940 28568 11946 28580
rect 12158 28568 12164 28580
rect 12216 28608 12222 28620
rect 12621 28611 12679 28617
rect 12621 28608 12633 28611
rect 12216 28580 12633 28608
rect 12216 28568 12222 28580
rect 12621 28577 12633 28580
rect 12667 28577 12679 28611
rect 12621 28571 12679 28577
rect 15930 28568 15936 28620
rect 15988 28568 15994 28620
rect 16040 28608 16068 28648
rect 17862 28636 17868 28688
rect 17920 28636 17926 28688
rect 20272 28676 20300 28716
rect 20349 28713 20361 28747
rect 20395 28744 20407 28747
rect 21358 28744 21364 28756
rect 20395 28716 21364 28744
rect 20395 28713 20407 28716
rect 20349 28707 20407 28713
rect 21358 28704 21364 28716
rect 21416 28704 21422 28756
rect 22554 28704 22560 28756
rect 22612 28744 22618 28756
rect 22833 28747 22891 28753
rect 22833 28744 22845 28747
rect 22612 28716 22845 28744
rect 22612 28704 22618 28716
rect 22833 28713 22845 28716
rect 22879 28713 22891 28747
rect 22833 28707 22891 28713
rect 23382 28704 23388 28756
rect 23440 28704 23446 28756
rect 20438 28676 20444 28688
rect 19306 28648 20208 28676
rect 20272 28648 20444 28676
rect 16326 28611 16384 28617
rect 16326 28608 16338 28611
rect 16040 28580 16338 28608
rect 16326 28577 16338 28580
rect 16372 28577 16384 28611
rect 16326 28571 16384 28577
rect 16482 28568 16488 28620
rect 16540 28568 16546 28620
rect 17494 28608 17500 28620
rect 17236 28580 17500 28608
rect 6696 28512 8156 28540
rect 6696 28500 6702 28512
rect 8202 28500 8208 28552
rect 8260 28540 8266 28552
rect 8260 28519 12922 28540
rect 8260 28513 12937 28519
rect 8260 28512 12891 28513
rect 8260 28500 8266 28512
rect 12434 28472 12440 28484
rect 6196 28444 6316 28472
rect 4154 28376 4752 28404
rect 3973 28367 4031 28373
rect 4890 28364 4896 28416
rect 4948 28404 4954 28416
rect 5077 28407 5135 28413
rect 5077 28404 5089 28407
rect 4948 28376 5089 28404
rect 4948 28364 4954 28376
rect 5077 28373 5089 28376
rect 5123 28373 5135 28407
rect 6288 28404 6316 28444
rect 7208 28444 12440 28472
rect 7208 28404 7236 28444
rect 12434 28432 12440 28444
rect 12492 28432 12498 28484
rect 12879 28479 12891 28512
rect 12925 28479 12937 28513
rect 15286 28500 15292 28552
rect 15344 28500 15350 28552
rect 15473 28543 15531 28549
rect 15473 28509 15485 28543
rect 15519 28540 15531 28543
rect 15654 28540 15660 28552
rect 15519 28512 15660 28540
rect 15519 28509 15531 28512
rect 15473 28503 15531 28509
rect 15654 28500 15660 28512
rect 15712 28500 15718 28552
rect 16206 28500 16212 28552
rect 16264 28500 16270 28552
rect 17236 28549 17264 28580
rect 17494 28568 17500 28580
rect 17552 28568 17558 28620
rect 18138 28568 18144 28620
rect 18196 28568 18202 28620
rect 18598 28568 18604 28620
rect 18656 28608 18662 28620
rect 19306 28608 19334 28648
rect 20180 28608 20208 28648
rect 20438 28636 20444 28648
rect 20496 28636 20502 28688
rect 22186 28676 22192 28688
rect 22112 28648 22192 28676
rect 18656 28580 19334 28608
rect 19812 28580 20024 28608
rect 20180 28580 20760 28608
rect 18656 28568 18662 28580
rect 19812 28552 19840 28580
rect 17221 28543 17279 28549
rect 17221 28509 17233 28543
rect 17267 28509 17279 28543
rect 17221 28503 17279 28509
rect 17405 28543 17463 28549
rect 17405 28509 17417 28543
rect 17451 28509 17463 28543
rect 17405 28503 17463 28509
rect 12879 28473 12937 28479
rect 6288 28376 7236 28404
rect 5077 28367 5135 28373
rect 7282 28364 7288 28416
rect 7340 28364 7346 28416
rect 8018 28364 8024 28416
rect 8076 28404 8082 28416
rect 12618 28404 12624 28416
rect 8076 28376 12624 28404
rect 8076 28364 8082 28376
rect 12618 28364 12624 28376
rect 12676 28364 12682 28416
rect 12710 28364 12716 28416
rect 12768 28404 12774 28416
rect 12894 28404 12922 28473
rect 17420 28472 17448 28503
rect 18230 28500 18236 28552
rect 18288 28549 18294 28552
rect 18288 28543 18316 28549
rect 18304 28509 18316 28543
rect 18288 28503 18316 28509
rect 18288 28500 18294 28503
rect 18414 28500 18420 28552
rect 18472 28500 18478 28552
rect 19794 28500 19800 28552
rect 19852 28500 19858 28552
rect 19886 28500 19892 28552
rect 19944 28500 19950 28552
rect 19996 28549 20024 28580
rect 19981 28543 20039 28549
rect 19981 28509 19993 28543
rect 20027 28509 20039 28543
rect 19981 28503 20039 28509
rect 20165 28543 20223 28549
rect 20165 28509 20177 28543
rect 20211 28509 20223 28543
rect 20165 28503 20223 28509
rect 20180 28472 20208 28503
rect 20438 28500 20444 28552
rect 20496 28540 20502 28552
rect 20533 28543 20591 28549
rect 20533 28540 20545 28543
rect 20496 28512 20545 28540
rect 20496 28500 20502 28512
rect 20533 28509 20545 28512
rect 20579 28509 20591 28543
rect 20533 28503 20591 28509
rect 20622 28500 20628 28552
rect 20680 28500 20686 28552
rect 20732 28540 20760 28580
rect 22112 28540 22140 28648
rect 22186 28636 22192 28648
rect 22244 28636 22250 28688
rect 22373 28679 22431 28685
rect 22373 28645 22385 28679
rect 22419 28676 22431 28679
rect 23842 28676 23848 28688
rect 22419 28648 23848 28676
rect 22419 28645 22431 28648
rect 22373 28639 22431 28645
rect 23842 28636 23848 28648
rect 23900 28636 23906 28688
rect 22204 28580 22416 28608
rect 22204 28549 22232 28580
rect 22388 28552 22416 28580
rect 22462 28568 22468 28620
rect 22520 28568 22526 28620
rect 20732 28512 22140 28540
rect 22189 28543 22247 28549
rect 22189 28509 22201 28543
rect 22235 28509 22247 28543
rect 22189 28503 22247 28509
rect 22281 28543 22339 28549
rect 22281 28509 22293 28543
rect 22327 28509 22339 28543
rect 22281 28503 22339 28509
rect 17052 28444 17448 28472
rect 19720 28444 20208 28472
rect 20892 28475 20950 28481
rect 13262 28404 13268 28416
rect 12768 28376 13268 28404
rect 12768 28364 12774 28376
rect 13262 28364 13268 28376
rect 13320 28364 13326 28416
rect 13633 28407 13691 28413
rect 13633 28373 13645 28407
rect 13679 28404 13691 28407
rect 13906 28404 13912 28416
rect 13679 28376 13912 28404
rect 13679 28373 13691 28376
rect 13633 28367 13691 28373
rect 13906 28364 13912 28376
rect 13964 28364 13970 28416
rect 16206 28364 16212 28416
rect 16264 28404 16270 28416
rect 16482 28404 16488 28416
rect 16264 28376 16488 28404
rect 16264 28364 16270 28376
rect 16482 28364 16488 28376
rect 16540 28364 16546 28416
rect 16574 28364 16580 28416
rect 16632 28404 16638 28416
rect 17052 28404 17080 28444
rect 16632 28376 17080 28404
rect 17129 28407 17187 28413
rect 16632 28364 16638 28376
rect 17129 28373 17141 28407
rect 17175 28404 17187 28407
rect 18414 28404 18420 28416
rect 17175 28376 18420 28404
rect 17175 28373 17187 28376
rect 17129 28367 17187 28373
rect 18414 28364 18420 28376
rect 18472 28364 18478 28416
rect 18874 28364 18880 28416
rect 18932 28404 18938 28416
rect 19242 28404 19248 28416
rect 18932 28376 19248 28404
rect 18932 28364 18938 28376
rect 19242 28364 19248 28376
rect 19300 28364 19306 28416
rect 19720 28413 19748 28444
rect 20892 28441 20904 28475
rect 20938 28441 20950 28475
rect 22296 28472 22324 28503
rect 22370 28500 22376 28552
rect 22428 28500 22434 28552
rect 22554 28500 22560 28552
rect 22612 28500 22618 28552
rect 23017 28543 23075 28549
rect 23017 28509 23029 28543
rect 23063 28509 23075 28543
rect 23017 28503 23075 28509
rect 22649 28475 22707 28481
rect 22649 28472 22661 28475
rect 22296 28444 22661 28472
rect 20892 28435 20950 28441
rect 22649 28441 22661 28444
rect 22695 28441 22707 28475
rect 22649 28435 22707 28441
rect 19705 28407 19763 28413
rect 19705 28373 19717 28407
rect 19751 28373 19763 28407
rect 19705 28367 19763 28373
rect 20070 28364 20076 28416
rect 20128 28364 20134 28416
rect 20530 28364 20536 28416
rect 20588 28404 20594 28416
rect 20907 28404 20935 28435
rect 20588 28376 20935 28404
rect 22005 28407 22063 28413
rect 20588 28364 20594 28376
rect 22005 28373 22017 28407
rect 22051 28404 22063 28407
rect 23032 28404 23060 28503
rect 23290 28500 23296 28552
rect 23348 28500 23354 28552
rect 23569 28543 23627 28549
rect 23569 28509 23581 28543
rect 23615 28509 23627 28543
rect 23569 28503 23627 28509
rect 23584 28472 23612 28503
rect 23658 28500 23664 28552
rect 23716 28540 23722 28552
rect 23845 28543 23903 28549
rect 23845 28540 23857 28543
rect 23716 28512 23857 28540
rect 23716 28500 23722 28512
rect 23845 28509 23857 28512
rect 23891 28509 23903 28543
rect 23845 28503 23903 28509
rect 23934 28500 23940 28552
rect 23992 28500 23998 28552
rect 23124 28444 23612 28472
rect 23124 28413 23152 28444
rect 22051 28376 23060 28404
rect 23109 28407 23167 28413
rect 22051 28373 22063 28376
rect 22005 28367 22063 28373
rect 23109 28373 23121 28407
rect 23155 28373 23167 28407
rect 23109 28367 23167 28373
rect 23658 28364 23664 28416
rect 23716 28364 23722 28416
rect 24118 28364 24124 28416
rect 24176 28364 24182 28416
rect 1104 28314 25000 28336
rect 1104 28262 6884 28314
rect 6936 28262 6948 28314
rect 7000 28262 7012 28314
rect 7064 28262 7076 28314
rect 7128 28262 7140 28314
rect 7192 28262 12818 28314
rect 12870 28262 12882 28314
rect 12934 28262 12946 28314
rect 12998 28262 13010 28314
rect 13062 28262 13074 28314
rect 13126 28262 18752 28314
rect 18804 28262 18816 28314
rect 18868 28262 18880 28314
rect 18932 28262 18944 28314
rect 18996 28262 19008 28314
rect 19060 28262 24686 28314
rect 24738 28262 24750 28314
rect 24802 28262 24814 28314
rect 24866 28262 24878 28314
rect 24930 28262 24942 28314
rect 24994 28262 25000 28314
rect 1104 28240 25000 28262
rect 2038 28160 2044 28212
rect 2096 28200 2102 28212
rect 2409 28203 2467 28209
rect 2409 28200 2421 28203
rect 2096 28172 2421 28200
rect 2096 28160 2102 28172
rect 2409 28169 2421 28172
rect 2455 28169 2467 28203
rect 2409 28163 2467 28169
rect 3510 28160 3516 28212
rect 3568 28160 3574 28212
rect 4065 28203 4123 28209
rect 4065 28169 4077 28203
rect 4111 28200 4123 28203
rect 4338 28200 4344 28212
rect 4111 28172 4344 28200
rect 4111 28169 4123 28172
rect 4065 28163 4123 28169
rect 4338 28160 4344 28172
rect 4396 28160 4402 28212
rect 4614 28160 4620 28212
rect 4672 28160 4678 28212
rect 5721 28203 5779 28209
rect 4908 28172 5672 28200
rect 2222 28092 2228 28144
rect 2280 28132 2286 28144
rect 3050 28132 3056 28144
rect 2280 28104 3056 28132
rect 2280 28092 2286 28104
rect 3050 28092 3056 28104
rect 3108 28092 3114 28144
rect 3528 28132 3556 28160
rect 4908 28132 4936 28172
rect 3528 28104 4936 28132
rect 5166 28092 5172 28144
rect 5224 28132 5230 28144
rect 5353 28135 5411 28141
rect 5353 28132 5365 28135
rect 5224 28104 5365 28132
rect 5224 28092 5230 28104
rect 5353 28101 5365 28104
rect 5399 28101 5411 28135
rect 5644 28132 5672 28172
rect 5721 28169 5733 28203
rect 5767 28200 5779 28203
rect 6546 28200 6552 28212
rect 5767 28172 6552 28200
rect 5767 28169 5779 28172
rect 5721 28163 5779 28169
rect 6546 28160 6552 28172
rect 6604 28160 6610 28212
rect 10962 28200 10968 28212
rect 7116 28172 10968 28200
rect 7116 28132 7144 28172
rect 5644 28104 7144 28132
rect 5353 28095 5411 28101
rect 7374 28092 7380 28144
rect 7432 28092 7438 28144
rect 1671 28067 1729 28073
rect 1671 28033 1683 28067
rect 1717 28064 1729 28067
rect 1762 28064 1768 28076
rect 1717 28036 1768 28064
rect 1717 28033 1729 28036
rect 1671 28027 1729 28033
rect 1762 28024 1768 28036
rect 1820 28064 1826 28076
rect 2498 28064 2504 28076
rect 1820 28036 2504 28064
rect 1820 28024 1826 28036
rect 2498 28024 2504 28036
rect 2556 28024 2562 28076
rect 2774 28024 2780 28076
rect 2832 28024 2838 28076
rect 3068 28064 3096 28092
rect 3295 28067 3353 28073
rect 3295 28064 3307 28067
rect 3068 28036 3307 28064
rect 3295 28033 3307 28036
rect 3341 28033 3353 28067
rect 4893 28067 4951 28073
rect 4893 28064 4905 28067
rect 3295 28027 3353 28033
rect 4356 28036 4905 28064
rect 1394 27956 1400 28008
rect 1452 27956 1458 28008
rect 2130 27956 2136 28008
rect 2188 27996 2194 28008
rect 2406 27996 2412 28008
rect 2188 27968 2412 27996
rect 2188 27956 2194 27968
rect 2406 27956 2412 27968
rect 2464 27956 2470 28008
rect 3053 27999 3111 28005
rect 3053 27996 3065 27999
rect 2746 27968 3065 27996
rect 2590 27928 2596 27940
rect 2148 27900 2596 27928
rect 2148 27872 2176 27900
rect 2590 27888 2596 27900
rect 2648 27888 2654 27940
rect 2130 27820 2136 27872
rect 2188 27820 2194 27872
rect 2314 27820 2320 27872
rect 2372 27860 2378 27872
rect 2746 27860 2774 27968
rect 3053 27965 3065 27968
rect 3099 27965 3111 27999
rect 3053 27959 3111 27965
rect 4356 27928 4384 28036
rect 4893 28033 4905 28036
rect 4939 28033 4951 28067
rect 4893 28027 4951 28033
rect 4985 28067 5043 28073
rect 4985 28033 4997 28067
rect 5031 28064 5043 28067
rect 5902 28064 5908 28076
rect 5031 28036 5908 28064
rect 5031 28033 5043 28036
rect 4985 28027 5043 28033
rect 5902 28024 5908 28036
rect 5960 28024 5966 28076
rect 7392 28064 7420 28092
rect 7300 28036 7420 28064
rect 7484 28064 7512 28172
rect 10962 28160 10968 28172
rect 11020 28160 11026 28212
rect 11057 28203 11115 28209
rect 11057 28169 11069 28203
rect 11103 28169 11115 28203
rect 11057 28163 11115 28169
rect 8662 28092 8668 28144
rect 8720 28132 8726 28144
rect 8720 28104 10088 28132
rect 8720 28092 8726 28104
rect 7543 28067 7601 28073
rect 7543 28064 7555 28067
rect 7484 28036 7555 28064
rect 5074 27956 5080 28008
rect 5132 27956 5138 28008
rect 6638 27956 6644 28008
rect 6696 27996 6702 28008
rect 7300 28005 7328 28036
rect 7543 28033 7555 28036
rect 7589 28033 7601 28067
rect 7543 28027 7601 28033
rect 8202 28024 8208 28076
rect 8260 28064 8266 28076
rect 8907 28067 8965 28073
rect 8907 28064 8919 28067
rect 8260 28036 8919 28064
rect 8260 28024 8266 28036
rect 8907 28033 8919 28036
rect 8953 28033 8965 28067
rect 8907 28027 8965 28033
rect 10060 28005 10088 28104
rect 10594 28092 10600 28144
rect 10652 28092 10658 28144
rect 10319 28067 10377 28073
rect 10319 28033 10331 28067
rect 10365 28064 10377 28067
rect 10612 28064 10640 28092
rect 10365 28036 10640 28064
rect 11072 28064 11100 28163
rect 11238 28160 11244 28212
rect 11296 28200 11302 28212
rect 11793 28203 11851 28209
rect 11793 28200 11805 28203
rect 11296 28172 11805 28200
rect 11296 28160 11302 28172
rect 11793 28169 11805 28172
rect 11839 28169 11851 28203
rect 11793 28163 11851 28169
rect 12434 28160 12440 28212
rect 12492 28200 12498 28212
rect 15746 28200 15752 28212
rect 12492 28172 15752 28200
rect 12492 28160 12498 28172
rect 15746 28160 15752 28172
rect 15804 28160 15810 28212
rect 17681 28203 17739 28209
rect 17681 28169 17693 28203
rect 17727 28200 17739 28203
rect 17862 28200 17868 28212
rect 17727 28172 17868 28200
rect 17727 28169 17739 28172
rect 17681 28163 17739 28169
rect 17862 28160 17868 28172
rect 17920 28160 17926 28212
rect 18414 28160 18420 28212
rect 18472 28160 18478 28212
rect 19429 28203 19487 28209
rect 19429 28169 19441 28203
rect 19475 28200 19487 28203
rect 19886 28200 19892 28212
rect 19475 28172 19892 28200
rect 19475 28169 19487 28172
rect 19429 28163 19487 28169
rect 19886 28160 19892 28172
rect 19944 28160 19950 28212
rect 20530 28160 20536 28212
rect 20588 28160 20594 28212
rect 21634 28160 21640 28212
rect 21692 28200 21698 28212
rect 21913 28203 21971 28209
rect 21913 28200 21925 28203
rect 21692 28172 21925 28200
rect 21692 28160 21698 28172
rect 21913 28169 21925 28172
rect 21959 28169 21971 28203
rect 21913 28163 21971 28169
rect 22186 28160 22192 28212
rect 22244 28160 22250 28212
rect 23201 28203 23259 28209
rect 23201 28169 23213 28203
rect 23247 28200 23259 28203
rect 23566 28200 23572 28212
rect 23247 28172 23572 28200
rect 23247 28169 23259 28172
rect 23201 28163 23259 28169
rect 23566 28160 23572 28172
rect 23624 28160 23630 28212
rect 23658 28160 23664 28212
rect 23716 28200 23722 28212
rect 23716 28172 24164 28200
rect 23716 28160 23722 28172
rect 17034 28132 17040 28144
rect 16776 28104 17040 28132
rect 11514 28064 11520 28076
rect 11072 28036 11520 28064
rect 10365 28033 10377 28036
rect 10319 28027 10377 28033
rect 11514 28024 11520 28036
rect 11572 28024 11578 28076
rect 11606 28024 11612 28076
rect 11664 28064 11670 28076
rect 11664 28036 12434 28064
rect 11664 28024 11670 28036
rect 7285 27999 7343 28005
rect 7285 27996 7297 27999
rect 6696 27968 7297 27996
rect 6696 27956 6702 27968
rect 7285 27965 7297 27968
rect 7331 27965 7343 27999
rect 7285 27959 7343 27965
rect 8665 27999 8723 28005
rect 8665 27965 8677 27999
rect 8711 27965 8723 27999
rect 8665 27959 8723 27965
rect 10045 27999 10103 28005
rect 10045 27965 10057 27999
rect 10091 27965 10103 27999
rect 10045 27959 10103 27965
rect 4356 27900 4476 27928
rect 4448 27872 4476 27900
rect 5902 27888 5908 27940
rect 5960 27888 5966 27940
rect 2372 27832 2774 27860
rect 2961 27863 3019 27869
rect 2372 27820 2378 27832
rect 2961 27829 2973 27863
rect 3007 27860 3019 27863
rect 4246 27860 4252 27872
rect 3007 27832 4252 27860
rect 3007 27829 3019 27832
rect 2961 27823 3019 27829
rect 4246 27820 4252 27832
rect 4304 27820 4310 27872
rect 4430 27820 4436 27872
rect 4488 27820 4494 27872
rect 8294 27820 8300 27872
rect 8352 27820 8358 27872
rect 8680 27860 8708 27959
rect 9122 27860 9128 27872
rect 8680 27832 9128 27860
rect 9122 27820 9128 27832
rect 9180 27820 9186 27872
rect 9674 27820 9680 27872
rect 9732 27820 9738 27872
rect 10060 27860 10088 27959
rect 11790 27956 11796 28008
rect 11848 27956 11854 28008
rect 10318 27860 10324 27872
rect 10060 27832 10324 27860
rect 10318 27820 10324 27832
rect 10376 27820 10382 27872
rect 11238 27820 11244 27872
rect 11296 27860 11302 27872
rect 11609 27863 11667 27869
rect 11609 27860 11621 27863
rect 11296 27832 11621 27860
rect 11296 27820 11302 27832
rect 11609 27829 11621 27832
rect 11655 27829 11667 27863
rect 12406 27860 12434 28036
rect 14734 28024 14740 28076
rect 14792 28064 14798 28076
rect 15071 28067 15129 28073
rect 15071 28064 15083 28067
rect 14792 28036 15083 28064
rect 14792 28024 14798 28036
rect 15071 28033 15083 28036
rect 15117 28033 15129 28067
rect 15071 28027 15129 28033
rect 15930 28024 15936 28076
rect 15988 28024 15994 28076
rect 16669 28070 16727 28073
rect 16776 28070 16804 28104
rect 17034 28092 17040 28104
rect 17092 28092 17098 28144
rect 18294 28135 18352 28141
rect 18294 28101 18306 28135
rect 18340 28132 18352 28135
rect 18432 28132 18460 28160
rect 18690 28132 18696 28144
rect 18340 28104 18696 28132
rect 18340 28101 18352 28104
rect 18294 28095 18352 28101
rect 18690 28092 18696 28104
rect 18748 28092 18754 28144
rect 18782 28092 18788 28144
rect 18840 28132 18846 28144
rect 19610 28132 19616 28144
rect 18840 28104 19616 28132
rect 18840 28092 18846 28104
rect 19610 28092 19616 28104
rect 19668 28092 19674 28144
rect 16669 28067 16804 28070
rect 16669 28033 16681 28067
rect 16715 28042 16804 28067
rect 16715 28033 16727 28042
rect 16669 28027 16727 28033
rect 16850 28024 16856 28076
rect 16908 28064 16914 28076
rect 16943 28067 17001 28073
rect 16943 28064 16955 28067
rect 16908 28036 16955 28064
rect 16908 28024 16914 28036
rect 16943 28033 16955 28036
rect 16989 28033 17001 28067
rect 16943 28027 17001 28033
rect 19795 28067 19853 28073
rect 19795 28033 19807 28067
rect 19841 28064 19853 28067
rect 20254 28064 20260 28076
rect 19841 28036 20260 28064
rect 19841 28033 19853 28036
rect 19795 28027 19853 28033
rect 20254 28024 20260 28036
rect 20312 28024 20318 28076
rect 20548 28064 20576 28160
rect 22204 28132 22232 28160
rect 24136 28141 24164 28172
rect 24121 28135 24179 28141
rect 22204 28104 22692 28132
rect 21361 28067 21419 28073
rect 21361 28064 21373 28067
rect 20548 28036 21373 28064
rect 21361 28033 21373 28036
rect 21407 28033 21419 28067
rect 21361 28027 21419 28033
rect 22094 28024 22100 28076
rect 22152 28024 22158 28076
rect 22554 28064 22560 28076
rect 22296 28036 22560 28064
rect 14826 27956 14832 28008
rect 14884 27956 14890 28008
rect 15841 27931 15899 27937
rect 15841 27897 15853 27931
rect 15887 27928 15899 27931
rect 15948 27928 15976 28024
rect 18049 27999 18107 28005
rect 18049 27965 18061 27999
rect 18095 27965 18107 27999
rect 18049 27959 18107 27965
rect 15887 27900 15976 27928
rect 15887 27897 15899 27900
rect 15841 27891 15899 27897
rect 17862 27888 17868 27940
rect 17920 27928 17926 27940
rect 18064 27928 18092 27959
rect 19426 27956 19432 28008
rect 19484 27996 19490 28008
rect 19521 27999 19579 28005
rect 19521 27996 19533 27999
rect 19484 27968 19533 27996
rect 19484 27956 19490 27968
rect 19521 27965 19533 27968
rect 19567 27965 19579 27999
rect 19521 27959 19579 27965
rect 17920 27900 18092 27928
rect 21177 27931 21235 27937
rect 17920 27888 17926 27900
rect 21177 27897 21189 27931
rect 21223 27928 21235 27931
rect 22296 27928 22324 28036
rect 22554 28024 22560 28036
rect 22612 28024 22618 28076
rect 22664 28073 22692 28104
rect 24121 28101 24133 28135
rect 24167 28101 24179 28135
rect 24121 28095 24179 28101
rect 22649 28067 22707 28073
rect 22649 28033 22661 28067
rect 22695 28033 22707 28067
rect 22649 28027 22707 28033
rect 23385 28067 23443 28073
rect 23385 28033 23397 28067
rect 23431 28033 23443 28067
rect 23385 28027 23443 28033
rect 23400 27996 23428 28027
rect 23842 28024 23848 28076
rect 23900 28024 23906 28076
rect 22480 27968 23428 27996
rect 22480 27937 22508 27968
rect 21223 27900 22324 27928
rect 22465 27931 22523 27937
rect 21223 27897 21235 27900
rect 21177 27891 21235 27897
rect 22465 27897 22477 27931
rect 22511 27897 22523 27931
rect 22465 27891 22523 27897
rect 19334 27860 19340 27872
rect 12406 27832 19340 27860
rect 11609 27823 11667 27829
rect 19334 27820 19340 27832
rect 19392 27820 19398 27872
rect 19794 27820 19800 27872
rect 19852 27860 19858 27872
rect 20533 27863 20591 27869
rect 20533 27860 20545 27863
rect 19852 27832 20545 27860
rect 19852 27820 19858 27832
rect 20533 27829 20545 27832
rect 20579 27829 20591 27863
rect 20533 27823 20591 27829
rect 23658 27820 23664 27872
rect 23716 27820 23722 27872
rect 24394 27820 24400 27872
rect 24452 27820 24458 27872
rect 1104 27770 24840 27792
rect 1104 27718 3917 27770
rect 3969 27718 3981 27770
rect 4033 27718 4045 27770
rect 4097 27718 4109 27770
rect 4161 27718 4173 27770
rect 4225 27718 9851 27770
rect 9903 27718 9915 27770
rect 9967 27718 9979 27770
rect 10031 27718 10043 27770
rect 10095 27718 10107 27770
rect 10159 27718 15785 27770
rect 15837 27718 15849 27770
rect 15901 27718 15913 27770
rect 15965 27718 15977 27770
rect 16029 27718 16041 27770
rect 16093 27718 21719 27770
rect 21771 27718 21783 27770
rect 21835 27718 21847 27770
rect 21899 27718 21911 27770
rect 21963 27718 21975 27770
rect 22027 27718 24840 27770
rect 1104 27696 24840 27718
rect 1854 27616 1860 27668
rect 1912 27656 1918 27668
rect 3602 27656 3608 27668
rect 1912 27628 3608 27656
rect 1912 27616 1918 27628
rect 3602 27616 3608 27628
rect 3660 27616 3666 27668
rect 3694 27616 3700 27668
rect 3752 27656 3758 27668
rect 3752 27628 5396 27656
rect 3752 27616 3758 27628
rect 2866 27548 2872 27600
rect 2924 27588 2930 27600
rect 2961 27591 3019 27597
rect 2961 27588 2973 27591
rect 2924 27560 2973 27588
rect 2924 27548 2930 27560
rect 2961 27557 2973 27560
rect 3007 27557 3019 27591
rect 2961 27551 3019 27557
rect 3513 27591 3571 27597
rect 3513 27557 3525 27591
rect 3559 27588 3571 27591
rect 4614 27588 4620 27600
rect 3559 27560 4620 27588
rect 3559 27557 3571 27560
rect 3513 27551 3571 27557
rect 4614 27548 4620 27560
rect 4672 27548 4678 27600
rect 4154 27480 4160 27532
rect 4212 27520 4218 27532
rect 4338 27520 4344 27532
rect 4212 27492 4344 27520
rect 4212 27480 4218 27492
rect 4338 27480 4344 27492
rect 4396 27480 4402 27532
rect 5368 27520 5396 27628
rect 5534 27616 5540 27668
rect 5592 27656 5598 27668
rect 6086 27656 6092 27668
rect 5592 27628 6092 27656
rect 5592 27616 5598 27628
rect 6086 27616 6092 27628
rect 6144 27616 6150 27668
rect 11238 27616 11244 27668
rect 11296 27616 11302 27668
rect 11517 27659 11575 27665
rect 11517 27625 11529 27659
rect 11563 27656 11575 27659
rect 11790 27656 11796 27668
rect 11563 27628 11796 27656
rect 11563 27625 11575 27628
rect 11517 27619 11575 27625
rect 11790 27616 11796 27628
rect 11848 27616 11854 27668
rect 11992 27628 12570 27656
rect 5629 27591 5687 27597
rect 5629 27557 5641 27591
rect 5675 27588 5687 27591
rect 10597 27591 10655 27597
rect 5675 27560 6040 27588
rect 5675 27557 5687 27560
rect 5629 27551 5687 27557
rect 5902 27520 5908 27532
rect 5368 27492 5908 27520
rect 1394 27412 1400 27464
rect 1452 27412 1458 27464
rect 1671 27455 1729 27461
rect 1671 27452 1683 27455
rect 1596 27424 1683 27452
rect 1596 27396 1624 27424
rect 1671 27421 1683 27424
rect 1717 27421 1729 27455
rect 1671 27415 1729 27421
rect 2222 27412 2228 27464
rect 2280 27452 2286 27464
rect 2280 27448 2728 27452
rect 2769 27451 2827 27457
rect 2769 27448 2781 27451
rect 2280 27424 2781 27448
rect 2280 27412 2286 27424
rect 2700 27420 2781 27424
rect 2769 27417 2781 27420
rect 2815 27417 2827 27451
rect 2769 27411 2827 27417
rect 2958 27412 2964 27464
rect 3016 27452 3022 27464
rect 3053 27455 3111 27461
rect 3053 27452 3065 27455
rect 3016 27424 3065 27452
rect 3016 27412 3022 27424
rect 3053 27421 3065 27424
rect 3099 27421 3111 27455
rect 3053 27415 3111 27421
rect 3329 27455 3387 27461
rect 3329 27421 3341 27455
rect 3375 27421 3387 27455
rect 3329 27415 3387 27421
rect 1578 27344 1584 27396
rect 1636 27344 1642 27396
rect 3344 27384 3372 27415
rect 3786 27412 3792 27464
rect 3844 27412 3850 27464
rect 4617 27455 4675 27461
rect 4617 27421 4629 27455
rect 4663 27452 4675 27455
rect 4798 27452 4804 27464
rect 4663 27424 4804 27452
rect 4663 27421 4675 27424
rect 4617 27415 4675 27421
rect 4798 27412 4804 27424
rect 4856 27412 4862 27464
rect 4891 27455 4949 27461
rect 4891 27421 4903 27455
rect 4937 27452 4949 27455
rect 5368 27452 5396 27492
rect 5902 27480 5908 27492
rect 5960 27480 5966 27532
rect 6012 27506 6040 27560
rect 10597 27557 10609 27591
rect 10643 27588 10655 27591
rect 11992 27588 12020 27628
rect 10643 27560 12020 27588
rect 12542 27588 12570 27628
rect 14292 27628 14872 27656
rect 13538 27588 13544 27600
rect 12542 27560 13544 27588
rect 10643 27557 10655 27560
rect 10597 27551 10655 27557
rect 13538 27548 13544 27560
rect 13596 27548 13602 27600
rect 14292 27588 14320 27628
rect 13648 27560 14320 27588
rect 14844 27588 14872 27628
rect 17678 27616 17684 27668
rect 17736 27656 17742 27668
rect 22094 27656 22100 27668
rect 17736 27628 22100 27656
rect 17736 27616 17742 27628
rect 22094 27616 22100 27628
rect 22152 27616 22158 27668
rect 22296 27628 22782 27656
rect 14844 27560 17080 27588
rect 7834 27480 7840 27532
rect 7892 27520 7898 27532
rect 8202 27520 8208 27532
rect 7892 27492 8208 27520
rect 7892 27480 7898 27492
rect 8202 27480 8208 27492
rect 8260 27480 8266 27532
rect 9674 27480 9680 27532
rect 9732 27480 9738 27532
rect 10962 27480 10968 27532
rect 11020 27520 11026 27532
rect 11020 27492 11744 27520
rect 11020 27480 11026 27492
rect 4937 27424 5396 27452
rect 4937 27421 4949 27424
rect 4891 27415 4949 27421
rect 5442 27412 5448 27464
rect 5500 27452 5506 27464
rect 5500 27424 6224 27452
rect 5500 27412 5506 27424
rect 6196 27393 6224 27424
rect 6454 27412 6460 27464
rect 6512 27412 6518 27464
rect 6549 27455 6607 27461
rect 6549 27421 6561 27455
rect 6595 27452 6607 27455
rect 7282 27452 7288 27464
rect 6595 27424 7288 27452
rect 6595 27421 6607 27424
rect 6549 27415 6607 27421
rect 7282 27412 7288 27424
rect 7340 27412 7346 27464
rect 7558 27412 7564 27464
rect 7616 27452 7622 27464
rect 8018 27452 8024 27464
rect 7616 27424 8024 27452
rect 7616 27412 7622 27424
rect 8018 27412 8024 27424
rect 8076 27412 8082 27464
rect 9508 27424 10824 27452
rect 6181 27387 6239 27393
rect 2884 27356 3372 27384
rect 3896 27356 6132 27384
rect 2406 27276 2412 27328
rect 2464 27276 2470 27328
rect 2590 27276 2596 27328
rect 2648 27316 2654 27328
rect 2884 27316 2912 27356
rect 2648 27288 2912 27316
rect 3237 27319 3295 27325
rect 2648 27276 2654 27288
rect 3237 27285 3249 27319
rect 3283 27316 3295 27319
rect 3896 27316 3924 27356
rect 3283 27288 3924 27316
rect 3973 27319 4031 27325
rect 3283 27285 3295 27288
rect 3237 27279 3295 27285
rect 3973 27285 3985 27319
rect 4019 27316 4031 27319
rect 5442 27316 5448 27328
rect 4019 27288 5448 27316
rect 4019 27285 4031 27288
rect 3973 27279 4031 27285
rect 5442 27276 5448 27288
rect 5500 27276 5506 27328
rect 6104 27316 6132 27356
rect 6181 27353 6193 27387
rect 6227 27353 6239 27387
rect 6181 27347 6239 27353
rect 6914 27344 6920 27396
rect 6972 27344 6978 27396
rect 9508 27384 9536 27424
rect 7208 27356 9536 27384
rect 7208 27316 7236 27356
rect 9582 27344 9588 27396
rect 9640 27344 9646 27396
rect 9674 27344 9680 27396
rect 9732 27344 9738 27396
rect 10042 27344 10048 27396
rect 10100 27344 10106 27396
rect 10796 27384 10824 27424
rect 11146 27412 11152 27464
rect 11204 27412 11210 27464
rect 11425 27455 11483 27461
rect 11425 27421 11437 27455
rect 11471 27452 11483 27455
rect 11514 27452 11520 27464
rect 11471 27424 11520 27452
rect 11471 27421 11483 27424
rect 11425 27415 11483 27421
rect 11514 27412 11520 27424
rect 11572 27412 11578 27464
rect 11606 27412 11612 27464
rect 11664 27412 11670 27464
rect 11716 27452 11744 27492
rect 11882 27480 11888 27532
rect 11940 27480 11946 27532
rect 13170 27480 13176 27532
rect 13228 27520 13234 27532
rect 13648 27520 13676 27560
rect 17052 27532 17080 27560
rect 17310 27548 17316 27600
rect 17368 27588 17374 27600
rect 17368 27560 17632 27588
rect 17368 27548 17374 27560
rect 17604 27532 17632 27560
rect 18230 27548 18236 27600
rect 18288 27588 18294 27600
rect 18288 27560 20024 27588
rect 18288 27548 18294 27560
rect 13228 27492 13676 27520
rect 13228 27480 13234 27492
rect 17034 27480 17040 27532
rect 17092 27520 17098 27532
rect 17402 27520 17408 27532
rect 17092 27492 17408 27520
rect 17092 27480 17098 27492
rect 17402 27480 17408 27492
rect 17460 27480 17466 27532
rect 17586 27480 17592 27532
rect 17644 27480 17650 27532
rect 18690 27480 18696 27532
rect 18748 27520 18754 27532
rect 19429 27523 19487 27529
rect 18748 27492 18828 27520
rect 18748 27480 18754 27492
rect 12159 27455 12217 27461
rect 12159 27452 12171 27455
rect 11716 27424 12171 27452
rect 12159 27421 12171 27424
rect 12205 27452 12217 27455
rect 12526 27452 12532 27464
rect 12205 27424 12532 27452
rect 12205 27421 12217 27424
rect 12159 27415 12217 27421
rect 12526 27412 12532 27424
rect 12584 27412 12590 27464
rect 14182 27412 14188 27464
rect 14240 27452 14246 27464
rect 14366 27452 14372 27464
rect 14240 27424 14372 27452
rect 14240 27412 14246 27424
rect 14366 27412 14372 27424
rect 14424 27412 14430 27464
rect 14459 27455 14517 27461
rect 14459 27421 14471 27455
rect 14505 27452 14517 27455
rect 14826 27452 14832 27464
rect 14505 27424 14832 27452
rect 14505 27421 14517 27424
rect 14459 27415 14517 27421
rect 14826 27412 14832 27424
rect 14884 27412 14890 27464
rect 18800 27461 18828 27492
rect 19429 27489 19441 27523
rect 19475 27520 19487 27523
rect 19889 27523 19947 27529
rect 19889 27520 19901 27523
rect 19475 27492 19901 27520
rect 19475 27489 19487 27492
rect 19429 27483 19487 27489
rect 19889 27489 19901 27492
rect 19935 27489 19947 27523
rect 19889 27483 19947 27489
rect 18785 27455 18843 27461
rect 18785 27421 18797 27455
rect 18831 27421 18843 27455
rect 18785 27415 18843 27421
rect 19337 27455 19395 27461
rect 19337 27421 19349 27455
rect 19383 27421 19395 27455
rect 19337 27415 19395 27421
rect 14550 27384 14556 27396
rect 10796 27356 14556 27384
rect 14550 27344 14556 27356
rect 14608 27344 14614 27396
rect 19352 27384 19380 27415
rect 19794 27412 19800 27464
rect 19852 27412 19858 27464
rect 19996 27452 20024 27560
rect 20070 27480 20076 27532
rect 20128 27480 20134 27532
rect 22296 27452 22324 27628
rect 22754 27464 22782 27628
rect 23842 27616 23848 27668
rect 23900 27616 23906 27668
rect 23109 27591 23167 27597
rect 23109 27557 23121 27591
rect 23155 27588 23167 27591
rect 23860 27588 23888 27616
rect 23155 27560 23888 27588
rect 23155 27557 23167 27560
rect 23109 27551 23167 27557
rect 22649 27455 22707 27461
rect 22649 27452 22661 27455
rect 19996 27424 22324 27452
rect 22388 27424 22661 27452
rect 18616 27356 19380 27384
rect 6104 27288 7236 27316
rect 7285 27319 7343 27325
rect 7285 27285 7297 27319
rect 7331 27316 7343 27319
rect 7374 27316 7380 27328
rect 7331 27288 7380 27316
rect 7331 27285 7343 27288
rect 7285 27279 7343 27285
rect 7374 27276 7380 27288
rect 7432 27276 7438 27328
rect 7466 27276 7472 27328
rect 7524 27276 7530 27328
rect 7834 27276 7840 27328
rect 7892 27316 7898 27328
rect 8386 27316 8392 27328
rect 7892 27288 8392 27316
rect 7892 27276 7898 27288
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 9309 27319 9367 27325
rect 9309 27285 9321 27319
rect 9355 27316 9367 27319
rect 10318 27316 10324 27328
rect 9355 27288 10324 27316
rect 9355 27285 9367 27288
rect 9309 27279 9367 27285
rect 10318 27276 10324 27288
rect 10376 27276 10382 27328
rect 10410 27276 10416 27328
rect 10468 27276 10474 27328
rect 11882 27276 11888 27328
rect 11940 27316 11946 27328
rect 12342 27316 12348 27328
rect 11940 27288 12348 27316
rect 11940 27276 11946 27288
rect 12342 27276 12348 27288
rect 12400 27276 12406 27328
rect 12710 27276 12716 27328
rect 12768 27316 12774 27328
rect 12897 27319 12955 27325
rect 12897 27316 12909 27319
rect 12768 27288 12909 27316
rect 12768 27276 12774 27288
rect 12897 27285 12909 27288
rect 12943 27285 12955 27319
rect 12897 27279 12955 27285
rect 14734 27276 14740 27328
rect 14792 27316 14798 27328
rect 18616 27325 18644 27356
rect 20898 27344 20904 27396
rect 20956 27384 20962 27396
rect 22388 27384 22416 27424
rect 22649 27421 22661 27424
rect 22695 27421 22707 27455
rect 22649 27415 22707 27421
rect 22738 27412 22744 27464
rect 22796 27452 22802 27464
rect 23017 27455 23075 27461
rect 23017 27452 23029 27455
rect 22796 27424 23029 27452
rect 22796 27412 22802 27424
rect 23017 27421 23029 27424
rect 23063 27421 23075 27455
rect 23017 27415 23075 27421
rect 23293 27455 23351 27461
rect 23293 27421 23305 27455
rect 23339 27421 23351 27455
rect 23293 27415 23351 27421
rect 23385 27455 23443 27461
rect 23385 27421 23397 27455
rect 23431 27452 23443 27455
rect 23658 27452 23664 27464
rect 23431 27424 23664 27452
rect 23431 27421 23443 27424
rect 23385 27415 23443 27421
rect 23308 27384 23336 27415
rect 23658 27412 23664 27424
rect 23716 27412 23722 27464
rect 23750 27412 23756 27464
rect 23808 27452 23814 27464
rect 23845 27455 23903 27461
rect 23845 27452 23857 27455
rect 23808 27424 23857 27452
rect 23808 27412 23814 27424
rect 23845 27421 23857 27424
rect 23891 27421 23903 27455
rect 23845 27415 23903 27421
rect 20956 27356 22416 27384
rect 22480 27356 23336 27384
rect 24213 27387 24271 27393
rect 20956 27344 20962 27356
rect 15197 27319 15255 27325
rect 15197 27316 15209 27319
rect 14792 27288 15209 27316
rect 14792 27276 14798 27288
rect 15197 27285 15209 27288
rect 15243 27285 15255 27319
rect 15197 27279 15255 27285
rect 18601 27319 18659 27325
rect 18601 27285 18613 27319
rect 18647 27285 18659 27319
rect 18601 27279 18659 27285
rect 20073 27319 20131 27325
rect 20073 27285 20085 27319
rect 20119 27316 20131 27319
rect 21910 27316 21916 27328
rect 20119 27288 21916 27316
rect 20119 27285 20131 27288
rect 20073 27279 20131 27285
rect 21910 27276 21916 27288
rect 21968 27276 21974 27328
rect 22480 27325 22508 27356
rect 24213 27353 24225 27387
rect 24259 27384 24271 27387
rect 25130 27384 25136 27396
rect 24259 27356 25136 27384
rect 24259 27353 24271 27356
rect 24213 27347 24271 27353
rect 25130 27344 25136 27356
rect 25188 27344 25194 27396
rect 22465 27319 22523 27325
rect 22465 27285 22477 27319
rect 22511 27285 22523 27319
rect 22465 27279 22523 27285
rect 22830 27276 22836 27328
rect 22888 27276 22894 27328
rect 23566 27276 23572 27328
rect 23624 27276 23630 27328
rect 1104 27226 25000 27248
rect 1104 27174 6884 27226
rect 6936 27174 6948 27226
rect 7000 27174 7012 27226
rect 7064 27174 7076 27226
rect 7128 27174 7140 27226
rect 7192 27174 12818 27226
rect 12870 27174 12882 27226
rect 12934 27174 12946 27226
rect 12998 27174 13010 27226
rect 13062 27174 13074 27226
rect 13126 27174 18752 27226
rect 18804 27174 18816 27226
rect 18868 27174 18880 27226
rect 18932 27174 18944 27226
rect 18996 27174 19008 27226
rect 19060 27174 24686 27226
rect 24738 27174 24750 27226
rect 24802 27174 24814 27226
rect 24866 27174 24878 27226
rect 24930 27174 24942 27226
rect 24994 27174 25000 27226
rect 1104 27152 25000 27174
rect 1765 27115 1823 27121
rect 1765 27081 1777 27115
rect 1811 27112 1823 27115
rect 2130 27112 2136 27124
rect 1811 27084 2136 27112
rect 1811 27081 1823 27084
rect 1765 27075 1823 27081
rect 2130 27072 2136 27084
rect 2188 27072 2194 27124
rect 3050 27072 3056 27124
rect 3108 27072 3114 27124
rect 3697 27115 3755 27121
rect 3697 27081 3709 27115
rect 3743 27112 3755 27115
rect 3743 27084 9076 27112
rect 3743 27081 3755 27084
rect 3697 27075 3755 27081
rect 1302 27004 1308 27056
rect 1360 27044 1366 27056
rect 2869 27047 2927 27053
rect 1360 27016 2774 27044
rect 1360 27004 1366 27016
rect 474 26976 480 26988
rect 308 26948 480 26976
rect 308 26920 336 26948
rect 474 26936 480 26948
rect 532 26936 538 26988
rect 2038 26936 2044 26988
rect 2096 26936 2102 26988
rect 2130 26936 2136 26988
rect 2188 26936 2194 26988
rect 2498 26936 2504 26988
rect 2556 26936 2562 26988
rect 2746 26976 2774 27016
rect 2869 27013 2881 27047
rect 2915 27044 2927 27047
rect 4338 27044 4344 27056
rect 2915 27016 3740 27044
rect 2915 27013 2927 27016
rect 2869 27007 2927 27013
rect 3513 26979 3571 26985
rect 3513 26976 3525 26979
rect 2746 26948 3525 26976
rect 3513 26945 3525 26948
rect 3559 26945 3571 26979
rect 3513 26939 3571 26945
rect 290 26868 296 26920
rect 348 26868 354 26920
rect 2406 26868 2412 26920
rect 2464 26868 2470 26920
rect 1578 26772 1584 26784
rect 1044 26744 1584 26772
rect 14 26596 20 26648
rect 72 26636 78 26648
rect 842 26636 848 26648
rect 72 26608 848 26636
rect 72 26596 78 26608
rect 842 26596 848 26608
rect 900 26596 906 26648
rect 1044 26568 1072 26744
rect 1578 26732 1584 26744
rect 1636 26732 1642 26784
rect 3712 26772 3740 27016
rect 3804 27016 4344 27044
rect 3804 26985 3832 27016
rect 4338 27004 4344 27016
rect 4396 27044 4402 27056
rect 4522 27044 4528 27056
rect 4396 27016 4528 27044
rect 4396 27004 4402 27016
rect 4522 27004 4528 27016
rect 4580 27004 4586 27056
rect 4798 27004 4804 27056
rect 4856 27044 4862 27056
rect 6270 27044 6276 27056
rect 4856 27016 6276 27044
rect 4856 27004 4862 27016
rect 6270 27004 6276 27016
rect 6328 27004 6334 27056
rect 7558 27004 7564 27056
rect 7616 27044 7622 27056
rect 7745 27047 7803 27053
rect 7745 27044 7757 27047
rect 7616 27016 7757 27044
rect 7616 27004 7622 27016
rect 7745 27013 7757 27016
rect 7791 27013 7803 27047
rect 7745 27007 7803 27013
rect 7834 27004 7840 27056
rect 7892 27044 7898 27056
rect 8021 27047 8079 27053
rect 8021 27044 8033 27047
rect 7892 27016 8033 27044
rect 7892 27004 7898 27016
rect 8021 27013 8033 27016
rect 8067 27013 8079 27047
rect 8021 27007 8079 27013
rect 8113 27047 8171 27053
rect 8113 27013 8125 27047
rect 8159 27044 8171 27047
rect 8294 27044 8300 27056
rect 8159 27016 8300 27044
rect 8159 27013 8171 27016
rect 8113 27007 8171 27013
rect 8294 27004 8300 27016
rect 8352 27004 8358 27056
rect 8481 27047 8539 27053
rect 8481 27013 8493 27047
rect 8527 27044 8539 27047
rect 9048 27044 9076 27084
rect 9674 27072 9680 27124
rect 9732 27112 9738 27124
rect 10321 27115 10379 27121
rect 10321 27112 10333 27115
rect 9732 27084 10333 27112
rect 9732 27072 9738 27084
rect 10321 27081 10333 27084
rect 10367 27081 10379 27115
rect 10321 27075 10379 27081
rect 11146 27072 11152 27124
rect 11204 27072 11210 27124
rect 11606 27072 11612 27124
rect 11664 27072 11670 27124
rect 11885 27115 11943 27121
rect 11885 27081 11897 27115
rect 11931 27081 11943 27115
rect 11885 27075 11943 27081
rect 11054 27044 11060 27056
rect 8527 27016 8984 27044
rect 9048 27016 11060 27044
rect 8527 27013 8539 27016
rect 8481 27007 8539 27013
rect 3789 26979 3847 26985
rect 3789 26945 3801 26979
rect 3835 26945 3847 26979
rect 3789 26939 3847 26945
rect 4063 26979 4121 26985
rect 4063 26945 4075 26979
rect 4109 26976 4121 26979
rect 4154 26976 4160 26988
rect 4109 26948 4160 26976
rect 4109 26945 4121 26948
rect 4063 26939 4121 26945
rect 4154 26936 4160 26948
rect 4212 26976 4218 26988
rect 4614 26976 4620 26988
rect 4212 26948 4620 26976
rect 4212 26936 4218 26948
rect 4614 26936 4620 26948
rect 4672 26936 4678 26988
rect 8496 26976 8524 27007
rect 4724 26948 8524 26976
rect 4724 26772 4752 26948
rect 8846 26936 8852 26988
rect 8904 26985 8910 26988
rect 8904 26979 8921 26985
rect 8909 26945 8921 26979
rect 8956 26976 8984 27016
rect 11054 27004 11060 27016
rect 11112 27004 11118 27056
rect 11164 27044 11192 27072
rect 11900 27044 11928 27075
rect 12434 27072 12440 27124
rect 12492 27112 12498 27124
rect 15381 27115 15439 27121
rect 12492 27084 15240 27112
rect 12492 27072 12498 27084
rect 15212 27044 15240 27084
rect 15381 27081 15393 27115
rect 15427 27112 15439 27115
rect 18230 27112 18236 27124
rect 15427 27084 18236 27112
rect 15427 27081 15439 27084
rect 15381 27075 15439 27081
rect 18230 27072 18236 27084
rect 18288 27072 18294 27124
rect 21821 27115 21879 27121
rect 21821 27081 21833 27115
rect 21867 27081 21879 27115
rect 21821 27075 21879 27081
rect 20898 27044 20904 27056
rect 11164 27016 11928 27044
rect 11992 27016 13768 27044
rect 15212 27016 20904 27044
rect 9030 26976 9036 26988
rect 8956 26948 9036 26976
rect 8904 26939 8921 26945
rect 8904 26936 8910 26939
rect 9030 26936 9036 26948
rect 9088 26936 9094 26988
rect 9214 26936 9220 26988
rect 9272 26976 9278 26988
rect 9551 26979 9609 26985
rect 9551 26976 9563 26979
rect 9272 26948 9563 26976
rect 9272 26936 9278 26948
rect 9551 26945 9563 26948
rect 9597 26945 9609 26979
rect 9551 26939 9609 26945
rect 10134 26936 10140 26988
rect 10192 26936 10198 26988
rect 11606 26936 11612 26988
rect 11664 26976 11670 26988
rect 11793 26979 11851 26985
rect 11793 26976 11805 26979
rect 11664 26948 11805 26976
rect 11664 26936 11670 26948
rect 11793 26945 11805 26948
rect 11839 26945 11851 26979
rect 11793 26939 11851 26945
rect 8294 26868 8300 26920
rect 8352 26868 8358 26920
rect 9122 26868 9128 26920
rect 9180 26908 9186 26920
rect 9309 26911 9367 26917
rect 9309 26908 9321 26911
rect 9180 26880 9321 26908
rect 9180 26868 9186 26880
rect 9309 26877 9321 26880
rect 9355 26877 9367 26911
rect 9309 26871 9367 26877
rect 10152 26840 10180 26936
rect 10410 26868 10416 26920
rect 10468 26908 10474 26920
rect 11992 26908 12020 27016
rect 13740 26988 13768 27016
rect 20898 27004 20904 27016
rect 20956 27004 20962 27056
rect 21836 27044 21864 27075
rect 21910 27072 21916 27124
rect 21968 27112 21974 27124
rect 21968 27084 23980 27112
rect 21968 27072 21974 27084
rect 22640 27047 22698 27053
rect 21836 27016 22324 27044
rect 12066 26936 12072 26988
rect 12124 26936 12130 26988
rect 12342 26936 12348 26988
rect 12400 26976 12406 26988
rect 12435 26979 12493 26985
rect 12435 26976 12447 26979
rect 12400 26948 12447 26976
rect 12400 26936 12406 26948
rect 12435 26945 12447 26948
rect 12481 26976 12493 26979
rect 13630 26976 13636 26988
rect 12481 26948 13636 26976
rect 12481 26945 12493 26948
rect 12435 26939 12493 26945
rect 13630 26936 13636 26948
rect 13688 26936 13694 26988
rect 13722 26936 13728 26988
rect 13780 26936 13786 26988
rect 14550 26936 14556 26988
rect 14608 26985 14614 26988
rect 14608 26979 14636 26985
rect 14624 26945 14636 26979
rect 14608 26939 14636 26945
rect 14608 26936 14614 26939
rect 14734 26936 14740 26988
rect 14792 26936 14798 26988
rect 16943 26979 17001 26985
rect 16943 26945 16955 26979
rect 16989 26976 17001 26979
rect 17402 26976 17408 26988
rect 16989 26948 17408 26976
rect 16989 26945 17001 26948
rect 16943 26939 17001 26945
rect 17402 26936 17408 26948
rect 17460 26976 17466 26988
rect 19978 26976 19984 26988
rect 17460 26948 19984 26976
rect 17460 26936 17466 26948
rect 19978 26936 19984 26948
rect 20036 26936 20042 26988
rect 21358 26936 21364 26988
rect 21416 26976 21422 26988
rect 22005 26979 22063 26985
rect 22005 26976 22017 26979
rect 21416 26948 22017 26976
rect 21416 26936 21422 26948
rect 22005 26945 22017 26948
rect 22051 26945 22063 26979
rect 22005 26939 22063 26945
rect 22097 26979 22155 26985
rect 22097 26945 22109 26979
rect 22143 26976 22155 26979
rect 22186 26976 22192 26988
rect 22143 26948 22192 26976
rect 22143 26945 22155 26948
rect 22097 26939 22155 26945
rect 22186 26936 22192 26948
rect 22244 26936 22250 26988
rect 22296 26985 22324 27016
rect 22640 27013 22652 27047
rect 22686 27044 22698 27047
rect 22738 27044 22744 27056
rect 22686 27016 22744 27044
rect 22686 27013 22698 27016
rect 22640 27007 22698 27013
rect 22738 27004 22744 27016
rect 22796 27004 22802 27056
rect 23952 27053 23980 27084
rect 23937 27047 23995 27053
rect 23937 27013 23949 27047
rect 23983 27013 23995 27047
rect 23937 27007 23995 27013
rect 22281 26979 22339 26985
rect 22281 26945 22293 26979
rect 22327 26945 22339 26979
rect 22281 26939 22339 26945
rect 10468 26880 12020 26908
rect 10468 26868 10474 26880
rect 12158 26868 12164 26920
rect 12216 26868 12222 26920
rect 13538 26908 13544 26920
rect 13096 26880 13544 26908
rect 10152 26812 12296 26840
rect 12268 26784 12296 26812
rect 3712 26744 4752 26772
rect 4798 26732 4804 26784
rect 4856 26732 4862 26784
rect 9033 26775 9091 26781
rect 9033 26741 9045 26775
rect 9079 26772 9091 26775
rect 11054 26772 11060 26784
rect 9079 26744 11060 26772
rect 9079 26741 9091 26744
rect 9033 26735 9091 26741
rect 11054 26732 11060 26744
rect 11112 26732 11118 26784
rect 12250 26732 12256 26784
rect 12308 26732 12314 26784
rect 12434 26732 12440 26784
rect 12492 26772 12498 26784
rect 13096 26772 13124 26880
rect 13538 26868 13544 26880
rect 13596 26868 13602 26920
rect 13906 26868 13912 26920
rect 13964 26908 13970 26920
rect 14185 26911 14243 26917
rect 14185 26908 14197 26911
rect 13964 26880 14197 26908
rect 13964 26868 13970 26880
rect 14185 26877 14197 26880
rect 14231 26877 14243 26911
rect 14461 26911 14519 26917
rect 14461 26908 14473 26911
rect 14185 26871 14243 26877
rect 14292 26880 14473 26908
rect 12492 26744 13124 26772
rect 12492 26732 12498 26744
rect 13170 26732 13176 26784
rect 13228 26732 13234 26784
rect 14182 26732 14188 26784
rect 14240 26772 14246 26784
rect 14292 26772 14320 26880
rect 14461 26877 14473 26880
rect 14507 26877 14519 26911
rect 14461 26871 14519 26877
rect 16669 26911 16727 26917
rect 16669 26877 16681 26911
rect 16715 26877 16727 26911
rect 16669 26871 16727 26877
rect 16684 26840 16712 26871
rect 20070 26868 20076 26920
rect 20128 26908 20134 26920
rect 20622 26908 20628 26920
rect 20128 26880 20628 26908
rect 20128 26868 20134 26880
rect 20622 26868 20628 26880
rect 20680 26908 20686 26920
rect 22373 26911 22431 26917
rect 22373 26908 22385 26911
rect 20680 26880 22385 26908
rect 20680 26868 20686 26880
rect 22373 26877 22385 26880
rect 22419 26877 22431 26911
rect 22373 26871 22431 26877
rect 16592 26812 16712 26840
rect 14240 26744 14320 26772
rect 14240 26732 14246 26744
rect 14458 26732 14464 26784
rect 14516 26772 14522 26784
rect 14734 26772 14740 26784
rect 14516 26744 14740 26772
rect 14516 26732 14522 26744
rect 14734 26732 14740 26744
rect 14792 26772 14798 26784
rect 16592 26772 16620 26812
rect 19242 26800 19248 26852
rect 19300 26840 19306 26852
rect 19300 26812 22416 26840
rect 19300 26800 19306 26812
rect 14792 26744 16620 26772
rect 14792 26732 14798 26744
rect 16666 26732 16672 26784
rect 16724 26772 16730 26784
rect 17402 26772 17408 26784
rect 16724 26744 17408 26772
rect 16724 26732 16730 26744
rect 17402 26732 17408 26744
rect 17460 26732 17466 26784
rect 17678 26732 17684 26784
rect 17736 26732 17742 26784
rect 22186 26732 22192 26784
rect 22244 26732 22250 26784
rect 22388 26772 22416 26812
rect 23014 26772 23020 26784
rect 22388 26744 23020 26772
rect 23014 26732 23020 26744
rect 23072 26732 23078 26784
rect 23750 26732 23756 26784
rect 23808 26732 23814 26784
rect 24210 26732 24216 26784
rect 24268 26732 24274 26784
rect 1104 26682 24840 26704
rect 1104 26630 3917 26682
rect 3969 26630 3981 26682
rect 4033 26630 4045 26682
rect 4097 26630 4109 26682
rect 4161 26630 4173 26682
rect 4225 26630 9851 26682
rect 9903 26630 9915 26682
rect 9967 26630 9979 26682
rect 10031 26630 10043 26682
rect 10095 26630 10107 26682
rect 10159 26630 15785 26682
rect 15837 26630 15849 26682
rect 15901 26630 15913 26682
rect 15965 26630 15977 26682
rect 16029 26630 16041 26682
rect 16093 26630 21719 26682
rect 21771 26630 21783 26682
rect 21835 26630 21847 26682
rect 21899 26630 21911 26682
rect 21963 26630 21975 26682
rect 22027 26630 24840 26682
rect 1104 26608 24840 26630
rect 124 26540 1072 26568
rect 124 26512 152 26540
rect 1394 26528 1400 26580
rect 1452 26568 1458 26580
rect 1452 26540 1532 26568
rect 1452 26528 1458 26540
rect 106 26460 112 26512
rect 164 26460 170 26512
rect 1504 26432 1532 26540
rect 2130 26528 2136 26580
rect 2188 26568 2194 26580
rect 2777 26571 2835 26577
rect 2777 26568 2789 26571
rect 2188 26540 2789 26568
rect 2188 26528 2194 26540
rect 2777 26537 2789 26540
rect 2823 26537 2835 26571
rect 2777 26531 2835 26537
rect 2866 26528 2872 26580
rect 2924 26568 2930 26580
rect 2924 26540 4934 26568
rect 2924 26528 2930 26540
rect 1578 26460 1584 26512
rect 1636 26460 1642 26512
rect 4906 26500 4934 26540
rect 5442 26528 5448 26580
rect 5500 26568 5506 26580
rect 5500 26540 8248 26568
rect 5500 26528 5506 26540
rect 6454 26500 6460 26512
rect 4906 26472 6460 26500
rect 6454 26460 6460 26472
rect 6512 26500 6518 26512
rect 7190 26500 7196 26512
rect 6512 26472 7196 26500
rect 6512 26460 6518 26472
rect 7190 26460 7196 26472
rect 7248 26460 7254 26512
rect 8220 26500 8248 26540
rect 8294 26528 8300 26580
rect 8352 26528 8358 26580
rect 13078 26568 13084 26580
rect 8404 26540 13084 26568
rect 8404 26500 8432 26540
rect 13078 26528 13084 26540
rect 13136 26528 13142 26580
rect 13170 26528 13176 26580
rect 13228 26528 13234 26580
rect 13998 26528 14004 26580
rect 14056 26568 14062 26580
rect 15286 26568 15292 26580
rect 14056 26540 15292 26568
rect 14056 26528 14062 26540
rect 15286 26528 15292 26540
rect 15344 26528 15350 26580
rect 15470 26528 15476 26580
rect 15528 26568 15534 26580
rect 15838 26568 15844 26580
rect 15528 26540 15844 26568
rect 15528 26528 15534 26540
rect 15838 26528 15844 26540
rect 15896 26528 15902 26580
rect 17678 26528 17684 26580
rect 17736 26568 17742 26580
rect 17736 26540 17908 26568
rect 17736 26528 17742 26540
rect 8220 26472 8432 26500
rect 8662 26460 8668 26512
rect 8720 26500 8726 26512
rect 9214 26500 9220 26512
rect 8720 26472 9220 26500
rect 8720 26460 8726 26472
rect 9214 26460 9220 26472
rect 9272 26500 9278 26512
rect 11514 26500 11520 26512
rect 9272 26472 11520 26500
rect 9272 26460 9278 26472
rect 11514 26460 11520 26472
rect 11572 26460 11578 26512
rect 13188 26500 13216 26528
rect 14737 26503 14795 26509
rect 14737 26500 14749 26503
rect 13188 26472 14749 26500
rect 14737 26469 14749 26472
rect 14783 26469 14795 26503
rect 16574 26500 16580 26512
rect 14737 26463 14795 26469
rect 16040 26472 16580 26500
rect 1765 26435 1823 26441
rect 1765 26432 1777 26435
rect 1504 26404 1777 26432
rect 1394 26324 1400 26376
rect 1452 26324 1458 26376
rect 1596 26296 1624 26404
rect 1765 26401 1777 26404
rect 1811 26401 1823 26435
rect 1765 26395 1823 26401
rect 2774 26392 2780 26444
rect 2832 26432 2838 26444
rect 3326 26432 3332 26444
rect 2832 26404 3332 26432
rect 2832 26392 2838 26404
rect 3326 26392 3332 26404
rect 3384 26392 3390 26444
rect 4982 26392 4988 26444
rect 5040 26432 5046 26444
rect 5442 26432 5448 26444
rect 5040 26404 5448 26432
rect 5040 26392 5046 26404
rect 5442 26392 5448 26404
rect 5500 26392 5506 26444
rect 6638 26392 6644 26444
rect 6696 26432 6702 26444
rect 7285 26435 7343 26441
rect 7285 26432 7297 26435
rect 6696 26404 7297 26432
rect 6696 26392 6702 26404
rect 7285 26401 7297 26404
rect 7331 26401 7343 26435
rect 7285 26395 7343 26401
rect 12250 26392 12256 26444
rect 12308 26392 12314 26444
rect 13538 26392 13544 26444
rect 13596 26432 13602 26444
rect 14277 26435 14335 26441
rect 14277 26432 14289 26435
rect 13596 26404 14289 26432
rect 13596 26392 13602 26404
rect 14277 26401 14289 26404
rect 14323 26401 14335 26435
rect 14277 26395 14335 26401
rect 14366 26392 14372 26444
rect 14424 26432 14430 26444
rect 14424 26404 15056 26432
rect 14424 26392 14430 26404
rect 1670 26324 1676 26376
rect 1728 26364 1734 26376
rect 4249 26367 4307 26373
rect 1728 26337 2084 26364
rect 1728 26336 2035 26337
rect 1728 26324 1734 26336
rect 2023 26303 2035 26336
rect 2069 26306 2084 26337
rect 4249 26333 4261 26367
rect 4295 26364 4307 26367
rect 7559 26367 7617 26373
rect 4295 26336 4384 26364
rect 4540 26363 5396 26364
rect 4295 26333 4307 26336
rect 4249 26327 4307 26333
rect 4356 26308 4384 26336
rect 4523 26357 5396 26363
rect 4523 26323 4535 26357
rect 4569 26336 5396 26357
rect 4569 26323 4581 26336
rect 4523 26317 4581 26323
rect 2069 26303 2081 26306
rect 2023 26297 2081 26303
rect 1596 26268 1716 26296
rect 1688 26240 1716 26268
rect 4338 26256 4344 26308
rect 4396 26256 4402 26308
rect 5368 26240 5396 26336
rect 7559 26333 7571 26367
rect 7605 26364 7617 26367
rect 8018 26364 8024 26376
rect 7605 26336 8024 26364
rect 7605 26333 7617 26336
rect 7559 26327 7617 26333
rect 8018 26324 8024 26336
rect 8076 26364 8082 26376
rect 8570 26364 8576 26376
rect 8076 26336 8576 26364
rect 8076 26324 8082 26336
rect 8570 26324 8576 26336
rect 8628 26324 8634 26376
rect 11517 26367 11575 26373
rect 11517 26333 11529 26367
rect 11563 26333 11575 26367
rect 11517 26327 11575 26333
rect 11791 26367 11849 26373
rect 11791 26333 11803 26367
rect 11837 26364 11849 26367
rect 11882 26364 11888 26376
rect 11837 26336 11888 26364
rect 11837 26333 11849 26336
rect 11791 26327 11849 26333
rect 7190 26256 7196 26308
rect 7248 26296 7254 26308
rect 7742 26296 7748 26308
rect 7248 26268 7748 26296
rect 7248 26256 7254 26268
rect 7742 26256 7748 26268
rect 7800 26256 7806 26308
rect 7834 26256 7840 26308
rect 7892 26296 7898 26308
rect 9122 26296 9128 26308
rect 7892 26268 9128 26296
rect 7892 26256 7898 26268
rect 9122 26256 9128 26268
rect 9180 26256 9186 26308
rect 11532 26296 11560 26327
rect 11882 26324 11888 26336
rect 11940 26324 11946 26376
rect 12158 26324 12164 26376
rect 12216 26324 12222 26376
rect 12176 26296 12204 26324
rect 11532 26268 12204 26296
rect 12268 26296 12296 26392
rect 14093 26367 14151 26373
rect 14093 26333 14105 26367
rect 14139 26364 14151 26367
rect 14458 26364 14464 26376
rect 14139 26336 14464 26364
rect 14139 26333 14151 26336
rect 14093 26327 14151 26333
rect 14458 26324 14464 26336
rect 14516 26324 14522 26376
rect 15028 26373 15056 26404
rect 15286 26392 15292 26444
rect 15344 26392 15350 26444
rect 15470 26392 15476 26444
rect 15528 26432 15534 26444
rect 16040 26441 16068 26472
rect 16574 26460 16580 26472
rect 16632 26460 16638 26512
rect 16025 26435 16083 26441
rect 16025 26432 16037 26435
rect 15528 26404 16037 26432
rect 15528 26392 15534 26404
rect 16025 26401 16037 26404
rect 16071 26401 16083 26435
rect 16025 26395 16083 26401
rect 16114 26392 16120 26444
rect 16172 26432 16178 26444
rect 16209 26435 16267 26441
rect 16209 26432 16221 26435
rect 16172 26404 16221 26432
rect 16172 26392 16178 26404
rect 16209 26401 16221 26404
rect 16255 26432 16267 26435
rect 16298 26432 16304 26444
rect 16255 26404 16304 26432
rect 16255 26401 16267 26404
rect 16209 26395 16267 26401
rect 16298 26392 16304 26404
rect 16356 26392 16362 26444
rect 16666 26392 16672 26444
rect 16724 26392 16730 26444
rect 16758 26392 16764 26444
rect 16816 26432 16822 26444
rect 16945 26435 17003 26441
rect 16945 26432 16957 26435
rect 16816 26404 16957 26432
rect 16816 26392 16822 26404
rect 16945 26401 16957 26404
rect 16991 26401 17003 26435
rect 16945 26395 17003 26401
rect 17221 26435 17279 26441
rect 17221 26401 17233 26435
rect 17267 26432 17279 26435
rect 17880 26432 17908 26540
rect 21358 26528 21364 26580
rect 21416 26528 21422 26580
rect 21468 26540 22140 26568
rect 18049 26503 18107 26509
rect 18049 26469 18061 26503
rect 18095 26469 18107 26503
rect 18049 26463 18107 26469
rect 17267 26404 17908 26432
rect 18064 26432 18092 26463
rect 18064 26404 18460 26432
rect 17267 26401 17279 26404
rect 17221 26395 17279 26401
rect 15013 26367 15071 26373
rect 15013 26333 15025 26367
rect 15059 26333 15071 26367
rect 15013 26327 15071 26333
rect 15102 26324 15108 26376
rect 15160 26373 15166 26376
rect 15160 26367 15188 26373
rect 15176 26333 15188 26367
rect 15160 26327 15188 26333
rect 15160 26324 15166 26327
rect 17034 26324 17040 26376
rect 17092 26373 17098 26376
rect 17092 26367 17120 26373
rect 17108 26333 17120 26367
rect 17092 26327 17120 26333
rect 17092 26324 17098 26327
rect 17862 26324 17868 26376
rect 17920 26364 17926 26376
rect 18432 26373 18460 26404
rect 21082 26392 21088 26444
rect 21140 26432 21146 26444
rect 21468 26441 21496 26540
rect 21453 26435 21511 26441
rect 21453 26432 21465 26435
rect 21140 26404 21465 26432
rect 21140 26392 21146 26404
rect 21453 26401 21465 26404
rect 21499 26401 21511 26435
rect 22112 26432 22140 26540
rect 22278 26528 22284 26580
rect 22336 26568 22342 26580
rect 22465 26571 22523 26577
rect 22465 26568 22477 26571
rect 22336 26540 22477 26568
rect 22336 26528 22342 26540
rect 22465 26537 22477 26540
rect 22511 26537 22523 26571
rect 22465 26531 22523 26537
rect 22462 26432 22468 26444
rect 22112 26404 22468 26432
rect 21453 26395 21511 26401
rect 22462 26392 22468 26404
rect 22520 26432 22526 26444
rect 22833 26435 22891 26441
rect 22833 26432 22845 26435
rect 22520 26404 22845 26432
rect 22520 26392 22526 26404
rect 22833 26401 22845 26404
rect 22879 26401 22891 26435
rect 22833 26395 22891 26401
rect 18233 26367 18291 26373
rect 18233 26364 18245 26367
rect 17920 26336 18245 26364
rect 17920 26324 17926 26336
rect 18233 26333 18245 26336
rect 18279 26333 18291 26367
rect 18233 26327 18291 26333
rect 18417 26367 18475 26373
rect 18417 26333 18429 26367
rect 18463 26333 18475 26367
rect 18417 26327 18475 26333
rect 19981 26367 20039 26373
rect 19981 26333 19993 26367
rect 20027 26364 20039 26367
rect 20070 26364 20076 26376
rect 20027 26336 20076 26364
rect 20027 26333 20039 26336
rect 19981 26327 20039 26333
rect 20070 26324 20076 26336
rect 20128 26324 20134 26376
rect 21695 26367 21753 26373
rect 21695 26364 21707 26367
rect 21560 26336 21707 26364
rect 20254 26305 20260 26308
rect 15933 26299 15991 26305
rect 12268 26268 14320 26296
rect 1670 26188 1676 26240
rect 1728 26188 1734 26240
rect 4522 26188 4528 26240
rect 4580 26228 4586 26240
rect 5261 26231 5319 26237
rect 5261 26228 5273 26231
rect 4580 26200 5273 26228
rect 4580 26188 4586 26200
rect 5261 26197 5273 26200
rect 5307 26197 5319 26231
rect 5261 26191 5319 26197
rect 5350 26188 5356 26240
rect 5408 26188 5414 26240
rect 6270 26188 6276 26240
rect 6328 26228 6334 26240
rect 12434 26228 12440 26240
rect 6328 26200 12440 26228
rect 6328 26188 6334 26200
rect 12434 26188 12440 26200
rect 12492 26188 12498 26240
rect 12526 26188 12532 26240
rect 12584 26188 12590 26240
rect 14292 26228 14320 26268
rect 15933 26265 15945 26299
rect 15979 26296 15991 26299
rect 20226 26299 20260 26305
rect 20226 26296 20238 26299
rect 15979 26268 16252 26296
rect 15979 26265 15991 26268
rect 15933 26259 15991 26265
rect 15102 26228 15108 26240
rect 14292 26200 15108 26228
rect 15102 26188 15108 26200
rect 15160 26188 15166 26240
rect 16224 26228 16252 26268
rect 17696 26268 20238 26296
rect 17696 26228 17724 26268
rect 20226 26265 20238 26268
rect 20226 26259 20260 26265
rect 20254 26256 20260 26259
rect 20312 26256 20318 26308
rect 21358 26256 21364 26308
rect 21416 26296 21422 26308
rect 21560 26296 21588 26336
rect 21695 26333 21707 26336
rect 21741 26333 21753 26367
rect 23106 26364 23112 26376
rect 23067 26336 23112 26364
rect 21695 26327 21753 26333
rect 23106 26324 23112 26336
rect 23164 26324 23170 26376
rect 21416 26268 21588 26296
rect 21416 26256 21422 26268
rect 16224 26200 17724 26228
rect 18506 26188 18512 26240
rect 18564 26188 18570 26240
rect 23842 26188 23848 26240
rect 23900 26188 23906 26240
rect 1104 26138 25000 26160
rect 1104 26086 6884 26138
rect 6936 26086 6948 26138
rect 7000 26086 7012 26138
rect 7064 26086 7076 26138
rect 7128 26086 7140 26138
rect 7192 26086 12818 26138
rect 12870 26086 12882 26138
rect 12934 26086 12946 26138
rect 12998 26086 13010 26138
rect 13062 26086 13074 26138
rect 13126 26086 18752 26138
rect 18804 26086 18816 26138
rect 18868 26086 18880 26138
rect 18932 26086 18944 26138
rect 18996 26086 19008 26138
rect 19060 26086 24686 26138
rect 24738 26086 24750 26138
rect 24802 26086 24814 26138
rect 24866 26086 24878 26138
rect 24930 26086 24942 26138
rect 24994 26086 25000 26138
rect 1104 26064 25000 26086
rect 934 25984 940 26036
rect 992 26024 998 26036
rect 992 25996 1992 26024
rect 992 25984 998 25996
rect 842 25916 848 25968
rect 900 25956 906 25968
rect 900 25928 1900 25956
rect 900 25916 906 25928
rect 1397 25891 1455 25897
rect 1397 25857 1409 25891
rect 1443 25888 1455 25891
rect 1486 25888 1492 25900
rect 1443 25860 1492 25888
rect 1443 25857 1455 25860
rect 1397 25851 1455 25857
rect 1486 25848 1492 25860
rect 1544 25848 1550 25900
rect 1872 25897 1900 25928
rect 1964 25897 1992 25996
rect 2130 25984 2136 26036
rect 2188 25984 2194 26036
rect 2682 25984 2688 26036
rect 2740 25984 2746 26036
rect 5445 26027 5503 26033
rect 3804 25996 4934 26024
rect 3804 25900 3832 25996
rect 4062 25916 4068 25968
rect 4120 25916 4126 25968
rect 4157 25959 4215 25965
rect 4157 25925 4169 25959
rect 4203 25956 4215 25959
rect 4246 25956 4252 25968
rect 4203 25928 4252 25956
rect 4203 25925 4215 25928
rect 4157 25919 4215 25925
rect 4246 25916 4252 25928
rect 4304 25916 4310 25968
rect 4522 25916 4528 25968
rect 4580 25916 4586 25968
rect 4906 25965 4934 25996
rect 5445 25993 5457 26027
rect 5491 25993 5503 26027
rect 5445 25987 5503 25993
rect 4893 25959 4951 25965
rect 4893 25925 4905 25959
rect 4939 25925 4951 25959
rect 4893 25919 4951 25925
rect 5261 25959 5319 25965
rect 5261 25925 5273 25959
rect 5307 25956 5319 25959
rect 5460 25956 5488 25987
rect 6546 25984 6552 26036
rect 6604 26024 6610 26036
rect 7650 26024 7656 26036
rect 6604 25996 7656 26024
rect 6604 25984 6610 25996
rect 7650 25984 7656 25996
rect 7708 25984 7714 26036
rect 8110 25984 8116 26036
rect 8168 26024 8174 26036
rect 9490 26024 9496 26036
rect 8168 25996 9496 26024
rect 8168 25984 8174 25996
rect 9490 25984 9496 25996
rect 9548 25984 9554 26036
rect 9766 25984 9772 26036
rect 9824 26024 9830 26036
rect 10686 26024 10692 26036
rect 9824 25996 10692 26024
rect 9824 25984 9830 25996
rect 10686 25984 10692 25996
rect 10744 25984 10750 26036
rect 11514 25984 11520 26036
rect 11572 26024 11578 26036
rect 14826 26024 14832 26036
rect 11572 25996 14832 26024
rect 11572 25984 11578 25996
rect 14826 25984 14832 25996
rect 14884 25984 14890 26036
rect 16209 26027 16267 26033
rect 16209 25993 16221 26027
rect 16255 26024 16267 26027
rect 16666 26024 16672 26036
rect 16255 25996 16672 26024
rect 16255 25993 16267 25996
rect 16209 25987 16267 25993
rect 16666 25984 16672 25996
rect 16724 25984 16730 26036
rect 18969 26027 19027 26033
rect 18969 25993 18981 26027
rect 19015 26024 19027 26027
rect 19015 25996 19932 26024
rect 19015 25993 19027 25996
rect 18969 25987 19027 25993
rect 15194 25956 15200 25968
rect 5307 25928 5396 25956
rect 5460 25928 15200 25956
rect 5307 25925 5319 25928
rect 5261 25919 5319 25925
rect 1857 25891 1915 25897
rect 1857 25857 1869 25891
rect 1903 25857 1915 25891
rect 1857 25851 1915 25857
rect 1949 25891 2007 25897
rect 1949 25857 1961 25891
rect 1995 25857 2007 25891
rect 1949 25851 2007 25857
rect 2222 25848 2228 25900
rect 2280 25848 2286 25900
rect 2498 25848 2504 25900
rect 2556 25848 2562 25900
rect 3786 25848 3792 25900
rect 3844 25848 3850 25900
rect 4080 25888 4108 25916
rect 4433 25891 4491 25897
rect 4433 25888 4445 25891
rect 4080 25860 4445 25888
rect 4433 25857 4445 25860
rect 4479 25857 4491 25891
rect 4433 25851 4491 25857
rect 5074 25848 5080 25900
rect 5132 25888 5138 25900
rect 5368 25888 5396 25928
rect 15194 25916 15200 25928
rect 15252 25916 15258 25968
rect 15378 25916 15384 25968
rect 15436 25916 15442 25968
rect 17862 25965 17868 25968
rect 17856 25956 17868 25965
rect 17823 25928 17868 25956
rect 17856 25919 17868 25928
rect 17862 25916 17868 25919
rect 17920 25916 17926 25968
rect 18506 25916 18512 25968
rect 18564 25956 18570 25968
rect 18564 25928 19196 25956
rect 18564 25916 18570 25928
rect 5442 25888 5448 25900
rect 5132 25860 5304 25888
rect 5368 25860 5448 25888
rect 5132 25848 5138 25860
rect 4798 25780 4804 25832
rect 4856 25780 4862 25832
rect 5276 25820 5304 25860
rect 5442 25848 5448 25860
rect 5500 25848 5506 25900
rect 7835 25891 7893 25897
rect 7835 25857 7847 25891
rect 7881 25888 7893 25891
rect 10134 25888 10140 25900
rect 7881 25860 9168 25888
rect 7881 25857 7893 25860
rect 7835 25851 7893 25857
rect 5626 25820 5632 25832
rect 5276 25792 5632 25820
rect 5626 25780 5632 25792
rect 5684 25780 5690 25832
rect 7561 25823 7619 25829
rect 7561 25789 7573 25823
rect 7607 25789 7619 25823
rect 7561 25783 7619 25789
rect 2406 25712 2412 25764
rect 2464 25712 2470 25764
rect 1578 25644 1584 25696
rect 1636 25644 1642 25696
rect 1673 25687 1731 25693
rect 1673 25653 1685 25687
rect 1719 25684 1731 25687
rect 2222 25684 2228 25696
rect 1719 25656 2228 25684
rect 1719 25653 1731 25656
rect 1673 25647 1731 25653
rect 2222 25644 2228 25656
rect 2280 25644 2286 25696
rect 2314 25644 2320 25696
rect 2372 25684 2378 25696
rect 2866 25684 2872 25696
rect 2372 25656 2872 25684
rect 2372 25644 2378 25656
rect 2866 25644 2872 25656
rect 2924 25644 2930 25696
rect 6086 25644 6092 25696
rect 6144 25684 6150 25696
rect 6733 25687 6791 25693
rect 6733 25684 6745 25687
rect 6144 25656 6745 25684
rect 6144 25644 6150 25656
rect 6733 25653 6745 25656
rect 6779 25653 6791 25687
rect 7576 25684 7604 25783
rect 7834 25684 7840 25696
rect 7576 25656 7840 25684
rect 6733 25647 6791 25653
rect 7834 25644 7840 25656
rect 7892 25644 7898 25696
rect 8018 25644 8024 25696
rect 8076 25684 8082 25696
rect 8573 25687 8631 25693
rect 8573 25684 8585 25687
rect 8076 25656 8585 25684
rect 8076 25644 8082 25656
rect 8573 25653 8585 25656
rect 8619 25653 8631 25687
rect 9140 25684 9168 25860
rect 9968 25860 10140 25888
rect 9214 25780 9220 25832
rect 9272 25820 9278 25832
rect 9968 25829 9996 25860
rect 10134 25848 10140 25860
rect 10192 25848 10198 25900
rect 10227 25891 10285 25897
rect 10227 25857 10239 25891
rect 10273 25888 10285 25891
rect 11974 25888 11980 25900
rect 10273 25860 11980 25888
rect 10273 25857 10285 25860
rect 10227 25851 10285 25857
rect 11974 25848 11980 25860
rect 12032 25848 12038 25900
rect 15396 25888 15424 25916
rect 19168 25897 19196 25928
rect 19904 25897 19932 25996
rect 20254 25984 20260 26036
rect 20312 25984 20318 26036
rect 22830 25984 22836 26036
rect 22888 25984 22894 26036
rect 23842 25984 23848 26036
rect 23900 25984 23906 26036
rect 15471 25891 15529 25897
rect 15471 25888 15483 25891
rect 15396 25860 15483 25888
rect 15471 25857 15483 25860
rect 15517 25857 15529 25891
rect 19061 25891 19119 25897
rect 19061 25888 19073 25891
rect 15471 25851 15529 25857
rect 18616 25860 19073 25888
rect 9953 25823 10011 25829
rect 9953 25820 9965 25823
rect 9272 25792 9965 25820
rect 9272 25780 9278 25792
rect 9953 25789 9965 25792
rect 9999 25789 10011 25823
rect 9953 25783 10011 25789
rect 14734 25780 14740 25832
rect 14792 25820 14798 25832
rect 15197 25823 15255 25829
rect 15197 25820 15209 25823
rect 14792 25792 15209 25820
rect 14792 25780 14798 25792
rect 15197 25789 15209 25792
rect 15243 25789 15255 25823
rect 15197 25783 15255 25789
rect 17589 25823 17647 25829
rect 17589 25789 17601 25823
rect 17635 25789 17647 25823
rect 17589 25783 17647 25789
rect 10796 25724 11928 25752
rect 10796 25684 10824 25724
rect 11900 25696 11928 25724
rect 9140 25656 10824 25684
rect 8573 25647 8631 25653
rect 10870 25644 10876 25696
rect 10928 25684 10934 25696
rect 10965 25687 11023 25693
rect 10965 25684 10977 25687
rect 10928 25656 10977 25684
rect 10928 25644 10934 25656
rect 10965 25653 10977 25656
rect 11011 25653 11023 25687
rect 10965 25647 11023 25653
rect 11882 25644 11888 25696
rect 11940 25644 11946 25696
rect 13262 25644 13268 25696
rect 13320 25684 13326 25696
rect 15654 25684 15660 25696
rect 13320 25656 15660 25684
rect 13320 25644 13326 25656
rect 15654 25644 15660 25656
rect 15712 25644 15718 25696
rect 17604 25684 17632 25783
rect 18616 25696 18644 25860
rect 19061 25857 19073 25860
rect 19107 25857 19119 25891
rect 19061 25851 19119 25857
rect 19153 25891 19211 25897
rect 19153 25857 19165 25891
rect 19199 25857 19211 25891
rect 19429 25891 19487 25897
rect 19429 25888 19441 25891
rect 19153 25851 19211 25857
rect 19260 25860 19441 25888
rect 19076 25820 19104 25851
rect 19260 25820 19288 25860
rect 19429 25857 19441 25860
rect 19475 25857 19487 25891
rect 19429 25851 19487 25857
rect 19613 25891 19671 25897
rect 19613 25857 19625 25891
rect 19659 25888 19671 25891
rect 19889 25891 19947 25897
rect 19659 25860 19748 25888
rect 19659 25857 19671 25860
rect 19613 25851 19671 25857
rect 19076 25792 19288 25820
rect 19337 25823 19395 25829
rect 19337 25789 19349 25823
rect 19383 25820 19395 25823
rect 19521 25823 19579 25829
rect 19521 25820 19533 25823
rect 19383 25792 19533 25820
rect 19383 25789 19395 25792
rect 19337 25783 19395 25789
rect 19521 25789 19533 25792
rect 19567 25789 19579 25823
rect 19521 25783 19579 25789
rect 19720 25761 19748 25860
rect 19889 25857 19901 25891
rect 19935 25857 19947 25891
rect 20272 25888 20300 25984
rect 20625 25891 20683 25897
rect 20625 25888 20637 25891
rect 20272 25860 20637 25888
rect 19889 25851 19947 25857
rect 20625 25857 20637 25860
rect 20671 25857 20683 25891
rect 20625 25851 20683 25857
rect 21085 25891 21143 25897
rect 21085 25857 21097 25891
rect 21131 25857 21143 25891
rect 21085 25851 21143 25857
rect 21821 25891 21879 25897
rect 21821 25857 21833 25891
rect 21867 25888 21879 25891
rect 22278 25888 22284 25900
rect 21867 25860 22284 25888
rect 21867 25857 21879 25860
rect 21821 25851 21879 25857
rect 21100 25820 21128 25851
rect 22278 25848 22284 25860
rect 22336 25848 22342 25900
rect 22848 25888 22876 25984
rect 23860 25956 23888 25984
rect 23216 25928 23888 25956
rect 23216 25897 23244 25928
rect 22925 25891 22983 25897
rect 22925 25888 22937 25891
rect 22848 25860 22937 25888
rect 22925 25857 22937 25860
rect 22971 25857 22983 25891
rect 22925 25851 22983 25857
rect 23201 25891 23259 25897
rect 23201 25857 23213 25891
rect 23247 25857 23259 25891
rect 23201 25851 23259 25857
rect 23382 25848 23388 25900
rect 23440 25848 23446 25900
rect 23661 25891 23719 25897
rect 23661 25857 23673 25891
rect 23707 25888 23719 25891
rect 23860 25888 23888 25928
rect 23934 25916 23940 25968
rect 23992 25956 23998 25968
rect 24121 25959 24179 25965
rect 24121 25956 24133 25959
rect 23992 25928 24133 25956
rect 23992 25916 23998 25928
rect 24121 25925 24133 25928
rect 24167 25925 24179 25959
rect 24121 25919 24179 25925
rect 23707 25860 23888 25888
rect 23707 25857 23719 25860
rect 23661 25851 23719 25857
rect 20456 25792 21128 25820
rect 22097 25823 22155 25829
rect 20456 25761 20484 25792
rect 22097 25789 22109 25823
rect 22143 25820 22155 25823
rect 22186 25820 22192 25832
rect 22143 25792 22192 25820
rect 22143 25789 22155 25792
rect 22097 25783 22155 25789
rect 22186 25780 22192 25792
rect 22244 25780 22250 25832
rect 23293 25823 23351 25829
rect 23293 25789 23305 25823
rect 23339 25820 23351 25823
rect 23937 25823 23995 25829
rect 23937 25820 23949 25823
rect 23339 25792 23949 25820
rect 23339 25789 23351 25792
rect 23293 25783 23351 25789
rect 23937 25789 23949 25792
rect 23983 25789 23995 25823
rect 23937 25783 23995 25789
rect 25130 25780 25136 25832
rect 25188 25820 25194 25832
rect 25314 25820 25320 25832
rect 25188 25792 25320 25820
rect 25188 25780 25194 25792
rect 25314 25780 25320 25792
rect 25372 25780 25378 25832
rect 19705 25755 19763 25761
rect 19705 25721 19717 25755
rect 19751 25721 19763 25755
rect 19705 25715 19763 25721
rect 20441 25755 20499 25761
rect 20441 25721 20453 25755
rect 20487 25721 20499 25755
rect 20441 25715 20499 25721
rect 23017 25755 23075 25761
rect 23017 25721 23029 25755
rect 23063 25752 23075 25755
rect 23753 25755 23811 25761
rect 23753 25752 23765 25755
rect 23063 25724 23765 25752
rect 23063 25721 23075 25724
rect 23017 25715 23075 25721
rect 23753 25721 23765 25724
rect 23799 25721 23811 25755
rect 23753 25715 23811 25721
rect 17954 25684 17960 25696
rect 17604 25656 17960 25684
rect 17954 25644 17960 25656
rect 18012 25684 18018 25696
rect 18506 25684 18512 25696
rect 18012 25656 18512 25684
rect 18012 25644 18018 25656
rect 18506 25644 18512 25656
rect 18564 25644 18570 25696
rect 18598 25644 18604 25696
rect 18656 25644 18662 25696
rect 19242 25644 19248 25696
rect 19300 25644 19306 25696
rect 21177 25687 21235 25693
rect 21177 25653 21189 25687
rect 21223 25684 21235 25687
rect 21913 25687 21971 25693
rect 21913 25684 21925 25687
rect 21223 25656 21925 25684
rect 21223 25653 21235 25656
rect 21177 25647 21235 25653
rect 21913 25653 21925 25656
rect 21959 25653 21971 25687
rect 21913 25647 21971 25653
rect 22005 25687 22063 25693
rect 22005 25653 22017 25687
rect 22051 25684 22063 25687
rect 22554 25684 22560 25696
rect 22051 25656 22560 25684
rect 22051 25653 22063 25656
rect 22005 25647 22063 25653
rect 22554 25644 22560 25656
rect 22612 25644 22618 25696
rect 23842 25644 23848 25696
rect 23900 25644 23906 25696
rect 24394 25644 24400 25696
rect 24452 25644 24458 25696
rect 1104 25594 24840 25616
rect 1104 25542 3917 25594
rect 3969 25542 3981 25594
rect 4033 25542 4045 25594
rect 4097 25542 4109 25594
rect 4161 25542 4173 25594
rect 4225 25542 9851 25594
rect 9903 25542 9915 25594
rect 9967 25542 9979 25594
rect 10031 25542 10043 25594
rect 10095 25542 10107 25594
rect 10159 25542 15785 25594
rect 15837 25542 15849 25594
rect 15901 25542 15913 25594
rect 15965 25542 15977 25594
rect 16029 25542 16041 25594
rect 16093 25542 21719 25594
rect 21771 25542 21783 25594
rect 21835 25542 21847 25594
rect 21899 25542 21911 25594
rect 21963 25542 21975 25594
rect 22027 25542 24840 25594
rect 1104 25520 24840 25542
rect 1578 25440 1584 25492
rect 1636 25480 1642 25492
rect 6270 25480 6276 25492
rect 1636 25452 6276 25480
rect 1636 25440 1642 25452
rect 6270 25440 6276 25452
rect 6328 25440 6334 25492
rect 7466 25440 7472 25492
rect 7524 25480 7530 25492
rect 11517 25483 11575 25489
rect 7524 25452 11284 25480
rect 7524 25440 7530 25452
rect 2130 25372 2136 25424
rect 2188 25372 2194 25424
rect 2314 25372 2320 25424
rect 2372 25372 2378 25424
rect 5721 25415 5779 25421
rect 5721 25381 5733 25415
rect 5767 25381 5779 25415
rect 5721 25375 5779 25381
rect 9876 25384 10456 25412
rect 1397 25279 1455 25285
rect 1397 25245 1409 25279
rect 1443 25245 1455 25279
rect 1397 25239 1455 25245
rect 934 25100 940 25152
rect 992 25140 998 25152
rect 1412 25140 1440 25239
rect 1670 25236 1676 25288
rect 1728 25236 1734 25288
rect 1946 25236 1952 25288
rect 2004 25236 2010 25288
rect 2332 25285 2360 25372
rect 3234 25304 3240 25356
rect 3292 25344 3298 25356
rect 3602 25344 3608 25356
rect 3292 25316 3608 25344
rect 3292 25304 3298 25316
rect 3602 25304 3608 25316
rect 3660 25304 3666 25356
rect 4338 25304 4344 25356
rect 4396 25344 4402 25356
rect 4709 25347 4767 25353
rect 4709 25344 4721 25347
rect 4396 25316 4721 25344
rect 4396 25304 4402 25316
rect 4709 25313 4721 25316
rect 4755 25313 4767 25347
rect 5736 25344 5764 25375
rect 9876 25353 9904 25384
rect 10428 25356 10456 25384
rect 9861 25347 9919 25353
rect 5736 25316 6118 25344
rect 4709 25307 4767 25313
rect 9861 25313 9873 25347
rect 9907 25313 9919 25347
rect 9861 25307 9919 25313
rect 10042 25304 10048 25356
rect 10100 25344 10106 25356
rect 10321 25347 10379 25353
rect 10321 25344 10333 25347
rect 10100 25316 10333 25344
rect 10100 25304 10106 25316
rect 10321 25313 10333 25316
rect 10367 25313 10379 25347
rect 10321 25307 10379 25313
rect 10410 25304 10416 25356
rect 10468 25304 10474 25356
rect 10686 25304 10692 25356
rect 10744 25353 10750 25356
rect 10744 25347 10772 25353
rect 10760 25313 10772 25347
rect 10744 25307 10772 25313
rect 10744 25304 10750 25307
rect 10870 25304 10876 25356
rect 10928 25304 10934 25356
rect 11256 25344 11284 25452
rect 11517 25449 11529 25483
rect 11563 25480 11575 25483
rect 12066 25480 12072 25492
rect 11563 25452 12072 25480
rect 11563 25449 11575 25452
rect 11517 25443 11575 25449
rect 12066 25440 12072 25452
rect 12124 25440 12130 25492
rect 15194 25440 15200 25492
rect 15252 25480 15258 25492
rect 15252 25452 18552 25480
rect 15252 25440 15258 25452
rect 12526 25372 12532 25424
rect 12584 25372 12590 25424
rect 18524 25412 18552 25452
rect 18598 25440 18604 25492
rect 18656 25440 18662 25492
rect 19242 25440 19248 25492
rect 19300 25480 19306 25492
rect 19300 25452 22094 25480
rect 19300 25440 19306 25452
rect 19886 25412 19892 25424
rect 13464 25384 14872 25412
rect 18524 25384 19892 25412
rect 11606 25344 11612 25356
rect 11256 25316 11612 25344
rect 11606 25304 11612 25316
rect 11664 25344 11670 25356
rect 11885 25347 11943 25353
rect 11885 25344 11897 25347
rect 11664 25316 11897 25344
rect 11664 25304 11670 25316
rect 11885 25313 11897 25316
rect 11931 25313 11943 25347
rect 12805 25347 12863 25353
rect 12805 25344 12817 25347
rect 11885 25307 11943 25313
rect 12268 25316 12817 25344
rect 12268 25288 12296 25316
rect 12805 25313 12817 25316
rect 12851 25344 12863 25347
rect 13464 25344 13492 25384
rect 12851 25316 13492 25344
rect 12851 25313 12863 25316
rect 12805 25307 12863 25313
rect 13722 25304 13728 25356
rect 13780 25304 13786 25356
rect 14093 25347 14151 25353
rect 14093 25313 14105 25347
rect 14139 25344 14151 25347
rect 14458 25344 14464 25356
rect 14139 25316 14464 25344
rect 14139 25313 14151 25316
rect 14093 25307 14151 25313
rect 14458 25304 14464 25316
rect 14516 25304 14522 25356
rect 14642 25304 14648 25356
rect 14700 25344 14706 25356
rect 14737 25347 14795 25353
rect 14737 25344 14749 25347
rect 14700 25316 14749 25344
rect 14700 25304 14706 25316
rect 14737 25313 14749 25316
rect 14783 25313 14795 25347
rect 14844 25344 14872 25384
rect 19886 25372 19892 25384
rect 19944 25372 19950 25424
rect 20162 25372 20168 25424
rect 20220 25412 20226 25424
rect 21082 25412 21088 25424
rect 20220 25384 21088 25412
rect 20220 25372 20226 25384
rect 21082 25372 21088 25384
rect 21140 25372 21146 25424
rect 22066 25412 22094 25452
rect 23382 25440 23388 25492
rect 23440 25480 23446 25492
rect 23477 25483 23535 25489
rect 23477 25480 23489 25483
rect 23440 25452 23489 25480
rect 23440 25440 23446 25452
rect 23477 25449 23489 25452
rect 23523 25449 23535 25483
rect 23477 25443 23535 25449
rect 25866 25440 25872 25492
rect 25924 25440 25930 25492
rect 25884 25412 25912 25440
rect 22066 25384 25912 25412
rect 15013 25347 15071 25353
rect 15013 25344 15025 25347
rect 14844 25316 15025 25344
rect 14737 25307 14795 25313
rect 15013 25313 15025 25316
rect 15059 25313 15071 25347
rect 15013 25307 15071 25313
rect 15102 25304 15108 25356
rect 15160 25353 15166 25356
rect 15160 25347 15188 25353
rect 15176 25313 15188 25347
rect 15160 25307 15188 25313
rect 15160 25304 15166 25307
rect 15286 25304 15292 25356
rect 15344 25304 15350 25356
rect 16298 25304 16304 25356
rect 16356 25344 16362 25356
rect 16574 25344 16580 25356
rect 16356 25316 16580 25344
rect 16356 25304 16362 25316
rect 16574 25304 16580 25316
rect 16632 25304 16638 25356
rect 23474 25304 23480 25356
rect 23532 25344 23538 25356
rect 23934 25344 23940 25356
rect 23532 25316 23940 25344
rect 23532 25304 23538 25316
rect 23934 25304 23940 25316
rect 23992 25304 23998 25356
rect 2317 25279 2375 25285
rect 2317 25245 2329 25279
rect 2363 25245 2375 25279
rect 2317 25239 2375 25245
rect 2591 25279 2649 25285
rect 2591 25245 2603 25279
rect 2637 25276 2649 25279
rect 2682 25276 2688 25288
rect 2637 25248 2688 25276
rect 2637 25245 2649 25248
rect 2591 25239 2649 25245
rect 2682 25236 2688 25248
rect 2740 25236 2746 25288
rect 3050 25236 3056 25288
rect 3108 25276 3114 25288
rect 4951 25279 5009 25285
rect 4951 25276 4963 25279
rect 3108 25272 4660 25276
rect 4816 25272 4963 25276
rect 3108 25248 4963 25272
rect 3108 25236 3114 25248
rect 4632 25244 4844 25248
rect 4951 25245 4963 25248
rect 4997 25276 5009 25279
rect 4997 25248 5212 25276
rect 4997 25245 5009 25248
rect 4951 25239 5009 25245
rect 5184 25220 5212 25248
rect 5626 25236 5632 25288
rect 5684 25276 5690 25288
rect 9677 25279 9735 25285
rect 9677 25276 9689 25279
rect 5684 25248 9689 25276
rect 5684 25236 5690 25248
rect 9677 25245 9689 25248
rect 9723 25245 9735 25279
rect 9677 25239 9735 25245
rect 1872 25180 4936 25208
rect 992 25112 1440 25140
rect 992 25100 998 25112
rect 1578 25100 1584 25152
rect 1636 25100 1642 25152
rect 1872 25149 1900 25180
rect 4908 25152 4936 25180
rect 5166 25168 5172 25220
rect 5224 25168 5230 25220
rect 6086 25168 6092 25220
rect 6144 25208 6150 25220
rect 6549 25211 6607 25217
rect 6549 25208 6561 25211
rect 6144 25180 6561 25208
rect 6144 25168 6150 25180
rect 6549 25177 6561 25180
rect 6595 25177 6607 25211
rect 6549 25171 6607 25177
rect 6641 25211 6699 25217
rect 6641 25177 6653 25211
rect 6687 25208 6699 25211
rect 7009 25211 7067 25217
rect 6687 25180 6868 25208
rect 6687 25177 6699 25180
rect 6641 25171 6699 25177
rect 1857 25143 1915 25149
rect 1857 25109 1869 25143
rect 1903 25109 1915 25143
rect 1857 25103 1915 25109
rect 3326 25100 3332 25152
rect 3384 25100 3390 25152
rect 4890 25100 4896 25152
rect 4948 25100 4954 25152
rect 6270 25100 6276 25152
rect 6328 25140 6334 25152
rect 6454 25140 6460 25152
rect 6328 25112 6460 25140
rect 6328 25100 6334 25112
rect 6454 25100 6460 25112
rect 6512 25100 6518 25152
rect 6840 25140 6868 25180
rect 7009 25177 7021 25211
rect 7055 25208 7067 25211
rect 7190 25208 7196 25220
rect 7055 25180 7196 25208
rect 7055 25177 7067 25180
rect 7009 25171 7067 25177
rect 7190 25168 7196 25180
rect 7248 25168 7254 25220
rect 7374 25168 7380 25220
rect 7432 25168 7438 25220
rect 7282 25140 7288 25152
rect 6840 25112 7288 25140
rect 7282 25100 7288 25112
rect 7340 25100 7346 25152
rect 7558 25100 7564 25152
rect 7616 25100 7622 25152
rect 9692 25140 9720 25239
rect 10594 25236 10600 25288
rect 10652 25236 10658 25288
rect 12069 25279 12127 25285
rect 12069 25245 12081 25279
rect 12115 25245 12127 25279
rect 12069 25239 12127 25245
rect 11974 25140 11980 25152
rect 9692 25112 11980 25140
rect 11974 25100 11980 25112
rect 12032 25140 12038 25152
rect 12084 25140 12112 25239
rect 12250 25236 12256 25288
rect 12308 25236 12314 25288
rect 12894 25236 12900 25288
rect 12952 25285 12958 25288
rect 12952 25279 12980 25285
rect 12968 25245 12980 25279
rect 12952 25239 12980 25245
rect 12952 25236 12958 25239
rect 13078 25236 13084 25288
rect 13136 25236 13142 25288
rect 13740 25276 13768 25304
rect 14277 25279 14335 25285
rect 14277 25276 14289 25279
rect 13740 25248 14289 25276
rect 14277 25245 14289 25248
rect 14323 25245 14335 25279
rect 14277 25239 14335 25245
rect 17494 25236 17500 25288
rect 17552 25276 17558 25288
rect 17589 25279 17647 25285
rect 17589 25276 17601 25279
rect 17552 25248 17601 25276
rect 17552 25236 17558 25248
rect 17589 25245 17601 25248
rect 17635 25245 17647 25279
rect 17589 25239 17647 25245
rect 17863 25279 17921 25285
rect 17863 25245 17875 25279
rect 17909 25276 17921 25279
rect 17909 25248 18092 25276
rect 17909 25245 17921 25248
rect 17863 25239 17921 25245
rect 17954 25208 17960 25220
rect 15856 25180 17960 25208
rect 12032 25112 12112 25140
rect 12032 25100 12038 25112
rect 12434 25100 12440 25152
rect 12492 25140 12498 25152
rect 12618 25140 12624 25152
rect 12492 25112 12624 25140
rect 12492 25100 12498 25112
rect 12618 25100 12624 25112
rect 12676 25140 12682 25152
rect 12894 25140 12900 25152
rect 12676 25112 12900 25140
rect 12676 25100 12682 25112
rect 12894 25100 12900 25112
rect 12952 25100 12958 25152
rect 13725 25143 13783 25149
rect 13725 25109 13737 25143
rect 13771 25140 13783 25143
rect 15856 25140 15884 25180
rect 17954 25168 17960 25180
rect 18012 25168 18018 25220
rect 13771 25112 15884 25140
rect 13771 25109 13783 25112
rect 13725 25103 13783 25109
rect 15930 25100 15936 25152
rect 15988 25100 15994 25152
rect 16574 25100 16580 25152
rect 16632 25140 16638 25152
rect 18064 25140 18092 25248
rect 19978 25236 19984 25288
rect 20036 25276 20042 25288
rect 20257 25279 20315 25285
rect 20257 25276 20269 25279
rect 20036 25248 20269 25276
rect 20036 25236 20042 25248
rect 20257 25245 20269 25248
rect 20303 25245 20315 25279
rect 20257 25239 20315 25245
rect 20349 25279 20407 25285
rect 20349 25245 20361 25279
rect 20395 25276 20407 25279
rect 20438 25276 20444 25288
rect 20395 25248 20444 25276
rect 20395 25245 20407 25248
rect 20349 25239 20407 25245
rect 20438 25236 20444 25248
rect 20496 25236 20502 25288
rect 20533 25279 20591 25285
rect 20533 25245 20545 25279
rect 20579 25245 20591 25279
rect 20533 25239 20591 25245
rect 23661 25279 23719 25285
rect 23661 25245 23673 25279
rect 23707 25276 23719 25279
rect 23750 25276 23756 25288
rect 23707 25248 23756 25276
rect 23707 25245 23719 25248
rect 23661 25239 23719 25245
rect 20548 25208 20576 25239
rect 23750 25236 23756 25248
rect 23808 25236 23814 25288
rect 20088 25180 20576 25208
rect 20088 25149 20116 25180
rect 21174 25168 21180 25220
rect 21232 25208 21238 25220
rect 23845 25211 23903 25217
rect 23845 25208 23857 25211
rect 21232 25180 23857 25208
rect 21232 25168 21238 25180
rect 23845 25177 23857 25180
rect 23891 25177 23903 25211
rect 23845 25171 23903 25177
rect 16632 25112 18092 25140
rect 20073 25143 20131 25149
rect 16632 25100 16638 25112
rect 20073 25109 20085 25143
rect 20119 25109 20131 25143
rect 20073 25103 20131 25109
rect 20346 25100 20352 25152
rect 20404 25140 20410 25152
rect 20441 25143 20499 25149
rect 20441 25140 20453 25143
rect 20404 25112 20453 25140
rect 20404 25100 20410 25112
rect 20441 25109 20453 25112
rect 20487 25109 20499 25143
rect 20441 25103 20499 25109
rect 24118 25100 24124 25152
rect 24176 25100 24182 25152
rect 1104 25050 25000 25072
rect 290 24964 296 25016
rect 348 25004 354 25016
rect 658 25004 664 25016
rect 348 24976 664 25004
rect 348 24964 354 24976
rect 658 24964 664 24976
rect 716 24964 722 25016
rect 1104 24998 6884 25050
rect 6936 24998 6948 25050
rect 7000 24998 7012 25050
rect 7064 24998 7076 25050
rect 7128 24998 7140 25050
rect 7192 24998 12818 25050
rect 12870 24998 12882 25050
rect 12934 24998 12946 25050
rect 12998 24998 13010 25050
rect 13062 24998 13074 25050
rect 13126 24998 18752 25050
rect 18804 24998 18816 25050
rect 18868 24998 18880 25050
rect 18932 24998 18944 25050
rect 18996 24998 19008 25050
rect 19060 24998 24686 25050
rect 24738 24998 24750 25050
rect 24802 24998 24814 25050
rect 24866 24998 24878 25050
rect 24930 24998 24942 25050
rect 24994 24998 25000 25050
rect 1104 24976 25000 24998
rect 1578 24896 1584 24948
rect 1636 24936 1642 24948
rect 1854 24936 1860 24948
rect 1636 24908 1860 24936
rect 1636 24896 1642 24908
rect 1854 24896 1860 24908
rect 1912 24896 1918 24948
rect 2222 24896 2228 24948
rect 2280 24936 2286 24948
rect 3786 24936 3792 24948
rect 2280 24908 3792 24936
rect 2280 24896 2286 24908
rect 3786 24896 3792 24908
rect 3844 24936 3850 24948
rect 4525 24939 4583 24945
rect 4525 24936 4537 24939
rect 3844 24908 4537 24936
rect 3844 24896 3850 24908
rect 4525 24905 4537 24908
rect 4571 24905 4583 24939
rect 4525 24899 4583 24905
rect 7282 24896 7288 24948
rect 7340 24936 7346 24948
rect 7377 24939 7435 24945
rect 7377 24936 7389 24939
rect 7340 24908 7389 24936
rect 7340 24896 7346 24908
rect 7377 24905 7389 24908
rect 7423 24905 7435 24939
rect 9309 24939 9367 24945
rect 7377 24899 7435 24905
rect 8312 24908 9242 24936
rect 106 24828 112 24880
rect 164 24868 170 24880
rect 3050 24868 3056 24880
rect 164 24840 3056 24868
rect 164 24828 170 24840
rect 3050 24828 3056 24840
rect 3108 24828 3114 24880
rect 3418 24828 3424 24880
rect 3476 24828 3482 24880
rect 4157 24871 4215 24877
rect 3620 24840 3924 24868
rect 1394 24760 1400 24812
rect 1452 24760 1458 24812
rect 1671 24803 1729 24809
rect 1671 24769 1683 24803
rect 1717 24800 1729 24803
rect 2222 24800 2228 24812
rect 1717 24772 2228 24800
rect 1717 24769 1729 24772
rect 1671 24763 1729 24769
rect 2222 24760 2228 24772
rect 2280 24760 2286 24812
rect 2777 24803 2835 24809
rect 2777 24769 2789 24803
rect 2823 24769 2835 24803
rect 3620 24800 3648 24840
rect 2777 24763 2835 24769
rect 2976 24772 3648 24800
rect 2792 24664 2820 24763
rect 2976 24673 3004 24772
rect 3694 24760 3700 24812
rect 3752 24760 3758 24812
rect 3786 24760 3792 24812
rect 3844 24760 3850 24812
rect 3896 24800 3924 24840
rect 4157 24837 4169 24871
rect 4203 24868 4215 24871
rect 4246 24868 4252 24880
rect 4203 24840 4252 24868
rect 4203 24837 4215 24840
rect 4157 24831 4215 24837
rect 4246 24828 4252 24840
rect 4304 24828 4310 24880
rect 4338 24828 4344 24880
rect 4396 24868 4402 24880
rect 8312 24877 8340 24908
rect 8021 24871 8079 24877
rect 4396 24840 5856 24868
rect 4396 24828 4402 24840
rect 5442 24800 5448 24812
rect 3896 24772 5448 24800
rect 5442 24760 5448 24772
rect 5500 24760 5506 24812
rect 3326 24692 3332 24744
rect 3384 24692 3390 24744
rect 5828 24732 5856 24840
rect 8021 24837 8033 24871
rect 8067 24868 8079 24871
rect 8297 24871 8355 24877
rect 8067 24840 8156 24868
rect 8067 24837 8079 24840
rect 8021 24831 8079 24837
rect 5902 24760 5908 24812
rect 5960 24800 5966 24812
rect 6607 24803 6665 24809
rect 6607 24800 6619 24803
rect 5960 24772 6619 24800
rect 5960 24760 5966 24772
rect 6607 24769 6619 24772
rect 6653 24769 6665 24803
rect 8128 24800 8156 24840
rect 8297 24837 8309 24871
rect 8343 24837 8355 24871
rect 8297 24831 8355 24837
rect 9125 24871 9183 24877
rect 9125 24837 9137 24871
rect 9171 24837 9183 24871
rect 9214 24868 9242 24908
rect 9309 24905 9321 24939
rect 9355 24936 9367 24939
rect 10502 24936 10508 24948
rect 9355 24908 10508 24936
rect 9355 24905 9367 24908
rect 9309 24899 9367 24905
rect 10502 24896 10508 24908
rect 10560 24896 10566 24948
rect 10594 24896 10600 24948
rect 10652 24936 10658 24948
rect 12250 24936 12256 24948
rect 10652 24908 12256 24936
rect 10652 24896 10658 24908
rect 12250 24896 12256 24908
rect 12308 24896 12314 24948
rect 13170 24896 13176 24948
rect 13228 24896 13234 24948
rect 15930 24896 15936 24948
rect 15988 24896 15994 24948
rect 19889 24939 19947 24945
rect 19889 24905 19901 24939
rect 19935 24936 19947 24939
rect 19978 24936 19984 24948
rect 19935 24908 19984 24936
rect 19935 24905 19947 24908
rect 19889 24899 19947 24905
rect 19978 24896 19984 24908
rect 20036 24896 20042 24948
rect 20254 24936 20260 24948
rect 20070 24908 20260 24936
rect 9214 24840 9720 24868
rect 9125 24831 9183 24837
rect 8202 24800 8208 24812
rect 8128 24772 8208 24800
rect 6607 24763 6665 24769
rect 8202 24760 8208 24772
rect 8260 24760 8266 24812
rect 8386 24760 8392 24812
rect 8444 24760 8450 24812
rect 8757 24803 8815 24809
rect 8757 24769 8769 24803
rect 8803 24800 8815 24803
rect 8938 24800 8944 24812
rect 8803 24772 8944 24800
rect 8803 24769 8815 24772
rect 8757 24763 8815 24769
rect 8938 24760 8944 24772
rect 8996 24760 9002 24812
rect 8024 24744 8076 24750
rect 9140 24744 9168 24831
rect 9692 24800 9720 24840
rect 9692 24772 9904 24800
rect 6365 24735 6423 24741
rect 6365 24732 6377 24735
rect 5828 24704 6377 24732
rect 6365 24701 6377 24704
rect 6411 24701 6423 24735
rect 6365 24695 6423 24701
rect 2056 24636 2820 24664
rect 2961 24667 3019 24673
rect 1302 24556 1308 24608
rect 1360 24596 1366 24608
rect 2056 24596 2084 24636
rect 2961 24633 2973 24667
rect 3007 24633 3019 24667
rect 2961 24627 3019 24633
rect 4706 24624 4712 24676
rect 4764 24624 4770 24676
rect 5350 24624 5356 24676
rect 5408 24664 5414 24676
rect 6086 24664 6092 24676
rect 5408 24636 6092 24664
rect 5408 24624 5414 24636
rect 6086 24624 6092 24636
rect 6144 24624 6150 24676
rect 1360 24568 2084 24596
rect 1360 24556 1366 24568
rect 2406 24556 2412 24608
rect 2464 24556 2470 24608
rect 6380 24596 6408 24695
rect 9122 24692 9128 24744
rect 9180 24692 9186 24744
rect 9490 24692 9496 24744
rect 9548 24692 9554 24744
rect 9674 24692 9680 24744
rect 9732 24692 9738 24744
rect 8024 24686 8076 24692
rect 9876 24664 9904 24772
rect 10502 24760 10508 24812
rect 10560 24809 10566 24812
rect 10560 24803 10588 24809
rect 10576 24769 10588 24803
rect 10560 24763 10588 24769
rect 10689 24803 10747 24809
rect 10689 24769 10701 24803
rect 10735 24769 10747 24803
rect 10689 24763 10747 24769
rect 11333 24803 11391 24809
rect 11333 24769 11345 24803
rect 11379 24800 11391 24803
rect 11514 24800 11520 24812
rect 11379 24772 11520 24800
rect 11379 24769 11391 24772
rect 11333 24763 11391 24769
rect 10560 24760 10566 24763
rect 10042 24692 10048 24744
rect 10100 24732 10106 24744
rect 10137 24735 10195 24741
rect 10137 24732 10149 24735
rect 10100 24704 10149 24732
rect 10100 24692 10106 24704
rect 10137 24701 10149 24704
rect 10183 24701 10195 24735
rect 10410 24732 10416 24744
rect 10137 24695 10195 24701
rect 10242 24704 10416 24732
rect 10242 24664 10270 24704
rect 10410 24692 10416 24704
rect 10468 24692 10474 24744
rect 10704 24732 10732 24763
rect 11514 24760 11520 24772
rect 11572 24760 11578 24812
rect 12435 24803 12493 24809
rect 12435 24769 12447 24803
rect 12481 24800 12493 24803
rect 13262 24800 13268 24812
rect 12481 24772 13268 24800
rect 12481 24769 12493 24772
rect 12435 24763 12493 24769
rect 13262 24760 13268 24772
rect 13320 24760 13326 24812
rect 14826 24760 14832 24812
rect 14884 24800 14890 24812
rect 15470 24800 15476 24812
rect 14884 24772 15476 24800
rect 14884 24760 14890 24772
rect 15470 24760 15476 24772
rect 15528 24760 15534 24812
rect 15948 24800 15976 24896
rect 17954 24828 17960 24880
rect 18012 24828 18018 24880
rect 19242 24828 19248 24880
rect 19300 24868 19306 24880
rect 20070 24868 20098 24908
rect 20254 24896 20260 24908
rect 20312 24896 20318 24948
rect 19300 24840 20098 24868
rect 21560 24840 23888 24868
rect 19300 24828 19306 24840
rect 16393 24803 16451 24809
rect 16393 24800 16405 24803
rect 15948 24772 16405 24800
rect 16393 24769 16405 24772
rect 16439 24769 16451 24803
rect 16393 24763 16451 24769
rect 17497 24803 17555 24809
rect 17497 24769 17509 24803
rect 17543 24769 17555 24803
rect 17972 24800 18000 24828
rect 18782 24809 18788 24812
rect 18765 24803 18788 24809
rect 18765 24800 18777 24803
rect 17972 24772 18777 24800
rect 17497 24763 17555 24769
rect 18765 24769 18777 24772
rect 18765 24763 18788 24769
rect 10870 24732 10876 24744
rect 10704 24704 10876 24732
rect 10870 24692 10876 24704
rect 10928 24692 10934 24744
rect 12158 24692 12164 24744
rect 12216 24692 12222 24744
rect 16114 24692 16120 24744
rect 16172 24732 16178 24744
rect 17512 24732 17540 24763
rect 18782 24760 18788 24763
rect 18840 24760 18846 24812
rect 19981 24803 20039 24809
rect 19981 24769 19993 24803
rect 20027 24800 20039 24803
rect 20162 24800 20168 24812
rect 20027 24772 20168 24800
rect 20027 24769 20039 24772
rect 19981 24763 20039 24769
rect 16172 24704 17540 24732
rect 16172 24692 16178 24704
rect 18506 24692 18512 24744
rect 18564 24692 18570 24744
rect 9876 24636 10270 24664
rect 14550 24624 14556 24676
rect 14608 24664 14614 24676
rect 14918 24664 14924 24676
rect 14608 24636 14924 24664
rect 14608 24624 14614 24636
rect 14918 24624 14924 24636
rect 14976 24664 14982 24676
rect 16850 24664 16856 24676
rect 14976 24636 16856 24664
rect 14976 24624 14982 24636
rect 16850 24624 16856 24636
rect 16908 24624 16914 24676
rect 17494 24624 17500 24676
rect 17552 24664 17558 24676
rect 19996 24664 20024 24763
rect 20162 24760 20168 24772
rect 20220 24760 20226 24812
rect 20254 24760 20260 24812
rect 20312 24800 20318 24812
rect 20312 24772 20355 24800
rect 20312 24760 20318 24772
rect 20990 24760 20996 24812
rect 21048 24800 21054 24812
rect 21560 24800 21588 24840
rect 21048 24772 21588 24800
rect 21048 24760 21054 24772
rect 21634 24760 21640 24812
rect 21692 24800 21698 24812
rect 22097 24803 22155 24809
rect 22097 24800 22109 24803
rect 21692 24772 22109 24800
rect 21692 24760 21698 24772
rect 22097 24769 22109 24772
rect 22143 24769 22155 24803
rect 22741 24803 22799 24809
rect 22741 24800 22753 24803
rect 22097 24763 22155 24769
rect 22296 24772 22753 24800
rect 22296 24676 22324 24772
rect 22741 24769 22753 24772
rect 22787 24769 22799 24803
rect 22741 24763 22799 24769
rect 23198 24760 23204 24812
rect 23256 24760 23262 24812
rect 23293 24803 23351 24809
rect 23293 24769 23305 24803
rect 23339 24800 23351 24803
rect 23382 24800 23388 24812
rect 23339 24772 23388 24800
rect 23339 24769 23351 24772
rect 23293 24763 23351 24769
rect 23382 24760 23388 24772
rect 23440 24760 23446 24812
rect 23474 24760 23480 24812
rect 23532 24800 23538 24812
rect 23569 24803 23627 24809
rect 23569 24800 23581 24803
rect 23532 24772 23581 24800
rect 23532 24760 23538 24772
rect 23569 24769 23581 24772
rect 23615 24769 23627 24803
rect 23569 24763 23627 24769
rect 23753 24803 23811 24809
rect 23753 24769 23765 24803
rect 23799 24769 23811 24803
rect 23860 24800 23888 24840
rect 24121 24803 24179 24809
rect 24121 24800 24133 24803
rect 23860 24772 24133 24800
rect 23753 24763 23811 24769
rect 24121 24769 24133 24772
rect 24167 24769 24179 24803
rect 24121 24763 24179 24769
rect 23768 24732 23796 24763
rect 23492 24704 23796 24732
rect 17552 24636 17908 24664
rect 17552 24624 17558 24636
rect 6730 24596 6736 24608
rect 6380 24568 6736 24596
rect 6730 24556 6736 24568
rect 6788 24556 6794 24608
rect 10686 24556 10692 24608
rect 10744 24596 10750 24608
rect 10870 24596 10876 24608
rect 10744 24568 10876 24596
rect 10744 24556 10750 24568
rect 10870 24556 10876 24568
rect 10928 24596 10934 24608
rect 12986 24596 12992 24608
rect 10928 24568 12992 24596
rect 10928 24556 10934 24568
rect 12986 24556 12992 24568
rect 13044 24556 13050 24608
rect 14182 24556 14188 24608
rect 14240 24596 14246 24608
rect 15102 24596 15108 24608
rect 14240 24568 15108 24596
rect 14240 24556 14246 24568
rect 15102 24556 15108 24568
rect 15160 24556 15166 24608
rect 16206 24556 16212 24608
rect 16264 24556 16270 24608
rect 17313 24599 17371 24605
rect 17313 24565 17325 24599
rect 17359 24596 17371 24599
rect 17770 24596 17776 24608
rect 17359 24568 17776 24596
rect 17359 24565 17371 24568
rect 17313 24559 17371 24565
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 17880 24596 17908 24636
rect 19904 24636 20024 24664
rect 19904 24596 19932 24636
rect 22278 24624 22284 24676
rect 22336 24624 22342 24676
rect 23017 24667 23075 24673
rect 23017 24633 23029 24667
rect 23063 24664 23075 24667
rect 23492 24664 23520 24704
rect 23063 24636 23520 24664
rect 23063 24633 23075 24636
rect 23017 24627 23075 24633
rect 17880 24568 19932 24596
rect 19978 24556 19984 24608
rect 20036 24596 20042 24608
rect 20438 24596 20444 24608
rect 20036 24568 20444 24596
rect 20036 24556 20042 24568
rect 20438 24556 20444 24568
rect 20496 24596 20502 24608
rect 20993 24599 21051 24605
rect 20993 24596 21005 24599
rect 20496 24568 21005 24596
rect 20496 24556 20502 24568
rect 20993 24565 21005 24568
rect 21039 24565 21051 24599
rect 20993 24559 21051 24565
rect 21913 24599 21971 24605
rect 21913 24565 21925 24599
rect 21959 24596 21971 24599
rect 22370 24596 22376 24608
rect 21959 24568 22376 24596
rect 21959 24565 21971 24568
rect 21913 24559 21971 24565
rect 22370 24556 22376 24568
rect 22428 24556 22434 24608
rect 22557 24599 22615 24605
rect 22557 24565 22569 24599
rect 22603 24596 22615 24599
rect 22922 24596 22928 24608
rect 22603 24568 22928 24596
rect 22603 24565 22615 24568
rect 22557 24559 22615 24565
rect 22922 24556 22928 24568
rect 22980 24556 22986 24608
rect 23477 24599 23535 24605
rect 23477 24565 23489 24599
rect 23523 24596 23535 24599
rect 23566 24596 23572 24608
rect 23523 24568 23572 24596
rect 23523 24565 23535 24568
rect 23477 24559 23535 24565
rect 23566 24556 23572 24568
rect 23624 24556 23630 24608
rect 23658 24556 23664 24608
rect 23716 24556 23722 24608
rect 24394 24556 24400 24608
rect 24452 24556 24458 24608
rect 382 24488 388 24540
rect 440 24488 446 24540
rect 1104 24506 24840 24528
rect 400 24336 428 24488
rect 1104 24454 3917 24506
rect 3969 24454 3981 24506
rect 4033 24454 4045 24506
rect 4097 24454 4109 24506
rect 4161 24454 4173 24506
rect 4225 24454 9851 24506
rect 9903 24454 9915 24506
rect 9967 24454 9979 24506
rect 10031 24454 10043 24506
rect 10095 24454 10107 24506
rect 10159 24454 15785 24506
rect 15837 24454 15849 24506
rect 15901 24454 15913 24506
rect 15965 24454 15977 24506
rect 16029 24454 16041 24506
rect 16093 24454 21719 24506
rect 21771 24454 21783 24506
rect 21835 24454 21847 24506
rect 21899 24454 21911 24506
rect 21963 24454 21975 24506
rect 22027 24454 24840 24506
rect 1104 24432 24840 24454
rect 3050 24352 3056 24404
rect 3108 24352 3114 24404
rect 3142 24352 3148 24404
rect 3200 24392 3206 24404
rect 3694 24392 3700 24404
rect 3200 24364 3700 24392
rect 3200 24352 3206 24364
rect 3694 24352 3700 24364
rect 3752 24352 3758 24404
rect 3786 24352 3792 24404
rect 3844 24392 3850 24404
rect 4801 24395 4859 24401
rect 4801 24392 4813 24395
rect 3844 24364 4813 24392
rect 3844 24352 3850 24364
rect 4801 24361 4813 24364
rect 4847 24361 4859 24395
rect 8570 24392 8576 24404
rect 4801 24355 4859 24361
rect 8496 24364 8576 24392
rect 382 24284 388 24336
rect 440 24284 446 24336
rect 2406 24216 2412 24268
rect 2464 24216 2470 24268
rect 2866 24216 2872 24268
rect 2924 24256 2930 24268
rect 3789 24259 3847 24265
rect 3789 24256 3801 24259
rect 2924 24228 3801 24256
rect 2924 24216 2930 24228
rect 3789 24225 3801 24228
rect 3835 24225 3847 24259
rect 3789 24219 3847 24225
rect 2222 24148 2228 24200
rect 2280 24188 2286 24200
rect 4063 24191 4121 24197
rect 2280 24160 3924 24188
rect 2280 24148 2286 24160
rect 1765 24123 1823 24129
rect 1765 24089 1777 24123
rect 1811 24120 1823 24123
rect 1854 24120 1860 24132
rect 1811 24092 1860 24120
rect 1811 24089 1823 24092
rect 1765 24083 1823 24089
rect 1854 24080 1860 24092
rect 1912 24080 1918 24132
rect 2041 24123 2099 24129
rect 2041 24089 2053 24123
rect 2087 24089 2099 24123
rect 2041 24083 2099 24089
rect 2056 24052 2084 24083
rect 2130 24080 2136 24132
rect 2188 24080 2194 24132
rect 2501 24123 2559 24129
rect 2501 24089 2513 24123
rect 2547 24120 2559 24123
rect 2958 24120 2964 24132
rect 2547 24092 2964 24120
rect 2547 24089 2559 24092
rect 2501 24083 2559 24089
rect 2958 24080 2964 24092
rect 3016 24080 3022 24132
rect 3896 24120 3924 24160
rect 4063 24157 4075 24191
rect 4109 24188 4121 24191
rect 4154 24188 4160 24200
rect 4109 24160 4160 24188
rect 4109 24157 4121 24160
rect 4063 24151 4121 24157
rect 4154 24148 4160 24160
rect 4212 24188 4218 24200
rect 6454 24188 6460 24200
rect 4212 24160 6460 24188
rect 4212 24148 4218 24160
rect 6454 24148 6460 24160
rect 6512 24148 6518 24200
rect 8496 24188 8524 24364
rect 8570 24352 8576 24364
rect 8628 24352 8634 24404
rect 9490 24352 9496 24404
rect 9548 24392 9554 24404
rect 9548 24364 9904 24392
rect 9548 24352 9554 24364
rect 9876 24324 9904 24364
rect 10226 24352 10232 24404
rect 10284 24352 10290 24404
rect 15933 24395 15991 24401
rect 12360 24364 13216 24392
rect 12360 24324 12388 24364
rect 9876 24296 12388 24324
rect 8570 24216 8576 24268
rect 8628 24256 8634 24268
rect 9214 24256 9220 24268
rect 8628 24228 9220 24256
rect 8628 24216 8634 24228
rect 9214 24216 9220 24228
rect 9272 24216 9278 24268
rect 11606 24216 11612 24268
rect 11664 24216 11670 24268
rect 11793 24259 11851 24265
rect 11793 24225 11805 24259
rect 11839 24256 11851 24259
rect 11974 24256 11980 24268
rect 11839 24228 11980 24256
rect 11839 24225 11851 24228
rect 11793 24219 11851 24225
rect 11974 24216 11980 24228
rect 12032 24216 12038 24268
rect 12250 24216 12256 24268
rect 12308 24216 12314 24268
rect 12360 24256 12388 24296
rect 13188 24268 13216 24364
rect 15933 24361 15945 24395
rect 15979 24392 15991 24395
rect 16114 24392 16120 24404
rect 15979 24364 16120 24392
rect 15979 24361 15991 24364
rect 15933 24355 15991 24361
rect 16114 24352 16120 24364
rect 16172 24352 16178 24404
rect 16206 24352 16212 24404
rect 16264 24352 16270 24404
rect 17494 24352 17500 24404
rect 17552 24392 17558 24404
rect 17552 24364 17724 24392
rect 17552 24352 17558 24364
rect 14642 24284 14648 24336
rect 14700 24324 14706 24336
rect 14737 24327 14795 24333
rect 14737 24324 14749 24327
rect 14700 24296 14749 24324
rect 14700 24284 14706 24296
rect 14737 24293 14749 24296
rect 14783 24293 14795 24327
rect 14737 24287 14795 24293
rect 12667 24259 12725 24265
rect 12360 24228 12572 24256
rect 12544 24197 12572 24228
rect 12667 24225 12679 24259
rect 12713 24256 12725 24259
rect 12986 24256 12992 24268
rect 12713 24228 12992 24256
rect 12713 24225 12725 24228
rect 12667 24219 12725 24225
rect 12986 24216 12992 24228
rect 13044 24216 13050 24268
rect 13170 24216 13176 24268
rect 13228 24256 13234 24268
rect 14093 24259 14151 24265
rect 14093 24256 14105 24259
rect 13228 24228 14105 24256
rect 13228 24216 13234 24228
rect 14093 24225 14105 24228
rect 14139 24225 14151 24259
rect 14093 24219 14151 24225
rect 14277 24259 14335 24265
rect 14277 24225 14289 24259
rect 14323 24256 14335 24259
rect 14366 24256 14372 24268
rect 14323 24228 14372 24256
rect 14323 24225 14335 24228
rect 14277 24219 14335 24225
rect 9491 24191 9549 24197
rect 9491 24188 9503 24191
rect 8496 24160 9503 24188
rect 9491 24157 9503 24160
rect 9537 24188 9549 24191
rect 12529 24191 12587 24197
rect 9537 24160 11744 24188
rect 9537 24157 9549 24160
rect 9491 24151 9549 24157
rect 11716 24132 11744 24160
rect 12529 24157 12541 24191
rect 12575 24157 12587 24191
rect 12529 24151 12587 24157
rect 12802 24148 12808 24200
rect 12860 24148 12866 24200
rect 13722 24148 13728 24200
rect 13780 24188 13786 24200
rect 14182 24188 14188 24200
rect 13780 24160 14188 24188
rect 13780 24148 13786 24160
rect 14182 24148 14188 24160
rect 14240 24148 14246 24200
rect 6914 24120 6920 24132
rect 3896 24092 6920 24120
rect 6914 24080 6920 24092
rect 6972 24080 6978 24132
rect 7650 24080 7656 24132
rect 7708 24120 7714 24132
rect 9766 24120 9772 24132
rect 7708 24092 9772 24120
rect 7708 24080 7714 24092
rect 9766 24080 9772 24092
rect 9824 24080 9830 24132
rect 11698 24080 11704 24132
rect 11756 24080 11762 24132
rect 14292 24120 14320 24219
rect 14366 24216 14372 24228
rect 14424 24216 14430 24268
rect 14826 24216 14832 24268
rect 14884 24256 14890 24268
rect 15013 24259 15071 24265
rect 15013 24256 15025 24259
rect 14884 24228 15025 24256
rect 14884 24216 14890 24228
rect 15013 24225 15025 24228
rect 15059 24225 15071 24259
rect 15013 24219 15071 24225
rect 15102 24216 15108 24268
rect 15160 24265 15166 24268
rect 15160 24259 15188 24265
rect 15176 24225 15188 24259
rect 15160 24219 15188 24225
rect 15160 24216 15166 24219
rect 15286 24216 15292 24268
rect 15344 24216 15350 24268
rect 16224 24256 16252 24352
rect 16224 24228 16804 24256
rect 16298 24148 16304 24200
rect 16356 24188 16362 24200
rect 16776 24197 16804 24228
rect 16850 24216 16856 24268
rect 16908 24256 16914 24268
rect 17037 24259 17095 24265
rect 17037 24256 17049 24259
rect 16908 24228 17049 24256
rect 16908 24216 16914 24228
rect 17037 24225 17049 24228
rect 17083 24225 17095 24259
rect 17037 24219 17095 24225
rect 16577 24191 16635 24197
rect 16577 24188 16589 24191
rect 16356 24160 16589 24188
rect 16356 24148 16362 24160
rect 16577 24157 16589 24160
rect 16623 24157 16635 24191
rect 16577 24151 16635 24157
rect 16761 24191 16819 24197
rect 16761 24157 16773 24191
rect 16807 24157 16819 24191
rect 16761 24151 16819 24157
rect 17311 24191 17369 24197
rect 17311 24157 17323 24191
rect 17357 24188 17369 24191
rect 17696 24188 17724 24364
rect 20346 24352 20352 24404
rect 20404 24352 20410 24404
rect 21358 24352 21364 24404
rect 21416 24352 21422 24404
rect 21634 24352 21640 24404
rect 21692 24392 21698 24404
rect 21729 24395 21787 24401
rect 21729 24392 21741 24395
rect 21692 24364 21741 24392
rect 21692 24352 21698 24364
rect 21729 24361 21741 24364
rect 21775 24361 21787 24395
rect 21729 24355 21787 24361
rect 22922 24352 22928 24404
rect 22980 24352 22986 24404
rect 23198 24352 23204 24404
rect 23256 24392 23262 24404
rect 23385 24395 23443 24401
rect 23385 24392 23397 24395
rect 23256 24364 23397 24392
rect 23256 24352 23262 24364
rect 23385 24361 23397 24364
rect 23431 24361 23443 24395
rect 23385 24355 23443 24361
rect 23566 24352 23572 24404
rect 23624 24392 23630 24404
rect 25774 24392 25780 24404
rect 23624 24364 25780 24392
rect 23624 24352 23630 24364
rect 25774 24352 25780 24364
rect 25832 24352 25838 24404
rect 20162 24324 20168 24336
rect 17357 24160 17724 24188
rect 17788 24296 20168 24324
rect 17357 24157 17369 24160
rect 17311 24151 17369 24157
rect 17788 24120 17816 24296
rect 20162 24284 20168 24296
rect 20220 24284 20226 24336
rect 19797 24259 19855 24265
rect 19797 24225 19809 24259
rect 19843 24256 19855 24259
rect 20073 24259 20131 24265
rect 20073 24256 20085 24259
rect 19843 24228 20085 24256
rect 19843 24225 19855 24228
rect 19797 24219 19855 24225
rect 20073 24225 20085 24228
rect 20119 24225 20131 24259
rect 20073 24219 20131 24225
rect 20257 24259 20315 24265
rect 20257 24225 20269 24259
rect 20303 24256 20315 24259
rect 20364 24256 20392 24352
rect 20303 24228 20392 24256
rect 21376 24256 21404 24352
rect 22940 24324 22968 24352
rect 22940 24296 23520 24324
rect 21376 24228 22140 24256
rect 20303 24225 20315 24228
rect 20257 24219 20315 24225
rect 17954 24148 17960 24200
rect 18012 24188 18018 24200
rect 18322 24188 18328 24200
rect 18012 24160 18328 24188
rect 18012 24148 18018 24160
rect 18322 24148 18328 24160
rect 18380 24148 18386 24200
rect 18782 24148 18788 24200
rect 18840 24188 18846 24200
rect 19429 24191 19487 24197
rect 19429 24188 19441 24191
rect 18840 24160 19441 24188
rect 18840 24148 18846 24160
rect 19429 24157 19441 24160
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24157 19763 24191
rect 19705 24151 19763 24157
rect 19720 24120 19748 24151
rect 19886 24148 19892 24200
rect 19944 24148 19950 24200
rect 19978 24148 19984 24200
rect 20036 24148 20042 24200
rect 20162 24148 20168 24200
rect 20220 24188 20226 24200
rect 20349 24191 20407 24197
rect 20349 24188 20361 24191
rect 20220 24160 20361 24188
rect 20220 24148 20226 24160
rect 20349 24157 20361 24160
rect 20395 24188 20407 24191
rect 22005 24191 22063 24197
rect 22005 24188 22017 24191
rect 20395 24160 22017 24188
rect 20395 24157 20407 24160
rect 20349 24151 20407 24157
rect 22005 24157 22017 24160
rect 22051 24157 22063 24191
rect 22112 24188 22140 24228
rect 22278 24197 22284 24200
rect 22261 24191 22284 24197
rect 22261 24188 22273 24191
rect 22112 24160 22273 24188
rect 22005 24151 22063 24157
rect 22261 24157 22273 24160
rect 22261 24151 22284 24157
rect 22278 24148 22284 24151
rect 22336 24148 22342 24200
rect 23492 24197 23520 24296
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24157 23535 24191
rect 23477 24151 23535 24157
rect 23934 24148 23940 24200
rect 23992 24148 23998 24200
rect 13372 24092 14320 24120
rect 16776 24092 17816 24120
rect 19260 24092 19748 24120
rect 19904 24120 19932 24148
rect 20622 24129 20628 24132
rect 20594 24123 20628 24129
rect 20594 24120 20606 24123
rect 19904 24092 20606 24120
rect 2222 24052 2228 24064
rect 2056 24024 2228 24052
rect 2222 24012 2228 24024
rect 2280 24012 2286 24064
rect 2869 24055 2927 24061
rect 2869 24021 2881 24055
rect 2915 24052 2927 24055
rect 3234 24052 3240 24064
rect 2915 24024 3240 24052
rect 2915 24021 2927 24024
rect 2869 24015 2927 24021
rect 3234 24012 3240 24024
rect 3292 24012 3298 24064
rect 9674 24012 9680 24064
rect 9732 24052 9738 24064
rect 10594 24052 10600 24064
rect 9732 24024 10600 24052
rect 9732 24012 9738 24024
rect 10594 24012 10600 24024
rect 10652 24052 10658 24064
rect 13372 24052 13400 24092
rect 10652 24024 13400 24052
rect 13449 24055 13507 24061
rect 10652 24012 10658 24024
rect 13449 24021 13461 24055
rect 13495 24052 13507 24055
rect 16776 24052 16804 24092
rect 13495 24024 16804 24052
rect 13495 24021 13507 24024
rect 13449 24015 13507 24021
rect 16850 24012 16856 24064
rect 16908 24012 16914 24064
rect 18046 24012 18052 24064
rect 18104 24012 18110 24064
rect 19260 24061 19288 24092
rect 20594 24089 20606 24092
rect 20594 24083 20628 24089
rect 20622 24080 20628 24083
rect 20680 24080 20686 24132
rect 21174 24080 21180 24132
rect 21232 24080 21238 24132
rect 19245 24055 19303 24061
rect 19245 24021 19257 24055
rect 19291 24021 19303 24055
rect 19245 24015 19303 24021
rect 20257 24055 20315 24061
rect 20257 24021 20269 24055
rect 20303 24052 20315 24055
rect 21192 24052 21220 24080
rect 20303 24024 21220 24052
rect 20303 24021 20315 24024
rect 20257 24015 20315 24021
rect 23566 24012 23572 24064
rect 23624 24012 23630 24064
rect 24118 24012 24124 24064
rect 24176 24012 24182 24064
rect 1104 23962 25000 23984
rect 1104 23910 6884 23962
rect 6936 23910 6948 23962
rect 7000 23910 7012 23962
rect 7064 23910 7076 23962
rect 7128 23910 7140 23962
rect 7192 23910 12818 23962
rect 12870 23910 12882 23962
rect 12934 23910 12946 23962
rect 12998 23910 13010 23962
rect 13062 23910 13074 23962
rect 13126 23910 18752 23962
rect 18804 23910 18816 23962
rect 18868 23910 18880 23962
rect 18932 23910 18944 23962
rect 18996 23910 19008 23962
rect 19060 23910 24686 23962
rect 24738 23910 24750 23962
rect 24802 23910 24814 23962
rect 24866 23910 24878 23962
rect 24930 23910 24942 23962
rect 24994 23910 25000 23962
rect 1104 23888 25000 23910
rect 2130 23808 2136 23860
rect 2188 23848 2194 23860
rect 2777 23851 2835 23857
rect 2777 23848 2789 23851
rect 2188 23820 2789 23848
rect 2188 23808 2194 23820
rect 2777 23817 2789 23820
rect 2823 23817 2835 23851
rect 2777 23811 2835 23817
rect 3418 23808 3424 23860
rect 3476 23808 3482 23860
rect 3510 23808 3516 23860
rect 3568 23848 3574 23860
rect 3605 23851 3663 23857
rect 3605 23848 3617 23851
rect 3568 23820 3617 23848
rect 3568 23808 3574 23820
rect 3605 23817 3617 23820
rect 3651 23817 3663 23851
rect 4982 23848 4988 23860
rect 3605 23811 3663 23817
rect 4540 23820 4988 23848
rect 1302 23740 1308 23792
rect 1360 23780 1366 23792
rect 3436 23780 3464 23808
rect 1360 23752 2774 23780
rect 3436 23752 3556 23780
rect 1360 23740 1366 23752
rect 1486 23672 1492 23724
rect 1544 23672 1550 23724
rect 1670 23672 1676 23724
rect 1728 23712 1734 23724
rect 1765 23715 1823 23721
rect 1765 23712 1777 23715
rect 1728 23684 1777 23712
rect 1728 23672 1734 23684
rect 1765 23681 1777 23684
rect 1811 23681 1823 23715
rect 1765 23675 1823 23681
rect 2039 23715 2097 23721
rect 2039 23681 2051 23715
rect 2085 23712 2097 23715
rect 2590 23712 2596 23724
rect 2085 23684 2596 23712
rect 2085 23681 2097 23684
rect 2039 23675 2097 23681
rect 2590 23672 2596 23684
rect 2648 23672 2654 23724
rect 2746 23712 2774 23752
rect 3145 23715 3203 23721
rect 3145 23712 3157 23715
rect 2746 23684 3157 23712
rect 3145 23681 3157 23684
rect 3191 23681 3203 23715
rect 3145 23675 3203 23681
rect 3418 23672 3424 23724
rect 3476 23672 3482 23724
rect 1394 23604 1400 23656
rect 1452 23644 1458 23656
rect 1688 23644 1716 23672
rect 1452 23616 1716 23644
rect 3528 23644 3556 23752
rect 4540 23724 4568 23820
rect 4982 23808 4988 23820
rect 5040 23808 5046 23860
rect 5074 23808 5080 23860
rect 5132 23848 5138 23860
rect 5350 23848 5356 23860
rect 5132 23820 5356 23848
rect 5132 23808 5138 23820
rect 5350 23808 5356 23820
rect 5408 23808 5414 23860
rect 8386 23808 8392 23860
rect 8444 23848 8450 23860
rect 9125 23851 9183 23857
rect 9125 23848 9137 23851
rect 8444 23820 9137 23848
rect 8444 23808 8450 23820
rect 9125 23817 9137 23820
rect 9171 23817 9183 23851
rect 9125 23811 9183 23817
rect 12250 23808 12256 23860
rect 12308 23848 12314 23860
rect 12529 23851 12587 23857
rect 12529 23848 12541 23851
rect 12308 23820 12541 23848
rect 12308 23808 12314 23820
rect 12529 23817 12541 23820
rect 12575 23817 12587 23851
rect 12529 23811 12587 23817
rect 13446 23808 13452 23860
rect 13504 23808 13510 23860
rect 14918 23808 14924 23860
rect 14976 23848 14982 23860
rect 16574 23848 16580 23860
rect 14976 23820 16580 23848
rect 14976 23808 14982 23820
rect 16574 23808 16580 23820
rect 16632 23808 16638 23860
rect 16850 23808 16856 23860
rect 16908 23848 16914 23860
rect 16908 23820 18184 23848
rect 16908 23808 16914 23820
rect 8938 23780 8944 23792
rect 7760 23752 8944 23780
rect 4246 23672 4252 23724
rect 4304 23712 4310 23724
rect 4341 23715 4399 23721
rect 4341 23712 4353 23715
rect 4304 23684 4353 23712
rect 4304 23672 4310 23684
rect 4341 23681 4353 23684
rect 4387 23681 4399 23715
rect 4341 23675 4399 23681
rect 4522 23672 4528 23724
rect 4580 23672 4586 23724
rect 5258 23672 5264 23724
rect 5316 23672 5322 23724
rect 5378 23647 5436 23653
rect 5378 23644 5390 23647
rect 3528 23616 5390 23644
rect 1452 23604 1458 23616
rect 5378 23613 5390 23616
rect 5424 23613 5436 23647
rect 5378 23607 5436 23613
rect 5534 23604 5540 23656
rect 5592 23604 5598 23656
rect 1673 23579 1731 23585
rect 1673 23545 1685 23579
rect 1719 23545 1731 23579
rect 1673 23539 1731 23545
rect 1688 23508 1716 23539
rect 4982 23536 4988 23588
rect 5040 23536 5046 23588
rect 7760 23576 7788 23752
rect 8938 23740 8944 23752
rect 8996 23780 9002 23792
rect 13464 23780 13492 23808
rect 8996 23752 11284 23780
rect 8996 23740 9002 23752
rect 11256 23724 11284 23752
rect 11532 23752 12478 23780
rect 13464 23752 16954 23780
rect 8387 23715 8445 23721
rect 8387 23681 8399 23715
rect 8433 23712 8445 23715
rect 8433 23684 9674 23712
rect 8433 23681 8445 23684
rect 8387 23675 8445 23681
rect 7834 23604 7840 23656
rect 7892 23644 7898 23656
rect 8018 23644 8024 23656
rect 7892 23616 8024 23644
rect 7892 23604 7898 23616
rect 8018 23604 8024 23616
rect 8076 23644 8082 23656
rect 8113 23647 8171 23653
rect 8113 23644 8125 23647
rect 8076 23616 8125 23644
rect 8076 23604 8082 23616
rect 8113 23613 8125 23616
rect 8159 23613 8171 23647
rect 8113 23607 8171 23613
rect 6104 23548 7788 23576
rect 2774 23508 2780 23520
rect 1688 23480 2780 23508
rect 2774 23468 2780 23480
rect 2832 23468 2838 23520
rect 3329 23511 3387 23517
rect 3329 23477 3341 23511
rect 3375 23508 3387 23511
rect 6104 23508 6132 23548
rect 3375 23480 6132 23508
rect 3375 23477 3387 23480
rect 3329 23471 3387 23477
rect 6178 23468 6184 23520
rect 6236 23468 6242 23520
rect 9646 23508 9674 23684
rect 11238 23672 11244 23724
rect 11296 23672 11302 23724
rect 11532 23721 11560 23752
rect 11517 23715 11575 23721
rect 11517 23712 11529 23715
rect 11348 23684 11529 23712
rect 11054 23604 11060 23656
rect 11112 23644 11118 23656
rect 11348 23644 11376 23684
rect 11517 23681 11529 23684
rect 11563 23681 11575 23715
rect 11517 23675 11575 23681
rect 11698 23672 11704 23724
rect 11756 23712 11762 23724
rect 11791 23715 11849 23721
rect 11791 23712 11803 23715
rect 11756 23684 11803 23712
rect 11756 23672 11762 23684
rect 11791 23681 11803 23684
rect 11837 23712 11849 23715
rect 12342 23712 12348 23724
rect 11837 23684 12348 23712
rect 11837 23681 11849 23684
rect 11791 23675 11849 23681
rect 12342 23672 12348 23684
rect 12400 23672 12406 23724
rect 11112 23616 11376 23644
rect 12450 23644 12478 23752
rect 16926 23751 16954 23752
rect 16926 23745 16985 23751
rect 13630 23672 13636 23724
rect 13688 23712 13694 23724
rect 15286 23721 15292 23724
rect 15255 23715 15292 23721
rect 15255 23712 15267 23715
rect 13688 23684 15267 23712
rect 13688 23672 13694 23684
rect 15255 23681 15267 23684
rect 15255 23675 15292 23681
rect 15286 23672 15292 23675
rect 15344 23672 15350 23724
rect 16926 23714 16939 23745
rect 16927 23711 16939 23714
rect 16973 23711 16985 23745
rect 16927 23705 16985 23711
rect 18046 23672 18052 23724
rect 18104 23672 18110 23724
rect 18156 23712 18184 23820
rect 20622 23808 20628 23860
rect 20680 23808 20686 23860
rect 20809 23851 20867 23857
rect 20809 23817 20821 23851
rect 20855 23817 20867 23851
rect 20809 23811 20867 23817
rect 18233 23715 18291 23721
rect 18233 23712 18245 23715
rect 18156 23684 18245 23712
rect 18233 23681 18245 23684
rect 18279 23681 18291 23715
rect 18233 23675 18291 23681
rect 18598 23672 18604 23724
rect 18656 23672 18662 23724
rect 20640 23712 20668 23808
rect 20824 23780 20852 23811
rect 23474 23808 23480 23860
rect 23532 23808 23538 23860
rect 23106 23780 23112 23792
rect 20824 23752 21496 23780
rect 21468 23721 21496 23752
rect 21560 23752 23112 23780
rect 20993 23715 21051 23721
rect 20993 23712 21005 23715
rect 20640 23684 21005 23712
rect 20993 23681 21005 23684
rect 21039 23681 21051 23715
rect 20993 23675 21051 23681
rect 21453 23715 21511 23721
rect 21453 23681 21465 23715
rect 21499 23681 21511 23715
rect 21453 23675 21511 23681
rect 14642 23644 14648 23656
rect 12450 23616 14648 23644
rect 11112 23604 11118 23616
rect 14642 23604 14648 23616
rect 14700 23644 14706 23656
rect 15013 23647 15071 23653
rect 15013 23644 15025 23647
rect 14700 23616 15025 23644
rect 14700 23604 14706 23616
rect 15013 23613 15025 23616
rect 15059 23613 15071 23647
rect 16669 23647 16727 23653
rect 16669 23644 16681 23647
rect 15013 23607 15071 23613
rect 15672 23616 16681 23644
rect 13262 23508 13268 23520
rect 9646 23480 13268 23508
rect 13262 23468 13268 23480
rect 13320 23508 13326 23520
rect 13630 23508 13636 23520
rect 13320 23480 13636 23508
rect 13320 23468 13326 23480
rect 13630 23468 13636 23480
rect 13688 23468 13694 23520
rect 15028 23508 15056 23607
rect 15672 23508 15700 23616
rect 16669 23613 16681 23616
rect 16715 23613 16727 23647
rect 16669 23607 16727 23613
rect 17494 23604 17500 23656
rect 17552 23644 17558 23656
rect 21560 23644 21588 23752
rect 23106 23740 23112 23752
rect 23164 23740 23170 23792
rect 21821 23715 21879 23721
rect 21821 23712 21833 23715
rect 17552 23616 21588 23644
rect 21652 23684 21833 23712
rect 17552 23604 17558 23616
rect 21652 23588 21680 23684
rect 21821 23681 21833 23684
rect 21867 23712 21879 23715
rect 22189 23715 22247 23721
rect 22189 23712 22201 23715
rect 21867 23684 22201 23712
rect 21867 23681 21879 23684
rect 21821 23675 21879 23681
rect 22189 23681 22201 23684
rect 22235 23681 22247 23715
rect 22189 23675 22247 23681
rect 22370 23672 22376 23724
rect 22428 23672 22434 23724
rect 22462 23672 22468 23724
rect 22520 23672 22526 23724
rect 22739 23715 22797 23721
rect 22739 23681 22751 23715
rect 22785 23712 22797 23715
rect 22830 23712 22836 23724
rect 22785 23684 22836 23712
rect 22785 23681 22797 23684
rect 22739 23675 22797 23681
rect 22830 23672 22836 23684
rect 22888 23672 22894 23724
rect 24026 23672 24032 23724
rect 24084 23712 24090 23724
rect 24121 23715 24179 23721
rect 24121 23712 24133 23715
rect 24084 23684 24133 23712
rect 24084 23672 24090 23684
rect 24121 23681 24133 23684
rect 24167 23681 24179 23715
rect 24121 23675 24179 23681
rect 22097 23647 22155 23653
rect 22097 23613 22109 23647
rect 22143 23644 22155 23647
rect 22281 23647 22339 23653
rect 22281 23644 22293 23647
rect 22143 23616 22293 23644
rect 22143 23613 22155 23616
rect 22097 23607 22155 23613
rect 22281 23613 22293 23616
rect 22327 23613 22339 23647
rect 22281 23607 22339 23613
rect 18322 23536 18328 23588
rect 18380 23536 18386 23588
rect 19794 23536 19800 23588
rect 19852 23536 19858 23588
rect 21634 23536 21640 23588
rect 21692 23536 21698 23588
rect 15028 23480 15700 23508
rect 16025 23511 16083 23517
rect 16025 23477 16037 23511
rect 16071 23508 16083 23511
rect 16114 23508 16120 23520
rect 16071 23480 16120 23508
rect 16071 23477 16083 23480
rect 16025 23471 16083 23477
rect 16114 23468 16120 23480
rect 16172 23468 16178 23520
rect 16574 23468 16580 23520
rect 16632 23508 16638 23520
rect 17681 23511 17739 23517
rect 17681 23508 17693 23511
rect 16632 23480 17693 23508
rect 16632 23468 16638 23480
rect 17681 23477 17693 23480
rect 17727 23477 17739 23511
rect 17681 23471 17739 23477
rect 18782 23468 18788 23520
rect 18840 23508 18846 23520
rect 19812 23508 19840 23536
rect 18840 23480 19840 23508
rect 21545 23511 21603 23517
rect 18840 23468 18846 23480
rect 21545 23477 21557 23511
rect 21591 23508 21603 23511
rect 21913 23511 21971 23517
rect 21913 23508 21925 23511
rect 21591 23480 21925 23508
rect 21591 23477 21603 23480
rect 21545 23471 21603 23477
rect 21913 23477 21925 23480
rect 21959 23477 21971 23511
rect 21913 23471 21971 23477
rect 22005 23511 22063 23517
rect 22005 23477 22017 23511
rect 22051 23508 22063 23511
rect 23934 23508 23940 23520
rect 22051 23480 23940 23508
rect 22051 23477 22063 23480
rect 22005 23471 22063 23477
rect 23934 23468 23940 23480
rect 23992 23468 23998 23520
rect 24394 23468 24400 23520
rect 24452 23468 24458 23520
rect 1104 23418 24840 23440
rect 1104 23366 3917 23418
rect 3969 23366 3981 23418
rect 4033 23366 4045 23418
rect 4097 23366 4109 23418
rect 4161 23366 4173 23418
rect 4225 23366 9851 23418
rect 9903 23366 9915 23418
rect 9967 23366 9979 23418
rect 10031 23366 10043 23418
rect 10095 23366 10107 23418
rect 10159 23366 15785 23418
rect 15837 23366 15849 23418
rect 15901 23366 15913 23418
rect 15965 23366 15977 23418
rect 16029 23366 16041 23418
rect 16093 23366 21719 23418
rect 21771 23366 21783 23418
rect 21835 23366 21847 23418
rect 21899 23366 21911 23418
rect 21963 23366 21975 23418
rect 22027 23366 24840 23418
rect 1104 23344 24840 23366
rect 2498 23264 2504 23316
rect 2556 23304 2562 23316
rect 2556 23276 5488 23304
rect 2556 23264 2562 23276
rect 1394 23128 1400 23180
rect 1452 23128 1458 23180
rect 3068 23177 3096 23276
rect 5460 23236 5488 23276
rect 5534 23264 5540 23316
rect 5592 23304 5598 23316
rect 5813 23307 5871 23313
rect 5813 23304 5825 23307
rect 5592 23276 5825 23304
rect 5592 23264 5598 23276
rect 5813 23273 5825 23276
rect 5859 23273 5871 23307
rect 5813 23267 5871 23273
rect 6917 23307 6975 23313
rect 6917 23273 6929 23307
rect 6963 23304 6975 23307
rect 7190 23304 7196 23316
rect 6963 23276 7196 23304
rect 6963 23273 6975 23276
rect 6917 23267 6975 23273
rect 7190 23264 7196 23276
rect 7248 23264 7254 23316
rect 7300 23276 8708 23304
rect 7300 23236 7328 23276
rect 8680 23248 8708 23276
rect 9214 23264 9220 23316
rect 9272 23304 9278 23316
rect 17773 23307 17831 23313
rect 9272 23276 16988 23304
rect 9272 23264 9278 23276
rect 5460 23208 7328 23236
rect 8662 23196 8668 23248
rect 8720 23196 8726 23248
rect 12066 23196 12072 23248
rect 12124 23236 12130 23248
rect 12526 23236 12532 23248
rect 12124 23208 12532 23236
rect 12124 23196 12130 23208
rect 12526 23196 12532 23208
rect 12584 23196 12590 23248
rect 16025 23239 16083 23245
rect 16025 23205 16037 23239
rect 16071 23236 16083 23239
rect 16114 23236 16120 23248
rect 16071 23208 16120 23236
rect 16071 23205 16083 23208
rect 16025 23199 16083 23205
rect 16114 23196 16120 23208
rect 16172 23196 16178 23248
rect 16960 23236 16988 23276
rect 17773 23273 17785 23307
rect 17819 23304 17831 23307
rect 18598 23304 18604 23316
rect 17819 23276 18604 23304
rect 17819 23273 17831 23276
rect 17773 23267 17831 23273
rect 18598 23264 18604 23276
rect 18656 23264 18662 23316
rect 19334 23264 19340 23316
rect 19392 23304 19398 23316
rect 19392 23276 21588 23304
rect 19392 23264 19398 23276
rect 21560 23236 21588 23276
rect 21634 23264 21640 23316
rect 21692 23304 21698 23316
rect 21913 23307 21971 23313
rect 21913 23304 21925 23307
rect 21692 23276 21925 23304
rect 21692 23264 21698 23276
rect 21913 23273 21925 23276
rect 21959 23273 21971 23307
rect 21913 23267 21971 23273
rect 23474 23264 23480 23316
rect 23532 23264 23538 23316
rect 23566 23264 23572 23316
rect 23624 23304 23630 23316
rect 23937 23307 23995 23313
rect 23937 23304 23949 23307
rect 23624 23276 23949 23304
rect 23624 23264 23630 23276
rect 23937 23273 23949 23276
rect 23983 23273 23995 23307
rect 23937 23267 23995 23273
rect 24026 23264 24032 23316
rect 24084 23264 24090 23316
rect 22738 23236 22744 23248
rect 16960 23208 20484 23236
rect 21560 23208 22744 23236
rect 3053 23171 3111 23177
rect 3053 23137 3065 23171
rect 3099 23137 3111 23171
rect 3053 23131 3111 23137
rect 6730 23128 6736 23180
rect 6788 23168 6794 23180
rect 7377 23171 7435 23177
rect 7377 23168 7389 23171
rect 6788 23140 6960 23168
rect 6788 23128 6794 23140
rect 1671 23103 1729 23109
rect 1671 23069 1683 23103
rect 1717 23100 1729 23103
rect 2682 23100 2688 23112
rect 1717 23072 2688 23100
rect 1717 23069 1729 23072
rect 1671 23063 1729 23069
rect 2682 23060 2688 23072
rect 2740 23060 2746 23112
rect 2777 23103 2835 23109
rect 2777 23069 2789 23103
rect 2823 23069 2835 23103
rect 2777 23063 2835 23069
rect 4801 23103 4859 23109
rect 4801 23069 4813 23103
rect 4847 23069 4859 23103
rect 4801 23063 4859 23069
rect 5075 23103 5133 23109
rect 5075 23069 5087 23103
rect 5121 23100 5133 23103
rect 5442 23100 5448 23112
rect 5121 23072 5448 23100
rect 5121 23069 5133 23072
rect 5075 23063 5133 23069
rect 1302 22992 1308 23044
rect 1360 23032 1366 23044
rect 2792 23032 2820 23063
rect 1360 23004 2820 23032
rect 1360 22992 1366 23004
rect 4338 22992 4344 23044
rect 4396 23032 4402 23044
rect 4816 23032 4844 23063
rect 5442 23060 5448 23072
rect 5500 23060 5506 23112
rect 6178 23060 6184 23112
rect 6236 23100 6242 23112
rect 6641 23103 6699 23109
rect 6641 23100 6653 23103
rect 6236 23072 6653 23100
rect 6236 23060 6242 23072
rect 6641 23069 6653 23072
rect 6687 23069 6699 23103
rect 6641 23063 6699 23069
rect 6825 23103 6883 23109
rect 6825 23069 6837 23103
rect 6871 23069 6883 23103
rect 6825 23063 6883 23069
rect 6840 23032 6868 23063
rect 4396 23004 6224 23032
rect 4396 22992 4402 23004
rect 6196 22976 6224 23004
rect 6472 23004 6868 23032
rect 6932 23032 6960 23140
rect 7208 23140 7389 23168
rect 7098 23060 7104 23112
rect 7156 23060 7162 23112
rect 7208 23032 7236 23140
rect 7377 23137 7389 23140
rect 7423 23137 7435 23171
rect 7377 23131 7435 23137
rect 11698 23128 11704 23180
rect 11756 23168 11762 23180
rect 13538 23168 13544 23180
rect 11756 23140 13544 23168
rect 11756 23128 11762 23140
rect 13538 23128 13544 23140
rect 13596 23128 13602 23180
rect 13906 23128 13912 23180
rect 13964 23168 13970 23180
rect 15381 23171 15439 23177
rect 15381 23168 15393 23171
rect 13964 23140 15393 23168
rect 13964 23128 13970 23140
rect 15381 23137 15393 23140
rect 15427 23137 15439 23171
rect 16418 23171 16476 23177
rect 16418 23168 16430 23171
rect 15381 23131 15439 23137
rect 15470 23140 16430 23168
rect 7285 23103 7343 23109
rect 7285 23069 7297 23103
rect 7331 23094 7343 23103
rect 7331 23069 7512 23094
rect 7285 23066 7512 23069
rect 7285 23063 7343 23066
rect 6932 23004 7236 23032
rect 7484 23032 7512 23066
rect 7558 23060 7564 23112
rect 7616 23100 7622 23112
rect 7651 23103 7709 23109
rect 7651 23100 7663 23103
rect 7616 23072 7663 23100
rect 7616 23060 7622 23072
rect 7651 23069 7663 23072
rect 7697 23100 7709 23103
rect 7697 23072 8616 23100
rect 7697 23069 7709 23072
rect 7651 23063 7709 23069
rect 7484 23004 7604 23032
rect 2406 22924 2412 22976
rect 2464 22924 2470 22976
rect 4614 22924 4620 22976
rect 4672 22964 4678 22976
rect 5442 22964 5448 22976
rect 4672 22936 5448 22964
rect 4672 22924 4678 22936
rect 5442 22924 5448 22936
rect 5500 22924 5506 22976
rect 6178 22924 6184 22976
rect 6236 22924 6242 22976
rect 6472 22973 6500 23004
rect 7576 22976 7604 23004
rect 8294 22992 8300 23044
rect 8352 23032 8358 23044
rect 8588 23032 8616 23072
rect 9122 23060 9128 23112
rect 9180 23060 9186 23112
rect 9766 23060 9772 23112
rect 9824 23100 9830 23112
rect 9953 23103 10011 23109
rect 9953 23100 9965 23103
rect 9824 23072 9965 23100
rect 9824 23060 9830 23072
rect 9953 23069 9965 23072
rect 9999 23069 10011 23103
rect 9953 23063 10011 23069
rect 10134 23060 10140 23112
rect 10192 23100 10198 23112
rect 10227 23103 10285 23109
rect 10227 23100 10239 23103
rect 10192 23072 10239 23100
rect 10192 23060 10198 23072
rect 10227 23069 10239 23072
rect 10273 23069 10285 23103
rect 10227 23063 10285 23069
rect 14826 23060 14832 23112
rect 14884 23100 14890 23112
rect 15010 23100 15016 23112
rect 14884 23072 15016 23100
rect 14884 23060 14890 23072
rect 15010 23060 15016 23072
rect 15068 23100 15074 23112
rect 15470 23100 15498 23140
rect 16418 23137 16430 23140
rect 16464 23137 16476 23171
rect 16418 23131 16476 23137
rect 20456 23112 20484 23208
rect 22738 23196 22744 23208
rect 22796 23196 22802 23248
rect 20901 23171 20959 23177
rect 20901 23168 20913 23171
rect 20732 23140 20913 23168
rect 15068 23072 15498 23100
rect 15565 23103 15623 23109
rect 15068 23060 15074 23072
rect 15565 23069 15577 23103
rect 15611 23069 15623 23103
rect 15565 23063 15623 23069
rect 8352 23004 8524 23032
rect 8588 23004 11100 23032
rect 8352 22992 8358 23004
rect 6457 22967 6515 22973
rect 6457 22933 6469 22967
rect 6503 22933 6515 22967
rect 6457 22927 6515 22933
rect 7285 22967 7343 22973
rect 7285 22933 7297 22967
rect 7331 22964 7343 22967
rect 7466 22964 7472 22976
rect 7331 22936 7472 22964
rect 7331 22933 7343 22936
rect 7285 22927 7343 22933
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 7558 22924 7564 22976
rect 7616 22924 7622 22976
rect 8386 22924 8392 22976
rect 8444 22924 8450 22976
rect 8496 22964 8524 23004
rect 9766 22964 9772 22976
rect 8496 22936 9772 22964
rect 9766 22924 9772 22936
rect 9824 22924 9830 22976
rect 10962 22924 10968 22976
rect 11020 22924 11026 22976
rect 11072 22964 11100 23004
rect 11330 22992 11336 23044
rect 11388 23032 11394 23044
rect 12434 23032 12440 23044
rect 11388 23004 12440 23032
rect 11388 22992 11394 23004
rect 12434 22992 12440 23004
rect 12492 22992 12498 23044
rect 15194 22992 15200 23044
rect 15252 23032 15258 23044
rect 15580 23032 15608 23063
rect 16298 23060 16304 23112
rect 16356 23060 16362 23112
rect 16574 23060 16580 23112
rect 16632 23060 16638 23112
rect 17681 23103 17739 23109
rect 17681 23069 17693 23103
rect 17727 23069 17739 23103
rect 17681 23063 17739 23069
rect 15252 23004 15608 23032
rect 17696 23032 17724 23063
rect 17770 23060 17776 23112
rect 17828 23100 17834 23112
rect 17865 23103 17923 23109
rect 17865 23100 17877 23103
rect 17828 23072 17877 23100
rect 17828 23060 17834 23072
rect 17865 23069 17877 23072
rect 17911 23069 17923 23103
rect 17865 23063 17923 23069
rect 18046 23060 18052 23112
rect 18104 23060 18110 23112
rect 20438 23060 20444 23112
rect 20496 23060 20502 23112
rect 18064 23032 18092 23060
rect 17696 23004 18092 23032
rect 15252 22992 15258 23004
rect 19518 22992 19524 23044
rect 19576 23032 19582 23044
rect 20622 23032 20628 23044
rect 19576 23004 20628 23032
rect 19576 22992 19582 23004
rect 20622 22992 20628 23004
rect 20680 22992 20686 23044
rect 20732 23032 20760 23140
rect 20901 23137 20913 23140
rect 20947 23137 20959 23171
rect 20901 23131 20959 23137
rect 22462 23128 22468 23180
rect 22520 23128 22526 23180
rect 23492 23168 23520 23264
rect 23658 23196 23664 23248
rect 23716 23236 23722 23248
rect 23716 23208 24164 23236
rect 23716 23196 23722 23208
rect 24136 23177 24164 23208
rect 24121 23171 24179 23177
rect 23492 23140 23888 23168
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 21143 23103 21201 23109
rect 21143 23100 21155 23103
rect 20864 23072 21155 23100
rect 20864 23060 20870 23072
rect 21143 23069 21155 23072
rect 21189 23069 21201 23103
rect 21143 23063 21201 23069
rect 22480 23032 22508 23128
rect 23382 23060 23388 23112
rect 23440 23060 23446 23112
rect 23860 23109 23888 23140
rect 24121 23137 24133 23171
rect 24167 23137 24179 23171
rect 24121 23131 24179 23137
rect 23477 23103 23535 23109
rect 23477 23069 23489 23103
rect 23523 23069 23535 23103
rect 23477 23063 23535 23069
rect 23845 23103 23903 23109
rect 23845 23069 23857 23103
rect 23891 23069 23903 23103
rect 23845 23063 23903 23069
rect 20732 23004 22508 23032
rect 22554 22992 22560 23044
rect 22612 23032 22618 23044
rect 23492 23032 23520 23063
rect 22612 23004 23520 23032
rect 22612 22992 22618 23004
rect 13354 22964 13360 22976
rect 11072 22936 13360 22964
rect 13354 22924 13360 22936
rect 13412 22924 13418 22976
rect 17221 22967 17279 22973
rect 17221 22933 17233 22967
rect 17267 22964 17279 22967
rect 20898 22964 20904 22976
rect 17267 22936 20904 22964
rect 17267 22933 17279 22936
rect 17221 22927 17279 22933
rect 20898 22924 20904 22936
rect 20956 22924 20962 22976
rect 23198 22924 23204 22976
rect 23256 22924 23262 22976
rect 23658 22924 23664 22976
rect 23716 22924 23722 22976
rect 1104 22874 25000 22896
rect 1104 22822 6884 22874
rect 6936 22822 6948 22874
rect 7000 22822 7012 22874
rect 7064 22822 7076 22874
rect 7128 22822 7140 22874
rect 7192 22822 12818 22874
rect 12870 22822 12882 22874
rect 12934 22822 12946 22874
rect 12998 22822 13010 22874
rect 13062 22822 13074 22874
rect 13126 22822 18752 22874
rect 18804 22822 18816 22874
rect 18868 22822 18880 22874
rect 18932 22822 18944 22874
rect 18996 22822 19008 22874
rect 19060 22822 24686 22874
rect 24738 22822 24750 22874
rect 24802 22822 24814 22874
rect 24866 22822 24878 22874
rect 24930 22822 24942 22874
rect 24994 22822 25000 22874
rect 1104 22800 25000 22822
rect 1210 22720 1216 22772
rect 1268 22760 1274 22772
rect 9033 22763 9091 22769
rect 9033 22760 9045 22763
rect 1268 22732 9045 22760
rect 1268 22720 1274 22732
rect 9033 22729 9045 22732
rect 9079 22729 9091 22763
rect 9033 22723 9091 22729
rect 9122 22720 9128 22772
rect 9180 22720 9186 22772
rect 9214 22720 9220 22772
rect 9272 22720 9278 22772
rect 9953 22763 10011 22769
rect 9953 22729 9965 22763
rect 9999 22760 10011 22763
rect 9999 22732 11744 22760
rect 9999 22729 10011 22732
rect 9953 22723 10011 22729
rect 4246 22692 4252 22704
rect 2700 22664 4252 22692
rect 1671 22637 1729 22643
rect 1394 22584 1400 22636
rect 1452 22584 1458 22636
rect 1671 22603 1683 22637
rect 1717 22624 1729 22637
rect 2700 22624 2728 22664
rect 4246 22652 4252 22664
rect 4304 22652 4310 22704
rect 7929 22695 7987 22701
rect 7929 22692 7941 22695
rect 6104 22664 7941 22692
rect 1717 22603 2728 22624
rect 1671 22597 2728 22603
rect 1686 22596 2728 22597
rect 2774 22584 2780 22636
rect 2832 22584 2838 22636
rect 3142 22584 3148 22636
rect 3200 22584 3206 22636
rect 3789 22627 3847 22633
rect 3789 22593 3801 22627
rect 3835 22624 3847 22627
rect 4062 22624 4068 22636
rect 3835 22596 4068 22624
rect 3835 22593 3847 22596
rect 3789 22587 3847 22593
rect 4062 22584 4068 22596
rect 4120 22584 4126 22636
rect 4341 22627 4399 22633
rect 4341 22593 4353 22627
rect 4387 22624 4399 22627
rect 4430 22624 4436 22636
rect 4387 22596 4436 22624
rect 4387 22593 4399 22596
rect 4341 22587 4399 22593
rect 4430 22584 4436 22596
rect 4488 22624 4494 22636
rect 4488 22596 4752 22624
rect 4488 22584 4494 22596
rect 3160 22556 3188 22584
rect 4246 22556 4252 22568
rect 3160 22528 4252 22556
rect 4246 22516 4252 22528
rect 4304 22556 4310 22568
rect 4525 22559 4583 22565
rect 4525 22556 4537 22559
rect 4304 22528 4537 22556
rect 4304 22516 4310 22528
rect 4525 22525 4537 22528
rect 4571 22525 4583 22559
rect 4525 22519 4583 22525
rect 2958 22448 2964 22500
rect 3016 22448 3022 22500
rect 4724 22488 4752 22596
rect 5350 22584 5356 22636
rect 5408 22633 5414 22636
rect 5408 22627 5436 22633
rect 5424 22593 5436 22627
rect 5408 22587 5436 22593
rect 5408 22584 5414 22587
rect 4890 22516 4896 22568
rect 4948 22516 4954 22568
rect 4982 22516 4988 22568
rect 5040 22516 5046 22568
rect 5261 22559 5319 22565
rect 5261 22556 5273 22559
rect 5090 22528 5273 22556
rect 4798 22488 4804 22500
rect 4724 22460 4804 22488
rect 4798 22448 4804 22460
rect 4856 22448 4862 22500
rect 4908 22488 4936 22516
rect 5090 22488 5118 22528
rect 5261 22525 5273 22528
rect 5307 22525 5319 22559
rect 5261 22519 5319 22525
rect 5534 22516 5540 22568
rect 5592 22516 5598 22568
rect 4908 22460 5118 22488
rect 2406 22380 2412 22432
rect 2464 22380 2470 22432
rect 3970 22380 3976 22432
rect 4028 22380 4034 22432
rect 5534 22380 5540 22432
rect 5592 22420 5598 22432
rect 6104 22420 6132 22664
rect 7929 22661 7941 22664
rect 7975 22661 7987 22695
rect 7929 22655 7987 22661
rect 8205 22695 8263 22701
rect 8205 22661 8217 22695
rect 8251 22692 8263 22695
rect 9140 22692 9168 22720
rect 8251 22664 9168 22692
rect 8251 22661 8263 22664
rect 8205 22655 8263 22661
rect 10226 22652 10232 22704
rect 10284 22652 10290 22704
rect 10321 22695 10379 22701
rect 10321 22661 10333 22695
rect 10367 22692 10379 22695
rect 10962 22692 10968 22704
rect 10367 22664 10968 22692
rect 10367 22661 10379 22664
rect 10321 22655 10379 22661
rect 10962 22652 10968 22664
rect 11020 22652 11026 22704
rect 11057 22695 11115 22701
rect 11057 22661 11069 22695
rect 11103 22692 11115 22695
rect 11146 22692 11152 22704
rect 11103 22664 11152 22692
rect 11103 22661 11115 22664
rect 11057 22655 11115 22661
rect 11146 22652 11152 22664
rect 11204 22652 11210 22704
rect 11716 22692 11744 22732
rect 13262 22720 13268 22772
rect 13320 22720 13326 22772
rect 13814 22720 13820 22772
rect 13872 22720 13878 22772
rect 16666 22720 16672 22772
rect 16724 22760 16730 22772
rect 17034 22760 17040 22772
rect 16724 22732 17040 22760
rect 16724 22720 16730 22732
rect 17034 22720 17040 22732
rect 17092 22720 17098 22772
rect 19889 22763 19947 22769
rect 19889 22729 19901 22763
rect 19935 22729 19947 22763
rect 19889 22723 19947 22729
rect 13280 22692 13308 22720
rect 11716 22664 13308 22692
rect 6639 22627 6697 22633
rect 6639 22593 6651 22627
rect 6685 22624 6697 22627
rect 7834 22624 7840 22636
rect 6685 22596 7840 22624
rect 6685 22593 6697 22596
rect 6639 22587 6697 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 8294 22584 8300 22636
rect 8352 22584 8358 22636
rect 8662 22584 8668 22636
rect 8720 22584 8726 22636
rect 9122 22584 9128 22636
rect 9180 22624 9186 22636
rect 10410 22624 10416 22636
rect 9180 22596 10416 22624
rect 9180 22584 9186 22596
rect 10410 22584 10416 22596
rect 10468 22584 10474 22636
rect 10686 22584 10692 22636
rect 10744 22584 10750 22636
rect 11716 22633 11744 22664
rect 11701 22627 11759 22633
rect 11701 22593 11713 22627
rect 11747 22593 11759 22627
rect 11701 22587 11759 22593
rect 11882 22584 11888 22636
rect 11940 22584 11946 22636
rect 11974 22584 11980 22636
rect 12032 22624 12038 22636
rect 12955 22627 13013 22633
rect 12955 22624 12967 22627
rect 12032 22596 12967 22624
rect 12032 22584 12038 22596
rect 12955 22593 12967 22596
rect 13001 22593 13013 22627
rect 13832 22624 13860 22720
rect 18230 22652 18236 22704
rect 18288 22692 18294 22704
rect 18386 22695 18444 22701
rect 18386 22692 18398 22695
rect 18288 22664 18398 22692
rect 18288 22652 18294 22664
rect 18386 22661 18398 22664
rect 18432 22661 18444 22695
rect 19904 22692 19932 22723
rect 23198 22720 23204 22772
rect 23256 22720 23262 22772
rect 23661 22763 23719 22769
rect 23661 22729 23673 22763
rect 23707 22760 23719 22763
rect 23750 22760 23756 22772
rect 23707 22732 23756 22760
rect 23707 22729 23719 22732
rect 23661 22723 23719 22729
rect 23750 22720 23756 22732
rect 23808 22720 23814 22772
rect 19904 22664 20392 22692
rect 18386 22655 18444 22661
rect 14427 22627 14485 22633
rect 14427 22624 14439 22627
rect 13832 22596 14439 22624
rect 12955 22587 13013 22593
rect 14427 22593 14439 22596
rect 14473 22593 14485 22627
rect 14427 22587 14485 22593
rect 15654 22584 15660 22636
rect 15712 22624 15718 22636
rect 16298 22624 16304 22636
rect 15712 22596 16304 22624
rect 15712 22584 15718 22596
rect 16298 22584 16304 22596
rect 16356 22624 16362 22636
rect 19242 22624 19248 22636
rect 16356 22596 19248 22624
rect 16356 22584 16362 22596
rect 19242 22584 19248 22596
rect 19300 22584 19306 22636
rect 19610 22584 19616 22636
rect 19668 22584 19674 22636
rect 20364 22633 20392 22664
rect 20438 22652 20444 22704
rect 20496 22692 20502 22704
rect 21266 22692 21272 22704
rect 20496 22664 21272 22692
rect 20496 22652 20502 22664
rect 21266 22652 21272 22664
rect 21324 22652 21330 22704
rect 23216 22692 23244 22720
rect 23216 22664 23888 22692
rect 20073 22627 20131 22633
rect 20073 22593 20085 22627
rect 20119 22593 20131 22627
rect 20073 22587 20131 22593
rect 20165 22627 20223 22633
rect 20165 22593 20177 22627
rect 20211 22593 20223 22627
rect 20165 22587 20223 22593
rect 20349 22627 20407 22633
rect 20349 22593 20361 22627
rect 20395 22593 20407 22627
rect 20349 22587 20407 22593
rect 23385 22627 23443 22633
rect 23385 22593 23397 22627
rect 23431 22593 23443 22627
rect 23385 22587 23443 22593
rect 6178 22516 6184 22568
rect 6236 22556 6242 22568
rect 6365 22559 6423 22565
rect 6365 22556 6377 22559
rect 6236 22528 6377 22556
rect 6236 22516 6242 22528
rect 6365 22525 6377 22528
rect 6411 22525 6423 22559
rect 6365 22519 6423 22525
rect 5592 22392 6132 22420
rect 5592 22380 5598 22392
rect 6178 22380 6184 22432
rect 6236 22380 6242 22432
rect 6380 22420 6408 22519
rect 8386 22516 8392 22568
rect 8444 22516 8450 22568
rect 10502 22516 10508 22568
rect 10560 22516 10566 22568
rect 11241 22491 11299 22497
rect 11241 22457 11253 22491
rect 11287 22488 11299 22491
rect 11330 22488 11336 22500
rect 11287 22460 11336 22488
rect 11287 22457 11299 22460
rect 11241 22451 11299 22457
rect 11330 22448 11336 22460
rect 11388 22488 11394 22500
rect 11900 22488 11928 22584
rect 12710 22516 12716 22568
rect 12768 22516 12774 22568
rect 14185 22559 14243 22565
rect 14185 22525 14197 22559
rect 14231 22525 14243 22559
rect 14185 22519 14243 22525
rect 18141 22559 18199 22565
rect 18141 22525 18153 22559
rect 18187 22525 18199 22559
rect 20088 22556 20116 22587
rect 18141 22519 18199 22525
rect 19536 22528 20116 22556
rect 11388 22460 11928 22488
rect 11388 22448 11394 22460
rect 6638 22420 6644 22432
rect 6380 22392 6644 22420
rect 6638 22380 6644 22392
rect 6696 22380 6702 22432
rect 7190 22380 7196 22432
rect 7248 22420 7254 22432
rect 7374 22420 7380 22432
rect 7248 22392 7380 22420
rect 7248 22380 7254 22392
rect 7374 22380 7380 22392
rect 7432 22380 7438 22432
rect 9398 22380 9404 22432
rect 9456 22420 9462 22432
rect 9766 22420 9772 22432
rect 9456 22392 9772 22420
rect 9456 22380 9462 22392
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 11882 22380 11888 22432
rect 11940 22380 11946 22432
rect 13722 22380 13728 22432
rect 13780 22380 13786 22432
rect 14200 22420 14228 22519
rect 14642 22420 14648 22432
rect 14200 22392 14648 22420
rect 14642 22380 14648 22392
rect 14700 22380 14706 22432
rect 15102 22380 15108 22432
rect 15160 22420 15166 22432
rect 15197 22423 15255 22429
rect 15197 22420 15209 22423
rect 15160 22392 15209 22420
rect 15160 22380 15166 22392
rect 15197 22389 15209 22392
rect 15243 22389 15255 22423
rect 15197 22383 15255 22389
rect 15378 22380 15384 22432
rect 15436 22420 15442 22432
rect 15749 22423 15807 22429
rect 15749 22420 15761 22423
rect 15436 22392 15761 22420
rect 15436 22380 15442 22392
rect 15749 22389 15761 22392
rect 15795 22389 15807 22423
rect 18156 22420 18184 22519
rect 19536 22497 19564 22528
rect 19521 22491 19579 22497
rect 19521 22457 19533 22491
rect 19567 22457 19579 22491
rect 19521 22451 19579 22457
rect 19886 22448 19892 22500
rect 19944 22488 19950 22500
rect 20180 22488 20208 22587
rect 23400 22556 23428 22587
rect 23566 22584 23572 22636
rect 23624 22584 23630 22636
rect 23860 22633 23888 22664
rect 23845 22627 23903 22633
rect 23845 22593 23857 22627
rect 23891 22593 23903 22627
rect 23845 22587 23903 22593
rect 24121 22627 24179 22633
rect 24121 22593 24133 22627
rect 24167 22593 24179 22627
rect 24121 22587 24179 22593
rect 23658 22556 23664 22568
rect 23400 22528 23664 22556
rect 23658 22516 23664 22528
rect 23716 22516 23722 22568
rect 19944 22460 20208 22488
rect 19944 22448 19950 22460
rect 20622 22448 20628 22500
rect 20680 22488 20686 22500
rect 24136 22488 24164 22587
rect 20680 22460 24164 22488
rect 20680 22448 20686 22460
rect 18506 22420 18512 22432
rect 18156 22392 18512 22420
rect 15749 22383 15807 22389
rect 18506 22380 18512 22392
rect 18564 22420 18570 22432
rect 19242 22420 19248 22432
rect 18564 22392 19248 22420
rect 18564 22380 18570 22392
rect 19242 22380 19248 22392
rect 19300 22380 19306 22432
rect 19702 22380 19708 22432
rect 19760 22380 19766 22432
rect 20254 22380 20260 22432
rect 20312 22380 20318 22432
rect 23474 22380 23480 22432
rect 23532 22380 23538 22432
rect 24394 22380 24400 22432
rect 24452 22380 24458 22432
rect 1104 22330 24840 22352
rect 1104 22278 3917 22330
rect 3969 22278 3981 22330
rect 4033 22278 4045 22330
rect 4097 22278 4109 22330
rect 4161 22278 4173 22330
rect 4225 22278 9851 22330
rect 9903 22278 9915 22330
rect 9967 22278 9979 22330
rect 10031 22278 10043 22330
rect 10095 22278 10107 22330
rect 10159 22278 15785 22330
rect 15837 22278 15849 22330
rect 15901 22278 15913 22330
rect 15965 22278 15977 22330
rect 16029 22278 16041 22330
rect 16093 22278 21719 22330
rect 21771 22278 21783 22330
rect 21835 22278 21847 22330
rect 21899 22278 21911 22330
rect 21963 22278 21975 22330
rect 22027 22278 24840 22330
rect 1104 22256 24840 22278
rect 14 22176 20 22228
rect 72 22216 78 22228
rect 1302 22216 1308 22228
rect 72 22188 1308 22216
rect 72 22176 78 22188
rect 1302 22176 1308 22188
rect 1360 22176 1366 22228
rect 2774 22176 2780 22228
rect 2832 22216 2838 22228
rect 2869 22219 2927 22225
rect 2869 22216 2881 22219
rect 2832 22188 2881 22216
rect 2832 22176 2838 22188
rect 2869 22185 2881 22188
rect 2915 22185 2927 22219
rect 4338 22216 4344 22228
rect 2869 22179 2927 22185
rect 3896 22188 4344 22216
rect 3896 22092 3924 22188
rect 4338 22176 4344 22188
rect 4396 22176 4402 22228
rect 4893 22219 4951 22225
rect 4893 22185 4905 22219
rect 4939 22216 4951 22219
rect 4982 22216 4988 22228
rect 4939 22188 4988 22216
rect 4939 22185 4951 22188
rect 4893 22179 4951 22185
rect 4982 22176 4988 22188
rect 5040 22176 5046 22228
rect 5166 22176 5172 22228
rect 5224 22216 5230 22228
rect 5224 22188 7512 22216
rect 5224 22176 5230 22188
rect 7374 22108 7380 22160
rect 7432 22108 7438 22160
rect 2314 22040 2320 22092
rect 2372 22040 2378 22092
rect 3878 22040 3884 22092
rect 3936 22040 3942 22092
rect 4890 22040 4896 22092
rect 4948 22080 4954 22092
rect 5534 22080 5540 22092
rect 4948 22052 5540 22080
rect 4948 22040 4954 22052
rect 5534 22040 5540 22052
rect 5592 22040 5598 22092
rect 5994 22080 6000 22092
rect 5644 22052 6000 22080
rect 5644 22024 5672 22052
rect 5994 22040 6000 22052
rect 6052 22040 6058 22092
rect 7190 22040 7196 22092
rect 7248 22040 7254 22092
rect 7484 22080 7512 22188
rect 7558 22176 7564 22228
rect 7616 22176 7622 22228
rect 7666 22188 10180 22216
rect 7666 22080 7694 22188
rect 10152 22148 10180 22188
rect 10502 22176 10508 22228
rect 10560 22176 10566 22228
rect 11974 22216 11980 22228
rect 10612 22188 11980 22216
rect 10612 22148 10640 22188
rect 11974 22176 11980 22188
rect 12032 22176 12038 22228
rect 12710 22176 12716 22228
rect 12768 22176 12774 22228
rect 13924 22188 19334 22216
rect 10152 22120 10640 22148
rect 11054 22108 11060 22160
rect 11112 22108 11118 22160
rect 12728 22148 12756 22176
rect 12636 22120 12756 22148
rect 7484 22052 7694 22080
rect 8570 22040 8576 22092
rect 8628 22080 8634 22092
rect 9214 22080 9220 22092
rect 8628 22052 9220 22080
rect 8628 22040 8634 22052
rect 9214 22040 9220 22052
rect 9272 22040 9278 22092
rect 9398 22040 9404 22092
rect 9456 22080 9462 22092
rect 9493 22083 9551 22089
rect 9493 22080 9505 22083
rect 9456 22052 9505 22080
rect 9456 22040 9462 22052
rect 9493 22049 9505 22052
rect 9539 22049 9551 22083
rect 9493 22043 9551 22049
rect 11072 22080 11100 22108
rect 12636 22089 12664 22120
rect 11241 22083 11299 22089
rect 11241 22080 11253 22083
rect 11072 22052 11253 22080
rect 1949 22015 2007 22021
rect 1949 21981 1961 22015
rect 1995 22012 2007 22015
rect 2406 22012 2412 22024
rect 1995 21984 2412 22012
rect 1995 21981 2007 21984
rect 1949 21975 2007 21981
rect 2406 21972 2412 21984
rect 2464 21972 2470 22024
rect 4139 21985 4197 21991
rect 1854 21904 1860 21956
rect 1912 21904 1918 21956
rect 2038 21904 2044 21956
rect 2096 21904 2102 21956
rect 2317 21947 2375 21953
rect 2317 21913 2329 21947
rect 2363 21944 2375 21947
rect 2685 21947 2743 21953
rect 2363 21916 2452 21944
rect 2363 21913 2375 21916
rect 2317 21907 2375 21913
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 2056 21876 2084 21904
rect 2424 21888 2452 21916
rect 2685 21913 2697 21947
rect 2731 21944 2743 21947
rect 3602 21944 3608 21956
rect 2731 21916 3608 21944
rect 2731 21913 2743 21916
rect 2685 21907 2743 21913
rect 3602 21904 3608 21916
rect 3660 21904 3666 21956
rect 4139 21951 4151 21985
rect 4185 21982 4197 21985
rect 4185 21951 4200 21982
rect 5626 21972 5632 22024
rect 5684 21972 5690 22024
rect 7101 22015 7159 22021
rect 7101 21981 7113 22015
rect 7147 22012 7159 22015
rect 7282 22012 7288 22024
rect 7147 21984 7288 22012
rect 7147 21981 7159 21984
rect 7101 21975 7159 21981
rect 7282 21972 7288 21984
rect 7340 21972 7346 22024
rect 7466 21972 7472 22024
rect 7524 21972 7530 22024
rect 7745 22015 7803 22021
rect 7745 21981 7757 22015
rect 7791 21981 7803 22015
rect 7745 21975 7803 21981
rect 4139 21945 4200 21951
rect 4172 21944 4200 21945
rect 4430 21944 4436 21956
rect 4172 21916 4436 21944
rect 4430 21904 4436 21916
rect 4488 21944 4494 21956
rect 5994 21944 6000 21956
rect 4488 21916 6000 21944
rect 4488 21904 4494 21916
rect 5994 21904 6000 21916
rect 6052 21904 6058 21956
rect 6178 21904 6184 21956
rect 6236 21944 6242 21956
rect 7760 21944 7788 21975
rect 8662 21972 8668 22024
rect 8720 22012 8726 22024
rect 9306 22012 9312 22024
rect 8720 21984 9312 22012
rect 8720 21972 8726 21984
rect 9306 21972 9312 21984
rect 9364 21972 9370 22024
rect 9767 22015 9825 22021
rect 9767 21981 9779 22015
rect 9813 22012 9825 22015
rect 10226 22012 10232 22024
rect 9813 21984 10232 22012
rect 9813 21981 9825 21984
rect 9767 21975 9825 21981
rect 10226 21972 10232 21984
rect 10284 22012 10290 22024
rect 10410 22012 10416 22024
rect 10284 21984 10416 22012
rect 10284 21972 10290 21984
rect 10410 21972 10416 21984
rect 10468 21972 10474 22024
rect 6236 21916 7788 21944
rect 6236 21904 6242 21916
rect 8202 21904 8208 21956
rect 8260 21944 8266 21956
rect 11072 21944 11100 22052
rect 11241 22049 11253 22052
rect 11287 22049 11299 22083
rect 11241 22043 11299 22049
rect 12621 22083 12679 22089
rect 12621 22049 12633 22083
rect 12667 22049 12679 22083
rect 12621 22043 12679 22049
rect 11499 21985 11557 21991
rect 11499 21951 11511 21985
rect 11545 21982 11557 21985
rect 11545 21956 11560 21982
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 12863 22015 12921 22021
rect 12863 22012 12875 22015
rect 12492 21984 12875 22012
rect 12492 21972 12498 21984
rect 12863 21981 12875 21984
rect 12909 22012 12921 22015
rect 13924 22012 13952 22188
rect 15102 22108 15108 22160
rect 15160 22108 15166 22160
rect 17862 22108 17868 22160
rect 17920 22148 17926 22160
rect 18414 22148 18420 22160
rect 17920 22120 18420 22148
rect 17920 22108 17926 22120
rect 18414 22108 18420 22120
rect 18472 22108 18478 22160
rect 15378 22040 15384 22092
rect 15436 22040 15442 22092
rect 15519 22083 15577 22089
rect 15519 22049 15531 22083
rect 15565 22080 15577 22083
rect 16022 22080 16028 22092
rect 15565 22052 16028 22080
rect 15565 22049 15577 22052
rect 15519 22043 15577 22049
rect 16022 22040 16028 22052
rect 16080 22040 16086 22092
rect 19306 22080 19334 22188
rect 19702 22176 19708 22228
rect 19760 22216 19766 22228
rect 19797 22219 19855 22225
rect 19797 22216 19809 22219
rect 19760 22188 19809 22216
rect 19760 22176 19766 22188
rect 19797 22185 19809 22188
rect 19843 22185 19855 22219
rect 19797 22179 19855 22185
rect 20254 22176 20260 22228
rect 20312 22176 20318 22228
rect 21275 22188 21956 22216
rect 20272 22148 20300 22176
rect 19996 22120 20300 22148
rect 19886 22080 19892 22092
rect 19306 22052 19564 22080
rect 19536 22024 19564 22052
rect 19720 22052 19892 22080
rect 12909 21984 13952 22012
rect 14461 22015 14519 22021
rect 12909 21981 12921 21984
rect 12863 21975 12921 21981
rect 14461 21981 14473 22015
rect 14507 21981 14519 22015
rect 14461 21975 14519 21981
rect 14645 22015 14703 22021
rect 14645 21981 14657 22015
rect 14691 21981 14703 22015
rect 14645 21975 14703 21981
rect 11499 21945 11520 21951
rect 8260 21916 11100 21944
rect 8260 21904 8266 21916
rect 11514 21904 11520 21945
rect 11572 21904 11578 21956
rect 14476 21944 14504 21975
rect 11624 21916 14504 21944
rect 1627 21848 2084 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 2406 21836 2412 21888
rect 2464 21836 2470 21888
rect 2958 21836 2964 21888
rect 3016 21876 3022 21888
rect 11624 21876 11652 21916
rect 12176 21888 12204 21916
rect 3016 21848 11652 21876
rect 3016 21836 3022 21848
rect 12158 21836 12164 21888
rect 12216 21836 12222 21888
rect 12250 21836 12256 21888
rect 12308 21836 12314 21888
rect 13538 21836 13544 21888
rect 13596 21876 13602 21888
rect 13633 21879 13691 21885
rect 13633 21876 13645 21879
rect 13596 21848 13645 21876
rect 13596 21836 13602 21848
rect 13633 21845 13645 21848
rect 13679 21845 13691 21879
rect 13633 21839 13691 21845
rect 13814 21836 13820 21888
rect 13872 21876 13878 21888
rect 14660 21876 14688 21975
rect 15654 21972 15660 22024
rect 15712 21972 15718 22024
rect 17310 21972 17316 22024
rect 17368 22012 17374 22024
rect 17678 22012 17684 22024
rect 17368 21984 17684 22012
rect 17368 21972 17374 21984
rect 17678 21972 17684 21984
rect 17736 21972 17742 22024
rect 18230 21972 18236 22024
rect 18288 22012 18294 22024
rect 18877 22015 18935 22021
rect 18877 22012 18889 22015
rect 18288 21984 18889 22012
rect 18288 21972 18294 21984
rect 18877 21981 18889 21984
rect 18923 21981 18935 22015
rect 18877 21975 18935 21981
rect 19518 21972 19524 22024
rect 19576 21972 19582 22024
rect 19720 22021 19748 22052
rect 19886 22040 19892 22052
rect 19944 22040 19950 22092
rect 19996 22089 20024 22120
rect 19981 22083 20039 22089
rect 19981 22049 19993 22083
rect 20027 22049 20039 22083
rect 19981 22043 20039 22049
rect 20162 22040 20168 22092
rect 20220 22080 20226 22092
rect 20257 22083 20315 22089
rect 20257 22080 20269 22083
rect 20220 22052 20269 22080
rect 20220 22040 20226 22052
rect 20257 22049 20269 22052
rect 20303 22049 20315 22083
rect 20257 22043 20315 22049
rect 19705 22015 19763 22021
rect 19705 21981 19717 22015
rect 19751 21981 19763 22015
rect 20272 22012 20300 22043
rect 21275 22012 21303 22188
rect 21637 22151 21695 22157
rect 21637 22117 21649 22151
rect 21683 22117 21695 22151
rect 21637 22111 21695 22117
rect 20272 21984 21303 22012
rect 21652 22012 21680 22111
rect 21818 22108 21824 22160
rect 21876 22108 21882 22160
rect 21928 22080 21956 22188
rect 21928 22052 22324 22080
rect 22296 22024 22324 22052
rect 22005 22015 22063 22021
rect 22005 22012 22017 22015
rect 21652 21984 22017 22012
rect 19705 21975 19763 21981
rect 22005 21981 22017 21984
rect 22051 21981 22063 22015
rect 22005 21975 22063 21981
rect 22278 21972 22284 22024
rect 22336 22012 22342 22024
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 22336 21984 22385 22012
rect 22336 21972 22342 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 23937 22015 23995 22021
rect 23937 21981 23949 22015
rect 23983 22012 23995 22015
rect 25682 22012 25688 22024
rect 23983 21984 25688 22012
rect 23983 21981 23995 21984
rect 23937 21975 23995 21981
rect 25682 21972 25688 21984
rect 25740 21972 25746 22024
rect 20530 21953 20536 21956
rect 20524 21944 20536 21953
rect 16316 21916 20116 21944
rect 20491 21916 20536 21944
rect 16316 21885 16344 21916
rect 13872 21848 14688 21876
rect 16301 21879 16359 21885
rect 13872 21836 13878 21848
rect 16301 21845 16313 21879
rect 16347 21845 16359 21879
rect 16301 21839 16359 21845
rect 18693 21879 18751 21885
rect 18693 21845 18705 21879
rect 18739 21876 18751 21879
rect 19610 21876 19616 21888
rect 18739 21848 19616 21876
rect 18739 21845 18751 21848
rect 18693 21839 18751 21845
rect 19610 21836 19616 21848
rect 19668 21836 19674 21888
rect 19978 21836 19984 21888
rect 20036 21836 20042 21888
rect 20088 21876 20116 21916
rect 20524 21907 20536 21916
rect 20530 21904 20536 21907
rect 20588 21904 20594 21956
rect 22646 21953 22652 21956
rect 22618 21947 22652 21953
rect 22618 21944 22630 21947
rect 22066 21916 22630 21944
rect 22066 21876 22094 21916
rect 22618 21913 22630 21916
rect 22618 21907 22652 21913
rect 22646 21904 22652 21907
rect 22704 21904 22710 21956
rect 20088 21848 22094 21876
rect 23750 21836 23756 21888
rect 23808 21836 23814 21888
rect 24118 21836 24124 21888
rect 24176 21836 24182 21888
rect 1104 21786 25000 21808
rect 1104 21734 6884 21786
rect 6936 21734 6948 21786
rect 7000 21734 7012 21786
rect 7064 21734 7076 21786
rect 7128 21734 7140 21786
rect 7192 21734 12818 21786
rect 12870 21734 12882 21786
rect 12934 21734 12946 21786
rect 12998 21734 13010 21786
rect 13062 21734 13074 21786
rect 13126 21734 18752 21786
rect 18804 21734 18816 21786
rect 18868 21734 18880 21786
rect 18932 21734 18944 21786
rect 18996 21734 19008 21786
rect 19060 21734 24686 21786
rect 24738 21734 24750 21786
rect 24802 21734 24814 21786
rect 24866 21734 24878 21786
rect 24930 21734 24942 21786
rect 24994 21734 25000 21786
rect 1104 21712 25000 21734
rect 1857 21675 1915 21681
rect 1857 21641 1869 21675
rect 1903 21672 1915 21675
rect 3878 21672 3884 21684
rect 1903 21644 2176 21672
rect 1903 21641 1915 21644
rect 1857 21635 1915 21641
rect 2148 21616 2176 21644
rect 2240 21644 3884 21672
rect 1026 21564 1032 21616
rect 1084 21604 1090 21616
rect 1084 21576 1992 21604
rect 1084 21564 1090 21576
rect 1394 21496 1400 21548
rect 1452 21496 1458 21548
rect 1964 21545 1992 21576
rect 2130 21564 2136 21616
rect 2188 21564 2194 21616
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21505 1731 21539
rect 1673 21499 1731 21505
rect 1949 21539 2007 21545
rect 1949 21505 1961 21539
rect 1995 21505 2007 21539
rect 1949 21499 2007 21505
rect 842 21428 848 21480
rect 900 21468 906 21480
rect 1688 21468 1716 21499
rect 2038 21496 2044 21548
rect 2096 21536 2102 21548
rect 2240 21545 2268 21644
rect 3878 21632 3884 21644
rect 3936 21632 3942 21684
rect 6730 21632 6736 21684
rect 6788 21672 6794 21684
rect 8202 21672 8208 21684
rect 6788 21644 8208 21672
rect 6788 21632 6794 21644
rect 8202 21632 8208 21644
rect 8260 21632 8266 21684
rect 8386 21632 8392 21684
rect 8444 21672 8450 21684
rect 9217 21675 9275 21681
rect 9217 21672 9229 21675
rect 8444 21644 9229 21672
rect 8444 21632 8450 21644
rect 9217 21641 9229 21644
rect 9263 21641 9275 21675
rect 9217 21635 9275 21641
rect 12158 21632 12164 21684
rect 12216 21672 12222 21684
rect 13173 21675 13231 21681
rect 13173 21672 13185 21675
rect 12216 21644 13185 21672
rect 12216 21632 12222 21644
rect 13173 21641 13185 21644
rect 13219 21641 13231 21675
rect 13173 21635 13231 21641
rect 13464 21644 13676 21672
rect 2590 21564 2596 21616
rect 2648 21604 2654 21616
rect 2648 21576 4016 21604
rect 2648 21564 2654 21576
rect 2225 21539 2283 21545
rect 2225 21536 2237 21539
rect 2096 21508 2237 21536
rect 2096 21496 2102 21508
rect 2225 21505 2237 21508
rect 2271 21505 2283 21539
rect 2225 21499 2283 21505
rect 2498 21496 2504 21548
rect 2556 21536 2562 21548
rect 3050 21536 3056 21548
rect 2556 21508 3056 21536
rect 2556 21496 2562 21508
rect 3050 21496 3056 21508
rect 3108 21536 3114 21548
rect 3108 21508 3464 21536
rect 3108 21496 3114 21508
rect 900 21440 1716 21468
rect 900 21428 906 21440
rect 1581 21403 1639 21409
rect 1581 21369 1593 21403
rect 1627 21400 1639 21403
rect 1627 21372 2360 21400
rect 1627 21369 1639 21372
rect 1581 21363 1639 21369
rect 2332 21344 2360 21372
rect 2130 21292 2136 21344
rect 2188 21292 2194 21344
rect 2314 21292 2320 21344
rect 2372 21292 2378 21344
rect 3234 21292 3240 21344
rect 3292 21292 3298 21344
rect 3436 21332 3464 21508
rect 3786 21496 3792 21548
rect 3844 21536 3850 21548
rect 3879 21539 3937 21545
rect 3879 21536 3891 21539
rect 3844 21508 3891 21536
rect 3844 21496 3850 21508
rect 3879 21505 3891 21508
rect 3925 21505 3937 21539
rect 3988 21536 4016 21576
rect 4246 21564 4252 21616
rect 4304 21604 4310 21616
rect 7650 21604 7656 21616
rect 4304 21576 7656 21604
rect 4304 21564 4310 21576
rect 7650 21564 7656 21576
rect 7708 21564 7714 21616
rect 6883 21539 6941 21545
rect 6883 21536 6895 21539
rect 3988 21508 6895 21536
rect 3879 21499 3937 21505
rect 6883 21505 6895 21508
rect 6929 21505 6941 21539
rect 6883 21499 6941 21505
rect 7558 21496 7564 21548
rect 7616 21536 7622 21548
rect 7742 21536 7748 21548
rect 7616 21508 7748 21536
rect 7616 21496 7622 21508
rect 7742 21496 7748 21508
rect 7800 21496 7806 21548
rect 8220 21545 8248 21632
rect 8570 21564 8576 21616
rect 8628 21604 8634 21616
rect 13464 21604 13492 21644
rect 8628 21576 13492 21604
rect 8628 21564 8634 21576
rect 13538 21564 13544 21616
rect 13596 21564 13602 21616
rect 8479 21549 8537 21555
rect 8205 21539 8263 21545
rect 8205 21505 8217 21539
rect 8251 21505 8263 21539
rect 8205 21499 8263 21505
rect 8386 21496 8392 21548
rect 8444 21536 8450 21548
rect 8479 21546 8491 21549
rect 8478 21536 8491 21546
rect 8444 21515 8491 21536
rect 8525 21515 8537 21549
rect 8444 21509 8537 21515
rect 8444 21508 8506 21509
rect 8444 21496 8450 21508
rect 9306 21496 9312 21548
rect 9364 21536 9370 21548
rect 11440 21536 11652 21546
rect 11791 21539 11849 21545
rect 11791 21536 11803 21539
rect 9364 21518 11803 21536
rect 9364 21508 11468 21518
rect 11624 21508 11803 21518
rect 9364 21496 9370 21508
rect 11791 21505 11803 21508
rect 11837 21536 11849 21539
rect 12342 21536 12348 21548
rect 11837 21508 12348 21536
rect 11837 21505 11849 21508
rect 11791 21499 11849 21505
rect 12342 21496 12348 21508
rect 12400 21496 12406 21548
rect 13262 21496 13268 21548
rect 13320 21536 13326 21548
rect 13449 21539 13507 21545
rect 13449 21536 13461 21539
rect 13320 21508 13461 21536
rect 13320 21496 13326 21508
rect 13449 21505 13461 21508
rect 13495 21505 13507 21539
rect 13648 21536 13676 21644
rect 14182 21632 14188 21684
rect 14240 21672 14246 21684
rect 14277 21675 14335 21681
rect 14277 21672 14289 21675
rect 14240 21644 14289 21672
rect 14240 21632 14246 21644
rect 14277 21641 14289 21644
rect 14323 21641 14335 21675
rect 14277 21635 14335 21641
rect 15654 21632 15660 21684
rect 15712 21672 15718 21684
rect 15749 21675 15807 21681
rect 15749 21672 15761 21675
rect 15712 21644 15761 21672
rect 15712 21632 15718 21644
rect 15749 21641 15761 21644
rect 15795 21641 15807 21675
rect 15749 21635 15807 21641
rect 19886 21632 19892 21684
rect 19944 21632 19950 21684
rect 19978 21632 19984 21684
rect 20036 21672 20042 21684
rect 20990 21672 20996 21684
rect 20036 21644 20996 21672
rect 20036 21632 20042 21644
rect 20990 21632 20996 21644
rect 21048 21632 21054 21684
rect 21560 21644 22508 21672
rect 13814 21536 13820 21548
rect 13648 21508 13820 21536
rect 13449 21499 13507 21505
rect 13814 21496 13820 21508
rect 13872 21536 13878 21548
rect 13909 21539 13967 21545
rect 13909 21536 13921 21539
rect 13872 21508 13921 21536
rect 13872 21496 13878 21508
rect 13909 21505 13921 21508
rect 13955 21505 13967 21539
rect 13909 21499 13967 21505
rect 13998 21496 14004 21548
rect 14056 21536 14062 21548
rect 14200 21536 14228 21632
rect 14056 21508 14228 21536
rect 14056 21496 14062 21508
rect 14918 21496 14924 21548
rect 14976 21536 14982 21548
rect 15011 21539 15069 21545
rect 15011 21536 15023 21539
rect 14976 21508 15023 21536
rect 14976 21496 14982 21508
rect 15011 21505 15023 21508
rect 15057 21505 15069 21539
rect 15011 21499 15069 21505
rect 16666 21496 16672 21548
rect 16724 21496 16730 21548
rect 17678 21496 17684 21548
rect 17736 21545 17742 21548
rect 17736 21539 17764 21545
rect 17752 21505 17764 21539
rect 19119 21539 19177 21545
rect 19119 21536 19131 21539
rect 17736 21499 17764 21505
rect 18708 21508 19131 21536
rect 17736 21496 17742 21499
rect 3510 21428 3516 21480
rect 3568 21468 3574 21480
rect 3605 21471 3663 21477
rect 3605 21468 3617 21471
rect 3568 21440 3617 21468
rect 3568 21428 3574 21440
rect 3605 21437 3617 21440
rect 3651 21437 3663 21471
rect 6178 21468 6184 21480
rect 3605 21431 3663 21437
rect 4264 21440 6184 21468
rect 4264 21332 4292 21440
rect 6178 21428 6184 21440
rect 6236 21428 6242 21480
rect 6638 21428 6644 21480
rect 6696 21428 6702 21480
rect 11054 21428 11060 21480
rect 11112 21468 11118 21480
rect 11517 21471 11575 21477
rect 11517 21468 11529 21471
rect 11112 21440 11529 21468
rect 11112 21428 11118 21440
rect 11517 21437 11529 21440
rect 11563 21437 11575 21471
rect 11517 21431 11575 21437
rect 13722 21428 13728 21480
rect 13780 21428 13786 21480
rect 14734 21428 14740 21480
rect 14792 21428 14798 21480
rect 16390 21428 16396 21480
rect 16448 21468 16454 21480
rect 16850 21468 16856 21480
rect 16448 21440 16856 21468
rect 16448 21428 16454 21440
rect 16850 21428 16856 21440
rect 16908 21428 16914 21480
rect 17589 21471 17647 21477
rect 17589 21468 17601 21471
rect 16960 21440 17601 21468
rect 4430 21360 4436 21412
rect 4488 21400 4494 21412
rect 16960 21400 16988 21440
rect 17589 21437 17601 21440
rect 17635 21437 17647 21471
rect 17589 21431 17647 21437
rect 17862 21428 17868 21480
rect 17920 21428 17926 21480
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 18598 21468 18604 21480
rect 18104 21440 18604 21468
rect 18104 21428 18110 21440
rect 18598 21428 18604 21440
rect 18656 21428 18662 21480
rect 4488 21372 6776 21400
rect 4488 21360 4494 21372
rect 3436 21304 4292 21332
rect 4522 21292 4528 21344
rect 4580 21332 4586 21344
rect 4617 21335 4675 21341
rect 4617 21332 4629 21335
rect 4580 21304 4629 21332
rect 4580 21292 4586 21304
rect 4617 21301 4629 21304
rect 4663 21301 4675 21335
rect 6748 21332 6776 21372
rect 7576 21372 8340 21400
rect 7576 21332 7604 21372
rect 6748 21304 7604 21332
rect 4617 21295 4675 21301
rect 7650 21292 7656 21344
rect 7708 21292 7714 21344
rect 8312 21332 8340 21372
rect 16500 21372 16988 21400
rect 17313 21403 17371 21409
rect 16500 21344 16528 21372
rect 17313 21369 17325 21403
rect 17359 21369 17371 21403
rect 18708 21400 18736 21508
rect 19119 21505 19131 21508
rect 19165 21505 19177 21539
rect 19119 21499 19177 21505
rect 20530 21496 20536 21548
rect 20588 21536 20594 21548
rect 20993 21539 21051 21545
rect 20993 21536 21005 21539
rect 20588 21508 21005 21536
rect 20588 21496 20594 21508
rect 20993 21505 21005 21508
rect 21039 21505 21051 21539
rect 20993 21499 21051 21505
rect 21453 21539 21511 21545
rect 21453 21505 21465 21539
rect 21499 21505 21511 21539
rect 21453 21499 21511 21505
rect 18877 21471 18935 21477
rect 18877 21437 18889 21471
rect 18923 21437 18935 21471
rect 21468 21468 21496 21499
rect 18877 21431 18935 21437
rect 20824 21440 21496 21468
rect 17313 21363 17371 21369
rect 18248 21372 18736 21400
rect 9030 21332 9036 21344
rect 8312 21304 9036 21332
rect 9030 21292 9036 21304
rect 9088 21292 9094 21344
rect 12526 21292 12532 21344
rect 12584 21292 12590 21344
rect 14461 21335 14519 21341
rect 14461 21301 14473 21335
rect 14507 21332 14519 21335
rect 15102 21332 15108 21344
rect 14507 21304 15108 21332
rect 14507 21301 14519 21304
rect 14461 21295 14519 21301
rect 15102 21292 15108 21304
rect 15160 21292 15166 21344
rect 15654 21292 15660 21344
rect 15712 21332 15718 21344
rect 16482 21332 16488 21344
rect 15712 21304 16488 21332
rect 15712 21292 15718 21304
rect 16482 21292 16488 21304
rect 16540 21292 16546 21344
rect 17034 21292 17040 21344
rect 17092 21332 17098 21344
rect 17328 21332 17356 21363
rect 17092 21304 17356 21332
rect 17092 21292 17098 21304
rect 17678 21292 17684 21344
rect 17736 21332 17742 21344
rect 18248 21332 18276 21372
rect 17736 21304 18276 21332
rect 17736 21292 17742 21304
rect 18506 21292 18512 21344
rect 18564 21292 18570 21344
rect 18892 21332 18920 21431
rect 20824 21409 20852 21440
rect 20809 21403 20867 21409
rect 20809 21369 20821 21403
rect 20855 21369 20867 21403
rect 21174 21400 21180 21412
rect 20809 21363 20867 21369
rect 21100 21372 21180 21400
rect 19886 21332 19892 21344
rect 18892 21304 19892 21332
rect 19886 21292 19892 21304
rect 19944 21332 19950 21344
rect 21100 21332 21128 21372
rect 21174 21360 21180 21372
rect 21232 21400 21238 21412
rect 21560 21400 21588 21644
rect 21910 21564 21916 21616
rect 21968 21604 21974 21616
rect 21968 21576 22416 21604
rect 21968 21564 21974 21576
rect 21821 21539 21879 21545
rect 21821 21505 21833 21539
rect 21867 21536 21879 21539
rect 22002 21536 22008 21548
rect 21867 21508 22008 21536
rect 21867 21505 21879 21508
rect 21821 21499 21879 21505
rect 22002 21496 22008 21508
rect 22060 21536 22066 21548
rect 22388 21545 22416 21576
rect 22480 21548 22508 21644
rect 22646 21632 22652 21684
rect 22704 21632 22710 21684
rect 23658 21632 23664 21684
rect 23716 21672 23722 21684
rect 23753 21675 23811 21681
rect 23753 21672 23765 21675
rect 23716 21644 23765 21672
rect 23716 21632 23722 21644
rect 23753 21641 23765 21644
rect 23799 21641 23811 21675
rect 23753 21635 23811 21641
rect 22189 21539 22247 21545
rect 22189 21536 22201 21539
rect 22060 21508 22201 21536
rect 22060 21496 22066 21508
rect 22189 21505 22201 21508
rect 22235 21505 22247 21539
rect 22189 21499 22247 21505
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 22462 21496 22468 21548
rect 22520 21496 22526 21548
rect 22664 21545 22692 21632
rect 22999 21569 23057 21575
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21505 22707 21539
rect 22999 21535 23011 21569
rect 23045 21566 23057 21569
rect 23045 21548 23060 21566
rect 22999 21529 23020 21535
rect 22649 21499 22707 21505
rect 23014 21496 23020 21529
rect 23072 21496 23078 21548
rect 23768 21536 23796 21635
rect 24121 21539 24179 21545
rect 24121 21536 24133 21539
rect 23768 21508 24133 21536
rect 24121 21505 24133 21508
rect 24167 21505 24179 21539
rect 24121 21499 24179 21505
rect 24486 21496 24492 21548
rect 24544 21536 24550 21548
rect 25314 21536 25320 21548
rect 24544 21508 25320 21536
rect 24544 21496 24550 21508
rect 25314 21496 25320 21508
rect 25372 21496 25378 21548
rect 22097 21471 22155 21477
rect 22097 21437 22109 21471
rect 22143 21468 22155 21471
rect 22281 21471 22339 21477
rect 22281 21468 22293 21471
rect 22143 21440 22293 21468
rect 22143 21437 22155 21440
rect 22097 21431 22155 21437
rect 22281 21437 22293 21440
rect 22327 21437 22339 21471
rect 22480 21468 22508 21496
rect 22741 21471 22799 21477
rect 22741 21468 22753 21471
rect 22480 21440 22753 21468
rect 22281 21431 22339 21437
rect 22741 21437 22753 21440
rect 22787 21437 22799 21471
rect 22741 21431 22799 21437
rect 23474 21428 23480 21480
rect 23532 21468 23538 21480
rect 24397 21471 24455 21477
rect 24397 21468 24409 21471
rect 23532 21440 24409 21468
rect 23532 21428 23538 21440
rect 24397 21437 24409 21440
rect 24443 21437 24455 21471
rect 24397 21431 24455 21437
rect 21232 21372 21588 21400
rect 22005 21403 22063 21409
rect 21232 21360 21238 21372
rect 22005 21369 22017 21403
rect 22051 21400 22063 21403
rect 22646 21400 22652 21412
rect 22051 21372 22652 21400
rect 22051 21369 22063 21372
rect 22005 21363 22063 21369
rect 22646 21360 22652 21372
rect 22704 21360 22710 21412
rect 24118 21360 24124 21412
rect 24176 21400 24182 21412
rect 24305 21403 24363 21409
rect 24305 21400 24317 21403
rect 24176 21372 24317 21400
rect 24176 21360 24182 21372
rect 24305 21369 24317 21372
rect 24351 21369 24363 21403
rect 24305 21363 24363 21369
rect 19944 21304 21128 21332
rect 21545 21335 21603 21341
rect 19944 21292 19950 21304
rect 21545 21301 21557 21335
rect 21591 21332 21603 21335
rect 21913 21335 21971 21341
rect 21913 21332 21925 21335
rect 21591 21304 21925 21332
rect 21591 21301 21603 21304
rect 21545 21295 21603 21301
rect 21913 21301 21925 21304
rect 21959 21301 21971 21335
rect 21913 21295 21971 21301
rect 22462 21292 22468 21344
rect 22520 21292 22526 21344
rect 24210 21292 24216 21344
rect 24268 21292 24274 21344
rect 1104 21242 24840 21264
rect 1104 21190 3917 21242
rect 3969 21190 3981 21242
rect 4033 21190 4045 21242
rect 4097 21190 4109 21242
rect 4161 21190 4173 21242
rect 4225 21190 9851 21242
rect 9903 21190 9915 21242
rect 9967 21190 9979 21242
rect 10031 21190 10043 21242
rect 10095 21190 10107 21242
rect 10159 21190 15785 21242
rect 15837 21190 15849 21242
rect 15901 21190 15913 21242
rect 15965 21190 15977 21242
rect 16029 21190 16041 21242
rect 16093 21190 21719 21242
rect 21771 21190 21783 21242
rect 21835 21190 21847 21242
rect 21899 21190 21911 21242
rect 21963 21190 21975 21242
rect 22027 21190 24840 21242
rect 1104 21168 24840 21190
rect 1581 21131 1639 21137
rect 1581 21097 1593 21131
rect 1627 21128 1639 21131
rect 1670 21128 1676 21140
rect 1627 21100 1676 21128
rect 1627 21097 1639 21100
rect 1581 21091 1639 21097
rect 1670 21088 1676 21100
rect 1728 21088 1734 21140
rect 1949 21131 2007 21137
rect 1949 21097 1961 21131
rect 1995 21128 2007 21131
rect 4430 21128 4436 21140
rect 1995 21100 4436 21128
rect 1995 21097 2007 21100
rect 1949 21091 2007 21097
rect 4430 21088 4436 21100
rect 4488 21088 4494 21140
rect 4982 21128 4988 21140
rect 4724 21100 4988 21128
rect 2038 21020 2044 21072
rect 2096 21060 2102 21072
rect 2096 21032 2176 21060
rect 2096 21020 2102 21032
rect 2148 21001 2176 21032
rect 2133 20995 2191 21001
rect 2133 20961 2145 20995
rect 2179 20961 2191 20995
rect 2133 20955 2191 20961
rect 2866 20952 2872 21004
rect 2924 20992 2930 21004
rect 3510 20992 3516 21004
rect 2924 20964 3516 20992
rect 2924 20952 2930 20964
rect 3510 20952 3516 20964
rect 3568 20992 3574 21004
rect 3694 20992 3700 21004
rect 3568 20964 3700 20992
rect 3568 20952 3574 20964
rect 3694 20952 3700 20964
rect 3752 20952 3758 21004
rect 4724 21001 4752 21100
rect 4982 21088 4988 21100
rect 5040 21088 5046 21140
rect 7101 21131 7159 21137
rect 7101 21097 7113 21131
rect 7147 21128 7159 21131
rect 7374 21128 7380 21140
rect 7147 21100 7380 21128
rect 7147 21097 7159 21100
rect 7101 21091 7159 21097
rect 7374 21088 7380 21100
rect 7432 21088 7438 21140
rect 9030 21088 9036 21140
rect 9088 21128 9094 21140
rect 11330 21128 11336 21140
rect 9088 21100 11336 21128
rect 9088 21088 9094 21100
rect 11330 21088 11336 21100
rect 11388 21128 11394 21140
rect 12526 21128 12532 21140
rect 11388 21100 11744 21128
rect 11388 21088 11394 21100
rect 7282 21060 7288 21072
rect 6932 21032 7288 21060
rect 4709 20995 4767 21001
rect 4709 20961 4721 20995
rect 4755 20961 4767 20995
rect 4709 20955 4767 20961
rect 934 20884 940 20936
rect 992 20924 998 20936
rect 1765 20927 1823 20933
rect 1765 20924 1777 20927
rect 992 20896 1777 20924
rect 992 20884 998 20896
rect 1765 20893 1777 20896
rect 1811 20893 1823 20927
rect 1765 20887 1823 20893
rect 2038 20884 2044 20936
rect 2096 20924 2102 20936
rect 2407 20927 2465 20933
rect 2407 20924 2419 20927
rect 2096 20896 2419 20924
rect 2096 20884 2102 20896
rect 2407 20893 2419 20896
rect 2453 20924 2465 20927
rect 3786 20924 3792 20936
rect 2453 20896 2636 20924
rect 2453 20893 2465 20896
rect 2407 20887 2465 20893
rect 2608 20868 2636 20896
rect 2700 20896 3792 20924
rect 2700 20868 2728 20896
rect 3786 20884 3792 20896
rect 3844 20884 3850 20936
rect 4983 20927 5041 20933
rect 4983 20893 4995 20927
rect 5029 20924 5041 20927
rect 6270 20924 6276 20936
rect 5029 20896 6276 20924
rect 5029 20893 5041 20896
rect 4983 20887 5041 20893
rect 6270 20884 6276 20896
rect 6328 20924 6334 20936
rect 6932 20924 6960 21032
rect 7282 21020 7288 21032
rect 7340 21020 7346 21072
rect 7650 20952 7656 21004
rect 7708 20952 7714 21004
rect 9214 20952 9220 21004
rect 9272 20992 9278 21004
rect 9401 20995 9459 21001
rect 9401 20992 9413 20995
rect 9272 20964 9413 20992
rect 9272 20952 9278 20964
rect 9401 20961 9413 20964
rect 9447 20961 9459 20995
rect 9401 20955 9459 20961
rect 11146 20952 11152 21004
rect 11204 20992 11210 21004
rect 11716 21001 11744 21100
rect 12176 21100 12532 21128
rect 12176 21069 12204 21100
rect 12526 21088 12532 21100
rect 12584 21088 12590 21140
rect 14734 21088 14740 21140
rect 14792 21128 14798 21140
rect 16666 21128 16672 21140
rect 14792 21100 16672 21128
rect 14792 21088 14798 21100
rect 16666 21088 16672 21100
rect 16724 21088 16730 21140
rect 18598 21088 18604 21140
rect 18656 21128 18662 21140
rect 18969 21131 19027 21137
rect 18969 21128 18981 21131
rect 18656 21100 18981 21128
rect 18656 21088 18662 21100
rect 18969 21097 18981 21100
rect 19015 21097 19027 21131
rect 18969 21091 19027 21097
rect 19058 21088 19064 21140
rect 19116 21128 19122 21140
rect 19116 21100 21864 21128
rect 19116 21088 19122 21100
rect 12161 21063 12219 21069
rect 12161 21029 12173 21063
rect 12207 21029 12219 21063
rect 12161 21023 12219 21029
rect 16025 21063 16083 21069
rect 16025 21029 16037 21063
rect 16071 21060 16083 21063
rect 17034 21060 17040 21072
rect 16071 21032 17040 21060
rect 16071 21029 16083 21032
rect 16025 21023 16083 21029
rect 17034 21020 17040 21032
rect 17092 21020 17098 21072
rect 18325 21063 18383 21069
rect 18325 21029 18337 21063
rect 18371 21060 18383 21063
rect 18371 21032 18920 21060
rect 18371 21029 18383 21032
rect 18325 21023 18383 21029
rect 11517 20995 11575 21001
rect 11517 20992 11529 20995
rect 11204 20964 11529 20992
rect 11204 20952 11210 20964
rect 11517 20961 11529 20964
rect 11563 20961 11575 20995
rect 11517 20955 11575 20961
rect 11701 20995 11759 21001
rect 11701 20961 11713 20995
rect 11747 20961 11759 20995
rect 11701 20955 11759 20961
rect 12250 20952 12256 21004
rect 12308 20992 12314 21004
rect 12308 20964 12756 20992
rect 12308 20952 12314 20964
rect 6328 20896 6960 20924
rect 6328 20884 6334 20896
rect 7282 20884 7288 20936
rect 7340 20924 7346 20936
rect 7340 20896 7420 20924
rect 7340 20884 7346 20896
rect 1486 20816 1492 20868
rect 1544 20816 1550 20868
rect 2590 20816 2596 20868
rect 2648 20816 2654 20868
rect 2682 20816 2688 20868
rect 2740 20816 2746 20868
rect 7392 20865 7420 20896
rect 7466 20884 7472 20936
rect 7524 20884 7530 20936
rect 7558 20884 7564 20936
rect 7616 20924 7622 20936
rect 8113 20927 8171 20933
rect 8113 20924 8125 20927
rect 7616 20896 8125 20924
rect 7616 20884 7622 20896
rect 8113 20893 8125 20896
rect 8159 20893 8171 20927
rect 9643 20927 9701 20933
rect 9643 20924 9655 20927
rect 8113 20887 8171 20893
rect 8312 20896 9655 20924
rect 7377 20859 7435 20865
rect 3528 20828 7052 20856
rect 3528 20800 3556 20828
rect 2130 20748 2136 20800
rect 2188 20788 2194 20800
rect 2498 20788 2504 20800
rect 2188 20760 2504 20788
rect 2188 20748 2194 20760
rect 2498 20748 2504 20760
rect 2556 20748 2562 20800
rect 3050 20748 3056 20800
rect 3108 20788 3114 20800
rect 3145 20791 3203 20797
rect 3145 20788 3157 20791
rect 3108 20760 3157 20788
rect 3108 20748 3114 20760
rect 3145 20757 3157 20760
rect 3191 20757 3203 20791
rect 3145 20751 3203 20757
rect 3510 20748 3516 20800
rect 3568 20748 3574 20800
rect 5442 20748 5448 20800
rect 5500 20788 5506 20800
rect 5721 20791 5779 20797
rect 5721 20788 5733 20791
rect 5500 20760 5733 20788
rect 5500 20748 5506 20760
rect 5721 20757 5733 20760
rect 5767 20757 5779 20791
rect 7024 20788 7052 20828
rect 7377 20825 7389 20859
rect 7423 20825 7435 20859
rect 7484 20856 7512 20884
rect 8312 20868 8340 20896
rect 9643 20893 9655 20896
rect 9689 20924 9701 20927
rect 9689 20896 11744 20924
rect 9689 20893 9701 20896
rect 9643 20887 9701 20893
rect 7653 20859 7711 20865
rect 7653 20856 7665 20859
rect 7484 20828 7665 20856
rect 7377 20819 7435 20825
rect 7653 20825 7665 20828
rect 7699 20825 7711 20859
rect 7653 20819 7711 20825
rect 7742 20816 7748 20868
rect 7800 20816 7806 20868
rect 8294 20816 8300 20868
rect 8352 20816 8358 20868
rect 8938 20856 8944 20868
rect 8496 20828 8944 20856
rect 8496 20797 8524 20828
rect 8938 20816 8944 20828
rect 8996 20816 9002 20868
rect 8481 20791 8539 20797
rect 8481 20788 8493 20791
rect 7024 20760 8493 20788
rect 5721 20751 5779 20757
rect 8481 20757 8493 20760
rect 8527 20757 8539 20791
rect 8481 20751 8539 20757
rect 8665 20791 8723 20797
rect 8665 20757 8677 20791
rect 8711 20788 8723 20791
rect 9030 20788 9036 20800
rect 8711 20760 9036 20788
rect 8711 20757 8723 20760
rect 8665 20751 8723 20757
rect 9030 20748 9036 20760
rect 9088 20748 9094 20800
rect 10410 20748 10416 20800
rect 10468 20748 10474 20800
rect 11716 20788 11744 20896
rect 12434 20884 12440 20936
rect 12492 20884 12498 20936
rect 12526 20884 12532 20936
rect 12584 20933 12590 20936
rect 12728 20933 12756 20964
rect 14550 20952 14556 21004
rect 14608 20992 14614 21004
rect 15010 20992 15016 21004
rect 14608 20964 15016 20992
rect 14608 20952 14614 20964
rect 15010 20952 15016 20964
rect 15068 20952 15074 21004
rect 18230 20992 18236 21004
rect 15672 20964 18236 20992
rect 12584 20927 12612 20933
rect 12600 20893 12612 20927
rect 12584 20887 12612 20893
rect 12713 20927 12771 20933
rect 12713 20893 12725 20927
rect 12759 20893 12771 20927
rect 15672 20924 15700 20964
rect 18230 20952 18236 20964
rect 18288 20952 18294 21004
rect 18432 20964 18828 20992
rect 15302 20903 15700 20924
rect 15271 20897 15700 20903
rect 15271 20894 15283 20897
rect 12713 20887 12771 20893
rect 12584 20884 12590 20887
rect 15212 20866 15283 20894
rect 15212 20856 15240 20866
rect 15271 20863 15283 20866
rect 15317 20896 15700 20897
rect 16393 20927 16451 20933
rect 15317 20866 15330 20896
rect 16393 20893 16405 20927
rect 16439 20893 16451 20927
rect 16393 20887 16451 20893
rect 16577 20927 16635 20933
rect 16577 20893 16589 20927
rect 16623 20924 16635 20927
rect 16758 20924 16764 20936
rect 16623 20896 16764 20924
rect 16623 20893 16635 20896
rect 16577 20887 16635 20893
rect 15317 20863 15329 20866
rect 15271 20857 15329 20863
rect 13280 20828 15240 20856
rect 13280 20788 13308 20828
rect 15562 20816 15568 20868
rect 15620 20856 15626 20868
rect 16408 20856 16436 20887
rect 16758 20884 16764 20896
rect 16816 20884 16822 20936
rect 17310 20884 17316 20936
rect 17368 20884 17374 20936
rect 17402 20884 17408 20936
rect 17460 20933 17466 20936
rect 17460 20927 17488 20933
rect 17476 20893 17488 20927
rect 17460 20887 17488 20893
rect 17460 20884 17466 20887
rect 17586 20884 17592 20936
rect 17644 20884 17650 20936
rect 18432 20924 18460 20964
rect 18248 20896 18460 20924
rect 18248 20865 18276 20896
rect 18506 20884 18512 20936
rect 18564 20929 18570 20936
rect 18800 20933 18828 20964
rect 18892 20933 18920 21032
rect 19518 21020 19524 21072
rect 19576 21060 19582 21072
rect 19978 21060 19984 21072
rect 19576 21032 19984 21060
rect 19576 21020 19582 21032
rect 19978 21020 19984 21032
rect 20036 21020 20042 21072
rect 21836 21060 21864 21100
rect 22094 21088 22100 21140
rect 22152 21128 22158 21140
rect 22189 21131 22247 21137
rect 22189 21128 22201 21131
rect 22152 21100 22201 21128
rect 22152 21088 22158 21100
rect 22189 21097 22201 21100
rect 22235 21097 22247 21131
rect 22189 21091 22247 21097
rect 22462 21088 22468 21140
rect 22520 21088 22526 21140
rect 22646 21088 22652 21140
rect 22704 21088 22710 21140
rect 23385 21131 23443 21137
rect 23385 21097 23397 21131
rect 23431 21128 23443 21131
rect 24210 21128 24216 21140
rect 23431 21100 24216 21128
rect 23431 21097 23443 21100
rect 23385 21091 23443 21097
rect 24210 21088 24216 21100
rect 24268 21088 24274 21140
rect 21836 21032 22094 21060
rect 18966 20952 18972 21004
rect 19024 20992 19030 21004
rect 19024 20964 20024 20992
rect 19024 20952 19030 20964
rect 18564 20884 18575 20929
rect 18785 20927 18843 20933
rect 18785 20893 18797 20927
rect 18831 20893 18843 20927
rect 18785 20887 18843 20893
rect 18877 20927 18935 20933
rect 18877 20893 18889 20927
rect 18923 20893 18935 20927
rect 19889 20927 19947 20933
rect 19889 20924 19901 20927
rect 18877 20887 18935 20893
rect 19628 20896 19901 20924
rect 18517 20883 18575 20884
rect 15620 20828 16436 20856
rect 18233 20859 18291 20865
rect 15620 20816 15626 20828
rect 18233 20825 18245 20859
rect 18279 20825 18291 20859
rect 18233 20819 18291 20825
rect 11716 20760 13308 20788
rect 13357 20791 13415 20797
rect 13357 20757 13369 20791
rect 13403 20788 13415 20791
rect 18506 20788 18512 20800
rect 13403 20760 18512 20788
rect 13403 20757 13415 20760
rect 13357 20751 13415 20757
rect 18506 20748 18512 20760
rect 18564 20748 18570 20800
rect 18601 20791 18659 20797
rect 18601 20757 18613 20791
rect 18647 20788 18659 20791
rect 19426 20788 19432 20800
rect 18647 20760 19432 20788
rect 18647 20757 18659 20760
rect 18601 20751 18659 20757
rect 19426 20748 19432 20760
rect 19484 20748 19490 20800
rect 19518 20748 19524 20800
rect 19576 20788 19582 20800
rect 19628 20788 19656 20896
rect 19889 20893 19901 20896
rect 19935 20893 19947 20927
rect 19889 20887 19947 20893
rect 19996 20856 20024 20964
rect 21174 20952 21180 21004
rect 21232 20952 21238 21004
rect 21419 20927 21477 20933
rect 21419 20924 21431 20927
rect 21275 20896 21431 20924
rect 21275 20856 21303 20896
rect 21419 20893 21431 20896
rect 21465 20893 21477 20927
rect 21419 20887 21477 20893
rect 19996 20828 21303 20856
rect 22066 20856 22094 21032
rect 22480 20924 22508 21088
rect 22664 20992 22692 21088
rect 22664 20964 23704 20992
rect 23676 20933 23704 20964
rect 23293 20927 23351 20933
rect 23293 20924 23305 20927
rect 22480 20896 23305 20924
rect 23293 20893 23305 20896
rect 23339 20893 23351 20927
rect 23293 20887 23351 20893
rect 23661 20927 23719 20933
rect 23661 20893 23673 20927
rect 23707 20893 23719 20927
rect 23661 20887 23719 20893
rect 22830 20856 22836 20868
rect 22066 20828 22836 20856
rect 22830 20816 22836 20828
rect 22888 20816 22894 20868
rect 19576 20760 19656 20788
rect 19576 20748 19582 20760
rect 19702 20748 19708 20800
rect 19760 20748 19766 20800
rect 23934 20748 23940 20800
rect 23992 20748 23998 20800
rect 1104 20698 25000 20720
rect 1104 20646 6884 20698
rect 6936 20646 6948 20698
rect 7000 20646 7012 20698
rect 7064 20646 7076 20698
rect 7128 20646 7140 20698
rect 7192 20646 12818 20698
rect 12870 20646 12882 20698
rect 12934 20646 12946 20698
rect 12998 20646 13010 20698
rect 13062 20646 13074 20698
rect 13126 20646 18752 20698
rect 18804 20646 18816 20698
rect 18868 20646 18880 20698
rect 18932 20646 18944 20698
rect 18996 20646 19008 20698
rect 19060 20646 24686 20698
rect 24738 20646 24750 20698
rect 24802 20646 24814 20698
rect 24866 20646 24878 20698
rect 24930 20646 24942 20698
rect 24994 20646 25000 20698
rect 1104 20624 25000 20646
rect 1210 20544 1216 20596
rect 1268 20584 1274 20596
rect 1627 20587 1685 20593
rect 1627 20584 1639 20587
rect 1268 20556 1639 20584
rect 1268 20544 1274 20556
rect 1627 20553 1639 20556
rect 1673 20553 1685 20587
rect 1627 20547 1685 20553
rect 2501 20587 2559 20593
rect 2501 20553 2513 20587
rect 2547 20553 2559 20587
rect 2501 20547 2559 20553
rect 2516 20516 2544 20547
rect 2590 20544 2596 20596
rect 2648 20584 2654 20596
rect 4801 20587 4859 20593
rect 4801 20584 4813 20587
rect 2648 20556 4813 20584
rect 2648 20544 2654 20556
rect 4801 20553 4813 20556
rect 4847 20584 4859 20587
rect 7374 20584 7380 20596
rect 4847 20556 7380 20584
rect 4847 20553 4859 20556
rect 4801 20547 4859 20553
rect 7374 20544 7380 20556
rect 7432 20544 7438 20596
rect 7742 20544 7748 20596
rect 7800 20584 7806 20596
rect 8573 20587 8631 20593
rect 8573 20584 8585 20587
rect 7800 20556 8585 20584
rect 7800 20544 7806 20556
rect 8573 20553 8585 20556
rect 8619 20553 8631 20587
rect 8573 20547 8631 20553
rect 9401 20587 9459 20593
rect 9401 20553 9413 20587
rect 9447 20584 9459 20587
rect 10318 20584 10324 20596
rect 9447 20556 10324 20584
rect 9447 20553 9459 20556
rect 9401 20547 9459 20553
rect 10318 20544 10324 20556
rect 10376 20584 10382 20596
rect 10778 20584 10784 20596
rect 10376 20556 10784 20584
rect 10376 20544 10382 20556
rect 10778 20544 10784 20556
rect 10836 20544 10842 20596
rect 11514 20544 11520 20596
rect 11572 20584 11578 20596
rect 12066 20584 12072 20596
rect 11572 20556 12072 20584
rect 11572 20544 11578 20556
rect 12066 20544 12072 20556
rect 12124 20544 12130 20596
rect 12434 20544 12440 20596
rect 12492 20544 12498 20596
rect 16482 20544 16488 20596
rect 16540 20584 16546 20596
rect 17494 20584 17500 20596
rect 16540 20556 17500 20584
rect 16540 20544 16546 20556
rect 17494 20544 17500 20556
rect 17552 20544 17558 20596
rect 17586 20544 17592 20596
rect 17644 20584 17650 20596
rect 17862 20584 17868 20596
rect 17644 20556 17868 20584
rect 17644 20544 17650 20556
rect 17862 20544 17868 20556
rect 17920 20584 17926 20596
rect 18049 20587 18107 20593
rect 18049 20584 18061 20587
rect 17920 20556 18061 20584
rect 17920 20544 17926 20556
rect 18049 20553 18061 20556
rect 18095 20553 18107 20587
rect 18049 20547 18107 20553
rect 18506 20544 18512 20596
rect 18564 20584 18570 20596
rect 19518 20584 19524 20596
rect 18564 20556 19524 20584
rect 18564 20544 18570 20556
rect 2774 20516 2780 20528
rect 2516 20488 2780 20516
rect 2774 20476 2780 20488
rect 2832 20476 2838 20528
rect 2869 20519 2927 20525
rect 2869 20485 2881 20519
rect 2915 20485 2927 20519
rect 2869 20479 2927 20485
rect 1394 20408 1400 20460
rect 1452 20408 1458 20460
rect 2317 20451 2375 20457
rect 2317 20448 2329 20451
rect 1504 20420 2329 20448
rect 1210 20340 1216 20392
rect 1268 20380 1274 20392
rect 1504 20380 1532 20420
rect 2317 20417 2329 20420
rect 2363 20417 2375 20451
rect 2884 20448 2912 20479
rect 3326 20476 3332 20528
rect 3384 20516 3390 20528
rect 3605 20519 3663 20525
rect 3605 20516 3617 20519
rect 3384 20488 3617 20516
rect 3384 20476 3390 20488
rect 3605 20485 3617 20488
rect 3651 20485 3663 20519
rect 3605 20479 3663 20485
rect 3973 20519 4031 20525
rect 3973 20485 3985 20519
rect 4019 20516 4031 20519
rect 4246 20516 4252 20528
rect 4019 20488 4252 20516
rect 4019 20485 4031 20488
rect 3973 20479 4031 20485
rect 4246 20476 4252 20488
rect 4304 20476 4310 20528
rect 4614 20476 4620 20528
rect 4672 20516 4678 20528
rect 5905 20519 5963 20525
rect 5905 20516 5917 20519
rect 4672 20488 5917 20516
rect 4672 20476 4678 20488
rect 5368 20460 5396 20488
rect 5905 20485 5917 20488
rect 5951 20485 5963 20519
rect 5905 20479 5963 20485
rect 6178 20476 6184 20528
rect 6236 20516 6242 20528
rect 9769 20519 9827 20525
rect 6236 20488 7602 20516
rect 6236 20476 6242 20488
rect 2958 20448 2964 20460
rect 2884 20420 2964 20448
rect 2317 20411 2375 20417
rect 2958 20408 2964 20420
rect 3016 20408 3022 20460
rect 3142 20408 3148 20460
rect 3200 20408 3206 20460
rect 3234 20408 3240 20460
rect 3292 20408 3298 20460
rect 4706 20408 4712 20460
rect 4764 20448 4770 20460
rect 4890 20448 4896 20460
rect 4764 20420 4896 20448
rect 4764 20408 4770 20420
rect 4890 20408 4896 20420
rect 4948 20448 4954 20460
rect 5077 20451 5135 20457
rect 5077 20448 5089 20451
rect 4948 20420 5089 20448
rect 4948 20408 4954 20420
rect 5077 20417 5089 20420
rect 5123 20417 5135 20451
rect 5077 20411 5135 20417
rect 5166 20408 5172 20460
rect 5224 20408 5230 20460
rect 5350 20408 5356 20460
rect 5408 20408 5414 20460
rect 5537 20451 5595 20457
rect 5537 20417 5549 20451
rect 5583 20448 5595 20451
rect 6638 20448 6644 20460
rect 5583 20420 6644 20448
rect 5583 20417 5595 20420
rect 5537 20411 5595 20417
rect 6638 20408 6644 20420
rect 6696 20448 6702 20460
rect 7466 20448 7472 20460
rect 6696 20420 7472 20448
rect 6696 20408 6702 20420
rect 7466 20408 7472 20420
rect 7524 20408 7530 20460
rect 7574 20448 7602 20488
rect 9769 20485 9781 20519
rect 9815 20516 9827 20519
rect 10410 20516 10416 20528
rect 9815 20488 10416 20516
rect 9815 20485 9827 20488
rect 9769 20479 9827 20485
rect 10410 20476 10416 20488
rect 10468 20476 10474 20528
rect 10502 20476 10508 20528
rect 10560 20516 10566 20528
rect 12452 20516 12480 20544
rect 10560 20488 11652 20516
rect 12452 20488 12756 20516
rect 10560 20476 10566 20488
rect 7803 20451 7861 20457
rect 7803 20448 7815 20451
rect 7574 20420 7815 20448
rect 7803 20417 7815 20420
rect 7849 20417 7861 20451
rect 7803 20411 7861 20417
rect 9030 20408 9036 20460
rect 9088 20448 9094 20460
rect 9582 20448 9588 20460
rect 9088 20420 9588 20448
rect 9088 20408 9094 20420
rect 9582 20408 9588 20420
rect 9640 20408 9646 20460
rect 9674 20408 9680 20460
rect 9732 20408 9738 20460
rect 10137 20451 10195 20457
rect 10137 20417 10149 20451
rect 10183 20448 10195 20451
rect 10962 20448 10968 20460
rect 10183 20420 10968 20448
rect 10183 20417 10195 20420
rect 10137 20411 10195 20417
rect 10962 20408 10968 20420
rect 11020 20408 11026 20460
rect 11624 20448 11652 20488
rect 12728 20457 12756 20488
rect 15286 20476 15292 20528
rect 15344 20516 15350 20528
rect 19444 20525 19472 20556
rect 19518 20544 19524 20556
rect 19576 20544 19582 20596
rect 22738 20544 22744 20596
rect 22796 20544 22802 20596
rect 23109 20587 23167 20593
rect 23109 20553 23121 20587
rect 23155 20584 23167 20587
rect 23566 20584 23572 20596
rect 23155 20556 23572 20584
rect 23155 20553 23167 20556
rect 23109 20547 23167 20553
rect 23566 20544 23572 20556
rect 23624 20544 23630 20596
rect 24305 20587 24363 20593
rect 24305 20553 24317 20587
rect 24351 20584 24363 20587
rect 24394 20584 24400 20596
rect 24351 20556 24400 20584
rect 24351 20553 24363 20556
rect 24305 20547 24363 20553
rect 24394 20544 24400 20556
rect 24452 20544 24458 20596
rect 19409 20519 19472 20525
rect 15344 20488 17322 20516
rect 15344 20476 15350 20488
rect 12713 20451 12771 20457
rect 11624 20420 12434 20448
rect 1268 20352 1532 20380
rect 1268 20340 1274 20352
rect 3050 20340 3056 20392
rect 3108 20340 3114 20392
rect 5442 20340 5448 20392
rect 5500 20340 5506 20392
rect 5902 20340 5908 20392
rect 5960 20380 5966 20392
rect 6730 20380 6736 20392
rect 5960 20352 6736 20380
rect 5960 20340 5966 20352
rect 6730 20340 6736 20352
rect 6788 20380 6794 20392
rect 7561 20383 7619 20389
rect 7561 20380 7573 20383
rect 6788 20352 7573 20380
rect 6788 20340 6794 20352
rect 7561 20349 7573 20352
rect 7607 20349 7619 20383
rect 12158 20380 12164 20392
rect 10442 20352 12164 20380
rect 7561 20343 7619 20349
rect 12158 20340 12164 20352
rect 12216 20340 12222 20392
rect 12406 20380 12434 20420
rect 12713 20417 12725 20451
rect 12759 20417 12771 20451
rect 12713 20411 12771 20417
rect 13998 20408 14004 20460
rect 14056 20408 14062 20460
rect 14366 20408 14372 20460
rect 14424 20448 14430 20460
rect 15010 20448 15016 20460
rect 14424 20420 15016 20448
rect 14424 20408 14430 20420
rect 15010 20408 15016 20420
rect 15068 20448 15074 20460
rect 17034 20448 17040 20460
rect 15068 20420 17040 20448
rect 15068 20408 15074 20420
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 17294 20457 17322 20488
rect 17696 20488 19380 20516
rect 17279 20451 17337 20457
rect 17279 20417 17291 20451
rect 17325 20417 17337 20451
rect 17279 20411 17337 20417
rect 13538 20380 13544 20392
rect 12406 20352 13544 20380
rect 13538 20340 13544 20352
rect 13596 20380 13602 20392
rect 14016 20380 14044 20408
rect 15286 20380 15292 20392
rect 13596 20352 14044 20380
rect 14476 20352 15292 20380
rect 13596 20340 13602 20352
rect 10962 20272 10968 20324
rect 11020 20312 11026 20324
rect 11974 20312 11980 20324
rect 11020 20284 11980 20312
rect 11020 20272 11026 20284
rect 11974 20272 11980 20284
rect 12032 20272 12038 20324
rect 12526 20272 12532 20324
rect 12584 20312 12590 20324
rect 14476 20312 14504 20352
rect 15286 20340 15292 20352
rect 15344 20340 15350 20392
rect 12584 20284 14504 20312
rect 12584 20272 12590 20284
rect 14550 20272 14556 20324
rect 14608 20312 14614 20324
rect 16942 20312 16948 20324
rect 14608 20284 16948 20312
rect 14608 20272 14614 20284
rect 16942 20272 16948 20284
rect 17000 20272 17006 20324
rect 4154 20204 4160 20256
rect 4212 20204 4218 20256
rect 6086 20204 6092 20256
rect 6144 20204 6150 20256
rect 6178 20204 6184 20256
rect 6236 20244 6242 20256
rect 7834 20244 7840 20256
rect 6236 20216 7840 20244
rect 6236 20204 6242 20216
rect 7834 20204 7840 20216
rect 7892 20204 7898 20256
rect 10686 20204 10692 20256
rect 10744 20204 10750 20256
rect 11514 20204 11520 20256
rect 11572 20244 11578 20256
rect 12710 20244 12716 20256
rect 11572 20216 12716 20244
rect 11572 20204 11578 20216
rect 12710 20204 12716 20216
rect 12768 20244 12774 20256
rect 17696 20244 17724 20488
rect 18506 20408 18512 20460
rect 18564 20408 18570 20460
rect 18598 20408 18604 20460
rect 18656 20408 18662 20460
rect 19153 20451 19211 20457
rect 19153 20417 19165 20451
rect 19199 20448 19211 20451
rect 19242 20448 19248 20460
rect 19199 20420 19248 20448
rect 19199 20417 19211 20420
rect 19153 20411 19211 20417
rect 19242 20408 19248 20420
rect 19300 20408 19306 20460
rect 19352 20448 19380 20488
rect 19409 20485 19421 20519
rect 19455 20488 19472 20519
rect 19536 20488 22094 20516
rect 19455 20485 19467 20488
rect 19409 20479 19467 20485
rect 19536 20448 19564 20488
rect 19352 20420 19564 20448
rect 19702 20408 19708 20460
rect 19760 20448 19766 20460
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 19760 20420 20637 20448
rect 19760 20408 19766 20420
rect 20625 20417 20637 20420
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 21085 20451 21143 20457
rect 21085 20417 21097 20451
rect 21131 20417 21143 20451
rect 21085 20411 21143 20417
rect 18785 20383 18843 20389
rect 18785 20349 18797 20383
rect 18831 20349 18843 20383
rect 21100 20380 21128 20411
rect 18785 20343 18843 20349
rect 20548 20352 21128 20380
rect 22066 20380 22094 20488
rect 22554 20408 22560 20460
rect 22612 20448 22618 20460
rect 22756 20448 22784 20544
rect 23750 20516 23756 20528
rect 23308 20488 23756 20516
rect 23308 20457 23336 20488
rect 23750 20476 23756 20488
rect 23808 20476 23814 20528
rect 23842 20476 23848 20528
rect 23900 20516 23906 20528
rect 24029 20519 24087 20525
rect 24029 20516 24041 20519
rect 23900 20488 24041 20516
rect 23900 20476 23906 20488
rect 24029 20485 24041 20488
rect 24075 20485 24087 20519
rect 24029 20479 24087 20485
rect 22833 20451 22891 20457
rect 22833 20448 22845 20451
rect 22612 20420 22845 20448
rect 22612 20408 22618 20420
rect 22833 20417 22845 20420
rect 22879 20417 22891 20451
rect 22833 20411 22891 20417
rect 23293 20451 23351 20457
rect 23293 20417 23305 20451
rect 23339 20417 23351 20451
rect 23293 20411 23351 20417
rect 23477 20451 23535 20457
rect 23477 20417 23489 20451
rect 23523 20448 23535 20451
rect 25866 20448 25872 20460
rect 23523 20420 25872 20448
rect 23523 20417 23535 20420
rect 23477 20411 23535 20417
rect 25866 20408 25872 20420
rect 25924 20408 25930 20460
rect 22066 20352 22876 20380
rect 18800 20312 18828 20343
rect 19058 20312 19064 20324
rect 18800 20284 19064 20312
rect 19058 20272 19064 20284
rect 19116 20272 19122 20324
rect 20548 20321 20576 20352
rect 20533 20315 20591 20321
rect 20533 20281 20545 20315
rect 20579 20281 20591 20315
rect 20533 20275 20591 20281
rect 22848 20256 22876 20352
rect 12768 20216 17724 20244
rect 18693 20247 18751 20253
rect 12768 20204 12774 20216
rect 18693 20213 18705 20247
rect 18739 20244 18751 20247
rect 20254 20244 20260 20256
rect 18739 20216 20260 20244
rect 18739 20213 18751 20216
rect 18693 20207 18751 20213
rect 20254 20204 20260 20216
rect 20312 20204 20318 20256
rect 20714 20204 20720 20256
rect 20772 20204 20778 20256
rect 20901 20247 20959 20253
rect 20901 20213 20913 20247
rect 20947 20244 20959 20247
rect 21358 20244 21364 20256
rect 20947 20216 21364 20244
rect 20947 20213 20959 20216
rect 20901 20207 20959 20213
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 22649 20247 22707 20253
rect 22649 20213 22661 20247
rect 22695 20244 22707 20247
rect 22738 20244 22744 20256
rect 22695 20216 22744 20244
rect 22695 20213 22707 20216
rect 22649 20207 22707 20213
rect 22738 20204 22744 20216
rect 22796 20204 22802 20256
rect 22830 20204 22836 20256
rect 22888 20204 22894 20256
rect 23750 20204 23756 20256
rect 23808 20204 23814 20256
rect 1104 20154 24840 20176
rect 1104 20102 3917 20154
rect 3969 20102 3981 20154
rect 4033 20102 4045 20154
rect 4097 20102 4109 20154
rect 4161 20102 4173 20154
rect 4225 20102 9851 20154
rect 9903 20102 9915 20154
rect 9967 20102 9979 20154
rect 10031 20102 10043 20154
rect 10095 20102 10107 20154
rect 10159 20102 15785 20154
rect 15837 20102 15849 20154
rect 15901 20102 15913 20154
rect 15965 20102 15977 20154
rect 16029 20102 16041 20154
rect 16093 20102 21719 20154
rect 21771 20102 21783 20154
rect 21835 20102 21847 20154
rect 21899 20102 21911 20154
rect 21963 20102 21975 20154
rect 22027 20102 24840 20154
rect 1104 20080 24840 20102
rect 1581 20043 1639 20049
rect 1581 20009 1593 20043
rect 1627 20040 1639 20043
rect 1762 20040 1768 20052
rect 1627 20012 1768 20040
rect 1627 20009 1639 20012
rect 1581 20003 1639 20009
rect 1762 20000 1768 20012
rect 1820 20000 1826 20052
rect 1946 20000 1952 20052
rect 2004 20040 2010 20052
rect 2004 20012 3464 20040
rect 2004 20000 2010 20012
rect 2682 19932 2688 19984
rect 2740 19932 2746 19984
rect 3436 19972 3464 20012
rect 3510 20000 3516 20052
rect 3568 20000 3574 20052
rect 5166 20000 5172 20052
rect 5224 20040 5230 20052
rect 6273 20043 6331 20049
rect 6273 20040 6285 20043
rect 5224 20012 6285 20040
rect 5224 20000 5230 20012
rect 6273 20009 6285 20012
rect 6319 20009 6331 20043
rect 6273 20003 6331 20009
rect 7558 20000 7564 20052
rect 7616 20040 7622 20052
rect 8018 20040 8024 20052
rect 7616 20012 8024 20040
rect 7616 20000 7622 20012
rect 8018 20000 8024 20012
rect 8076 20040 8082 20052
rect 8076 20012 10364 20040
rect 8076 20000 8082 20012
rect 4706 19972 4712 19984
rect 3436 19944 4712 19972
rect 4706 19932 4712 19944
rect 4764 19932 4770 19984
rect 2976 19876 3556 19904
rect 1397 19839 1455 19845
rect 1397 19805 1409 19839
rect 1443 19836 1455 19839
rect 1578 19836 1584 19848
rect 1443 19808 1584 19836
rect 1443 19805 1455 19808
rect 1397 19799 1455 19805
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 1670 19796 1676 19848
rect 1728 19796 1734 19848
rect 1947 19839 2005 19845
rect 1947 19805 1959 19839
rect 1993 19836 2005 19839
rect 2976 19836 3004 19876
rect 3528 19848 3556 19876
rect 4982 19864 4988 19916
rect 5040 19864 5046 19916
rect 9030 19864 9036 19916
rect 9088 19904 9094 19916
rect 9214 19904 9220 19916
rect 9088 19876 9220 19904
rect 9088 19864 9094 19876
rect 9214 19864 9220 19876
rect 9272 19904 9278 19916
rect 9398 19904 9404 19916
rect 9272 19876 9404 19904
rect 9272 19864 9278 19876
rect 9398 19864 9404 19876
rect 9456 19904 9462 19916
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 9456 19876 9689 19904
rect 9456 19864 9462 19876
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 9677 19867 9735 19873
rect 1993 19808 3004 19836
rect 3053 19839 3111 19845
rect 1993 19805 2005 19808
rect 1947 19799 2005 19805
rect 3053 19805 3065 19839
rect 3099 19805 3111 19839
rect 3053 19799 3111 19805
rect 1302 19728 1308 19780
rect 1360 19768 1366 19780
rect 3068 19768 3096 19799
rect 3326 19796 3332 19848
rect 3384 19796 3390 19848
rect 3510 19796 3516 19848
rect 3568 19796 3574 19848
rect 3786 19796 3792 19848
rect 3844 19796 3850 19848
rect 5000 19836 5028 19864
rect 5261 19839 5319 19845
rect 5261 19836 5273 19839
rect 5000 19808 5273 19836
rect 5261 19805 5273 19808
rect 5307 19805 5319 19839
rect 5261 19799 5319 19805
rect 5535 19839 5593 19845
rect 5535 19805 5547 19839
rect 5581 19836 5593 19839
rect 10336 19836 10364 20012
rect 10962 20000 10968 20052
rect 11020 20040 11026 20052
rect 11606 20040 11612 20052
rect 11020 20012 11612 20040
rect 11020 20000 11026 20012
rect 11606 20000 11612 20012
rect 11664 20000 11670 20052
rect 11974 20040 11980 20052
rect 11806 20012 11980 20040
rect 10689 19975 10747 19981
rect 10689 19941 10701 19975
rect 10735 19972 10747 19975
rect 11701 19975 11759 19981
rect 11701 19972 11713 19975
rect 10735 19944 11713 19972
rect 10735 19941 10747 19944
rect 10689 19935 10747 19941
rect 11701 19941 11713 19944
rect 11747 19941 11759 19975
rect 11701 19935 11759 19941
rect 11057 19907 11115 19913
rect 11057 19873 11069 19907
rect 11103 19904 11115 19907
rect 11146 19904 11152 19916
rect 11103 19876 11152 19904
rect 11103 19873 11115 19876
rect 11057 19867 11115 19873
rect 11146 19864 11152 19876
rect 11204 19864 11210 19916
rect 11241 19907 11299 19913
rect 11241 19873 11253 19907
rect 11287 19904 11299 19907
rect 11330 19904 11336 19916
rect 11287 19876 11336 19904
rect 11287 19873 11299 19876
rect 11241 19867 11299 19873
rect 11330 19864 11336 19876
rect 11388 19864 11394 19916
rect 11806 19904 11834 20012
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 12066 20000 12072 20052
rect 12124 20040 12130 20052
rect 14550 20040 14556 20052
rect 12124 20012 14556 20040
rect 12124 20000 12130 20012
rect 14550 20000 14556 20012
rect 14608 20000 14614 20052
rect 14734 20000 14740 20052
rect 14792 20040 14798 20052
rect 14792 20012 18368 20040
rect 14792 20000 14798 20012
rect 18340 19972 18368 20012
rect 18506 20000 18512 20052
rect 18564 20040 18570 20052
rect 18693 20043 18751 20049
rect 18693 20040 18705 20043
rect 18564 20012 18705 20040
rect 18564 20000 18570 20012
rect 18693 20009 18705 20012
rect 18739 20009 18751 20043
rect 18693 20003 18751 20009
rect 18340 19944 18552 19972
rect 12094 19907 12152 19913
rect 12094 19904 12106 19907
rect 11806 19876 12106 19904
rect 12094 19873 12106 19876
rect 12140 19873 12152 19907
rect 12094 19867 12152 19873
rect 14366 19864 14372 19916
rect 14424 19904 14430 19916
rect 14461 19907 14519 19913
rect 14461 19904 14473 19907
rect 14424 19876 14473 19904
rect 14424 19864 14430 19876
rect 14461 19873 14473 19876
rect 14507 19873 14519 19907
rect 14461 19867 14519 19873
rect 17034 19864 17040 19916
rect 17092 19904 17098 19916
rect 17681 19907 17739 19913
rect 17681 19904 17693 19907
rect 17092 19876 17693 19904
rect 17092 19864 17098 19876
rect 17681 19873 17693 19876
rect 17727 19873 17739 19907
rect 17681 19867 17739 19873
rect 5581 19808 5856 19836
rect 5581 19805 5593 19808
rect 5535 19799 5593 19805
rect 5350 19768 5356 19780
rect 1360 19740 3096 19768
rect 3160 19740 5356 19768
rect 1360 19728 1366 19740
rect 198 19660 204 19712
rect 256 19700 262 19712
rect 1578 19700 1584 19712
rect 256 19672 1584 19700
rect 256 19660 262 19672
rect 1578 19660 1584 19672
rect 1636 19660 1642 19712
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 3160 19700 3188 19740
rect 5350 19728 5356 19740
rect 5408 19728 5414 19780
rect 5828 19768 5856 19808
rect 7944 19808 9674 19836
rect 7650 19768 7656 19780
rect 5828 19740 7656 19768
rect 7650 19728 7656 19740
rect 7708 19768 7714 19780
rect 7944 19768 7972 19808
rect 7708 19740 7972 19768
rect 7708 19728 7714 19740
rect 8018 19728 8024 19780
rect 8076 19768 8082 19780
rect 9490 19768 9496 19780
rect 8076 19740 9496 19768
rect 8076 19728 8082 19740
rect 9490 19728 9496 19740
rect 9548 19728 9554 19780
rect 1728 19672 3188 19700
rect 3237 19703 3295 19709
rect 1728 19660 1734 19672
rect 3237 19669 3249 19703
rect 3283 19700 3295 19703
rect 3602 19700 3608 19712
rect 3283 19672 3608 19700
rect 3283 19669 3295 19672
rect 3237 19663 3295 19669
rect 3602 19660 3608 19672
rect 3660 19700 3666 19712
rect 3878 19700 3884 19712
rect 3660 19672 3884 19700
rect 3660 19660 3666 19672
rect 3878 19660 3884 19672
rect 3936 19660 3942 19712
rect 3973 19703 4031 19709
rect 3973 19669 3985 19703
rect 4019 19700 4031 19703
rect 8570 19700 8576 19712
rect 4019 19672 8576 19700
rect 4019 19669 4031 19672
rect 3973 19663 4031 19669
rect 8570 19660 8576 19672
rect 8628 19660 8634 19712
rect 8938 19660 8944 19712
rect 8996 19700 9002 19712
rect 9214 19700 9220 19712
rect 8996 19672 9220 19700
rect 8996 19660 9002 19672
rect 9214 19660 9220 19672
rect 9272 19660 9278 19712
rect 9646 19700 9674 19808
rect 9935 19809 9993 19815
rect 9935 19775 9947 19809
rect 9981 19806 9993 19809
rect 10336 19808 11192 19836
rect 9981 19780 9996 19806
rect 11164 19780 11192 19808
rect 11974 19796 11980 19848
rect 12032 19796 12038 19848
rect 12250 19796 12256 19848
rect 12308 19796 12314 19848
rect 13814 19796 13820 19848
rect 13872 19836 13878 19848
rect 13909 19839 13967 19845
rect 13909 19836 13921 19839
rect 13872 19808 13921 19836
rect 13872 19796 13878 19808
rect 13909 19805 13921 19808
rect 13955 19805 13967 19839
rect 14734 19836 14740 19848
rect 14695 19808 14740 19836
rect 13909 19799 13967 19805
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 16482 19836 16488 19848
rect 14844 19808 16488 19836
rect 9935 19769 9956 19775
rect 9950 19728 9956 19769
rect 10008 19768 10014 19780
rect 11054 19768 11060 19780
rect 10008 19740 11060 19768
rect 10008 19728 10014 19740
rect 11054 19728 11060 19740
rect 11112 19728 11118 19780
rect 11146 19728 11152 19780
rect 11204 19728 11210 19780
rect 13630 19728 13636 19780
rect 13688 19768 13694 19780
rect 14844 19768 14872 19808
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 17939 19809 17997 19815
rect 17939 19806 17951 19809
rect 13688 19740 14872 19768
rect 13688 19728 13694 19740
rect 14918 19728 14924 19780
rect 14976 19768 14982 19780
rect 17494 19768 17500 19780
rect 14976 19740 17500 19768
rect 14976 19728 14982 19740
rect 17494 19728 17500 19740
rect 17552 19768 17558 19780
rect 17938 19775 17951 19806
rect 17985 19775 17997 19809
rect 17938 19769 17997 19775
rect 17938 19768 17966 19769
rect 17552 19740 17966 19768
rect 18524 19768 18552 19944
rect 18708 19836 18736 20003
rect 19058 20000 19064 20052
rect 19116 20040 19122 20052
rect 19337 20043 19395 20049
rect 19337 20040 19349 20043
rect 19116 20012 19349 20040
rect 19116 20000 19122 20012
rect 19337 20009 19349 20012
rect 19383 20009 19395 20043
rect 19337 20003 19395 20009
rect 19886 20000 19892 20052
rect 19944 20040 19950 20052
rect 19944 20012 20668 20040
rect 19944 20000 19950 20012
rect 19904 19972 19932 20000
rect 19812 19944 19932 19972
rect 19812 19913 19840 19944
rect 19797 19907 19855 19913
rect 19797 19873 19809 19907
rect 19843 19873 19855 19907
rect 20640 19904 20668 20012
rect 20714 20000 20720 20052
rect 20772 20040 20778 20052
rect 21269 20043 21327 20049
rect 21269 20040 21281 20043
rect 20772 20012 21281 20040
rect 20772 20000 20778 20012
rect 21269 20009 21281 20012
rect 21315 20009 21327 20043
rect 21269 20003 21327 20009
rect 21358 20000 21364 20052
rect 21416 20000 21422 20052
rect 21542 20000 21548 20052
rect 21600 20040 21606 20052
rect 22005 20043 22063 20049
rect 22005 20040 22017 20043
rect 21600 20012 22017 20040
rect 21600 20000 21606 20012
rect 22005 20009 22017 20012
rect 22051 20009 22063 20043
rect 23842 20040 23848 20052
rect 22005 20003 22063 20009
rect 22204 20012 23848 20040
rect 20809 19975 20867 19981
rect 20809 19941 20821 19975
rect 20855 19941 20867 19975
rect 21376 19972 21404 20000
rect 22204 19972 22232 20012
rect 23842 20000 23848 20012
rect 23900 20000 23906 20052
rect 21376 19944 21772 19972
rect 20809 19935 20867 19941
rect 20714 19904 20720 19916
rect 20640 19876 20720 19904
rect 19797 19867 19855 19873
rect 20714 19864 20720 19876
rect 20772 19864 20778 19916
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 18708 19808 19257 19836
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 19426 19796 19432 19848
rect 19484 19796 19490 19848
rect 19610 19796 19616 19848
rect 19668 19796 19674 19848
rect 20824 19836 20852 19935
rect 21453 19907 21511 19913
rect 21453 19873 21465 19907
rect 21499 19904 21511 19907
rect 21637 19907 21695 19913
rect 21637 19904 21649 19907
rect 21499 19876 21649 19904
rect 21499 19873 21511 19876
rect 21453 19867 21511 19873
rect 21637 19873 21649 19876
rect 21683 19873 21695 19907
rect 21637 19867 21695 19873
rect 21744 19845 21772 19944
rect 22066 19944 22232 19972
rect 21177 19839 21235 19845
rect 21177 19836 21189 19839
rect 20055 19809 20113 19815
rect 19628 19768 19656 19796
rect 20055 19775 20067 19809
rect 20101 19806 20113 19809
rect 20824 19808 21189 19836
rect 20101 19775 20116 19806
rect 21177 19805 21189 19808
rect 21223 19836 21235 19839
rect 21545 19839 21603 19845
rect 21545 19836 21557 19839
rect 21223 19808 21557 19836
rect 21223 19805 21235 19808
rect 21177 19799 21235 19805
rect 21545 19805 21557 19808
rect 21591 19805 21603 19839
rect 21545 19799 21603 19805
rect 21729 19839 21787 19845
rect 21729 19805 21741 19839
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 21818 19796 21824 19848
rect 21876 19796 21882 19848
rect 20055 19769 20116 19775
rect 18524 19740 19656 19768
rect 20088 19768 20116 19769
rect 22066 19768 22094 19944
rect 22189 19839 22247 19845
rect 22189 19805 22201 19839
rect 22235 19836 22247 19839
rect 22278 19836 22284 19848
rect 22235 19808 22284 19836
rect 22235 19805 22247 19808
rect 22189 19799 22247 19805
rect 22278 19796 22284 19808
rect 22336 19836 22342 19848
rect 22336 19808 22692 19836
rect 22336 19796 22342 19808
rect 20088 19740 20208 19768
rect 17552 19728 17558 19740
rect 20180 19712 20208 19740
rect 21468 19740 22094 19768
rect 22456 19771 22514 19777
rect 12066 19700 12072 19712
rect 9646 19672 12072 19700
rect 12066 19660 12072 19672
rect 12124 19660 12130 19712
rect 12897 19703 12955 19709
rect 12897 19669 12909 19703
rect 12943 19700 12955 19703
rect 13170 19700 13176 19712
rect 12943 19672 13176 19700
rect 12943 19669 12955 19672
rect 12897 19663 12955 19669
rect 13170 19660 13176 19672
rect 13228 19660 13234 19712
rect 15470 19660 15476 19712
rect 15528 19660 15534 19712
rect 15746 19660 15752 19712
rect 15804 19700 15810 19712
rect 20070 19700 20076 19712
rect 15804 19672 20076 19700
rect 15804 19660 15810 19672
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 20162 19660 20168 19712
rect 20220 19660 20226 19712
rect 21468 19709 21496 19740
rect 22456 19737 22468 19771
rect 22502 19768 22514 19771
rect 22554 19768 22560 19780
rect 22502 19740 22560 19768
rect 22502 19737 22514 19740
rect 22456 19731 22514 19737
rect 22554 19728 22560 19740
rect 22612 19728 22618 19780
rect 22664 19712 22692 19808
rect 23290 19796 23296 19848
rect 23348 19836 23354 19848
rect 23845 19839 23903 19845
rect 23845 19836 23857 19839
rect 23348 19808 23857 19836
rect 23348 19796 23354 19808
rect 23845 19805 23857 19808
rect 23891 19805 23903 19839
rect 23845 19799 23903 19805
rect 24210 19728 24216 19780
rect 24268 19728 24274 19780
rect 21453 19703 21511 19709
rect 21453 19669 21465 19703
rect 21499 19669 21511 19703
rect 21453 19663 21511 19669
rect 22646 19660 22652 19712
rect 22704 19660 22710 19712
rect 23566 19660 23572 19712
rect 23624 19660 23630 19712
rect 1104 19610 25000 19632
rect 1104 19558 6884 19610
rect 6936 19558 6948 19610
rect 7000 19558 7012 19610
rect 7064 19558 7076 19610
rect 7128 19558 7140 19610
rect 7192 19558 12818 19610
rect 12870 19558 12882 19610
rect 12934 19558 12946 19610
rect 12998 19558 13010 19610
rect 13062 19558 13074 19610
rect 13126 19558 18752 19610
rect 18804 19558 18816 19610
rect 18868 19558 18880 19610
rect 18932 19558 18944 19610
rect 18996 19558 19008 19610
rect 19060 19558 24686 19610
rect 24738 19558 24750 19610
rect 24802 19558 24814 19610
rect 24866 19558 24878 19610
rect 24930 19558 24942 19610
rect 24994 19558 25000 19610
rect 1104 19536 25000 19558
rect 1302 19456 1308 19508
rect 1360 19496 1366 19508
rect 3786 19496 3792 19508
rect 1360 19468 3792 19496
rect 1360 19456 1366 19468
rect 3786 19456 3792 19468
rect 3844 19456 3850 19508
rect 3878 19456 3884 19508
rect 3936 19496 3942 19508
rect 6638 19496 6644 19508
rect 3936 19468 6644 19496
rect 3936 19456 3942 19468
rect 6638 19456 6644 19468
rect 6696 19456 6702 19508
rect 7558 19456 7564 19508
rect 7616 19456 7622 19508
rect 7650 19456 7656 19508
rect 7708 19456 7714 19508
rect 7742 19456 7748 19508
rect 7800 19496 7806 19508
rect 8481 19499 8539 19505
rect 8481 19496 8493 19499
rect 7800 19468 8493 19496
rect 7800 19456 7806 19468
rect 8481 19465 8493 19468
rect 8527 19465 8539 19499
rect 8481 19459 8539 19465
rect 9212 19456 9218 19508
rect 9270 19496 9276 19508
rect 9270 19468 9352 19496
rect 9270 19456 9276 19468
rect 3142 19428 3148 19440
rect 1412 19400 1808 19428
rect 1412 19369 1440 19400
rect 1780 19372 1808 19400
rect 2746 19400 3148 19428
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19329 1455 19363
rect 1397 19323 1455 19329
rect 1578 19320 1584 19372
rect 1636 19360 1642 19372
rect 1671 19363 1729 19369
rect 1671 19360 1683 19363
rect 1636 19332 1683 19360
rect 1636 19320 1642 19332
rect 1671 19329 1683 19332
rect 1717 19329 1729 19363
rect 1671 19323 1729 19329
rect 1762 19320 1768 19372
rect 1820 19320 1826 19372
rect 2746 19292 2774 19400
rect 3142 19388 3148 19400
rect 3200 19388 3206 19440
rect 7576 19428 7604 19456
rect 3252 19400 3832 19428
rect 2866 19320 2872 19372
rect 2924 19320 2930 19372
rect 3252 19360 3280 19400
rect 3068 19334 3280 19360
rect 2976 19332 3280 19334
rect 3419 19363 3477 19369
rect 2332 19264 2774 19292
rect 2976 19306 3096 19332
rect 3419 19329 3431 19363
rect 3465 19360 3477 19363
rect 3510 19360 3516 19372
rect 3465 19332 3516 19360
rect 3465 19329 3477 19332
rect 3419 19323 3477 19329
rect 3510 19320 3516 19332
rect 3568 19320 3574 19372
rect 2332 19168 2360 19264
rect 2314 19116 2320 19168
rect 2372 19116 2378 19168
rect 2406 19116 2412 19168
rect 2464 19116 2470 19168
rect 2976 19165 3004 19306
rect 3140 19295 3198 19301
rect 3140 19261 3152 19295
rect 3186 19261 3198 19295
rect 3140 19255 3198 19261
rect 3050 19184 3056 19236
rect 3108 19224 3114 19236
rect 3160 19224 3188 19255
rect 3108 19196 3188 19224
rect 3804 19224 3832 19400
rect 7484 19400 7604 19428
rect 5534 19252 5540 19304
rect 5592 19292 5598 19304
rect 7484 19301 7512 19400
rect 7668 19360 7696 19456
rect 7727 19363 7785 19369
rect 7727 19360 7739 19363
rect 7668 19332 7739 19360
rect 7727 19329 7739 19332
rect 7773 19329 7785 19363
rect 7727 19323 7785 19329
rect 8938 19320 8944 19372
rect 8996 19320 9002 19372
rect 9199 19363 9257 19369
rect 9199 19329 9211 19363
rect 9245 19360 9257 19363
rect 9324 19360 9352 19468
rect 9398 19456 9404 19508
rect 9456 19456 9462 19508
rect 9490 19456 9496 19508
rect 9548 19496 9554 19508
rect 9953 19499 10011 19505
rect 9548 19468 9674 19496
rect 9548 19456 9554 19468
rect 9245 19332 9352 19360
rect 9416 19360 9444 19456
rect 9646 19428 9674 19468
rect 9953 19465 9965 19499
rect 9999 19496 10011 19499
rect 12158 19496 12164 19508
rect 9999 19468 12164 19496
rect 9999 19465 10011 19468
rect 9953 19459 10011 19465
rect 12158 19456 12164 19468
rect 12216 19456 12222 19508
rect 12250 19456 12256 19508
rect 12308 19496 12314 19508
rect 12529 19499 12587 19505
rect 12529 19496 12541 19499
rect 12308 19468 12541 19496
rect 12308 19456 12314 19468
rect 12529 19465 12541 19468
rect 12575 19465 12587 19499
rect 12529 19459 12587 19465
rect 12894 19456 12900 19508
rect 12952 19496 12958 19508
rect 16850 19496 16856 19508
rect 12952 19468 16856 19496
rect 12952 19456 12958 19468
rect 9646 19400 11652 19428
rect 11514 19360 11520 19372
rect 9416 19332 11520 19360
rect 9245 19329 9257 19332
rect 9199 19323 9257 19329
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 11624 19360 11652 19400
rect 11775 19393 11833 19399
rect 11775 19390 11787 19393
rect 11774 19360 11787 19390
rect 11624 19359 11787 19360
rect 11821 19359 11833 19393
rect 12986 19388 12992 19440
rect 13044 19428 13050 19440
rect 13538 19428 13544 19440
rect 13044 19400 13544 19428
rect 13044 19388 13050 19400
rect 13538 19388 13544 19400
rect 13596 19388 13602 19440
rect 13722 19388 13728 19440
rect 13780 19388 13786 19440
rect 11624 19353 11833 19359
rect 11624 19332 11802 19353
rect 12526 19320 12532 19372
rect 12584 19360 12590 19372
rect 12710 19360 12716 19372
rect 12584 19332 12716 19360
rect 12584 19320 12590 19332
rect 12710 19320 12716 19332
rect 12768 19360 12774 19372
rect 12897 19363 12955 19369
rect 12897 19360 12909 19363
rect 12768 19332 12909 19360
rect 12768 19320 12774 19332
rect 12897 19329 12909 19332
rect 12943 19329 12955 19363
rect 12897 19323 12955 19329
rect 13171 19363 13229 19369
rect 13171 19329 13183 19363
rect 13217 19360 13229 19363
rect 13740 19360 13768 19388
rect 13217 19332 13768 19360
rect 14277 19363 14335 19369
rect 13217 19329 13229 19332
rect 13171 19323 13229 19329
rect 14277 19329 14289 19363
rect 14323 19360 14335 19363
rect 14323 19332 14412 19360
rect 14323 19329 14335 19332
rect 14277 19323 14335 19329
rect 7469 19295 7527 19301
rect 7469 19292 7481 19295
rect 5592 19264 7481 19292
rect 5592 19252 5598 19264
rect 7469 19261 7481 19264
rect 7515 19261 7527 19295
rect 7469 19255 7527 19261
rect 8846 19224 8852 19236
rect 3804 19196 7052 19224
rect 3108 19184 3114 19196
rect 2961 19159 3019 19165
rect 2961 19125 2973 19159
rect 3007 19125 3019 19159
rect 2961 19119 3019 19125
rect 3234 19116 3240 19168
rect 3292 19156 3298 19168
rect 4157 19159 4215 19165
rect 4157 19156 4169 19159
rect 3292 19128 4169 19156
rect 3292 19116 3298 19128
rect 4157 19125 4169 19128
rect 4203 19125 4215 19159
rect 7024 19156 7052 19196
rect 8128 19196 8852 19224
rect 8128 19156 8156 19196
rect 8846 19184 8852 19196
rect 8904 19184 8910 19236
rect 14384 19224 14412 19332
rect 14476 19301 14504 19468
rect 16850 19456 16856 19468
rect 16908 19456 16914 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 20864 19468 22692 19496
rect 20864 19456 20870 19468
rect 16482 19388 16488 19440
rect 16540 19428 16546 19440
rect 16540 19400 16954 19428
rect 16540 19388 16546 19400
rect 16926 19399 16954 19400
rect 16926 19393 16985 19399
rect 15470 19320 15476 19372
rect 15528 19320 15534 19372
rect 16926 19362 16939 19393
rect 16927 19359 16939 19362
rect 16973 19359 16985 19393
rect 16927 19353 16985 19359
rect 19610 19320 19616 19372
rect 19668 19360 19674 19372
rect 20438 19360 20444 19372
rect 19668 19332 20444 19360
rect 19668 19320 19674 19332
rect 20438 19320 20444 19332
rect 20496 19320 20502 19372
rect 21082 19320 21088 19372
rect 21140 19360 21146 19372
rect 21818 19360 21824 19372
rect 21140 19332 21824 19360
rect 21140 19320 21146 19332
rect 21818 19320 21824 19332
rect 21876 19320 21882 19372
rect 22370 19320 22376 19372
rect 22428 19360 22434 19372
rect 22465 19363 22523 19369
rect 22465 19360 22477 19363
rect 22428 19332 22477 19360
rect 22428 19320 22434 19332
rect 22465 19329 22477 19332
rect 22511 19329 22523 19363
rect 22664 19360 22692 19468
rect 24026 19388 24032 19440
rect 24084 19428 24090 19440
rect 24121 19431 24179 19437
rect 24121 19428 24133 19431
rect 24084 19400 24133 19428
rect 24084 19388 24090 19400
rect 24121 19397 24133 19400
rect 24167 19397 24179 19431
rect 24121 19391 24179 19397
rect 22739 19363 22797 19369
rect 22739 19360 22751 19363
rect 22664 19332 22751 19360
rect 22465 19323 22523 19329
rect 22739 19329 22751 19332
rect 22785 19360 22797 19363
rect 25866 19360 25872 19372
rect 22785 19332 25872 19360
rect 22785 19329 22797 19332
rect 22739 19323 22797 19329
rect 25866 19320 25872 19332
rect 25924 19320 25930 19372
rect 14461 19295 14519 19301
rect 14461 19261 14473 19295
rect 14507 19261 14519 19295
rect 14461 19255 14519 19261
rect 14826 19252 14832 19304
rect 14884 19252 14890 19304
rect 15194 19252 15200 19304
rect 15252 19252 15258 19304
rect 15286 19252 15292 19304
rect 15344 19301 15350 19304
rect 15344 19295 15372 19301
rect 15360 19261 15372 19295
rect 15344 19255 15372 19261
rect 15344 19252 15350 19255
rect 16666 19252 16672 19304
rect 16724 19252 16730 19304
rect 14844 19224 14872 19252
rect 13832 19196 14872 19224
rect 7024 19128 8156 19156
rect 4157 19119 4215 19125
rect 8570 19116 8576 19168
rect 8628 19156 8634 19168
rect 13832 19156 13860 19196
rect 14918 19184 14924 19236
rect 14976 19184 14982 19236
rect 15856 19196 16620 19224
rect 8628 19128 13860 19156
rect 13909 19159 13967 19165
rect 8628 19116 8634 19128
rect 13909 19125 13921 19159
rect 13955 19156 13967 19159
rect 13998 19156 14004 19168
rect 13955 19128 14004 19156
rect 13955 19125 13967 19128
rect 13909 19119 13967 19125
rect 13998 19116 14004 19128
rect 14056 19116 14062 19168
rect 14734 19116 14740 19168
rect 14792 19156 14798 19168
rect 15856 19156 15884 19196
rect 14792 19128 15884 19156
rect 14792 19116 14798 19128
rect 16114 19116 16120 19168
rect 16172 19116 16178 19168
rect 16482 19116 16488 19168
rect 16540 19116 16546 19168
rect 16592 19156 16620 19196
rect 17328 19196 18644 19224
rect 17328 19156 17356 19196
rect 18616 19168 18644 19196
rect 16592 19128 17356 19156
rect 17678 19116 17684 19168
rect 17736 19116 17742 19168
rect 18598 19116 18604 19168
rect 18656 19116 18662 19168
rect 23474 19116 23480 19168
rect 23532 19116 23538 19168
rect 24394 19116 24400 19168
rect 24452 19116 24458 19168
rect 1104 19066 24840 19088
rect 1104 19014 3917 19066
rect 3969 19014 3981 19066
rect 4033 19014 4045 19066
rect 4097 19014 4109 19066
rect 4161 19014 4173 19066
rect 4225 19014 9851 19066
rect 9903 19014 9915 19066
rect 9967 19014 9979 19066
rect 10031 19014 10043 19066
rect 10095 19014 10107 19066
rect 10159 19014 15785 19066
rect 15837 19014 15849 19066
rect 15901 19014 15913 19066
rect 15965 19014 15977 19066
rect 16029 19014 16041 19066
rect 16093 19014 21719 19066
rect 21771 19014 21783 19066
rect 21835 19014 21847 19066
rect 21899 19014 21911 19066
rect 21963 19014 21975 19066
rect 22027 19014 24840 19066
rect 1104 18992 24840 19014
rect 1486 18912 1492 18964
rect 1544 18952 1550 18964
rect 6638 18952 6644 18964
rect 1544 18924 6644 18952
rect 1544 18912 1550 18924
rect 6638 18912 6644 18924
rect 6696 18912 6702 18964
rect 8846 18912 8852 18964
rect 8904 18952 8910 18964
rect 10502 18952 10508 18964
rect 8904 18924 10508 18952
rect 8904 18912 8910 18924
rect 10502 18912 10508 18924
rect 10560 18912 10566 18964
rect 12360 18924 14872 18952
rect 1946 18844 1952 18896
rect 2004 18844 2010 18896
rect 6825 18887 6883 18893
rect 6825 18853 6837 18887
rect 6871 18853 6883 18887
rect 12360 18884 12388 18924
rect 6825 18847 6883 18853
rect 8496 18856 12388 18884
rect 934 18776 940 18828
rect 992 18816 998 18828
rect 2317 18819 2375 18825
rect 992 18788 1808 18816
rect 992 18776 998 18788
rect 750 18708 756 18760
rect 808 18748 814 18760
rect 1780 18757 1808 18788
rect 2317 18785 2329 18819
rect 2363 18785 2375 18819
rect 2317 18779 2375 18785
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 808 18720 1409 18748
rect 808 18708 814 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18717 1823 18751
rect 1765 18711 1823 18717
rect 1578 18572 1584 18624
rect 1636 18572 1642 18624
rect 2332 18612 2360 18779
rect 3694 18776 3700 18828
rect 3752 18816 3758 18828
rect 4249 18819 4307 18825
rect 4249 18816 4261 18819
rect 3752 18788 4261 18816
rect 3752 18776 3758 18788
rect 4249 18785 4261 18788
rect 4295 18785 4307 18819
rect 6840 18816 6868 18847
rect 6840 18788 7222 18816
rect 4249 18779 4307 18785
rect 4523 18751 4581 18757
rect 2575 18721 2633 18727
rect 2575 18687 2587 18721
rect 2621 18718 2633 18721
rect 2621 18692 2634 18718
rect 4523 18717 4535 18751
rect 4569 18748 4581 18751
rect 4614 18748 4620 18760
rect 4569 18720 4620 18748
rect 4569 18717 4581 18720
rect 4523 18711 4581 18717
rect 4614 18708 4620 18720
rect 4672 18708 4678 18760
rect 5534 18708 5540 18760
rect 5592 18748 5598 18760
rect 5813 18751 5871 18757
rect 5813 18748 5825 18751
rect 5592 18720 5825 18748
rect 5592 18708 5598 18720
rect 5813 18717 5825 18720
rect 5859 18717 5871 18751
rect 5813 18711 5871 18717
rect 6071 18721 6129 18727
rect 2575 18681 2596 18687
rect 2590 18640 2596 18681
rect 2648 18640 2654 18692
rect 3602 18680 3608 18692
rect 2700 18652 3608 18680
rect 2700 18612 2728 18652
rect 3602 18640 3608 18652
rect 3660 18640 3666 18692
rect 6071 18687 6083 18721
rect 6117 18718 6129 18721
rect 6117 18687 6130 18718
rect 7282 18708 7288 18760
rect 7340 18748 7346 18760
rect 7558 18748 7564 18760
rect 7340 18720 7564 18748
rect 7340 18708 7346 18720
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 7650 18708 7656 18760
rect 7708 18708 7714 18760
rect 7742 18708 7748 18760
rect 7800 18708 7806 18760
rect 8113 18751 8171 18757
rect 8113 18717 8125 18751
rect 8159 18748 8171 18751
rect 8202 18748 8208 18760
rect 8159 18720 8208 18748
rect 8159 18717 8171 18720
rect 8113 18711 8171 18717
rect 8202 18708 8208 18720
rect 8260 18748 8266 18760
rect 8496 18748 8524 18856
rect 9030 18776 9036 18828
rect 9088 18816 9094 18828
rect 10226 18816 10232 18828
rect 9088 18788 10232 18816
rect 9088 18776 9094 18788
rect 10226 18776 10232 18788
rect 10284 18776 10290 18828
rect 10962 18776 10968 18828
rect 11020 18816 11026 18828
rect 11020 18788 12158 18816
rect 11020 18776 11026 18788
rect 8260 18720 8524 18748
rect 8260 18708 8266 18720
rect 9582 18708 9588 18760
rect 9640 18748 9646 18760
rect 12130 18748 12158 18788
rect 12434 18776 12440 18828
rect 12492 18776 12498 18828
rect 14844 18816 14872 18924
rect 14918 18912 14924 18964
rect 14976 18952 14982 18964
rect 15105 18955 15163 18961
rect 15105 18952 15117 18955
rect 14976 18924 15117 18952
rect 14976 18912 14982 18924
rect 15105 18921 15117 18924
rect 15151 18921 15163 18955
rect 15105 18915 15163 18921
rect 15470 18912 15476 18964
rect 15528 18952 15534 18964
rect 16390 18952 16396 18964
rect 15528 18924 16396 18952
rect 15528 18912 15534 18924
rect 16390 18912 16396 18924
rect 16448 18912 16454 18964
rect 16482 18912 16488 18964
rect 16540 18912 16546 18964
rect 20990 18912 20996 18964
rect 21048 18952 21054 18964
rect 21048 18924 24256 18952
rect 21048 18912 21054 18924
rect 15286 18816 15292 18828
rect 14844 18788 15292 18816
rect 15286 18776 15292 18788
rect 15344 18816 15350 18828
rect 15749 18819 15807 18825
rect 15749 18816 15761 18819
rect 15344 18788 15761 18816
rect 15344 18776 15350 18788
rect 15749 18785 15761 18788
rect 15795 18785 15807 18819
rect 15749 18779 15807 18785
rect 16390 18776 16396 18828
rect 16448 18776 16454 18828
rect 16500 18816 16528 18912
rect 20533 18887 20591 18893
rect 20533 18853 20545 18887
rect 20579 18853 20591 18887
rect 20533 18847 20591 18853
rect 22925 18887 22983 18893
rect 22925 18853 22937 18887
rect 22971 18884 22983 18887
rect 23477 18887 23535 18893
rect 23477 18884 23489 18887
rect 22971 18856 23489 18884
rect 22971 18853 22983 18856
rect 22925 18847 22983 18853
rect 23477 18853 23489 18856
rect 23523 18853 23535 18887
rect 23477 18847 23535 18853
rect 16669 18819 16727 18825
rect 16669 18816 16681 18819
rect 16500 18788 16681 18816
rect 16669 18785 16681 18788
rect 16715 18785 16727 18819
rect 16669 18779 16727 18785
rect 16945 18819 17003 18825
rect 16945 18785 16957 18819
rect 16991 18816 17003 18819
rect 17678 18816 17684 18828
rect 16991 18788 17684 18816
rect 16991 18785 17003 18788
rect 16945 18779 17003 18785
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 20548 18816 20576 18847
rect 20548 18788 21312 18816
rect 12679 18751 12737 18757
rect 12679 18748 12691 18751
rect 9640 18720 11928 18748
rect 12130 18720 12691 18748
rect 9640 18708 9646 18720
rect 6071 18681 6130 18687
rect 6102 18680 6130 18681
rect 11054 18680 11060 18692
rect 6102 18652 6224 18680
rect 6196 18624 6224 18652
rect 8404 18652 11060 18680
rect 2332 18584 2728 18612
rect 2774 18572 2780 18624
rect 2832 18612 2838 18624
rect 3329 18615 3387 18621
rect 3329 18612 3341 18615
rect 2832 18584 3341 18612
rect 2832 18572 2838 18584
rect 3329 18581 3341 18584
rect 3375 18581 3387 18615
rect 3329 18575 3387 18581
rect 4338 18572 4344 18624
rect 4396 18612 4402 18624
rect 4982 18612 4988 18624
rect 4396 18584 4988 18612
rect 4396 18572 4402 18584
rect 4982 18572 4988 18584
rect 5040 18572 5046 18624
rect 5166 18572 5172 18624
rect 5224 18612 5230 18624
rect 5261 18615 5319 18621
rect 5261 18612 5273 18615
rect 5224 18584 5273 18612
rect 5224 18572 5230 18584
rect 5261 18581 5273 18584
rect 5307 18581 5319 18615
rect 5261 18575 5319 18581
rect 6178 18572 6184 18624
rect 6236 18572 6242 18624
rect 7377 18615 7435 18621
rect 7377 18581 7389 18615
rect 7423 18612 7435 18615
rect 8404 18612 8432 18652
rect 11054 18640 11060 18652
rect 11112 18640 11118 18692
rect 11900 18680 11928 18720
rect 12544 18692 12572 18720
rect 12679 18717 12691 18720
rect 12725 18717 12737 18751
rect 12679 18711 12737 18717
rect 14093 18751 14151 18757
rect 14093 18717 14105 18751
rect 14139 18717 14151 18751
rect 14093 18711 14151 18717
rect 14367 18751 14425 18757
rect 14367 18717 14379 18751
rect 14413 18748 14425 18751
rect 14734 18748 14740 18760
rect 14413 18720 14740 18748
rect 14413 18717 14425 18720
rect 14367 18711 14425 18717
rect 12066 18680 12072 18692
rect 11900 18652 12072 18680
rect 12066 18640 12072 18652
rect 12124 18640 12130 18692
rect 12526 18640 12532 18692
rect 12584 18640 12590 18692
rect 12894 18640 12900 18692
rect 12952 18640 12958 18692
rect 12986 18640 12992 18692
rect 13044 18680 13050 18692
rect 13722 18680 13728 18692
rect 13044 18652 13728 18680
rect 13044 18640 13050 18652
rect 13722 18640 13728 18652
rect 13780 18640 13786 18692
rect 14108 18680 14136 18711
rect 14734 18708 14740 18720
rect 14792 18708 14798 18760
rect 14826 18708 14832 18760
rect 14884 18748 14890 18760
rect 16850 18757 16856 18760
rect 15933 18751 15991 18757
rect 15933 18748 15945 18751
rect 14884 18720 15945 18748
rect 14884 18708 14890 18720
rect 15933 18717 15945 18720
rect 15979 18717 15991 18751
rect 15933 18711 15991 18717
rect 16807 18751 16856 18757
rect 16807 18717 16819 18751
rect 16853 18717 16856 18751
rect 16807 18711 16856 18717
rect 16850 18708 16856 18711
rect 16908 18708 16914 18760
rect 19610 18708 19616 18760
rect 19668 18708 19674 18760
rect 19794 18708 19800 18760
rect 19852 18708 19858 18760
rect 21284 18757 21312 18788
rect 23658 18776 23664 18828
rect 23716 18776 23722 18828
rect 20717 18751 20775 18757
rect 20717 18717 20729 18751
rect 20763 18717 20775 18751
rect 20717 18711 20775 18717
rect 21269 18751 21327 18757
rect 21269 18717 21281 18751
rect 21315 18717 21327 18751
rect 21269 18711 21327 18717
rect 14108 18652 14412 18680
rect 7423 18584 8432 18612
rect 8481 18615 8539 18621
rect 7423 18581 7435 18584
rect 7377 18575 7435 18581
rect 8481 18581 8493 18615
rect 8527 18612 8539 18615
rect 8570 18612 8576 18624
rect 8527 18584 8576 18612
rect 8527 18581 8539 18584
rect 8481 18575 8539 18581
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 8662 18572 8668 18624
rect 8720 18572 8726 18624
rect 9674 18572 9680 18624
rect 9732 18612 9738 18624
rect 11974 18612 11980 18624
rect 9732 18584 11980 18612
rect 9732 18572 9738 18584
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12434 18572 12440 18624
rect 12492 18612 12498 18624
rect 12912 18612 12940 18640
rect 14384 18624 14412 18652
rect 17678 18640 17684 18692
rect 17736 18680 17742 18692
rect 20346 18680 20352 18692
rect 17736 18652 20352 18680
rect 17736 18640 17742 18652
rect 20346 18640 20352 18652
rect 20404 18680 20410 18692
rect 20732 18680 20760 18711
rect 22738 18708 22744 18760
rect 22796 18748 22802 18760
rect 22833 18751 22891 18757
rect 22833 18748 22845 18751
rect 22796 18720 22845 18748
rect 22796 18708 22802 18720
rect 22833 18717 22845 18720
rect 22879 18717 22891 18751
rect 22833 18711 22891 18717
rect 23293 18751 23351 18757
rect 23293 18717 23305 18751
rect 23339 18717 23351 18751
rect 23293 18711 23351 18717
rect 23385 18751 23443 18757
rect 23385 18717 23397 18751
rect 23431 18748 23443 18751
rect 23474 18748 23480 18760
rect 23431 18720 23480 18748
rect 23431 18717 23443 18720
rect 23385 18711 23443 18717
rect 20404 18652 20760 18680
rect 23308 18680 23336 18711
rect 23474 18708 23480 18720
rect 23532 18708 23538 18760
rect 23566 18708 23572 18760
rect 23624 18708 23630 18760
rect 23845 18751 23903 18757
rect 23845 18717 23857 18751
rect 23891 18748 23903 18751
rect 24118 18748 24124 18760
rect 23891 18720 24124 18748
rect 23891 18717 23903 18720
rect 23845 18711 23903 18717
rect 24118 18708 24124 18720
rect 24176 18708 24182 18760
rect 23584 18680 23612 18708
rect 23308 18652 23612 18680
rect 20404 18640 20410 18652
rect 24228 18624 24256 18924
rect 12492 18584 12940 18612
rect 12492 18572 12498 18584
rect 13446 18572 13452 18624
rect 13504 18572 13510 18624
rect 14366 18572 14372 18624
rect 14424 18572 14430 18624
rect 15010 18572 15016 18624
rect 15068 18612 15074 18624
rect 16666 18612 16672 18624
rect 15068 18584 16672 18612
rect 15068 18572 15074 18584
rect 16666 18572 16672 18584
rect 16724 18612 16730 18624
rect 17494 18612 17500 18624
rect 16724 18584 17500 18612
rect 16724 18572 16730 18584
rect 17494 18572 17500 18584
rect 17552 18572 17558 18624
rect 17589 18615 17647 18621
rect 17589 18581 17601 18615
rect 17635 18612 17647 18615
rect 18046 18612 18052 18624
rect 17635 18584 18052 18612
rect 17635 18581 17647 18584
rect 17589 18575 17647 18581
rect 18046 18572 18052 18584
rect 18104 18572 18110 18624
rect 19702 18572 19708 18624
rect 19760 18572 19766 18624
rect 21361 18615 21419 18621
rect 21361 18581 21373 18615
rect 21407 18612 21419 18615
rect 21910 18612 21916 18624
rect 21407 18584 21916 18612
rect 21407 18581 21419 18584
rect 21361 18575 21419 18581
rect 21910 18572 21916 18584
rect 21968 18572 21974 18624
rect 23109 18615 23167 18621
rect 23109 18581 23121 18615
rect 23155 18612 23167 18615
rect 23474 18612 23480 18624
rect 23155 18584 23480 18612
rect 23155 18581 23167 18584
rect 23109 18575 23167 18581
rect 23474 18572 23480 18584
rect 23532 18572 23538 18624
rect 23566 18572 23572 18624
rect 23624 18612 23630 18624
rect 23661 18615 23719 18621
rect 23661 18612 23673 18615
rect 23624 18584 23673 18612
rect 23624 18572 23630 18584
rect 23661 18581 23673 18584
rect 23707 18581 23719 18615
rect 23661 18575 23719 18581
rect 24118 18572 24124 18624
rect 24176 18572 24182 18624
rect 24210 18572 24216 18624
rect 24268 18572 24274 18624
rect 1104 18522 25000 18544
rect 1104 18470 6884 18522
rect 6936 18470 6948 18522
rect 7000 18470 7012 18522
rect 7064 18470 7076 18522
rect 7128 18470 7140 18522
rect 7192 18470 12818 18522
rect 12870 18470 12882 18522
rect 12934 18470 12946 18522
rect 12998 18470 13010 18522
rect 13062 18470 13074 18522
rect 13126 18470 18752 18522
rect 18804 18470 18816 18522
rect 18868 18470 18880 18522
rect 18932 18470 18944 18522
rect 18996 18470 19008 18522
rect 19060 18470 24686 18522
rect 24738 18470 24750 18522
rect 24802 18470 24814 18522
rect 24866 18470 24878 18522
rect 24930 18470 24942 18522
rect 24994 18470 25000 18522
rect 1104 18448 25000 18470
rect 3510 18368 3516 18420
rect 3568 18408 3574 18420
rect 5813 18411 5871 18417
rect 5813 18408 5825 18411
rect 3568 18380 5825 18408
rect 3568 18368 3574 18380
rect 5813 18377 5825 18380
rect 5859 18377 5871 18411
rect 5813 18371 5871 18377
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 6546 18408 6552 18420
rect 5960 18380 6552 18408
rect 5960 18368 5966 18380
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 6730 18368 6736 18420
rect 6788 18408 6794 18420
rect 7837 18411 7895 18417
rect 6788 18380 7788 18408
rect 6788 18368 6794 18380
rect 750 18300 756 18352
rect 808 18340 814 18352
rect 1489 18343 1547 18349
rect 1489 18340 1501 18343
rect 808 18312 1501 18340
rect 808 18300 814 18312
rect 1489 18309 1501 18312
rect 1535 18309 1547 18343
rect 1489 18303 1547 18309
rect 1670 18300 1676 18352
rect 1728 18300 1734 18352
rect 2222 18340 2228 18352
rect 2056 18312 2228 18340
rect 1854 18232 1860 18284
rect 1912 18232 1918 18284
rect 1946 18232 1952 18284
rect 2004 18232 2010 18284
rect 1872 18136 1900 18232
rect 2056 18213 2084 18312
rect 2222 18300 2228 18312
rect 2280 18300 2286 18352
rect 6196 18312 6500 18340
rect 3234 18232 3240 18284
rect 3292 18232 3298 18284
rect 4338 18272 4344 18284
rect 3896 18244 4344 18272
rect 2041 18207 2099 18213
rect 2041 18173 2053 18207
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 2225 18207 2283 18213
rect 2225 18173 2237 18207
rect 2271 18204 2283 18207
rect 2314 18204 2320 18216
rect 2271 18176 2320 18204
rect 2271 18173 2283 18176
rect 2225 18167 2283 18173
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 2961 18207 3019 18213
rect 2961 18204 2973 18207
rect 2608 18176 2973 18204
rect 2608 18136 2636 18176
rect 2961 18173 2973 18176
rect 3007 18173 3019 18207
rect 2961 18167 3019 18173
rect 3099 18207 3157 18213
rect 3099 18173 3111 18207
rect 3145 18204 3157 18207
rect 3786 18204 3792 18216
rect 3145 18176 3792 18204
rect 3145 18173 3157 18176
rect 3099 18167 3157 18173
rect 3786 18164 3792 18176
rect 3844 18204 3850 18216
rect 3896 18204 3924 18244
rect 4338 18232 4344 18244
rect 4396 18232 4402 18284
rect 4982 18232 4988 18284
rect 5040 18281 5046 18284
rect 5040 18275 5068 18281
rect 5056 18241 5068 18275
rect 5040 18235 5068 18241
rect 5040 18232 5046 18235
rect 5166 18232 5172 18284
rect 5224 18232 5230 18284
rect 6196 18281 6224 18312
rect 6181 18275 6239 18281
rect 6181 18241 6193 18275
rect 6227 18241 6239 18275
rect 6472 18272 6500 18312
rect 6638 18300 6644 18352
rect 6696 18340 6702 18352
rect 6696 18312 7420 18340
rect 6696 18300 6702 18312
rect 6825 18275 6883 18281
rect 6825 18272 6837 18275
rect 6472 18244 6837 18272
rect 6181 18235 6239 18241
rect 6825 18241 6837 18244
rect 6871 18241 6883 18275
rect 6825 18235 6883 18241
rect 6914 18232 6920 18284
rect 6972 18232 6978 18284
rect 7282 18232 7288 18284
rect 7340 18232 7346 18284
rect 7392 18272 7420 18312
rect 7466 18300 7472 18352
rect 7524 18340 7530 18352
rect 7653 18343 7711 18349
rect 7653 18340 7665 18343
rect 7524 18312 7665 18340
rect 7524 18300 7530 18312
rect 7653 18309 7665 18312
rect 7699 18309 7711 18343
rect 7760 18340 7788 18380
rect 7837 18377 7849 18411
rect 7883 18408 7895 18411
rect 9677 18411 9735 18417
rect 7883 18380 9628 18408
rect 7883 18377 7895 18380
rect 7837 18371 7895 18377
rect 7760 18312 9352 18340
rect 7653 18303 7711 18309
rect 8939 18275 8997 18281
rect 7392 18244 7696 18272
rect 3844 18176 3924 18204
rect 3973 18207 4031 18213
rect 3844 18164 3850 18176
rect 3973 18173 3985 18207
rect 4019 18173 4031 18207
rect 3973 18167 4031 18173
rect 1872 18108 2636 18136
rect 2685 18139 2743 18145
rect 2685 18105 2697 18139
rect 2731 18136 2743 18139
rect 2774 18136 2780 18148
rect 2731 18108 2780 18136
rect 2731 18105 2743 18108
rect 2685 18099 2743 18105
rect 2774 18096 2780 18108
rect 2832 18096 2838 18148
rect 1765 18071 1823 18077
rect 1765 18037 1777 18071
rect 1811 18068 1823 18071
rect 3050 18068 3056 18080
rect 1811 18040 3056 18068
rect 1811 18037 1823 18040
rect 1765 18031 1823 18037
rect 3050 18028 3056 18040
rect 3108 18028 3114 18080
rect 3326 18028 3332 18080
rect 3384 18068 3390 18080
rect 3881 18071 3939 18077
rect 3881 18068 3893 18071
rect 3384 18040 3893 18068
rect 3384 18028 3390 18040
rect 3881 18037 3893 18040
rect 3927 18037 3939 18071
rect 3988 18068 4016 18167
rect 4154 18164 4160 18216
rect 4212 18164 4218 18216
rect 4522 18164 4528 18216
rect 4580 18204 4586 18216
rect 4617 18207 4675 18213
rect 4617 18204 4629 18207
rect 4580 18176 4629 18204
rect 4580 18164 4586 18176
rect 4617 18173 4629 18176
rect 4663 18173 4675 18207
rect 4617 18167 4675 18173
rect 4893 18207 4951 18213
rect 4893 18173 4905 18207
rect 4939 18204 4951 18207
rect 4939 18176 6316 18204
rect 4939 18173 4951 18176
rect 4893 18167 4951 18173
rect 6288 18136 6316 18176
rect 6730 18164 6736 18216
rect 6788 18164 6794 18216
rect 7668 18136 7696 18244
rect 8939 18241 8951 18275
rect 8985 18272 8997 18275
rect 9030 18272 9036 18284
rect 8985 18244 9036 18272
rect 8985 18241 8997 18244
rect 8939 18235 8997 18241
rect 9030 18232 9036 18244
rect 9088 18232 9094 18284
rect 7742 18164 7748 18216
rect 7800 18204 7806 18216
rect 8665 18207 8723 18213
rect 8665 18204 8677 18207
rect 7800 18176 8677 18204
rect 7800 18164 7806 18176
rect 8665 18173 8677 18176
rect 8711 18173 8723 18207
rect 8665 18167 8723 18173
rect 9324 18136 9352 18312
rect 9600 18204 9628 18380
rect 9677 18377 9689 18411
rect 9723 18377 9735 18411
rect 9677 18371 9735 18377
rect 9692 18284 9720 18371
rect 10226 18368 10232 18420
rect 10284 18408 10290 18420
rect 10594 18408 10600 18420
rect 10284 18380 10600 18408
rect 10284 18368 10290 18380
rect 10594 18368 10600 18380
rect 10652 18368 10658 18420
rect 13722 18408 13728 18420
rect 13002 18380 13728 18408
rect 11974 18300 11980 18352
rect 12032 18340 12038 18352
rect 12894 18340 12900 18352
rect 12032 18312 12900 18340
rect 12032 18300 12038 18312
rect 12894 18300 12900 18312
rect 12952 18300 12958 18352
rect 13002 18340 13030 18380
rect 13722 18368 13728 18380
rect 13780 18368 13786 18420
rect 15470 18368 15476 18420
rect 15528 18368 15534 18420
rect 16209 18411 16267 18417
rect 16209 18377 16221 18411
rect 16255 18408 16267 18411
rect 16390 18408 16396 18420
rect 16255 18380 16396 18408
rect 16255 18377 16267 18380
rect 16209 18371 16267 18377
rect 16390 18368 16396 18380
rect 16448 18368 16454 18420
rect 19337 18411 19395 18417
rect 19337 18377 19349 18411
rect 19383 18408 19395 18411
rect 19705 18411 19763 18417
rect 19383 18380 19656 18408
rect 19383 18377 19395 18380
rect 19337 18371 19395 18377
rect 13002 18312 13032 18340
rect 9674 18232 9680 18284
rect 9732 18232 9738 18284
rect 10594 18232 10600 18284
rect 10652 18232 10658 18284
rect 10962 18272 10968 18284
rect 10704 18244 10968 18272
rect 10704 18204 10732 18244
rect 10962 18232 10968 18244
rect 11020 18232 11026 18284
rect 11054 18232 11060 18284
rect 11112 18272 11118 18284
rect 12250 18272 12256 18284
rect 11112 18244 12256 18272
rect 11112 18232 11118 18244
rect 12250 18232 12256 18244
rect 12308 18272 12314 18284
rect 12618 18272 12624 18284
rect 12308 18244 12624 18272
rect 12308 18232 12314 18244
rect 12618 18232 12624 18244
rect 12676 18272 12682 18284
rect 12805 18276 12863 18281
rect 12728 18275 12863 18276
rect 12728 18272 12817 18275
rect 12676 18248 12817 18272
rect 12676 18244 12756 18248
rect 12676 18232 12682 18244
rect 12805 18241 12817 18248
rect 12851 18241 12863 18275
rect 12805 18235 12863 18241
rect 9600 18176 10732 18204
rect 12912 18204 12940 18300
rect 13004 18281 13032 18312
rect 15470 18311 15498 18368
rect 17972 18312 19380 18340
rect 15455 18305 15513 18311
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 13722 18232 13728 18284
rect 13780 18232 13786 18284
rect 13998 18232 14004 18284
rect 14056 18232 14062 18284
rect 15010 18232 15016 18284
rect 15068 18272 15074 18284
rect 15197 18275 15255 18281
rect 15197 18272 15209 18275
rect 15068 18244 15209 18272
rect 15068 18232 15074 18244
rect 15197 18241 15209 18244
rect 15243 18241 15255 18275
rect 15455 18271 15467 18305
rect 15501 18271 15513 18305
rect 17972 18281 18000 18312
rect 19352 18284 19380 18312
rect 15455 18265 15513 18271
rect 17957 18275 18015 18281
rect 15197 18235 15255 18241
rect 17957 18241 17969 18275
rect 18003 18241 18015 18275
rect 17957 18235 18015 18241
rect 18046 18232 18052 18284
rect 18104 18272 18110 18284
rect 18213 18275 18271 18281
rect 18213 18272 18225 18275
rect 18104 18244 18225 18272
rect 18104 18232 18110 18244
rect 18213 18241 18225 18244
rect 18259 18241 18271 18275
rect 18213 18235 18271 18241
rect 19334 18232 19340 18284
rect 19392 18232 19398 18284
rect 19426 18232 19432 18284
rect 19484 18232 19490 18284
rect 19628 18272 19656 18380
rect 19705 18377 19717 18411
rect 19751 18408 19763 18411
rect 19794 18408 19800 18420
rect 19751 18380 19800 18408
rect 19751 18377 19763 18380
rect 19705 18371 19763 18377
rect 19794 18368 19800 18380
rect 19852 18368 19858 18420
rect 22278 18368 22284 18420
rect 22336 18408 22342 18420
rect 22336 18380 22508 18408
rect 22336 18368 22342 18380
rect 20346 18349 20352 18352
rect 20329 18343 20352 18349
rect 20329 18309 20341 18343
rect 20329 18303 20352 18309
rect 20346 18300 20352 18303
rect 20404 18300 20410 18352
rect 22094 18300 22100 18352
rect 22152 18300 22158 18352
rect 19889 18275 19947 18281
rect 19889 18272 19901 18275
rect 19628 18244 19901 18272
rect 19889 18241 19901 18244
rect 19935 18241 19947 18275
rect 19889 18235 19947 18241
rect 21634 18232 21640 18284
rect 21692 18272 21698 18284
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 21692 18244 21833 18272
rect 21692 18232 21698 18244
rect 21821 18241 21833 18244
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 21910 18232 21916 18284
rect 21968 18232 21974 18284
rect 22480 18281 22508 18380
rect 23382 18368 23388 18420
rect 23440 18368 23446 18420
rect 23474 18368 23480 18420
rect 23532 18368 23538 18420
rect 23569 18411 23627 18417
rect 23569 18377 23581 18411
rect 23615 18408 23627 18411
rect 23658 18408 23664 18420
rect 23615 18380 23664 18408
rect 23615 18377 23627 18380
rect 23569 18371 23627 18377
rect 23658 18368 23664 18380
rect 23716 18368 23722 18420
rect 24394 18368 24400 18420
rect 24452 18368 24458 18420
rect 22756 18312 23336 18340
rect 22373 18275 22431 18281
rect 22373 18272 22385 18275
rect 22020 18244 22385 18272
rect 12912 18176 13400 18204
rect 12434 18136 12440 18148
rect 6288 18108 6408 18136
rect 7668 18108 7788 18136
rect 9324 18108 12440 18136
rect 6380 18080 6408 18108
rect 4890 18068 4896 18080
rect 3988 18040 4896 18068
rect 3881 18031 3939 18037
rect 4890 18028 4896 18040
rect 4948 18068 4954 18080
rect 5258 18068 5264 18080
rect 4948 18040 5264 18068
rect 4948 18028 4954 18040
rect 5258 18028 5264 18040
rect 5316 18028 5322 18080
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 5902 18068 5908 18080
rect 5592 18040 5908 18068
rect 5592 18028 5598 18040
rect 5902 18028 5908 18040
rect 5960 18028 5966 18080
rect 6362 18028 6368 18080
rect 6420 18028 6426 18080
rect 7760 18068 7788 18108
rect 12434 18096 12440 18108
rect 12492 18096 12498 18148
rect 13372 18136 13400 18176
rect 13446 18164 13452 18216
rect 13504 18164 13510 18216
rect 13842 18207 13900 18213
rect 13842 18204 13854 18207
rect 13556 18176 13854 18204
rect 13556 18136 13584 18176
rect 13842 18173 13854 18176
rect 13888 18173 13900 18207
rect 19352 18204 19380 18232
rect 20073 18207 20131 18213
rect 20073 18204 20085 18207
rect 19352 18176 20085 18204
rect 13842 18167 13900 18173
rect 20073 18173 20085 18176
rect 20119 18173 20131 18207
rect 22020 18204 22048 18244
rect 22373 18241 22385 18244
rect 22419 18241 22431 18275
rect 22373 18235 22431 18241
rect 22465 18275 22523 18281
rect 22465 18241 22477 18275
rect 22511 18241 22523 18275
rect 22465 18235 22523 18241
rect 22649 18275 22707 18281
rect 22649 18241 22661 18275
rect 22695 18241 22707 18275
rect 22649 18235 22707 18241
rect 20073 18167 20131 18173
rect 21468 18176 22048 18204
rect 22097 18207 22155 18213
rect 13372 18108 13584 18136
rect 14642 18096 14648 18148
rect 14700 18096 14706 18148
rect 17954 18136 17960 18148
rect 15856 18108 17960 18136
rect 10413 18071 10471 18077
rect 10413 18068 10425 18071
rect 7760 18040 10425 18068
rect 10413 18037 10425 18040
rect 10459 18037 10471 18071
rect 10413 18031 10471 18037
rect 10962 18028 10968 18080
rect 11020 18068 11026 18080
rect 11882 18068 11888 18080
rect 11020 18040 11888 18068
rect 11020 18028 11026 18040
rect 11882 18028 11888 18040
rect 11940 18028 11946 18080
rect 11974 18028 11980 18080
rect 12032 18028 12038 18080
rect 12342 18028 12348 18080
rect 12400 18068 12406 18080
rect 15856 18068 15884 18108
rect 17954 18096 17960 18108
rect 18012 18096 18018 18148
rect 21468 18145 21496 18176
rect 22097 18173 22109 18207
rect 22143 18204 22155 18207
rect 22557 18207 22615 18213
rect 22557 18204 22569 18207
rect 22143 18176 22569 18204
rect 22143 18173 22155 18176
rect 22097 18167 22155 18173
rect 22557 18173 22569 18176
rect 22603 18173 22615 18207
rect 22557 18167 22615 18173
rect 21453 18139 21511 18145
rect 19306 18108 19656 18136
rect 12400 18040 15884 18068
rect 12400 18028 12406 18040
rect 15930 18028 15936 18080
rect 15988 18068 15994 18080
rect 19306 18068 19334 18108
rect 15988 18040 19334 18068
rect 15988 18028 15994 18040
rect 19518 18028 19524 18080
rect 19576 18028 19582 18080
rect 19628 18068 19656 18108
rect 21453 18105 21465 18139
rect 21499 18105 21511 18139
rect 21453 18099 21511 18105
rect 22189 18139 22247 18145
rect 22189 18105 22201 18139
rect 22235 18136 22247 18139
rect 22664 18136 22692 18235
rect 22235 18108 22692 18136
rect 22235 18105 22247 18108
rect 22189 18099 22247 18105
rect 22756 18080 22784 18312
rect 23308 18281 23336 18312
rect 23400 18281 23428 18368
rect 22833 18275 22891 18281
rect 22833 18241 22845 18275
rect 22879 18272 22891 18275
rect 23293 18275 23351 18281
rect 22879 18244 23152 18272
rect 22879 18241 22891 18244
rect 22833 18235 22891 18241
rect 23124 18145 23152 18244
rect 23293 18241 23305 18275
rect 23339 18241 23351 18275
rect 23293 18235 23351 18241
rect 23385 18275 23443 18281
rect 23385 18241 23397 18275
rect 23431 18241 23443 18275
rect 23492 18272 23520 18368
rect 23569 18275 23627 18281
rect 23569 18272 23581 18275
rect 23492 18244 23581 18272
rect 23385 18235 23443 18241
rect 23569 18241 23581 18244
rect 23615 18241 23627 18275
rect 23569 18235 23627 18241
rect 23750 18232 23756 18284
rect 23808 18232 23814 18284
rect 24210 18232 24216 18284
rect 24268 18232 24274 18284
rect 23109 18139 23167 18145
rect 23109 18105 23121 18139
rect 23155 18105 23167 18139
rect 23109 18099 23167 18105
rect 22738 18068 22744 18080
rect 19628 18040 22744 18068
rect 22738 18028 22744 18040
rect 22796 18028 22802 18080
rect 22925 18071 22983 18077
rect 22925 18037 22937 18071
rect 22971 18068 22983 18071
rect 23934 18068 23940 18080
rect 22971 18040 23940 18068
rect 22971 18037 22983 18040
rect 22925 18031 22983 18037
rect 23934 18028 23940 18040
rect 23992 18028 23998 18080
rect 24026 18028 24032 18080
rect 24084 18028 24090 18080
rect 1104 17978 24840 18000
rect 1104 17926 3917 17978
rect 3969 17926 3981 17978
rect 4033 17926 4045 17978
rect 4097 17926 4109 17978
rect 4161 17926 4173 17978
rect 4225 17926 9851 17978
rect 9903 17926 9915 17978
rect 9967 17926 9979 17978
rect 10031 17926 10043 17978
rect 10095 17926 10107 17978
rect 10159 17926 15785 17978
rect 15837 17926 15849 17978
rect 15901 17926 15913 17978
rect 15965 17926 15977 17978
rect 16029 17926 16041 17978
rect 16093 17926 21719 17978
rect 21771 17926 21783 17978
rect 21835 17926 21847 17978
rect 21899 17926 21911 17978
rect 21963 17926 21975 17978
rect 22027 17926 24840 17978
rect 1104 17904 24840 17926
rect 3326 17864 3332 17876
rect 1596 17836 3332 17864
rect 1596 17669 1624 17836
rect 3326 17824 3332 17836
rect 3384 17824 3390 17876
rect 5445 17867 5503 17873
rect 5445 17833 5457 17867
rect 5491 17864 5503 17867
rect 6730 17864 6736 17876
rect 5491 17836 6736 17864
rect 5491 17833 5503 17836
rect 5445 17827 5503 17833
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 6825 17867 6883 17873
rect 6825 17833 6837 17867
rect 6871 17864 6883 17867
rect 6914 17864 6920 17876
rect 6871 17836 6920 17864
rect 6871 17833 6883 17836
rect 6825 17827 6883 17833
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 10686 17824 10692 17876
rect 10744 17864 10750 17876
rect 10873 17867 10931 17873
rect 10873 17864 10885 17867
rect 10744 17836 10885 17864
rect 10744 17824 10750 17836
rect 10873 17833 10885 17836
rect 10919 17833 10931 17867
rect 10873 17827 10931 17833
rect 12805 17867 12863 17873
rect 12805 17833 12817 17867
rect 12851 17864 12863 17867
rect 12894 17864 12900 17876
rect 12851 17836 12900 17864
rect 12851 17833 12863 17836
rect 12805 17827 12863 17833
rect 12894 17824 12900 17836
rect 12952 17824 12958 17876
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 17310 17864 17316 17876
rect 15252 17836 17316 17864
rect 15252 17824 15258 17836
rect 17310 17824 17316 17836
rect 17368 17824 17374 17876
rect 18046 17824 18052 17876
rect 18104 17824 18110 17876
rect 18417 17867 18475 17873
rect 18417 17833 18429 17867
rect 18463 17864 18475 17867
rect 19334 17864 19340 17876
rect 18463 17836 19340 17864
rect 18463 17833 18475 17836
rect 18417 17827 18475 17833
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 19610 17824 19616 17876
rect 19668 17864 19674 17876
rect 20257 17867 20315 17873
rect 20257 17864 20269 17867
rect 19668 17836 20269 17864
rect 19668 17824 19674 17836
rect 20257 17833 20269 17836
rect 20303 17833 20315 17867
rect 20257 17827 20315 17833
rect 21634 17824 21640 17876
rect 21692 17864 21698 17876
rect 21729 17867 21787 17873
rect 21729 17864 21741 17867
rect 21692 17836 21741 17864
rect 21692 17824 21698 17836
rect 21729 17833 21741 17836
rect 21775 17864 21787 17867
rect 22278 17864 22284 17876
rect 21775 17836 22284 17864
rect 21775 17833 21787 17836
rect 21729 17827 21787 17833
rect 22278 17824 22284 17836
rect 22336 17824 22342 17876
rect 1854 17756 1860 17808
rect 1912 17756 1918 17808
rect 2317 17799 2375 17805
rect 2317 17765 2329 17799
rect 2363 17796 2375 17799
rect 2406 17796 2412 17808
rect 2363 17768 2412 17796
rect 2363 17765 2375 17768
rect 2317 17759 2375 17765
rect 2406 17756 2412 17768
rect 2464 17756 2470 17808
rect 9674 17756 9680 17808
rect 9732 17756 9738 17808
rect 1872 17728 1900 17756
rect 2593 17731 2651 17737
rect 2593 17728 2605 17731
rect 1872 17700 2605 17728
rect 2593 17697 2605 17700
rect 2639 17697 2651 17731
rect 2593 17691 2651 17697
rect 2866 17688 2872 17740
rect 2924 17688 2930 17740
rect 7650 17688 7656 17740
rect 7708 17728 7714 17740
rect 9953 17731 10011 17737
rect 9953 17728 9965 17731
rect 7708 17700 9965 17728
rect 7708 17688 7714 17700
rect 9953 17697 9965 17700
rect 9999 17728 10011 17731
rect 9999 17700 11284 17728
rect 9999 17697 10011 17700
rect 9953 17691 10011 17697
rect 1581 17663 1639 17669
rect 1581 17629 1593 17663
rect 1627 17629 1639 17663
rect 1581 17623 1639 17629
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17629 1731 17663
rect 1673 17623 1731 17629
rect 1688 17592 1716 17623
rect 1762 17620 1768 17672
rect 1820 17660 1826 17672
rect 2774 17669 2780 17672
rect 1857 17663 1915 17669
rect 1857 17660 1869 17663
rect 1820 17632 1869 17660
rect 1820 17620 1826 17632
rect 1857 17629 1869 17632
rect 1903 17629 1915 17663
rect 1857 17623 1915 17629
rect 2731 17663 2780 17669
rect 2731 17629 2743 17663
rect 2777 17629 2780 17663
rect 2731 17623 2780 17629
rect 2774 17620 2780 17623
rect 2832 17620 2838 17672
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17629 4491 17663
rect 4433 17623 4491 17629
rect 4707 17663 4765 17669
rect 4707 17629 4719 17663
rect 4753 17660 4765 17663
rect 5166 17660 5172 17672
rect 4753 17632 5172 17660
rect 4753 17629 4765 17632
rect 4707 17623 4765 17629
rect 4448 17592 4476 17623
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 5810 17620 5816 17672
rect 5868 17620 5874 17672
rect 6086 17660 6092 17672
rect 6047 17632 6092 17660
rect 6086 17620 6092 17632
rect 6144 17660 6150 17672
rect 6454 17660 6460 17672
rect 6144 17632 6460 17660
rect 6144 17620 6150 17632
rect 6454 17620 6460 17632
rect 6512 17620 6518 17672
rect 9030 17620 9036 17672
rect 9088 17620 9094 17672
rect 10134 17669 10140 17672
rect 9217 17663 9275 17669
rect 9217 17629 9229 17663
rect 9263 17629 9275 17663
rect 9217 17623 9275 17629
rect 10091 17663 10140 17669
rect 10091 17629 10103 17663
rect 10137 17629 10140 17663
rect 10091 17623 10140 17629
rect 5828 17592 5856 17620
rect 1688 17564 1900 17592
rect 1397 17527 1455 17533
rect 1397 17493 1409 17527
rect 1443 17524 1455 17527
rect 1578 17524 1584 17536
rect 1443 17496 1584 17524
rect 1443 17493 1455 17496
rect 1397 17487 1455 17493
rect 1578 17484 1584 17496
rect 1636 17484 1642 17536
rect 1872 17524 1900 17564
rect 3436 17564 4384 17592
rect 4448 17564 5856 17592
rect 2222 17524 2228 17536
rect 1872 17496 2228 17524
rect 2222 17484 2228 17496
rect 2280 17524 2286 17536
rect 2406 17524 2412 17536
rect 2280 17496 2412 17524
rect 2280 17484 2286 17496
rect 2406 17484 2412 17496
rect 2464 17484 2470 17536
rect 2958 17484 2964 17536
rect 3016 17524 3022 17536
rect 3436 17524 3464 17564
rect 3016 17496 3464 17524
rect 3016 17484 3022 17496
rect 3510 17484 3516 17536
rect 3568 17484 3574 17536
rect 4356 17524 4384 17564
rect 9122 17524 9128 17536
rect 4356 17496 9128 17524
rect 9122 17484 9128 17496
rect 9180 17524 9186 17536
rect 9232 17524 9260 17623
rect 10134 17620 10140 17623
rect 10192 17620 10198 17672
rect 10226 17620 10232 17672
rect 10284 17620 10290 17672
rect 9180 17496 9260 17524
rect 11256 17524 11284 17700
rect 11698 17688 11704 17740
rect 11756 17688 11762 17740
rect 18064 17728 18092 17824
rect 19058 17756 19064 17808
rect 19116 17796 19122 17808
rect 19116 17768 19288 17796
rect 19116 17756 19122 17768
rect 19260 17737 19288 17768
rect 19245 17731 19303 17737
rect 18064 17700 18644 17728
rect 11793 17663 11851 17669
rect 11793 17629 11805 17663
rect 11839 17660 11851 17663
rect 11974 17660 11980 17672
rect 11839 17632 11980 17660
rect 11839 17629 11851 17632
rect 11793 17623 11851 17629
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 12250 17620 12256 17672
rect 12308 17620 12314 17672
rect 15194 17660 15200 17672
rect 12360 17632 15200 17660
rect 11514 17552 11520 17604
rect 11572 17552 11578 17604
rect 11882 17552 11888 17604
rect 11940 17552 11946 17604
rect 12360 17524 12388 17632
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 16945 17663 17003 17669
rect 16945 17629 16957 17663
rect 16991 17660 17003 17663
rect 17310 17660 17316 17672
rect 16991 17632 17316 17660
rect 16991 17629 17003 17632
rect 16945 17623 17003 17629
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 17954 17620 17960 17672
rect 18012 17660 18018 17672
rect 18616 17669 18644 17700
rect 19245 17697 19257 17731
rect 19291 17697 19303 17731
rect 19245 17691 19303 17697
rect 18233 17663 18291 17669
rect 18233 17660 18245 17663
rect 18012 17632 18245 17660
rect 18012 17620 18018 17632
rect 18233 17629 18245 17632
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 18601 17663 18659 17669
rect 18601 17629 18613 17663
rect 18647 17629 18659 17663
rect 18601 17623 18659 17629
rect 19519 17663 19577 17669
rect 19519 17629 19531 17663
rect 19565 17660 19577 17663
rect 19886 17660 19892 17672
rect 19565 17632 19892 17660
rect 19565 17629 19577 17632
rect 13446 17552 13452 17604
rect 13504 17592 13510 17604
rect 18984 17598 19334 17626
rect 19519 17623 19577 17629
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 20714 17620 20720 17672
rect 20772 17620 20778 17672
rect 20990 17669 20996 17672
rect 20959 17663 20996 17669
rect 20959 17629 20971 17663
rect 20959 17623 20996 17629
rect 20990 17620 20996 17623
rect 21048 17620 21054 17672
rect 22557 17663 22615 17669
rect 22557 17629 22569 17663
rect 22603 17629 22615 17663
rect 22557 17623 22615 17629
rect 18984 17592 19012 17598
rect 13504 17564 19012 17592
rect 19306 17592 19334 17598
rect 22572 17592 22600 17623
rect 22646 17620 22652 17672
rect 22704 17620 22710 17672
rect 22738 17620 22744 17672
rect 22796 17660 22802 17672
rect 22905 17663 22963 17669
rect 22905 17660 22917 17663
rect 22796 17632 22917 17660
rect 22796 17620 22802 17632
rect 22905 17629 22917 17632
rect 22951 17629 22963 17663
rect 22905 17623 22963 17629
rect 19306 17564 22508 17592
rect 22572 17564 22692 17592
rect 13504 17552 13510 17564
rect 11256 17496 12388 17524
rect 9180 17484 9186 17496
rect 12434 17484 12440 17536
rect 12492 17524 12498 17536
rect 12621 17527 12679 17533
rect 12621 17524 12633 17527
rect 12492 17496 12633 17524
rect 12492 17484 12498 17496
rect 12621 17493 12633 17496
rect 12667 17493 12679 17527
rect 12621 17487 12679 17493
rect 14642 17484 14648 17536
rect 14700 17524 14706 17536
rect 16574 17524 16580 17536
rect 14700 17496 16580 17524
rect 14700 17484 14706 17496
rect 16574 17484 16580 17496
rect 16632 17484 16638 17536
rect 16758 17484 16764 17536
rect 16816 17524 16822 17536
rect 17034 17524 17040 17536
rect 16816 17496 17040 17524
rect 16816 17484 16822 17496
rect 17034 17484 17040 17496
rect 17092 17484 17098 17536
rect 17126 17484 17132 17536
rect 17184 17484 17190 17536
rect 19058 17484 19064 17536
rect 19116 17524 19122 17536
rect 20714 17524 20720 17536
rect 19116 17496 20720 17524
rect 19116 17484 19122 17496
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 22370 17484 22376 17536
rect 22428 17484 22434 17536
rect 22480 17524 22508 17564
rect 22554 17524 22560 17536
rect 22480 17496 22560 17524
rect 22554 17484 22560 17496
rect 22612 17484 22618 17536
rect 22664 17524 22692 17564
rect 24029 17527 24087 17533
rect 24029 17524 24041 17527
rect 22664 17496 24041 17524
rect 24029 17493 24041 17496
rect 24075 17493 24087 17527
rect 24029 17487 24087 17493
rect 1104 17434 25000 17456
rect 1104 17382 6884 17434
rect 6936 17382 6948 17434
rect 7000 17382 7012 17434
rect 7064 17382 7076 17434
rect 7128 17382 7140 17434
rect 7192 17382 12818 17434
rect 12870 17382 12882 17434
rect 12934 17382 12946 17434
rect 12998 17382 13010 17434
rect 13062 17382 13074 17434
rect 13126 17382 18752 17434
rect 18804 17382 18816 17434
rect 18868 17382 18880 17434
rect 18932 17382 18944 17434
rect 18996 17382 19008 17434
rect 19060 17382 24686 17434
rect 24738 17382 24750 17434
rect 24802 17382 24814 17434
rect 24866 17382 24878 17434
rect 24930 17382 24942 17434
rect 24994 17382 25000 17434
rect 25498 17416 25504 17468
rect 25556 17416 25562 17468
rect 1104 17360 25000 17382
rect 934 17280 940 17332
rect 992 17320 998 17332
rect 1765 17323 1823 17329
rect 1765 17320 1777 17323
rect 992 17292 1777 17320
rect 992 17280 998 17292
rect 1765 17289 1777 17292
rect 1811 17289 1823 17323
rect 1765 17283 1823 17289
rect 1854 17280 1860 17332
rect 1912 17320 1918 17332
rect 2317 17323 2375 17329
rect 2317 17320 2329 17323
rect 1912 17292 2329 17320
rect 1912 17280 1918 17292
rect 2317 17289 2329 17292
rect 2363 17289 2375 17323
rect 3789 17323 3847 17329
rect 3789 17320 3801 17323
rect 2317 17283 2375 17289
rect 2746 17292 3801 17320
rect 1302 17212 1308 17264
rect 1360 17212 1366 17264
rect 1673 17255 1731 17261
rect 1673 17221 1685 17255
rect 1719 17252 1731 17255
rect 2746 17252 2774 17292
rect 3789 17289 3801 17292
rect 3835 17289 3847 17323
rect 3789 17283 3847 17289
rect 6270 17280 6276 17332
rect 6328 17320 6334 17332
rect 6546 17320 6552 17332
rect 6328 17292 6552 17320
rect 6328 17280 6334 17292
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 7742 17280 7748 17332
rect 7800 17320 7806 17332
rect 9214 17320 9220 17332
rect 7800 17292 9220 17320
rect 7800 17280 7806 17292
rect 9214 17280 9220 17292
rect 9272 17320 9278 17332
rect 9674 17320 9680 17332
rect 9272 17292 9536 17320
rect 9272 17280 9278 17292
rect 1719 17224 2774 17252
rect 1719 17221 1731 17224
rect 1673 17215 1731 17221
rect 3050 17212 3056 17264
rect 3108 17252 3114 17264
rect 3329 17255 3387 17261
rect 3329 17252 3341 17255
rect 3108 17224 3341 17252
rect 3108 17212 3114 17224
rect 3329 17221 3341 17224
rect 3375 17221 3387 17255
rect 3329 17215 3387 17221
rect 5902 17212 5908 17264
rect 5960 17252 5966 17264
rect 5960 17224 9444 17252
rect 5960 17212 5966 17224
rect 290 17076 296 17128
rect 348 17116 354 17128
rect 658 17116 664 17128
rect 348 17088 664 17116
rect 348 17076 354 17088
rect 658 17076 664 17088
rect 716 17076 722 17128
rect 1320 17116 1348 17212
rect 2222 17144 2228 17196
rect 2280 17144 2286 17196
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17184 2835 17187
rect 3973 17187 4031 17193
rect 2823 17156 3924 17184
rect 2823 17153 2835 17156
rect 2777 17147 2835 17153
rect 3896 17116 3924 17156
rect 3973 17153 3985 17187
rect 4019 17184 4031 17187
rect 6730 17184 6736 17196
rect 4019 17156 6736 17184
rect 4019 17153 4031 17156
rect 3973 17147 4031 17153
rect 6730 17144 6736 17156
rect 6788 17144 6794 17196
rect 7558 17144 7564 17196
rect 7616 17184 7622 17196
rect 7834 17184 7840 17196
rect 7616 17156 7840 17184
rect 7616 17144 7622 17156
rect 7834 17144 7840 17156
rect 7892 17184 7898 17196
rect 8263 17187 8321 17193
rect 8263 17184 8275 17187
rect 7892 17156 8275 17184
rect 7892 17144 7898 17156
rect 8263 17153 8275 17156
rect 8309 17153 8321 17187
rect 8263 17147 8321 17153
rect 5442 17116 5448 17128
rect 1320 17088 3464 17116
rect 3896 17088 5448 17116
rect 1302 17008 1308 17060
rect 1360 17048 1366 17060
rect 1360 17020 2774 17048
rect 1360 17008 1366 17020
rect 1762 16980 1768 16992
rect 768 16952 1768 16980
rect 768 16856 796 16952
rect 1762 16940 1768 16952
rect 1820 16940 1826 16992
rect 2746 16980 2774 17020
rect 3436 16989 3464 17088
rect 5442 17076 5448 17088
rect 5500 17076 5506 17128
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 7742 17116 7748 17128
rect 7248 17088 7748 17116
rect 7248 17076 7254 17088
rect 7742 17076 7748 17088
rect 7800 17116 7806 17128
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7800 17088 8033 17116
rect 7800 17076 7806 17088
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8021 17079 8079 17085
rect 2869 16983 2927 16989
rect 2869 16980 2881 16983
rect 2746 16952 2881 16980
rect 2869 16949 2881 16952
rect 2915 16949 2927 16983
rect 2869 16943 2927 16949
rect 3421 16983 3479 16989
rect 3421 16949 3433 16983
rect 3467 16949 3479 16983
rect 3421 16943 3479 16949
rect 8846 16940 8852 16992
rect 8904 16980 8910 16992
rect 9033 16983 9091 16989
rect 9033 16980 9045 16983
rect 8904 16952 9045 16980
rect 8904 16940 8910 16952
rect 9033 16949 9045 16952
rect 9079 16949 9091 16983
rect 9416 16980 9444 17224
rect 9508 17193 9536 17292
rect 9646 17280 9680 17320
rect 9732 17280 9738 17332
rect 10226 17280 10232 17332
rect 10284 17320 10290 17332
rect 10505 17323 10563 17329
rect 10505 17320 10517 17323
rect 10284 17292 10517 17320
rect 10284 17280 10290 17292
rect 10505 17289 10517 17292
rect 10551 17289 10563 17323
rect 10505 17283 10563 17289
rect 11882 17280 11888 17332
rect 11940 17320 11946 17332
rect 12713 17323 12771 17329
rect 12713 17320 12725 17323
rect 11940 17292 12725 17320
rect 11940 17280 11946 17292
rect 12713 17289 12725 17292
rect 12759 17289 12771 17323
rect 12713 17283 12771 17289
rect 13538 17280 13544 17332
rect 13596 17320 13602 17332
rect 20990 17320 20996 17332
rect 13596 17292 20996 17320
rect 13596 17280 13602 17292
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 22094 17280 22100 17332
rect 22152 17320 22158 17332
rect 23014 17320 23020 17332
rect 22152 17292 23020 17320
rect 22152 17280 22158 17292
rect 23014 17280 23020 17292
rect 23072 17280 23078 17332
rect 23750 17280 23756 17332
rect 23808 17320 23814 17332
rect 24489 17323 24547 17329
rect 24489 17320 24501 17323
rect 23808 17292 24501 17320
rect 23808 17280 23814 17292
rect 24489 17289 24501 17292
rect 24535 17289 24547 17323
rect 24489 17283 24547 17289
rect 9646 17264 9674 17280
rect 25516 17264 25544 17416
rect 9582 17212 9588 17264
rect 9640 17224 9674 17264
rect 9640 17212 9646 17224
rect 10318 17212 10324 17264
rect 10376 17212 10382 17264
rect 10980 17224 16712 17252
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17184 9551 17187
rect 9674 17184 9680 17196
rect 9539 17156 9680 17184
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 9674 17144 9680 17156
rect 9732 17144 9738 17196
rect 9767 17187 9825 17193
rect 9767 17153 9779 17187
rect 9813 17184 9825 17187
rect 10336 17184 10364 17212
rect 10980 17196 11008 17224
rect 9813 17156 10364 17184
rect 9813 17153 9825 17156
rect 9767 17147 9825 17153
rect 10962 17144 10968 17196
rect 11020 17144 11026 17196
rect 11974 17144 11980 17196
rect 12032 17184 12038 17196
rect 15028 17193 15056 17224
rect 15013 17187 15071 17193
rect 12032 17156 12075 17184
rect 12032 17144 12038 17156
rect 15013 17153 15025 17187
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 15287 17187 15345 17193
rect 15287 17153 15299 17187
rect 15333 17184 15345 17187
rect 16298 17184 16304 17196
rect 15333 17156 16304 17184
rect 15333 17153 15345 17156
rect 15287 17147 15345 17153
rect 16298 17144 16304 17156
rect 16356 17144 16362 17196
rect 16684 17193 16712 17224
rect 17494 17212 17500 17264
rect 17552 17252 17558 17264
rect 19610 17252 19616 17264
rect 17552 17224 19334 17252
rect 17552 17212 17558 17224
rect 16669 17187 16727 17193
rect 16669 17153 16681 17187
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 16943 17187 17001 17193
rect 16943 17153 16955 17187
rect 16989 17184 17001 17187
rect 18291 17187 18349 17193
rect 16989 17156 17356 17184
rect 16989 17153 17001 17156
rect 16943 17147 17001 17153
rect 10686 17076 10692 17128
rect 10744 17116 10750 17128
rect 11701 17119 11759 17125
rect 11701 17116 11713 17119
rect 10744 17088 11713 17116
rect 10744 17076 10750 17088
rect 11701 17085 11713 17088
rect 11747 17085 11759 17119
rect 11701 17079 11759 17085
rect 12618 17076 12624 17128
rect 12676 17116 12682 17128
rect 13630 17116 13636 17128
rect 12676 17088 13636 17116
rect 12676 17076 12682 17088
rect 13630 17076 13636 17088
rect 13688 17076 13694 17128
rect 12360 17020 14320 17048
rect 9582 16980 9588 16992
rect 9416 16952 9588 16980
rect 9033 16943 9091 16949
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 11974 16940 11980 16992
rect 12032 16980 12038 16992
rect 12360 16980 12388 17020
rect 12032 16952 12388 16980
rect 12032 16940 12038 16952
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 13814 16980 13820 16992
rect 12584 16952 13820 16980
rect 12584 16940 12590 16952
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 14182 16940 14188 16992
rect 14240 16940 14246 16992
rect 14292 16980 14320 17020
rect 14366 17008 14372 17060
rect 14424 17048 14430 17060
rect 14642 17048 14648 17060
rect 14424 17020 14648 17048
rect 14424 17008 14430 17020
rect 14642 17008 14648 17020
rect 14700 17008 14706 17060
rect 16390 17048 16396 17060
rect 15948 17020 16396 17048
rect 15378 16980 15384 16992
rect 14292 16952 15384 16980
rect 15378 16940 15384 16952
rect 15436 16980 15442 16992
rect 15948 16980 15976 17020
rect 16390 17008 16396 17020
rect 16448 17008 16454 17060
rect 15436 16952 15976 16980
rect 16025 16983 16083 16989
rect 15436 16940 15442 16952
rect 16025 16949 16037 16983
rect 16071 16980 16083 16983
rect 16114 16980 16120 16992
rect 16071 16952 16120 16980
rect 16071 16949 16083 16952
rect 16025 16943 16083 16949
rect 16114 16940 16120 16952
rect 16172 16940 16178 16992
rect 16298 16940 16304 16992
rect 16356 16980 16362 16992
rect 16684 16980 16712 17147
rect 16356 16952 16712 16980
rect 16356 16940 16362 16952
rect 17034 16940 17040 16992
rect 17092 16980 17098 16992
rect 17328 16980 17356 17156
rect 18291 17153 18303 17187
rect 18337 17184 18349 17187
rect 18690 17184 18696 17196
rect 18337 17156 18696 17184
rect 18337 17153 18349 17156
rect 18291 17147 18349 17153
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 17494 17076 17500 17128
rect 17552 17116 17558 17128
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 17552 17088 18061 17116
rect 17552 17076 17558 17088
rect 18049 17085 18061 17088
rect 18095 17085 18107 17119
rect 18049 17079 18107 17085
rect 17092 16952 17356 16980
rect 17092 16940 17098 16952
rect 17678 16940 17684 16992
rect 17736 16940 17742 16992
rect 18414 16940 18420 16992
rect 18472 16980 18478 16992
rect 19061 16983 19119 16989
rect 19061 16980 19073 16983
rect 18472 16952 19073 16980
rect 18472 16940 18478 16952
rect 19061 16949 19073 16952
rect 19107 16949 19119 16983
rect 19306 16980 19334 17224
rect 19444 17224 19616 17252
rect 19444 17193 19472 17224
rect 19610 17212 19616 17224
rect 19668 17212 19674 17264
rect 25498 17212 25504 17264
rect 25556 17212 25562 17264
rect 19429 17187 19487 17193
rect 19429 17153 19441 17187
rect 19475 17153 19487 17187
rect 19429 17147 19487 17153
rect 19518 17144 19524 17196
rect 19576 17144 19582 17196
rect 21266 17144 21272 17196
rect 21324 17184 21330 17196
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21324 17156 22017 17184
rect 21324 17144 21330 17156
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 22554 17144 22560 17196
rect 22612 17184 22618 17196
rect 23075 17187 23133 17193
rect 23075 17184 23087 17187
rect 22612 17156 23087 17184
rect 22612 17144 22618 17156
rect 23075 17153 23087 17156
rect 23121 17153 23133 17187
rect 24213 17187 24271 17193
rect 24213 17184 24225 17187
rect 23075 17147 23133 17153
rect 23860 17156 24225 17184
rect 19702 17076 19708 17128
rect 19760 17076 19766 17128
rect 20714 17076 20720 17128
rect 20772 17116 20778 17128
rect 21634 17116 21640 17128
rect 20772 17088 21640 17116
rect 20772 17076 20778 17088
rect 21634 17076 21640 17088
rect 21692 17116 21698 17128
rect 22833 17119 22891 17125
rect 22833 17116 22845 17119
rect 21692 17088 22845 17116
rect 21692 17076 21698 17088
rect 22833 17085 22845 17088
rect 22879 17085 22891 17119
rect 22833 17079 22891 17085
rect 19613 17051 19671 17057
rect 19613 17017 19625 17051
rect 19659 17048 19671 17051
rect 22738 17048 22744 17060
rect 19659 17020 22744 17048
rect 19659 17017 19671 17020
rect 19613 17011 19671 17017
rect 22738 17008 22744 17020
rect 22796 17008 22802 17060
rect 21542 16980 21548 16992
rect 19306 16952 21548 16980
rect 19061 16943 19119 16949
rect 21542 16940 21548 16952
rect 21600 16940 21606 16992
rect 21821 16983 21879 16989
rect 21821 16949 21833 16983
rect 21867 16980 21879 16983
rect 22462 16980 22468 16992
rect 21867 16952 22468 16980
rect 21867 16949 21879 16952
rect 21821 16943 21879 16949
rect 22462 16940 22468 16952
rect 22520 16940 22526 16992
rect 23290 16940 23296 16992
rect 23348 16980 23354 16992
rect 23860 16989 23888 17156
rect 24213 17153 24225 17156
rect 24259 17153 24271 17187
rect 24213 17147 24271 17153
rect 23934 17076 23940 17128
rect 23992 17116 23998 17128
rect 24305 17119 24363 17125
rect 24305 17116 24317 17119
rect 23992 17088 24317 17116
rect 23992 17076 23998 17088
rect 24305 17085 24317 17088
rect 24351 17085 24363 17119
rect 24305 17079 24363 17085
rect 24489 17119 24547 17125
rect 24489 17085 24501 17119
rect 24535 17085 24547 17119
rect 24489 17079 24547 17085
rect 23845 16983 23903 16989
rect 23845 16980 23857 16983
rect 23348 16952 23857 16980
rect 23348 16940 23354 16952
rect 23845 16949 23857 16952
rect 23891 16949 23903 16983
rect 24504 16980 24532 17079
rect 25038 17076 25044 17128
rect 25096 17116 25102 17128
rect 25406 17116 25412 17128
rect 25096 17088 25412 17116
rect 25096 17076 25102 17088
rect 25406 17076 25412 17088
rect 25464 17076 25470 17128
rect 24504 16952 24900 16980
rect 23845 16943 23903 16949
rect 1104 16890 24840 16912
rect 750 16804 756 16856
rect 808 16804 814 16856
rect 1104 16838 3917 16890
rect 3969 16838 3981 16890
rect 4033 16838 4045 16890
rect 4097 16838 4109 16890
rect 4161 16838 4173 16890
rect 4225 16838 9851 16890
rect 9903 16838 9915 16890
rect 9967 16838 9979 16890
rect 10031 16838 10043 16890
rect 10095 16838 10107 16890
rect 10159 16838 15785 16890
rect 15837 16838 15849 16890
rect 15901 16838 15913 16890
rect 15965 16838 15977 16890
rect 16029 16838 16041 16890
rect 16093 16838 21719 16890
rect 21771 16838 21783 16890
rect 21835 16838 21847 16890
rect 21899 16838 21911 16890
rect 21963 16838 21975 16890
rect 22027 16838 24840 16890
rect 1104 16816 24840 16838
rect 1302 16736 1308 16788
rect 1360 16776 1366 16788
rect 3237 16779 3295 16785
rect 3237 16776 3249 16779
rect 1360 16748 3249 16776
rect 1360 16736 1366 16748
rect 3237 16745 3249 16748
rect 3283 16745 3295 16779
rect 3237 16739 3295 16745
rect 3510 16736 3516 16788
rect 3568 16776 3574 16788
rect 8386 16776 8392 16788
rect 3568 16748 8392 16776
rect 3568 16736 3574 16748
rect 8386 16736 8392 16748
rect 8444 16736 8450 16788
rect 10796 16748 11468 16776
rect 1670 16668 1676 16720
rect 1728 16668 1734 16720
rect 8205 16711 8263 16717
rect 8205 16677 8217 16711
rect 8251 16708 8263 16711
rect 8294 16708 8300 16720
rect 8251 16680 8300 16708
rect 8251 16677 8263 16680
rect 8205 16671 8263 16677
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 1578 16532 1584 16584
rect 1636 16532 1642 16584
rect 1688 16581 1716 16668
rect 3694 16600 3700 16652
rect 3752 16640 3758 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 3752 16612 4077 16640
rect 3752 16600 3758 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 7190 16640 7196 16652
rect 4065 16603 4123 16609
rect 5276 16612 7196 16640
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16541 1731 16575
rect 1673 16535 1731 16541
rect 1947 16575 2005 16581
rect 1947 16541 1959 16575
rect 1993 16572 2005 16575
rect 2038 16572 2044 16584
rect 1993 16544 2044 16572
rect 1993 16541 2005 16544
rect 1947 16535 2005 16541
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 3145 16507 3203 16513
rect 3145 16504 3157 16507
rect 1412 16476 3157 16504
rect 1412 16445 1440 16476
rect 3145 16473 3157 16476
rect 3191 16473 3203 16507
rect 4080 16504 4108 16603
rect 4246 16532 4252 16584
rect 4304 16572 4310 16584
rect 4339 16575 4397 16581
rect 4339 16572 4351 16575
rect 4304 16544 4351 16572
rect 4304 16532 4310 16544
rect 4339 16541 4351 16544
rect 4385 16541 4397 16575
rect 4339 16535 4397 16541
rect 5276 16504 5304 16612
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 10318 16640 10324 16652
rect 9824 16612 10324 16640
rect 9824 16600 9830 16612
rect 10318 16600 10324 16612
rect 10376 16640 10382 16652
rect 10686 16640 10692 16652
rect 10376 16612 10692 16640
rect 10376 16600 10382 16612
rect 10686 16600 10692 16612
rect 10744 16640 10750 16652
rect 10796 16649 10824 16748
rect 10781 16643 10839 16649
rect 10781 16640 10793 16643
rect 10744 16612 10793 16640
rect 10744 16600 10750 16612
rect 10781 16609 10793 16612
rect 10827 16609 10839 16643
rect 11440 16640 11468 16748
rect 11698 16736 11704 16788
rect 11756 16776 11762 16788
rect 11793 16779 11851 16785
rect 11793 16776 11805 16779
rect 11756 16748 11805 16776
rect 11756 16736 11762 16748
rect 11793 16745 11805 16748
rect 11839 16745 11851 16779
rect 11793 16739 11851 16745
rect 12066 16736 12072 16788
rect 12124 16776 12130 16788
rect 13446 16776 13452 16788
rect 12124 16748 13452 16776
rect 12124 16736 12130 16748
rect 13446 16736 13452 16748
rect 13504 16736 13510 16788
rect 15654 16736 15660 16788
rect 15712 16736 15718 16788
rect 16114 16736 16120 16788
rect 16172 16736 16178 16788
rect 16666 16776 16672 16788
rect 16249 16748 16672 16776
rect 15672 16708 15700 16736
rect 15488 16680 15700 16708
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 11440 16612 12633 16640
rect 10781 16603 10839 16609
rect 5350 16532 5356 16584
rect 5408 16572 5414 16584
rect 7435 16575 7493 16581
rect 7435 16572 7447 16575
rect 5408 16544 7447 16572
rect 5408 16532 5414 16544
rect 7435 16541 7447 16544
rect 7481 16541 7493 16575
rect 7435 16535 7493 16541
rect 11039 16545 11097 16551
rect 4080 16476 5304 16504
rect 3145 16467 3203 16473
rect 5442 16464 5448 16516
rect 5500 16504 5506 16516
rect 9582 16504 9588 16516
rect 5500 16476 9588 16504
rect 5500 16464 5506 16476
rect 9582 16464 9588 16476
rect 9640 16464 9646 16516
rect 9766 16464 9772 16516
rect 9824 16504 9830 16516
rect 10226 16504 10232 16516
rect 9824 16476 10232 16504
rect 9824 16464 9830 16476
rect 10226 16464 10232 16476
rect 10284 16464 10290 16516
rect 10870 16464 10876 16516
rect 10928 16464 10934 16516
rect 11039 16511 11051 16545
rect 11085 16542 11097 16545
rect 11085 16511 11098 16542
rect 11039 16505 11098 16511
rect 11070 16504 11098 16505
rect 11070 16476 11836 16504
rect 1397 16439 1455 16445
rect 1397 16405 1409 16439
rect 1443 16405 1455 16439
rect 1397 16399 1455 16405
rect 2498 16396 2504 16448
rect 2556 16436 2562 16448
rect 2685 16439 2743 16445
rect 2685 16436 2697 16439
rect 2556 16408 2697 16436
rect 2556 16396 2562 16408
rect 2685 16405 2697 16408
rect 2731 16405 2743 16439
rect 2685 16399 2743 16405
rect 4982 16396 4988 16448
rect 5040 16436 5046 16448
rect 5077 16439 5135 16445
rect 5077 16436 5089 16439
rect 5040 16408 5089 16436
rect 5040 16396 5046 16408
rect 5077 16405 5089 16408
rect 5123 16405 5135 16439
rect 5077 16399 5135 16405
rect 7926 16396 7932 16448
rect 7984 16436 7990 16448
rect 8386 16436 8392 16448
rect 7984 16408 8392 16436
rect 7984 16396 7990 16408
rect 8386 16396 8392 16408
rect 8444 16396 8450 16448
rect 9398 16396 9404 16448
rect 9456 16436 9462 16448
rect 10888 16436 10916 16464
rect 11808 16448 11836 16476
rect 9456 16408 10916 16436
rect 9456 16396 9462 16408
rect 11790 16396 11796 16448
rect 11848 16396 11854 16448
rect 12452 16436 12480 16612
rect 12621 16609 12633 16612
rect 12667 16609 12679 16643
rect 12621 16603 12679 16609
rect 13354 16600 13360 16652
rect 13412 16600 13418 16652
rect 15488 16649 15516 16680
rect 15473 16643 15531 16649
rect 15473 16609 15485 16643
rect 15519 16609 15531 16643
rect 15473 16603 15531 16609
rect 15657 16643 15715 16649
rect 15657 16609 15669 16643
rect 15703 16640 15715 16643
rect 16022 16640 16028 16652
rect 15703 16612 16028 16640
rect 15703 16609 15715 16612
rect 15657 16603 15715 16609
rect 16022 16600 16028 16612
rect 16080 16600 16086 16652
rect 16132 16649 16160 16736
rect 16117 16643 16175 16649
rect 16117 16609 16129 16643
rect 16163 16609 16175 16643
rect 16249 16640 16277 16748
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 17310 16736 17316 16788
rect 17368 16736 17374 16788
rect 17678 16776 17684 16788
rect 17420 16748 17684 16776
rect 16510 16643 16568 16649
rect 16510 16640 16522 16643
rect 16249 16612 16522 16640
rect 16117 16603 16175 16609
rect 16510 16609 16522 16612
rect 16556 16609 16568 16643
rect 16510 16603 16568 16609
rect 16669 16643 16727 16649
rect 16669 16609 16681 16643
rect 16715 16640 16727 16643
rect 17420 16640 17448 16748
rect 17678 16736 17684 16748
rect 17736 16736 17742 16788
rect 22646 16776 22652 16788
rect 21008 16748 22652 16776
rect 18322 16668 18328 16720
rect 18380 16708 18386 16720
rect 18690 16708 18696 16720
rect 18380 16680 18696 16708
rect 18380 16668 18386 16680
rect 18690 16668 18696 16680
rect 18748 16668 18754 16720
rect 21008 16649 21036 16748
rect 22646 16736 22652 16748
rect 22704 16736 22710 16788
rect 22738 16736 22744 16788
rect 22796 16736 22802 16788
rect 23385 16779 23443 16785
rect 23385 16745 23397 16779
rect 23431 16776 23443 16779
rect 24872 16776 24900 16952
rect 23431 16748 24900 16776
rect 23431 16745 23443 16748
rect 23385 16739 23443 16745
rect 22370 16668 22376 16720
rect 22428 16668 22434 16720
rect 22756 16708 22784 16736
rect 22756 16680 23704 16708
rect 20993 16643 21051 16649
rect 20993 16640 21005 16643
rect 16715 16612 17448 16640
rect 20640 16612 21005 16640
rect 16715 16609 16727 16612
rect 16669 16603 16727 16609
rect 12526 16532 12532 16584
rect 12584 16572 12590 16584
rect 12895 16575 12953 16581
rect 12895 16572 12907 16575
rect 12584 16544 12907 16572
rect 12584 16532 12590 16544
rect 12895 16541 12907 16544
rect 12941 16572 12953 16575
rect 13372 16572 13400 16600
rect 12941 16544 13400 16572
rect 12941 16541 12953 16544
rect 12895 16535 12953 16541
rect 13446 16532 13452 16584
rect 13504 16572 13510 16584
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 13504 16544 14105 16572
rect 13504 16532 13510 16544
rect 14093 16541 14105 16544
rect 14139 16541 14151 16575
rect 14366 16572 14372 16584
rect 14327 16544 14372 16572
rect 14093 16535 14151 16541
rect 14366 16532 14372 16544
rect 14424 16532 14430 16584
rect 16390 16532 16396 16584
rect 16448 16532 16454 16584
rect 17310 16532 17316 16584
rect 17368 16572 17374 16584
rect 17405 16575 17463 16581
rect 17405 16572 17417 16575
rect 17368 16544 17417 16572
rect 17368 16532 17374 16544
rect 17405 16541 17417 16544
rect 17451 16572 17463 16575
rect 17451 16544 17540 16572
rect 17451 16541 17463 16544
rect 17405 16535 17463 16541
rect 17512 16516 17540 16544
rect 17663 16545 17721 16551
rect 13556 16476 15700 16504
rect 13556 16448 13584 16476
rect 13446 16436 13452 16448
rect 12452 16408 13452 16436
rect 13446 16396 13452 16408
rect 13504 16396 13510 16448
rect 13538 16396 13544 16448
rect 13596 16396 13602 16448
rect 13630 16396 13636 16448
rect 13688 16396 13694 16448
rect 14550 16396 14556 16448
rect 14608 16436 14614 16448
rect 15105 16439 15163 16445
rect 15105 16436 15117 16439
rect 14608 16408 15117 16436
rect 14608 16396 14614 16408
rect 15105 16405 15117 16408
rect 15151 16405 15163 16439
rect 15672 16436 15700 16476
rect 17494 16464 17500 16516
rect 17552 16464 17558 16516
rect 17663 16511 17675 16545
rect 17709 16511 17721 16545
rect 19242 16532 19248 16584
rect 19300 16572 19306 16584
rect 20640 16572 20668 16612
rect 20993 16609 21005 16612
rect 21039 16609 21051 16643
rect 22388 16640 22416 16668
rect 22388 16612 23520 16640
rect 20993 16603 21051 16609
rect 21266 16581 21272 16584
rect 21260 16572 21272 16581
rect 19300 16544 20668 16572
rect 21227 16544 21272 16572
rect 19300 16532 19306 16544
rect 21260 16535 21272 16544
rect 21266 16532 21272 16535
rect 21324 16532 21330 16584
rect 22462 16532 22468 16584
rect 22520 16532 22526 16584
rect 22925 16575 22983 16581
rect 22925 16572 22937 16575
rect 22664 16544 22937 16572
rect 17663 16505 17721 16511
rect 17678 16436 17706 16505
rect 22664 16504 22692 16544
rect 22925 16541 22937 16544
rect 22971 16541 22983 16575
rect 22925 16535 22983 16541
rect 23017 16575 23075 16581
rect 23017 16541 23029 16575
rect 23063 16572 23075 16575
rect 23106 16572 23112 16584
rect 23063 16544 23112 16572
rect 23063 16541 23075 16544
rect 23017 16535 23075 16541
rect 23106 16532 23112 16544
rect 23164 16532 23170 16584
rect 23201 16575 23259 16581
rect 23201 16541 23213 16575
rect 23247 16541 23259 16575
rect 23201 16535 23259 16541
rect 23216 16504 23244 16535
rect 23290 16532 23296 16584
rect 23348 16532 23354 16584
rect 23492 16581 23520 16612
rect 23676 16581 23704 16680
rect 23934 16600 23940 16652
rect 23992 16600 23998 16652
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16541 23719 16575
rect 23661 16535 23719 16541
rect 22388 16476 22692 16504
rect 22756 16476 23244 16504
rect 17862 16436 17868 16448
rect 15672 16408 17868 16436
rect 15105 16399 15163 16405
rect 17862 16396 17868 16408
rect 17920 16396 17926 16448
rect 18046 16396 18052 16448
rect 18104 16436 18110 16448
rect 22388 16445 22416 16476
rect 18417 16439 18475 16445
rect 18417 16436 18429 16439
rect 18104 16408 18429 16436
rect 18104 16396 18110 16408
rect 18417 16405 18429 16408
rect 18463 16405 18475 16439
rect 18417 16399 18475 16405
rect 22373 16439 22431 16445
rect 22373 16405 22385 16439
rect 22419 16405 22431 16439
rect 22373 16399 22431 16405
rect 22554 16396 22560 16448
rect 22612 16396 22618 16448
rect 22756 16445 22784 16476
rect 22741 16439 22799 16445
rect 22741 16405 22753 16439
rect 22787 16405 22799 16439
rect 22741 16399 22799 16405
rect 23201 16439 23259 16445
rect 23201 16405 23213 16439
rect 23247 16436 23259 16439
rect 23382 16436 23388 16448
rect 23247 16408 23388 16436
rect 23247 16405 23259 16408
rect 23201 16399 23259 16405
rect 23382 16396 23388 16408
rect 23440 16396 23446 16448
rect 1104 16346 25000 16368
rect 1104 16294 6884 16346
rect 6936 16294 6948 16346
rect 7000 16294 7012 16346
rect 7064 16294 7076 16346
rect 7128 16294 7140 16346
rect 7192 16294 12818 16346
rect 12870 16294 12882 16346
rect 12934 16294 12946 16346
rect 12998 16294 13010 16346
rect 13062 16294 13074 16346
rect 13126 16294 18752 16346
rect 18804 16294 18816 16346
rect 18868 16294 18880 16346
rect 18932 16294 18944 16346
rect 18996 16294 19008 16346
rect 19060 16294 24686 16346
rect 24738 16294 24750 16346
rect 24802 16294 24814 16346
rect 24866 16294 24878 16346
rect 24930 16294 24942 16346
rect 24994 16294 25000 16346
rect 1104 16272 25000 16294
rect 1578 16192 1584 16244
rect 1636 16232 1642 16244
rect 5629 16235 5687 16241
rect 5629 16232 5641 16235
rect 1636 16204 5641 16232
rect 1636 16192 1642 16204
rect 5629 16201 5641 16204
rect 5675 16201 5687 16235
rect 5629 16195 5687 16201
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 9493 16235 9551 16241
rect 9493 16232 9505 16235
rect 6788 16204 9505 16232
rect 6788 16192 6794 16204
rect 9493 16201 9505 16204
rect 9539 16201 9551 16235
rect 9493 16195 9551 16201
rect 9582 16192 9588 16244
rect 9640 16232 9646 16244
rect 10965 16235 11023 16241
rect 10965 16232 10977 16235
rect 9640 16204 10977 16232
rect 9640 16192 9646 16204
rect 10965 16201 10977 16204
rect 11011 16201 11023 16235
rect 10965 16195 11023 16201
rect 11422 16192 11428 16244
rect 11480 16232 11486 16244
rect 13633 16235 13691 16241
rect 13633 16232 13645 16235
rect 11480 16204 13645 16232
rect 11480 16192 11486 16204
rect 13633 16201 13645 16204
rect 13679 16232 13691 16235
rect 14090 16232 14096 16244
rect 13679 16204 14096 16232
rect 13679 16201 13691 16204
rect 13633 16195 13691 16201
rect 14090 16192 14096 16204
rect 14148 16192 14154 16244
rect 14921 16235 14979 16241
rect 14921 16201 14933 16235
rect 14967 16232 14979 16235
rect 18230 16232 18236 16244
rect 14967 16204 18236 16232
rect 14967 16201 14979 16204
rect 14921 16195 14979 16201
rect 1486 16124 1492 16176
rect 1544 16124 1550 16176
rect 2424 16136 3740 16164
rect 14 16056 20 16108
rect 72 16096 78 16108
rect 474 16096 480 16108
rect 72 16068 480 16096
rect 72 16056 78 16068
rect 474 16056 480 16068
rect 532 16056 538 16108
rect 2314 16056 2320 16108
rect 2372 16056 2378 16108
rect 2424 16105 2452 16136
rect 3712 16108 3740 16136
rect 5534 16124 5540 16176
rect 5592 16124 5598 16176
rect 9398 16124 9404 16176
rect 9456 16124 9462 16176
rect 13354 16164 13360 16176
rect 9508 16136 13360 16164
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16065 2467 16099
rect 2409 16059 2467 16065
rect 2682 16056 2688 16108
rect 2740 16056 2746 16108
rect 3694 16056 3700 16108
rect 3752 16056 3758 16108
rect 3786 16056 3792 16108
rect 3844 16056 3850 16108
rect 4798 16056 4804 16108
rect 4856 16105 4862 16108
rect 4856 16099 4884 16105
rect 4872 16065 4884 16099
rect 4856 16059 4884 16065
rect 4856 16056 4862 16059
rect 4982 16056 4988 16108
rect 5040 16056 5046 16108
rect 3973 16031 4031 16037
rect 3973 16028 3985 16031
rect 3344 16000 3985 16028
rect 1394 15852 1400 15904
rect 1452 15892 1458 15904
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 1452 15864 1593 15892
rect 1452 15852 1458 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 1581 15855 1639 15861
rect 2130 15852 2136 15904
rect 2188 15852 2194 15904
rect 2774 15852 2780 15904
rect 2832 15892 2838 15904
rect 3234 15892 3240 15904
rect 2832 15864 3240 15892
rect 2832 15852 2838 15864
rect 3234 15852 3240 15864
rect 3292 15892 3298 15904
rect 3344 15892 3372 16000
rect 3973 15997 3985 16000
rect 4019 15997 4031 16031
rect 3973 15991 4031 15997
rect 4706 15988 4712 16040
rect 4764 16028 4770 16040
rect 5552 16028 5580 16124
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 6546 16096 6552 16108
rect 5776 16068 6552 16096
rect 5776 16056 5782 16068
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 7653 16099 7711 16105
rect 7653 16065 7665 16099
rect 7699 16096 7711 16099
rect 7742 16096 7748 16108
rect 7699 16068 7748 16096
rect 7699 16065 7711 16068
rect 7653 16059 7711 16065
rect 7742 16056 7748 16068
rect 7800 16096 7806 16108
rect 7800 16068 7972 16096
rect 7800 16056 7806 16068
rect 7466 16028 7472 16040
rect 4764 16000 7472 16028
rect 4764 15988 4770 16000
rect 7466 15988 7472 16000
rect 7524 15988 7530 16040
rect 7837 16031 7895 16037
rect 7837 16028 7849 16031
rect 7668 16000 7849 16028
rect 3421 15963 3479 15969
rect 3421 15929 3433 15963
rect 3467 15960 3479 15963
rect 4433 15963 4491 15969
rect 4433 15960 4445 15963
rect 3467 15932 4445 15960
rect 3467 15929 3479 15932
rect 3421 15923 3479 15929
rect 4433 15929 4445 15932
rect 4479 15929 4491 15963
rect 4433 15923 4491 15929
rect 5626 15920 5632 15972
rect 5684 15960 5690 15972
rect 6914 15960 6920 15972
rect 5684 15932 6920 15960
rect 5684 15920 5690 15932
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7668 15904 7696 16000
rect 7837 15997 7849 16000
rect 7883 15997 7895 16031
rect 7944 16028 7972 16068
rect 8846 16056 8852 16108
rect 8904 16056 8910 16108
rect 8202 16028 8208 16040
rect 7944 16000 8208 16028
rect 7837 15991 7895 15997
rect 8202 15988 8208 16000
rect 8260 15988 8266 16040
rect 8294 15988 8300 16040
rect 8352 15988 8358 16040
rect 8754 16037 8760 16040
rect 8573 16031 8631 16037
rect 8573 16028 8585 16031
rect 8404 16000 8585 16028
rect 8404 15960 8432 16000
rect 8573 15997 8585 16000
rect 8619 15997 8631 16031
rect 8573 15991 8631 15997
rect 8711 16031 8760 16037
rect 8711 15997 8723 16031
rect 8757 15997 8760 16031
rect 8711 15991 8760 15997
rect 8754 15988 8760 15991
rect 8812 16028 8818 16040
rect 9416 16028 9444 16124
rect 8812 16000 9444 16028
rect 8812 15988 8818 16000
rect 7944 15932 8432 15960
rect 7944 15904 7972 15932
rect 3292 15864 3372 15892
rect 3292 15852 3298 15864
rect 4522 15852 4528 15904
rect 4580 15892 4586 15904
rect 7190 15892 7196 15904
rect 4580 15864 7196 15892
rect 4580 15852 4586 15864
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 7650 15852 7656 15904
rect 7708 15852 7714 15904
rect 7926 15852 7932 15904
rect 7984 15852 7990 15904
rect 8110 15852 8116 15904
rect 8168 15892 8174 15904
rect 9508 15892 9536 16136
rect 13354 16124 13360 16136
rect 13412 16124 13418 16176
rect 13909 16167 13967 16173
rect 13909 16133 13921 16167
rect 13955 16164 13967 16167
rect 14182 16164 14188 16176
rect 13955 16136 14188 16164
rect 13955 16133 13967 16136
rect 13909 16127 13967 16133
rect 14182 16124 14188 16136
rect 14240 16124 14246 16176
rect 14550 16164 14556 16176
rect 14292 16136 14556 16164
rect 9859 16099 9917 16105
rect 9859 16065 9871 16099
rect 9905 16096 9917 16099
rect 10502 16096 10508 16108
rect 9905 16068 10508 16096
rect 9905 16065 9917 16068
rect 9859 16059 9917 16065
rect 10502 16056 10508 16068
rect 10560 16056 10566 16108
rect 11146 16056 11152 16108
rect 11204 16056 11210 16108
rect 13538 16096 13544 16108
rect 13372 16068 13544 16096
rect 9582 15988 9588 16040
rect 9640 15988 9646 16040
rect 10520 16028 10548 16056
rect 13372 16028 13400 16068
rect 13538 16056 13544 16068
rect 13596 16056 13602 16108
rect 14001 16099 14059 16105
rect 14001 16065 14013 16099
rect 14047 16096 14059 16099
rect 14292 16096 14320 16136
rect 14550 16124 14556 16136
rect 14608 16124 14614 16176
rect 14734 16124 14740 16176
rect 14792 16124 14798 16176
rect 16942 16124 16948 16176
rect 17000 16164 17006 16176
rect 17000 16136 17172 16164
rect 17000 16124 17006 16136
rect 14047 16068 14320 16096
rect 14369 16099 14427 16105
rect 14047 16065 14059 16068
rect 14001 16059 14059 16065
rect 14369 16065 14381 16099
rect 14415 16096 14427 16099
rect 16206 16096 16212 16108
rect 14415 16068 16212 16096
rect 14415 16065 14427 16068
rect 14369 16059 14427 16065
rect 16206 16056 16212 16068
rect 16264 16096 16270 16108
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 16264 16068 17049 16096
rect 16264 16056 16270 16068
rect 17037 16065 17049 16068
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 10520 16000 13400 16028
rect 13636 16040 13688 16046
rect 17144 16028 17172 16136
rect 17236 16096 17264 16204
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 19794 16192 19800 16244
rect 19852 16232 19858 16244
rect 20070 16232 20076 16244
rect 19852 16204 20076 16232
rect 19852 16192 19858 16204
rect 20070 16192 20076 16204
rect 20128 16192 20134 16244
rect 20441 16235 20499 16241
rect 20441 16201 20453 16235
rect 20487 16201 20499 16235
rect 22278 16232 22284 16244
rect 20441 16195 20499 16201
rect 21091 16204 22284 16232
rect 19334 16173 19340 16176
rect 18877 16167 18935 16173
rect 18877 16133 18889 16167
rect 18923 16164 18935 16167
rect 19328 16164 19340 16173
rect 18923 16136 19340 16164
rect 18923 16133 18935 16136
rect 18877 16127 18935 16133
rect 19328 16127 19340 16136
rect 19334 16124 19340 16127
rect 19392 16124 19398 16176
rect 20456 16164 20484 16195
rect 20456 16136 21036 16164
rect 17236 16068 17356 16096
rect 17221 16031 17279 16037
rect 17221 16028 17233 16031
rect 17144 16000 17233 16028
rect 17221 15997 17233 16000
rect 17267 15997 17279 16031
rect 17328 16028 17356 16068
rect 17954 16056 17960 16108
rect 18012 16056 18018 16108
rect 19061 16099 19119 16105
rect 19061 16065 19073 16099
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 18074 16031 18132 16037
rect 18074 16028 18086 16031
rect 17328 16000 18086 16028
rect 17221 15991 17279 15997
rect 18074 15997 18086 16000
rect 18120 15997 18132 16031
rect 18074 15991 18132 15997
rect 18233 16031 18291 16037
rect 18233 15997 18245 16031
rect 18279 16028 18291 16031
rect 18414 16028 18420 16040
rect 18279 16000 18420 16028
rect 18279 15997 18291 16000
rect 18233 15991 18291 15997
rect 18414 15988 18420 16000
rect 18472 15988 18478 16040
rect 13636 15982 13688 15988
rect 17681 15963 17739 15969
rect 17681 15929 17693 15963
rect 17727 15929 17739 15963
rect 17681 15923 17739 15929
rect 8168 15864 9536 15892
rect 8168 15852 8174 15864
rect 10594 15852 10600 15904
rect 10652 15852 10658 15904
rect 17696 15892 17724 15923
rect 18046 15892 18052 15904
rect 17696 15864 18052 15892
rect 18046 15852 18052 15864
rect 18104 15852 18110 15904
rect 19076 15892 19104 16059
rect 20530 16056 20536 16108
rect 20588 16056 20594 16108
rect 21008 16105 21036 16136
rect 20993 16099 21051 16105
rect 20993 16065 21005 16099
rect 21039 16065 21051 16099
rect 20993 16059 21051 16065
rect 20070 15988 20076 16040
rect 20128 16028 20134 16040
rect 21091 16028 21119 16204
rect 22278 16192 22284 16204
rect 22336 16192 22342 16244
rect 23014 16192 23020 16244
rect 23072 16232 23078 16244
rect 24305 16235 24363 16241
rect 23072 16204 24072 16232
rect 23072 16192 23078 16204
rect 24044 16173 24072 16204
rect 24305 16201 24317 16235
rect 24351 16232 24363 16235
rect 24394 16232 24400 16244
rect 24351 16204 24400 16232
rect 24351 16201 24363 16204
rect 24305 16195 24363 16201
rect 24394 16192 24400 16204
rect 24452 16192 24458 16244
rect 24029 16167 24087 16173
rect 20128 16000 21119 16028
rect 21192 16136 22094 16164
rect 20128 15988 20134 16000
rect 21192 15960 21220 16136
rect 22066 16135 22094 16136
rect 22066 16129 22137 16135
rect 22066 16098 22091 16129
rect 22079 16095 22091 16098
rect 22125 16095 22137 16129
rect 24029 16133 24041 16167
rect 24075 16133 24087 16167
rect 24029 16127 24087 16133
rect 22079 16089 22137 16095
rect 23477 16099 23535 16105
rect 23477 16065 23489 16099
rect 23523 16096 23535 16099
rect 23842 16096 23848 16108
rect 23523 16068 23848 16096
rect 23523 16065 23535 16068
rect 23477 16059 23535 16065
rect 23842 16056 23848 16068
rect 23900 16056 23906 16108
rect 21634 15988 21640 16040
rect 21692 16028 21698 16040
rect 21821 16031 21879 16037
rect 21821 16028 21833 16031
rect 21692 16000 21833 16028
rect 21692 15988 21698 16000
rect 21821 15997 21833 16000
rect 21867 15997 21879 16031
rect 21821 15991 21879 15997
rect 23014 15988 23020 16040
rect 23072 16028 23078 16040
rect 24210 16028 24216 16040
rect 23072 16000 24216 16028
rect 23072 15988 23078 16000
rect 24210 15988 24216 16000
rect 24268 15988 24274 16040
rect 19996 15932 21220 15960
rect 19996 15904 20024 15932
rect 20732 15904 20760 15932
rect 19242 15892 19248 15904
rect 19076 15864 19248 15892
rect 19242 15852 19248 15864
rect 19300 15852 19306 15904
rect 19978 15852 19984 15904
rect 20036 15852 20042 15904
rect 20622 15852 20628 15904
rect 20680 15852 20686 15904
rect 20714 15852 20720 15904
rect 20772 15852 20778 15904
rect 20809 15895 20867 15901
rect 20809 15861 20821 15895
rect 20855 15892 20867 15895
rect 21358 15892 21364 15904
rect 20855 15864 21364 15892
rect 20855 15861 20867 15864
rect 20809 15855 20867 15861
rect 21358 15852 21364 15864
rect 21416 15852 21422 15904
rect 22833 15895 22891 15901
rect 22833 15861 22845 15895
rect 22879 15892 22891 15895
rect 23106 15892 23112 15904
rect 22879 15864 23112 15892
rect 22879 15861 22891 15864
rect 22833 15855 22891 15861
rect 23106 15852 23112 15864
rect 23164 15852 23170 15904
rect 23750 15852 23756 15904
rect 23808 15852 23814 15904
rect 1104 15802 24840 15824
rect 1104 15750 3917 15802
rect 3969 15750 3981 15802
rect 4033 15750 4045 15802
rect 4097 15750 4109 15802
rect 4161 15750 4173 15802
rect 4225 15750 9851 15802
rect 9903 15750 9915 15802
rect 9967 15750 9979 15802
rect 10031 15750 10043 15802
rect 10095 15750 10107 15802
rect 10159 15750 15785 15802
rect 15837 15750 15849 15802
rect 15901 15750 15913 15802
rect 15965 15750 15977 15802
rect 16029 15750 16041 15802
rect 16093 15750 21719 15802
rect 21771 15750 21783 15802
rect 21835 15750 21847 15802
rect 21899 15750 21911 15802
rect 21963 15750 21975 15802
rect 22027 15750 24840 15802
rect 1104 15728 24840 15750
rect 2038 15648 2044 15700
rect 2096 15688 2102 15700
rect 4522 15688 4528 15700
rect 2096 15660 4528 15688
rect 2096 15648 2102 15660
rect 4522 15648 4528 15660
rect 4580 15648 4586 15700
rect 4614 15648 4620 15700
rect 4672 15648 4678 15700
rect 8110 15688 8116 15700
rect 6748 15660 8116 15688
rect 1946 15620 1952 15632
rect 1688 15592 1952 15620
rect 1688 15348 1716 15592
rect 1946 15580 1952 15592
rect 2004 15620 2010 15632
rect 2409 15623 2467 15629
rect 2004 15592 2360 15620
rect 2004 15580 2010 15592
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15552 1823 15555
rect 2038 15552 2044 15564
rect 1811 15524 2044 15552
rect 1811 15521 1823 15524
rect 1765 15515 1823 15521
rect 2038 15512 2044 15524
rect 2096 15512 2102 15564
rect 2332 15552 2360 15592
rect 2409 15589 2421 15623
rect 2455 15620 2467 15623
rect 2498 15620 2504 15632
rect 2455 15592 2504 15620
rect 2455 15589 2467 15592
rect 2409 15583 2467 15589
rect 2498 15580 2504 15592
rect 2556 15580 2562 15632
rect 3418 15580 3424 15632
rect 3476 15620 3482 15632
rect 3789 15623 3847 15629
rect 3789 15620 3801 15623
rect 3476 15592 3801 15620
rect 3476 15580 3482 15592
rect 3789 15589 3801 15592
rect 3835 15589 3847 15623
rect 5442 15620 5448 15632
rect 3789 15583 3847 15589
rect 5276 15592 5448 15620
rect 2866 15561 2872 15564
rect 2685 15555 2743 15561
rect 2685 15552 2697 15555
rect 2332 15524 2697 15552
rect 2685 15521 2697 15524
rect 2731 15521 2743 15555
rect 2685 15515 2743 15521
rect 2823 15555 2872 15561
rect 2823 15521 2835 15555
rect 2869 15521 2872 15555
rect 2823 15515 2872 15521
rect 2866 15512 2872 15515
rect 2924 15552 2930 15564
rect 3326 15552 3332 15564
rect 2924 15524 3332 15552
rect 2924 15512 2930 15524
rect 3326 15512 3332 15524
rect 3384 15552 3390 15564
rect 5276 15552 5304 15592
rect 5442 15580 5448 15592
rect 5500 15580 5506 15632
rect 3384 15524 3556 15552
rect 3384 15512 3390 15524
rect 1946 15444 1952 15496
rect 2004 15444 2010 15496
rect 2958 15444 2964 15496
rect 3016 15444 3022 15496
rect 2590 15348 2596 15360
rect 1688 15320 2596 15348
rect 2590 15308 2596 15320
rect 2648 15308 2654 15360
rect 3528 15348 3556 15524
rect 3620 15524 5304 15552
rect 3620 15493 3648 15524
rect 5810 15512 5816 15564
rect 5868 15512 5874 15564
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15453 3663 15487
rect 3605 15447 3663 15453
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15484 4031 15487
rect 5258 15484 5264 15496
rect 4019 15456 5264 15484
rect 4019 15453 4031 15456
rect 3973 15447 4031 15453
rect 5258 15444 5264 15456
rect 5316 15444 5322 15496
rect 5460 15456 5856 15484
rect 4525 15419 4583 15425
rect 4525 15385 4537 15419
rect 4571 15416 4583 15419
rect 4614 15416 4620 15428
rect 4571 15388 4620 15416
rect 4571 15385 4583 15388
rect 4525 15379 4583 15385
rect 4614 15376 4620 15388
rect 4672 15376 4678 15428
rect 4706 15376 4712 15428
rect 4764 15376 4770 15428
rect 5077 15419 5135 15425
rect 5077 15385 5089 15419
rect 5123 15416 5135 15419
rect 5460 15416 5488 15456
rect 5828 15425 5856 15456
rect 5902 15444 5908 15496
rect 5960 15444 5966 15496
rect 5994 15444 6000 15496
rect 6052 15444 6058 15496
rect 5123 15388 5488 15416
rect 5813 15419 5871 15425
rect 5123 15385 5135 15388
rect 5077 15379 5135 15385
rect 5813 15385 5825 15419
rect 5859 15416 5871 15419
rect 6012 15416 6040 15444
rect 5859 15388 6040 15416
rect 5859 15385 5871 15388
rect 5813 15379 5871 15385
rect 6270 15376 6276 15428
rect 6328 15376 6334 15428
rect 6748 15416 6776 15660
rect 8110 15648 8116 15660
rect 8168 15648 8174 15700
rect 9214 15648 9220 15700
rect 9272 15688 9278 15700
rect 9582 15688 9588 15700
rect 9272 15660 9588 15688
rect 9272 15648 9278 15660
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 10594 15688 10600 15700
rect 10060 15660 10600 15688
rect 10060 15629 10088 15660
rect 10594 15648 10600 15660
rect 10652 15648 10658 15700
rect 11146 15648 11152 15700
rect 11204 15688 11210 15700
rect 11241 15691 11299 15697
rect 11241 15688 11253 15691
rect 11204 15660 11253 15688
rect 11204 15648 11210 15660
rect 11241 15657 11253 15660
rect 11287 15657 11299 15691
rect 17494 15688 17500 15700
rect 11241 15651 11299 15657
rect 11440 15660 17500 15688
rect 10045 15623 10103 15629
rect 10045 15589 10057 15623
rect 10091 15589 10103 15623
rect 10045 15583 10103 15589
rect 11440 15564 11468 15660
rect 17494 15648 17500 15660
rect 17552 15648 17558 15700
rect 19334 15648 19340 15700
rect 19392 15648 19398 15700
rect 19521 15691 19579 15697
rect 19521 15657 19533 15691
rect 19567 15688 19579 15691
rect 20530 15688 20536 15700
rect 19567 15660 20536 15688
rect 19567 15657 19579 15660
rect 19521 15651 19579 15657
rect 20530 15648 20536 15660
rect 20588 15648 20594 15700
rect 20622 15648 20628 15700
rect 20680 15688 20686 15700
rect 21269 15691 21327 15697
rect 21269 15688 21281 15691
rect 20680 15660 21281 15688
rect 20680 15648 20686 15660
rect 21269 15657 21281 15660
rect 21315 15657 21327 15691
rect 21269 15651 21327 15657
rect 21358 15648 21364 15700
rect 21416 15648 21422 15700
rect 22554 15648 22560 15700
rect 22612 15688 22618 15700
rect 23293 15691 23351 15697
rect 23293 15688 23305 15691
rect 22612 15660 23305 15688
rect 22612 15648 22618 15660
rect 23293 15657 23305 15660
rect 23339 15657 23351 15691
rect 23293 15651 23351 15657
rect 23382 15648 23388 15700
rect 23440 15648 23446 15700
rect 13354 15580 13360 15632
rect 13412 15580 13418 15632
rect 6822 15512 6828 15564
rect 6880 15512 6886 15564
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 7009 15555 7067 15561
rect 7009 15552 7021 15555
rect 6972 15524 7021 15552
rect 6972 15512 6978 15524
rect 7009 15521 7021 15524
rect 7055 15521 7067 15555
rect 7009 15515 7067 15521
rect 9401 15555 9459 15561
rect 9401 15521 9413 15555
rect 9447 15552 9459 15555
rect 10321 15555 10379 15561
rect 9447 15524 9812 15552
rect 9447 15521 9459 15524
rect 9401 15515 9459 15521
rect 6564 15388 6776 15416
rect 6840 15416 6868 15512
rect 9784 15496 9812 15524
rect 10321 15521 10333 15555
rect 10367 15552 10379 15555
rect 11238 15552 11244 15564
rect 10367 15524 11244 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 11422 15512 11428 15564
rect 11480 15512 11486 15564
rect 7190 15444 7196 15496
rect 7248 15484 7254 15496
rect 7283 15487 7341 15493
rect 7283 15484 7295 15487
rect 7248 15456 7295 15484
rect 7248 15444 7254 15456
rect 7283 15453 7295 15456
rect 7329 15453 7341 15487
rect 7283 15447 7341 15453
rect 7374 15444 7380 15496
rect 7432 15484 7438 15496
rect 7432 15456 8064 15484
rect 7432 15444 7438 15456
rect 7926 15416 7932 15428
rect 6840 15388 7932 15416
rect 4724 15348 4752 15376
rect 3528 15320 4752 15348
rect 5537 15351 5595 15357
rect 5537 15317 5549 15351
rect 5583 15348 5595 15351
rect 6564 15348 6592 15388
rect 5583 15320 6592 15348
rect 5583 15317 5595 15320
rect 5537 15311 5595 15317
rect 6638 15308 6644 15360
rect 6696 15308 6702 15360
rect 6840 15357 6868 15388
rect 7926 15376 7932 15388
rect 7984 15376 7990 15428
rect 8036 15416 8064 15456
rect 9582 15444 9588 15496
rect 9640 15444 9646 15496
rect 9766 15444 9772 15496
rect 9824 15444 9830 15496
rect 10410 15444 10416 15496
rect 10468 15493 10474 15496
rect 10468 15487 10496 15493
rect 10484 15453 10496 15487
rect 10468 15447 10496 15453
rect 10468 15444 10474 15447
rect 10594 15444 10600 15496
rect 10652 15444 10658 15496
rect 11793 15487 11851 15493
rect 11793 15453 11805 15487
rect 11839 15484 11851 15487
rect 11974 15484 11980 15496
rect 11839 15456 11980 15484
rect 11839 15453 11851 15456
rect 11793 15447 11851 15453
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 12067 15487 12125 15493
rect 12067 15453 12079 15487
rect 12113 15484 12125 15487
rect 12158 15484 12164 15496
rect 12113 15456 12164 15484
rect 12113 15453 12125 15456
rect 12067 15447 12125 15453
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 13173 15487 13231 15493
rect 13173 15453 13185 15487
rect 13219 15484 13231 15487
rect 13372 15484 13400 15580
rect 15194 15512 15200 15564
rect 15252 15552 15258 15564
rect 16390 15552 16396 15564
rect 15252 15524 16396 15552
rect 15252 15512 15258 15524
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 13219 15456 13400 15484
rect 13541 15487 13599 15493
rect 13219 15453 13231 15456
rect 13173 15447 13231 15453
rect 13541 15453 13553 15487
rect 13587 15484 13599 15487
rect 14458 15484 14464 15496
rect 13587 15456 14464 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 17310 15484 17316 15496
rect 14608 15456 17316 15484
rect 14608 15444 14614 15456
rect 17310 15444 17316 15456
rect 17368 15444 17374 15496
rect 19352 15484 19380 15648
rect 20809 15623 20867 15629
rect 20809 15589 20821 15623
rect 20855 15589 20867 15623
rect 21376 15620 21404 15648
rect 21376 15592 21772 15620
rect 20809 15583 20867 15589
rect 19518 15512 19524 15564
rect 19576 15552 19582 15564
rect 19794 15552 19800 15564
rect 19576 15524 19800 15552
rect 19576 15512 19582 15524
rect 19794 15512 19800 15524
rect 19852 15512 19858 15564
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 19352 15456 19717 15484
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 20824 15484 20852 15583
rect 21453 15555 21511 15561
rect 21453 15521 21465 15555
rect 21499 15552 21511 15555
rect 21637 15555 21695 15561
rect 21637 15552 21649 15555
rect 21499 15524 21649 15552
rect 21499 15521 21511 15524
rect 21453 15515 21511 15521
rect 21637 15521 21649 15524
rect 21683 15521 21695 15555
rect 21637 15515 21695 15521
rect 21744 15493 21772 15592
rect 23400 15552 23428 15648
rect 23477 15555 23535 15561
rect 23477 15552 23489 15555
rect 23400 15524 23489 15552
rect 23477 15521 23489 15524
rect 23523 15521 23535 15555
rect 23477 15515 23535 15521
rect 21177 15487 21235 15493
rect 21177 15484 21189 15487
rect 19705 15447 19763 15453
rect 20055 15457 20113 15463
rect 8036 15388 9628 15416
rect 6825 15351 6883 15357
rect 6825 15317 6837 15351
rect 6871 15317 6883 15351
rect 6825 15311 6883 15317
rect 7374 15308 7380 15360
rect 7432 15348 7438 15360
rect 8021 15351 8079 15357
rect 8021 15348 8033 15351
rect 7432 15320 8033 15348
rect 7432 15308 7438 15320
rect 8021 15317 8033 15320
rect 8067 15317 8079 15351
rect 9600 15348 9628 15388
rect 11072 15388 13768 15416
rect 11072 15348 11100 15388
rect 9600 15320 11100 15348
rect 8021 15311 8079 15317
rect 12066 15308 12072 15360
rect 12124 15348 12130 15360
rect 12805 15351 12863 15357
rect 12805 15348 12817 15351
rect 12124 15320 12817 15348
rect 12124 15308 12130 15320
rect 12805 15317 12817 15320
rect 12851 15317 12863 15351
rect 12805 15311 12863 15317
rect 13354 15308 13360 15360
rect 13412 15308 13418 15360
rect 13740 15357 13768 15388
rect 15194 15376 15200 15428
rect 15252 15416 15258 15428
rect 15562 15416 15568 15428
rect 15252 15388 15568 15416
rect 15252 15376 15258 15388
rect 15562 15376 15568 15388
rect 15620 15376 15626 15428
rect 20055 15423 20067 15457
rect 20101 15454 20113 15457
rect 20824 15456 21189 15484
rect 20101 15423 20116 15454
rect 21177 15453 21189 15456
rect 21223 15484 21235 15487
rect 21545 15487 21603 15493
rect 21545 15484 21557 15487
rect 21223 15456 21557 15484
rect 21223 15453 21235 15456
rect 21177 15447 21235 15453
rect 21545 15453 21557 15456
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 21729 15487 21787 15493
rect 21729 15453 21741 15487
rect 21775 15453 21787 15487
rect 21729 15447 21787 15453
rect 22646 15444 22652 15496
rect 22704 15444 22710 15496
rect 22925 15487 22983 15493
rect 22925 15453 22937 15487
rect 22971 15484 22983 15487
rect 23014 15484 23020 15496
rect 22971 15456 23020 15484
rect 22971 15453 22983 15456
rect 22925 15447 22983 15453
rect 23014 15444 23020 15456
rect 23072 15444 23078 15496
rect 23106 15444 23112 15496
rect 23164 15444 23170 15496
rect 23198 15444 23204 15496
rect 23256 15444 23262 15496
rect 23566 15444 23572 15496
rect 23624 15484 23630 15496
rect 23845 15487 23903 15493
rect 23845 15484 23857 15487
rect 23624 15456 23857 15484
rect 23624 15444 23630 15456
rect 23845 15453 23857 15456
rect 23891 15453 23903 15487
rect 23845 15447 23903 15453
rect 20055 15417 20116 15423
rect 20088 15416 20116 15417
rect 20438 15416 20444 15428
rect 20088 15388 20444 15416
rect 20438 15376 20444 15388
rect 20496 15376 20502 15428
rect 22741 15419 22799 15425
rect 22741 15385 22753 15419
rect 22787 15416 22799 15419
rect 23658 15416 23664 15428
rect 22787 15388 23664 15416
rect 22787 15385 22799 15388
rect 22741 15379 22799 15385
rect 23658 15376 23664 15388
rect 23716 15376 23722 15428
rect 13725 15351 13783 15357
rect 13725 15317 13737 15351
rect 13771 15317 13783 15351
rect 13725 15311 13783 15317
rect 15470 15308 15476 15360
rect 15528 15348 15534 15360
rect 16666 15348 16672 15360
rect 15528 15320 16672 15348
rect 15528 15308 15534 15320
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 21453 15351 21511 15357
rect 21453 15317 21465 15351
rect 21499 15348 21511 15351
rect 22462 15348 22468 15360
rect 21499 15320 22468 15348
rect 21499 15317 21511 15320
rect 21453 15311 21511 15317
rect 22462 15308 22468 15320
rect 22520 15308 22526 15360
rect 23109 15351 23167 15357
rect 23109 15317 23121 15351
rect 23155 15348 23167 15351
rect 23382 15348 23388 15360
rect 23155 15320 23388 15348
rect 23155 15317 23167 15320
rect 23109 15311 23167 15317
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 23474 15308 23480 15360
rect 23532 15308 23538 15360
rect 24118 15308 24124 15360
rect 24176 15308 24182 15360
rect 1104 15258 25000 15280
rect 1104 15206 6884 15258
rect 6936 15206 6948 15258
rect 7000 15206 7012 15258
rect 7064 15206 7076 15258
rect 7128 15206 7140 15258
rect 7192 15206 12818 15258
rect 12870 15206 12882 15258
rect 12934 15206 12946 15258
rect 12998 15206 13010 15258
rect 13062 15206 13074 15258
rect 13126 15206 18752 15258
rect 18804 15206 18816 15258
rect 18868 15206 18880 15258
rect 18932 15206 18944 15258
rect 18996 15206 19008 15258
rect 19060 15206 24686 15258
rect 24738 15206 24750 15258
rect 24802 15206 24814 15258
rect 24866 15206 24878 15258
rect 24930 15206 24942 15258
rect 24994 15206 25000 15258
rect 1104 15184 25000 15206
rect 1762 15104 1768 15156
rect 1820 15104 1826 15156
rect 2222 15104 2228 15156
rect 2280 15104 2286 15156
rect 2958 15104 2964 15156
rect 3016 15144 3022 15156
rect 3145 15147 3203 15153
rect 3145 15144 3157 15147
rect 3016 15116 3157 15144
rect 3016 15104 3022 15116
rect 3145 15113 3157 15116
rect 3191 15113 3203 15147
rect 3145 15107 3203 15113
rect 3694 15104 3700 15156
rect 3752 15104 3758 15156
rect 5810 15104 5816 15156
rect 5868 15144 5874 15156
rect 5905 15147 5963 15153
rect 5905 15144 5917 15147
rect 5868 15116 5917 15144
rect 5868 15104 5874 15116
rect 5905 15113 5917 15116
rect 5951 15113 5963 15147
rect 7650 15144 7656 15156
rect 5905 15107 5963 15113
rect 6932 15116 7656 15144
rect 1673 15079 1731 15085
rect 1673 15045 1685 15079
rect 1719 15076 1731 15079
rect 2130 15076 2136 15088
rect 1719 15048 2136 15076
rect 1719 15045 1731 15048
rect 1673 15039 1731 15045
rect 2130 15036 2136 15048
rect 2188 15036 2194 15088
rect 2240 15008 2268 15104
rect 3605 15079 3663 15085
rect 3605 15045 3617 15079
rect 3651 15076 3663 15079
rect 3651 15048 6868 15076
rect 3651 15045 3663 15048
rect 3605 15039 3663 15045
rect 2375 15011 2433 15017
rect 2375 15008 2387 15011
rect 2240 14980 2387 15008
rect 2375 14977 2387 14980
rect 2421 15008 2433 15011
rect 3786 15008 3792 15020
rect 2421 14980 3792 15008
rect 2421 14977 2433 14980
rect 2375 14971 2433 14977
rect 3786 14968 3792 14980
rect 3844 14968 3850 15020
rect 4522 14968 4528 15020
rect 4580 15008 4586 15020
rect 5135 15011 5193 15017
rect 5135 15008 5147 15011
rect 4580 14980 5147 15008
rect 4580 14968 4586 14980
rect 5135 14977 5147 14980
rect 5181 14977 5193 15011
rect 5135 14971 5193 14977
rect 1670 14900 1676 14952
rect 1728 14940 1734 14952
rect 2133 14943 2191 14949
rect 2133 14940 2145 14943
rect 1728 14912 2145 14940
rect 1728 14900 1734 14912
rect 2133 14909 2145 14912
rect 2179 14909 2191 14943
rect 2133 14903 2191 14909
rect 4706 14900 4712 14952
rect 4764 14940 4770 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4764 14912 4905 14940
rect 4764 14900 4770 14912
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 6730 14900 6736 14952
rect 6788 14900 6794 14952
rect 6840 14940 6868 15048
rect 6932 15017 6960 15116
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 9214 15104 9220 15156
rect 9272 15104 9278 15156
rect 10594 15104 10600 15156
rect 10652 15144 10658 15156
rect 10689 15147 10747 15153
rect 10689 15144 10701 15147
rect 10652 15116 10701 15144
rect 10652 15104 10658 15116
rect 10689 15113 10701 15116
rect 10735 15113 10747 15147
rect 10689 15107 10747 15113
rect 11514 15104 11520 15156
rect 11572 15144 11578 15156
rect 11701 15147 11759 15153
rect 11701 15144 11713 15147
rect 11572 15116 11713 15144
rect 11572 15104 11578 15116
rect 11701 15113 11713 15116
rect 11747 15113 11759 15147
rect 11701 15107 11759 15113
rect 11974 15104 11980 15156
rect 12032 15104 12038 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12805 15147 12863 15153
rect 12805 15144 12817 15147
rect 12492 15116 12817 15144
rect 12492 15104 12498 15116
rect 12805 15113 12817 15116
rect 12851 15113 12863 15147
rect 12805 15107 12863 15113
rect 12989 15147 13047 15153
rect 12989 15113 13001 15147
rect 13035 15144 13047 15147
rect 13538 15144 13544 15156
rect 13035 15116 13544 15144
rect 13035 15113 13047 15116
rect 12989 15107 13047 15113
rect 13538 15104 13544 15116
rect 13596 15104 13602 15156
rect 14918 15104 14924 15156
rect 14976 15144 14982 15156
rect 17402 15144 17408 15156
rect 14976 15116 17408 15144
rect 14976 15104 14982 15116
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 20162 15104 20168 15156
rect 20220 15144 20226 15156
rect 20622 15144 20628 15156
rect 20220 15116 20628 15144
rect 20220 15104 20226 15116
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 22373 15147 22431 15153
rect 22373 15113 22385 15147
rect 22419 15144 22431 15147
rect 23106 15144 23112 15156
rect 22419 15116 23112 15144
rect 22419 15113 22431 15116
rect 22373 15107 22431 15113
rect 23106 15104 23112 15116
rect 23164 15104 23170 15156
rect 23566 15144 23572 15156
rect 23308 15116 23572 15144
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 14977 6975 15011
rect 6917 14971 6975 14977
rect 7742 14968 7748 15020
rect 7800 15017 7806 15020
rect 7800 15011 7828 15017
rect 7816 14977 7828 15011
rect 9232 15008 9260 15104
rect 10870 15036 10876 15088
rect 10928 15076 10934 15088
rect 11992 15076 12020 15104
rect 10928 15048 12020 15076
rect 10928 15036 10934 15048
rect 12066 15036 12072 15088
rect 12124 15036 12130 15088
rect 14274 15076 14280 15088
rect 12406 15048 14280 15076
rect 9398 15008 9404 15020
rect 9232 14980 9404 15008
rect 7800 14971 7828 14977
rect 7800 14968 7806 14971
rect 9398 14968 9404 14980
rect 9456 15008 9462 15020
rect 9677 15011 9735 15017
rect 9677 15008 9689 15011
rect 9456 14980 9689 15008
rect 9456 14968 9462 14980
rect 9677 14977 9689 14980
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 9951 15011 10009 15017
rect 9951 14977 9963 15011
rect 9997 15008 10009 15011
rect 9997 14980 10362 15008
rect 9997 14977 10009 14980
rect 9951 14971 10009 14977
rect 7282 14940 7288 14952
rect 6840 14912 7288 14940
rect 7282 14900 7288 14912
rect 7340 14900 7346 14952
rect 7374 14900 7380 14952
rect 7432 14900 7438 14952
rect 7466 14900 7472 14952
rect 7524 14940 7530 14952
rect 7653 14943 7711 14949
rect 7653 14940 7665 14943
rect 7524 14912 7665 14940
rect 7524 14900 7530 14912
rect 7653 14909 7665 14912
rect 7699 14909 7711 14943
rect 7653 14903 7711 14909
rect 7926 14900 7932 14952
rect 7984 14900 7990 14952
rect 3694 14832 3700 14884
rect 3752 14872 3758 14884
rect 3970 14872 3976 14884
rect 3752 14844 3976 14872
rect 3752 14832 3758 14844
rect 3970 14832 3976 14844
rect 4028 14832 4034 14884
rect 6748 14872 6776 14900
rect 5736 14844 6776 14872
rect 2130 14764 2136 14816
rect 2188 14804 2194 14816
rect 5736 14804 5764 14844
rect 2188 14776 5764 14804
rect 2188 14764 2194 14776
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 8573 14807 8631 14813
rect 8573 14804 8585 14807
rect 5868 14776 8585 14804
rect 5868 14764 5874 14776
rect 8573 14773 8585 14776
rect 8619 14773 8631 14807
rect 8573 14767 8631 14773
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 10334 14804 10362 14980
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 12406 15008 12434 15048
rect 14274 15036 14280 15048
rect 14332 15036 14338 15088
rect 16574 15036 16580 15088
rect 16632 15036 16638 15088
rect 18248 15048 19288 15076
rect 12032 14980 12434 15008
rect 12483 15011 12541 15017
rect 12032 14968 12038 14980
rect 12483 14977 12495 15011
rect 12529 15008 12541 15011
rect 13170 15008 13176 15020
rect 12529 14980 13176 15008
rect 12529 14977 12541 14980
rect 12483 14971 12541 14977
rect 13170 14968 13176 14980
rect 13228 15008 13234 15020
rect 14369 15011 14427 15017
rect 14369 15008 14381 15011
rect 13228 14980 14381 15008
rect 13228 14968 13234 14980
rect 14369 14977 14381 14980
rect 14415 14977 14427 15011
rect 14369 14971 14427 14977
rect 11704 14952 11756 14958
rect 14185 14943 14243 14949
rect 14185 14909 14197 14943
rect 14231 14940 14243 14943
rect 14274 14940 14280 14952
rect 14231 14912 14280 14940
rect 14231 14909 14243 14912
rect 14185 14903 14243 14909
rect 14274 14900 14280 14912
rect 14332 14900 14338 14952
rect 14918 14900 14924 14952
rect 14976 14940 14982 14952
rect 15105 14943 15163 14949
rect 15105 14940 15117 14943
rect 14976 14912 15117 14940
rect 14976 14900 14982 14912
rect 15105 14909 15117 14912
rect 15151 14909 15163 14943
rect 15105 14903 15163 14909
rect 15194 14900 15200 14952
rect 15252 14949 15258 14952
rect 15252 14943 15280 14949
rect 15268 14909 15280 14943
rect 15252 14903 15280 14909
rect 15381 14943 15439 14949
rect 15381 14909 15393 14943
rect 15427 14940 15439 14943
rect 16206 14940 16212 14952
rect 15427 14912 16212 14940
rect 15427 14909 15439 14912
rect 15381 14903 15439 14909
rect 15252 14900 15258 14903
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 16592 14940 16620 15036
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 18248 15017 18276 15048
rect 19260 15020 19288 15048
rect 22922 15047 22928 15088
rect 22907 15041 22928 15047
rect 18233 15011 18291 15017
rect 18233 15008 18245 15011
rect 18012 14980 18245 15008
rect 18012 14968 18018 14980
rect 18233 14977 18245 14980
rect 18279 14977 18291 15011
rect 18489 15011 18547 15017
rect 18489 15008 18501 15011
rect 18233 14971 18291 14977
rect 18331 14980 18501 15008
rect 18331 14940 18359 14980
rect 18489 14977 18501 14980
rect 18535 15008 18547 15011
rect 18782 15008 18788 15020
rect 18535 14980 18788 15008
rect 18535 14977 18547 14980
rect 18489 14971 18547 14977
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 19242 14968 19248 15020
rect 19300 14968 19306 15020
rect 22554 14968 22560 15020
rect 22612 14968 22618 15020
rect 22907 15007 22919 15041
rect 22980 15036 22986 15088
rect 23014 15036 23020 15088
rect 23072 15076 23078 15088
rect 23308 15076 23336 15116
rect 23566 15104 23572 15116
rect 23624 15144 23630 15156
rect 23661 15147 23719 15153
rect 23661 15144 23673 15147
rect 23624 15116 23673 15144
rect 23624 15104 23630 15116
rect 23661 15113 23673 15116
rect 23707 15113 23719 15147
rect 23661 15107 23719 15113
rect 23072 15048 23336 15076
rect 23072 15036 23078 15048
rect 23474 15036 23480 15088
rect 23532 15076 23538 15088
rect 24121 15079 24179 15085
rect 24121 15076 24133 15079
rect 23532 15048 24133 15076
rect 23532 15036 23538 15048
rect 24121 15045 24133 15048
rect 24167 15045 24179 15079
rect 24121 15039 24179 15045
rect 22953 15010 22968 15036
rect 22953 15007 22965 15010
rect 22907 15001 22965 15007
rect 16592 14912 18359 14940
rect 21634 14900 21640 14952
rect 21692 14940 21698 14952
rect 22649 14943 22707 14949
rect 22649 14940 22661 14943
rect 21692 14912 22661 14940
rect 21692 14900 21698 14912
rect 22649 14909 22661 14912
rect 22695 14909 22707 14943
rect 22649 14903 22707 14909
rect 11704 14894 11756 14900
rect 14826 14832 14832 14884
rect 14884 14832 14890 14884
rect 10962 14804 10968 14816
rect 9732 14776 10968 14804
rect 9732 14764 9738 14776
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 14642 14764 14648 14816
rect 14700 14804 14706 14816
rect 14918 14804 14924 14816
rect 14700 14776 14924 14804
rect 14700 14764 14706 14776
rect 14918 14764 14924 14776
rect 14976 14764 14982 14816
rect 15194 14764 15200 14816
rect 15252 14804 15258 14816
rect 16025 14807 16083 14813
rect 16025 14804 16037 14807
rect 15252 14776 16037 14804
rect 15252 14764 15258 14776
rect 16025 14773 16037 14776
rect 16071 14773 16083 14807
rect 16025 14767 16083 14773
rect 19610 14764 19616 14816
rect 19668 14764 19674 14816
rect 24394 14764 24400 14816
rect 24452 14764 24458 14816
rect 1104 14714 24840 14736
rect 1104 14662 3917 14714
rect 3969 14662 3981 14714
rect 4033 14662 4045 14714
rect 4097 14662 4109 14714
rect 4161 14662 4173 14714
rect 4225 14662 9851 14714
rect 9903 14662 9915 14714
rect 9967 14662 9979 14714
rect 10031 14662 10043 14714
rect 10095 14662 10107 14714
rect 10159 14662 15785 14714
rect 15837 14662 15849 14714
rect 15901 14662 15913 14714
rect 15965 14662 15977 14714
rect 16029 14662 16041 14714
rect 16093 14662 21719 14714
rect 21771 14662 21783 14714
rect 21835 14662 21847 14714
rect 21899 14662 21911 14714
rect 21963 14662 21975 14714
rect 22027 14662 24840 14714
rect 1104 14640 24840 14662
rect 1578 14560 1584 14612
rect 1636 14560 1642 14612
rect 3053 14603 3111 14609
rect 3053 14569 3065 14603
rect 3099 14569 3111 14603
rect 5810 14600 5816 14612
rect 3053 14563 3111 14569
rect 3620 14572 5816 14600
rect 1302 14492 1308 14544
rect 1360 14532 1366 14544
rect 3068 14532 3096 14563
rect 1360 14504 3096 14532
rect 1360 14492 1366 14504
rect 3418 14464 3424 14476
rect 1504 14436 3424 14464
rect 1504 14405 1532 14436
rect 3418 14424 3424 14436
rect 3476 14424 3482 14476
rect 1489 14399 1547 14405
rect 1489 14365 1501 14399
rect 1535 14365 1547 14399
rect 1489 14359 1547 14365
rect 2222 14356 2228 14408
rect 2280 14356 2286 14408
rect 2498 14396 2504 14408
rect 2424 14368 2504 14396
rect 1302 14288 1308 14340
rect 1360 14328 1366 14340
rect 2424 14337 2452 14368
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 3620 14405 3648 14572
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 5902 14560 5908 14612
rect 5960 14600 5966 14612
rect 6549 14603 6607 14609
rect 6549 14600 6561 14603
rect 5960 14572 6561 14600
rect 5960 14560 5966 14572
rect 6549 14569 6561 14572
rect 6595 14569 6607 14603
rect 6549 14563 6607 14569
rect 7926 14560 7932 14612
rect 7984 14600 7990 14612
rect 8021 14603 8079 14609
rect 8021 14600 8033 14603
rect 7984 14572 8033 14600
rect 7984 14560 7990 14572
rect 8021 14569 8033 14572
rect 8067 14569 8079 14603
rect 8021 14563 8079 14569
rect 11698 14560 11704 14612
rect 11756 14600 11762 14612
rect 11793 14603 11851 14609
rect 11793 14600 11805 14603
rect 11756 14572 11805 14600
rect 11756 14560 11762 14572
rect 11793 14569 11805 14572
rect 11839 14569 11851 14603
rect 11793 14563 11851 14569
rect 14108 14572 14780 14600
rect 4154 14492 4160 14544
rect 4212 14492 4218 14544
rect 8386 14492 8392 14544
rect 8444 14532 8450 14544
rect 10134 14532 10140 14544
rect 8444 14504 10140 14532
rect 8444 14492 8450 14504
rect 10134 14492 10140 14504
rect 10192 14492 10198 14544
rect 4706 14424 4712 14476
rect 4764 14464 4770 14476
rect 5534 14464 5540 14476
rect 4764 14436 5540 14464
rect 4764 14424 4770 14436
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 6638 14424 6644 14476
rect 6696 14464 6702 14476
rect 6822 14464 6828 14476
rect 6696 14436 6828 14464
rect 6696 14424 6702 14436
rect 6822 14424 6828 14436
rect 6880 14464 6886 14476
rect 7009 14467 7067 14473
rect 7009 14464 7021 14467
rect 6880 14436 7021 14464
rect 6880 14424 6886 14436
rect 7009 14433 7021 14436
rect 7055 14433 7067 14467
rect 7009 14427 7067 14433
rect 12710 14424 12716 14476
rect 12768 14464 12774 14476
rect 14108 14473 14136 14572
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 12768 14436 14105 14464
rect 12768 14424 12774 14436
rect 14093 14433 14105 14436
rect 14139 14433 14151 14467
rect 14752 14464 14780 14572
rect 14826 14560 14832 14612
rect 14884 14600 14890 14612
rect 15105 14603 15163 14609
rect 15105 14600 15117 14603
rect 14884 14572 15117 14600
rect 14884 14560 14890 14572
rect 15105 14569 15117 14572
rect 15151 14569 15163 14603
rect 15105 14563 15163 14569
rect 16206 14560 16212 14612
rect 16264 14600 16270 14612
rect 16485 14603 16543 14609
rect 16485 14600 16497 14603
rect 16264 14572 16497 14600
rect 16264 14560 16270 14572
rect 16485 14569 16497 14572
rect 16531 14569 16543 14603
rect 16485 14563 16543 14569
rect 18230 14560 18236 14612
rect 18288 14600 18294 14612
rect 18288 14572 19840 14600
rect 18288 14560 18294 14572
rect 19812 14544 19840 14572
rect 20732 14572 22094 14600
rect 19334 14532 19340 14544
rect 17236 14504 19340 14532
rect 15473 14467 15531 14473
rect 15473 14464 15485 14467
rect 14752 14436 15485 14464
rect 14093 14427 14151 14433
rect 15473 14433 15485 14436
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 3605 14399 3663 14405
rect 3605 14365 3617 14399
rect 3651 14365 3663 14399
rect 3605 14359 3663 14365
rect 3786 14356 3792 14408
rect 3844 14396 3850 14408
rect 5779 14399 5837 14405
rect 5779 14396 5791 14399
rect 3844 14368 5791 14396
rect 3844 14356 3850 14368
rect 5779 14365 5791 14368
rect 5825 14396 5837 14399
rect 7251 14399 7309 14405
rect 7251 14396 7263 14399
rect 5825 14368 7263 14396
rect 5825 14365 5837 14368
rect 5779 14359 5837 14365
rect 7251 14365 7263 14368
rect 7297 14365 7309 14399
rect 7251 14359 7309 14365
rect 10781 14399 10839 14405
rect 10781 14365 10793 14399
rect 10827 14396 10839 14399
rect 10827 14368 10916 14396
rect 10827 14365 10839 14368
rect 10781 14359 10839 14365
rect 10888 14340 10916 14368
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 11790 14396 11796 14408
rect 11112 14368 11796 14396
rect 11112 14356 11118 14368
rect 11790 14356 11796 14368
rect 11848 14396 11854 14408
rect 14335 14399 14393 14405
rect 14335 14396 14347 14399
rect 11848 14368 14347 14396
rect 11848 14356 11854 14368
rect 14335 14365 14347 14368
rect 14381 14365 14393 14399
rect 17034 14396 17040 14408
rect 15746 14375 17040 14396
rect 14335 14359 14393 14365
rect 15731 14369 17040 14375
rect 2409 14331 2467 14337
rect 1360 14300 2176 14328
rect 1360 14288 1366 14300
rect 2038 14220 2044 14272
rect 2096 14220 2102 14272
rect 2148 14260 2176 14300
rect 2409 14297 2421 14331
rect 2455 14297 2467 14331
rect 2409 14291 2467 14297
rect 2958 14288 2964 14340
rect 3016 14288 3022 14340
rect 3881 14331 3939 14337
rect 3881 14297 3893 14331
rect 3927 14328 3939 14331
rect 3927 14300 3961 14328
rect 3927 14297 3939 14300
rect 3881 14291 3939 14297
rect 2501 14263 2559 14269
rect 2501 14260 2513 14263
rect 2148 14232 2513 14260
rect 2501 14229 2513 14232
rect 2547 14229 2559 14263
rect 2501 14223 2559 14229
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 3421 14263 3479 14269
rect 3421 14260 3433 14263
rect 2832 14232 3433 14260
rect 2832 14220 2838 14232
rect 3421 14229 3433 14232
rect 3467 14229 3479 14263
rect 3421 14223 3479 14229
rect 3510 14220 3516 14272
rect 3568 14260 3574 14272
rect 3896 14260 3924 14291
rect 4706 14288 4712 14340
rect 4764 14328 4770 14340
rect 7834 14328 7840 14340
rect 4764 14300 7840 14328
rect 4764 14288 4770 14300
rect 7834 14288 7840 14300
rect 7892 14288 7898 14340
rect 10870 14288 10876 14340
rect 10928 14288 10934 14340
rect 15731 14335 15743 14369
rect 15777 14368 17040 14369
rect 15777 14335 15789 14368
rect 17034 14356 17040 14368
rect 17092 14356 17098 14408
rect 15731 14329 15789 14335
rect 17236 14328 17264 14504
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 19794 14492 19800 14544
rect 19852 14492 19858 14544
rect 20732 14476 20760 14572
rect 18782 14424 18788 14476
rect 18840 14464 18846 14476
rect 18840 14436 18920 14464
rect 18840 14424 18846 14436
rect 18892 14405 18920 14436
rect 19242 14424 19248 14476
rect 19300 14464 19306 14476
rect 20714 14464 20720 14476
rect 19300 14436 20720 14464
rect 19300 14424 19306 14436
rect 20714 14424 20720 14436
rect 20772 14424 20778 14476
rect 22066 14464 22094 14572
rect 22554 14560 22560 14612
rect 22612 14600 22618 14612
rect 24213 14603 24271 14609
rect 24213 14600 24225 14603
rect 22612 14572 24225 14600
rect 22612 14560 22618 14572
rect 24213 14569 24225 14572
rect 24259 14569 24271 14603
rect 24213 14563 24271 14569
rect 22833 14467 22891 14473
rect 22833 14464 22845 14467
rect 22066 14436 22845 14464
rect 22833 14433 22845 14436
rect 22879 14433 22891 14467
rect 22833 14427 22891 14433
rect 18877 14399 18935 14405
rect 18877 14365 18889 14399
rect 18923 14365 18935 14399
rect 18877 14359 18935 14365
rect 19337 14399 19395 14405
rect 19337 14365 19349 14399
rect 19383 14365 19395 14399
rect 19337 14359 19395 14365
rect 19352 14328 19380 14359
rect 19610 14356 19616 14408
rect 19668 14396 19674 14408
rect 19981 14399 20039 14405
rect 19981 14396 19993 14399
rect 19668 14368 19993 14396
rect 19668 14356 19674 14368
rect 19981 14365 19993 14368
rect 20027 14365 20039 14399
rect 20984 14399 21042 14405
rect 20984 14396 20996 14399
rect 19981 14359 20039 14365
rect 20916 14368 20996 14396
rect 20916 14340 20944 14368
rect 20984 14365 20996 14368
rect 21030 14365 21042 14399
rect 20984 14359 21042 14365
rect 22186 14356 22192 14408
rect 22244 14356 22250 14408
rect 22649 14399 22707 14405
rect 22649 14365 22661 14399
rect 22695 14365 22707 14399
rect 22649 14359 22707 14365
rect 15856 14300 17264 14328
rect 18708 14300 19380 14328
rect 15856 14272 15884 14300
rect 4525 14263 4583 14269
rect 4525 14260 4537 14263
rect 3568 14232 4537 14260
rect 3568 14220 3574 14232
rect 4525 14229 4537 14232
rect 4571 14229 4583 14263
rect 4525 14223 4583 14229
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 10226 14260 10232 14272
rect 5592 14232 10232 14260
rect 5592 14220 5598 14232
rect 10226 14220 10232 14232
rect 10284 14260 10290 14272
rect 11146 14260 11152 14272
rect 10284 14232 11152 14260
rect 10284 14220 10290 14232
rect 11146 14220 11152 14232
rect 11204 14220 11210 14272
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14182 14260 14188 14272
rect 13872 14232 14188 14260
rect 13872 14220 13878 14232
rect 14182 14220 14188 14232
rect 14240 14260 14246 14272
rect 15838 14260 15844 14272
rect 14240 14232 15844 14260
rect 14240 14220 14246 14232
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 18708 14269 18736 14300
rect 19518 14288 19524 14340
rect 19576 14328 19582 14340
rect 19576 14300 20852 14328
rect 19576 14288 19582 14300
rect 18693 14263 18751 14269
rect 18693 14229 18705 14263
rect 18739 14229 18751 14263
rect 18693 14223 18751 14229
rect 19429 14263 19487 14269
rect 19429 14229 19441 14263
rect 19475 14260 19487 14263
rect 19702 14260 19708 14272
rect 19475 14232 19708 14260
rect 19475 14229 19487 14232
rect 19429 14223 19487 14229
rect 19702 14220 19708 14232
rect 19760 14220 19766 14272
rect 19797 14263 19855 14269
rect 19797 14229 19809 14263
rect 19843 14260 19855 14263
rect 20254 14260 20260 14272
rect 19843 14232 20260 14260
rect 19843 14229 19855 14232
rect 19797 14223 19855 14229
rect 20254 14220 20260 14232
rect 20312 14220 20318 14272
rect 20824 14260 20852 14300
rect 20898 14288 20904 14340
rect 20956 14288 20962 14340
rect 22664 14328 22692 14359
rect 23106 14337 23112 14340
rect 23100 14328 23112 14337
rect 22112 14300 22692 14328
rect 23067 14300 23112 14328
rect 21358 14260 21364 14272
rect 20824 14232 21364 14260
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 22112 14269 22140 14300
rect 23100 14291 23112 14300
rect 23106 14288 23112 14291
rect 23164 14288 23170 14340
rect 22097 14263 22155 14269
rect 22097 14229 22109 14263
rect 22143 14229 22155 14263
rect 22097 14223 22155 14229
rect 22278 14220 22284 14272
rect 22336 14220 22342 14272
rect 22465 14263 22523 14269
rect 22465 14229 22477 14263
rect 22511 14260 22523 14263
rect 23198 14260 23204 14272
rect 22511 14232 23204 14260
rect 22511 14229 22523 14232
rect 22465 14223 22523 14229
rect 23198 14220 23204 14232
rect 23256 14220 23262 14272
rect 1104 14170 25000 14192
rect 1104 14118 6884 14170
rect 6936 14118 6948 14170
rect 7000 14118 7012 14170
rect 7064 14118 7076 14170
rect 7128 14118 7140 14170
rect 7192 14118 12818 14170
rect 12870 14118 12882 14170
rect 12934 14118 12946 14170
rect 12998 14118 13010 14170
rect 13062 14118 13074 14170
rect 13126 14118 18752 14170
rect 18804 14118 18816 14170
rect 18868 14118 18880 14170
rect 18932 14118 18944 14170
rect 18996 14118 19008 14170
rect 19060 14118 24686 14170
rect 24738 14118 24750 14170
rect 24802 14118 24814 14170
rect 24866 14118 24878 14170
rect 24930 14118 24942 14170
rect 24994 14118 25000 14170
rect 1104 14096 25000 14118
rect 1394 14016 1400 14068
rect 1452 14056 1458 14068
rect 1765 14059 1823 14065
rect 1765 14056 1777 14059
rect 1452 14028 1777 14056
rect 1452 14016 1458 14028
rect 1765 14025 1777 14028
rect 1811 14025 1823 14059
rect 1765 14019 1823 14025
rect 2682 14016 2688 14068
rect 2740 14056 2746 14068
rect 3694 14056 3700 14068
rect 2740 14028 3700 14056
rect 2740 14016 2746 14028
rect 3694 14016 3700 14028
rect 3752 14056 3758 14068
rect 9214 14056 9220 14068
rect 3752 14028 9220 14056
rect 3752 14016 3758 14028
rect 1673 13991 1731 13997
rect 1673 13957 1685 13991
rect 1719 13957 1731 13991
rect 1673 13951 1731 13957
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 1688 13920 1716 13951
rect 1854 13948 1860 14000
rect 1912 13988 1918 14000
rect 2225 13991 2283 13997
rect 2225 13988 2237 13991
rect 1912 13960 2237 13988
rect 1912 13948 1918 13960
rect 2225 13957 2237 13960
rect 2271 13957 2283 13991
rect 2225 13951 2283 13957
rect 2700 13960 3832 13988
rect 2700 13929 2728 13960
rect 1452 13892 1716 13920
rect 2685 13923 2743 13929
rect 1452 13880 1458 13892
rect 2685 13889 2697 13923
rect 2731 13889 2743 13923
rect 2685 13883 2743 13889
rect 2959 13923 3017 13929
rect 2959 13889 2971 13923
rect 3005 13920 3017 13923
rect 3050 13920 3056 13932
rect 3005 13892 3056 13920
rect 3005 13889 3017 13892
rect 2959 13883 3017 13889
rect 3050 13880 3056 13892
rect 3108 13880 3114 13932
rect 3804 13864 3832 13960
rect 4338 13959 4366 14028
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 9401 14059 9459 14065
rect 9401 14025 9413 14059
rect 9447 14056 9459 14059
rect 9674 14056 9680 14068
rect 9447 14028 9680 14056
rect 9447 14025 9459 14028
rect 9401 14019 9459 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 9953 14059 10011 14065
rect 9953 14025 9965 14059
rect 9999 14025 10011 14059
rect 9953 14019 10011 14025
rect 4323 13953 4381 13959
rect 4323 13919 4335 13953
rect 4369 13919 4381 13953
rect 7374 13948 7380 14000
rect 7432 13988 7438 14000
rect 9968 13988 9996 14019
rect 10778 14016 10784 14068
rect 10836 14056 10842 14068
rect 13538 14056 13544 14068
rect 10836 14028 13544 14056
rect 10836 14016 10842 14028
rect 13538 14016 13544 14028
rect 13596 14016 13602 14068
rect 16298 14056 16304 14068
rect 15120 14028 16304 14056
rect 7432 13960 9996 13988
rect 12636 13960 14504 13988
rect 7432 13948 7438 13960
rect 4323 13913 4381 13919
rect 6638 13880 6644 13932
rect 6696 13920 6702 13932
rect 8386 13920 8392 13932
rect 6696 13892 8392 13920
rect 6696 13880 6702 13892
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 8662 13920 8668 13932
rect 8623 13892 8668 13920
rect 8662 13880 8668 13892
rect 8720 13920 8726 13932
rect 9490 13920 9496 13932
rect 8720 13892 9496 13920
rect 8720 13880 8726 13892
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 10778 13920 10784 13932
rect 9815 13892 10784 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 3786 13812 3792 13864
rect 3844 13852 3850 13864
rect 4065 13855 4123 13861
rect 4065 13852 4077 13855
rect 3844 13824 4077 13852
rect 3844 13812 3850 13824
rect 4065 13821 4077 13824
rect 4111 13821 4123 13855
rect 4065 13815 4123 13821
rect 9214 13812 9220 13864
rect 9272 13852 9278 13864
rect 12636 13852 12664 13960
rect 12987 13923 13045 13929
rect 12987 13889 12999 13923
rect 13033 13920 13045 13923
rect 13033 13892 13768 13920
rect 13033 13889 13045 13892
rect 12987 13883 13045 13889
rect 9272 13824 12664 13852
rect 9272 13812 9278 13824
rect 12710 13812 12716 13864
rect 12768 13812 12774 13864
rect 13740 13852 13768 13892
rect 13740 13824 14412 13852
rect 14384 13796 14412 13824
rect 1504 13756 2434 13784
rect 1394 13676 1400 13728
rect 1452 13716 1458 13728
rect 1504 13716 1532 13756
rect 1452 13688 1532 13716
rect 1452 13676 1458 13688
rect 2314 13676 2320 13728
rect 2372 13676 2378 13728
rect 2406 13716 2434 13756
rect 3344 13756 3830 13784
rect 2958 13716 2964 13728
rect 2406 13688 2964 13716
rect 2958 13676 2964 13688
rect 3016 13676 3022 13728
rect 3050 13676 3056 13728
rect 3108 13716 3114 13728
rect 3344 13716 3372 13756
rect 3108 13688 3372 13716
rect 3108 13676 3114 13688
rect 3694 13676 3700 13728
rect 3752 13676 3758 13728
rect 3802 13716 3830 13756
rect 4722 13756 6592 13784
rect 4722 13716 4750 13756
rect 6564 13728 6592 13756
rect 13648 13756 13860 13784
rect 3802 13688 4750 13716
rect 4982 13676 4988 13728
rect 5040 13716 5046 13728
rect 5077 13719 5135 13725
rect 5077 13716 5089 13719
rect 5040 13688 5089 13716
rect 5040 13676 5046 13688
rect 5077 13685 5089 13688
rect 5123 13685 5135 13719
rect 5077 13679 5135 13685
rect 6546 13676 6552 13728
rect 6604 13676 6610 13728
rect 6730 13676 6736 13728
rect 6788 13716 6794 13728
rect 13648 13716 13676 13756
rect 6788 13688 13676 13716
rect 6788 13676 6794 13688
rect 13722 13676 13728 13728
rect 13780 13676 13786 13728
rect 13832 13716 13860 13756
rect 14366 13744 14372 13796
rect 14424 13744 14430 13796
rect 14476 13784 14504 13960
rect 15120 13920 15148 14028
rect 16298 14016 16304 14028
rect 16356 14056 16362 14068
rect 19886 14056 19892 14068
rect 16356 14028 19892 14056
rect 16356 14016 16362 14028
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 21269 14059 21327 14065
rect 21269 14025 21281 14059
rect 21315 14056 21327 14059
rect 22186 14056 22192 14068
rect 21315 14028 22192 14056
rect 21315 14025 21327 14028
rect 21269 14019 21327 14025
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 23474 14016 23480 14068
rect 23532 14056 23538 14068
rect 23532 14028 24164 14056
rect 23532 14016 23538 14028
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 23014 13988 23020 14000
rect 15344 13960 23020 13988
rect 15344 13948 15350 13960
rect 23014 13948 23020 13960
rect 23072 13948 23078 14000
rect 15197 13923 15255 13929
rect 15197 13920 15209 13923
rect 15120 13892 15209 13920
rect 15197 13889 15209 13892
rect 15243 13889 15255 13923
rect 15197 13883 15255 13889
rect 15439 13923 15497 13929
rect 15439 13889 15451 13923
rect 15485 13920 15497 13923
rect 15838 13920 15844 13932
rect 15485 13892 15844 13920
rect 15485 13889 15497 13892
rect 15439 13883 15497 13889
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 16298 13880 16304 13932
rect 16356 13920 16362 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16356 13892 16681 13920
rect 16356 13880 16362 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 16943 13923 17001 13929
rect 16943 13889 16955 13923
rect 16989 13920 17001 13923
rect 17310 13920 17316 13932
rect 16989 13892 17316 13920
rect 16989 13889 17001 13892
rect 16943 13883 17001 13889
rect 17310 13880 17316 13892
rect 17368 13920 17374 13932
rect 17586 13920 17592 13932
rect 17368 13892 17592 13920
rect 17368 13880 17374 13892
rect 17586 13880 17592 13892
rect 17644 13880 17650 13932
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13920 18107 13923
rect 18230 13920 18236 13932
rect 18095 13892 18236 13920
rect 18095 13889 18107 13892
rect 18049 13883 18107 13889
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 18323 13923 18381 13929
rect 18323 13889 18335 13923
rect 18369 13920 18381 13923
rect 18690 13920 18696 13932
rect 18369 13892 18696 13920
rect 18369 13889 18381 13892
rect 18323 13883 18381 13889
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 19334 13880 19340 13932
rect 19392 13920 19398 13932
rect 19671 13923 19729 13929
rect 19671 13920 19683 13923
rect 19392 13892 19683 13920
rect 19392 13880 19398 13892
rect 19671 13889 19683 13892
rect 19717 13889 19729 13923
rect 19671 13883 19729 13889
rect 19794 13880 19800 13932
rect 19852 13920 19858 13932
rect 19852 13892 20668 13920
rect 19852 13880 19858 13892
rect 19426 13812 19432 13864
rect 19484 13812 19490 13864
rect 20640 13852 20668 13892
rect 20898 13880 20904 13932
rect 20956 13920 20962 13932
rect 21453 13923 21511 13929
rect 21453 13920 21465 13923
rect 20956 13892 21465 13920
rect 20956 13880 20962 13892
rect 21453 13889 21465 13892
rect 21499 13889 21511 13923
rect 21453 13883 21511 13889
rect 22095 13923 22153 13929
rect 22095 13889 22107 13923
rect 22141 13920 22153 13923
rect 22186 13920 22192 13932
rect 22141 13892 22192 13920
rect 22141 13889 22153 13892
rect 22095 13883 22153 13889
rect 22186 13880 22192 13892
rect 22244 13880 22250 13932
rect 22462 13880 22468 13932
rect 22520 13920 22526 13932
rect 23290 13920 23296 13932
rect 22520 13892 23296 13920
rect 22520 13880 22526 13892
rect 23290 13880 23296 13892
rect 23348 13880 23354 13932
rect 23385 13923 23443 13929
rect 23385 13889 23397 13923
rect 23431 13920 23443 13923
rect 23566 13920 23572 13932
rect 23431 13892 23572 13920
rect 23431 13889 23443 13892
rect 23385 13883 23443 13889
rect 23566 13880 23572 13892
rect 23624 13880 23630 13932
rect 23658 13880 23664 13932
rect 23716 13880 23722 13932
rect 24136 13929 24164 14028
rect 24121 13923 24179 13929
rect 24121 13889 24133 13923
rect 24167 13889 24179 13923
rect 24121 13883 24179 13889
rect 21634 13852 21640 13864
rect 20640 13824 21640 13852
rect 21634 13812 21640 13824
rect 21692 13852 21698 13864
rect 21821 13855 21879 13861
rect 21821 13852 21833 13855
rect 21692 13824 21833 13852
rect 21692 13812 21698 13824
rect 21821 13821 21833 13824
rect 21867 13821 21879 13855
rect 21821 13815 21879 13821
rect 15194 13784 15200 13796
rect 14476 13756 15200 13784
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 24029 13787 24087 13793
rect 24029 13784 24041 13787
rect 16132 13756 16344 13784
rect 16132 13716 16160 13756
rect 13832 13688 16160 13716
rect 16206 13676 16212 13728
rect 16264 13676 16270 13728
rect 16316 13716 16344 13756
rect 17328 13756 17816 13784
rect 17328 13716 17356 13756
rect 16316 13688 17356 13716
rect 17678 13676 17684 13728
rect 17736 13676 17742 13728
rect 17788 13716 17816 13756
rect 18708 13756 19196 13784
rect 18708 13716 18736 13756
rect 17788 13688 18736 13716
rect 19058 13676 19064 13728
rect 19116 13676 19122 13728
rect 19168 13716 19196 13756
rect 20088 13756 20576 13784
rect 20088 13716 20116 13756
rect 19168 13688 20116 13716
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 20441 13719 20499 13725
rect 20441 13716 20453 13719
rect 20220 13688 20453 13716
rect 20220 13676 20226 13688
rect 20441 13685 20453 13688
rect 20487 13685 20499 13719
rect 20548 13716 20576 13756
rect 22756 13756 24041 13784
rect 22756 13716 22784 13756
rect 24029 13753 24041 13756
rect 24075 13753 24087 13787
rect 24029 13747 24087 13753
rect 20548 13688 22784 13716
rect 22833 13719 22891 13725
rect 20441 13679 20499 13685
rect 22833 13685 22845 13719
rect 22879 13716 22891 13719
rect 22922 13716 22928 13728
rect 22879 13688 22928 13716
rect 22879 13685 22891 13688
rect 22833 13679 22891 13685
rect 22922 13676 22928 13688
rect 22980 13676 22986 13728
rect 1104 13626 24840 13648
rect 1104 13574 3917 13626
rect 3969 13574 3981 13626
rect 4033 13574 4045 13626
rect 4097 13574 4109 13626
rect 4161 13574 4173 13626
rect 4225 13574 9851 13626
rect 9903 13574 9915 13626
rect 9967 13574 9979 13626
rect 10031 13574 10043 13626
rect 10095 13574 10107 13626
rect 10159 13574 15785 13626
rect 15837 13574 15849 13626
rect 15901 13574 15913 13626
rect 15965 13574 15977 13626
rect 16029 13574 16041 13626
rect 16093 13574 21719 13626
rect 21771 13574 21783 13626
rect 21835 13574 21847 13626
rect 21899 13574 21911 13626
rect 21963 13574 21975 13626
rect 22027 13574 24840 13626
rect 1104 13552 24840 13574
rect 1762 13472 1768 13524
rect 1820 13472 1826 13524
rect 2222 13472 2228 13524
rect 2280 13512 2286 13524
rect 2280 13484 3464 13512
rect 2280 13472 2286 13484
rect 1578 13336 1584 13388
rect 1636 13376 1642 13388
rect 2225 13379 2283 13385
rect 2225 13376 2237 13379
rect 1636 13348 2237 13376
rect 1636 13336 1642 13348
rect 2225 13345 2237 13348
rect 2271 13345 2283 13379
rect 2225 13339 2283 13345
rect 3234 13336 3240 13388
rect 3292 13336 3298 13388
rect 3436 13376 3464 13484
rect 3510 13472 3516 13524
rect 3568 13512 3574 13524
rect 5905 13515 5963 13521
rect 5905 13512 5917 13515
rect 3568 13484 5917 13512
rect 3568 13472 3574 13484
rect 5905 13481 5917 13484
rect 5951 13481 5963 13515
rect 8938 13512 8944 13524
rect 5905 13475 5963 13481
rect 8404 13484 8944 13512
rect 3694 13404 3700 13456
rect 3752 13444 3758 13456
rect 4433 13447 4491 13453
rect 4433 13444 4445 13447
rect 3752 13416 4445 13444
rect 3752 13404 3758 13416
rect 4433 13413 4445 13416
rect 4479 13413 4491 13447
rect 4433 13407 4491 13413
rect 3789 13379 3847 13385
rect 3789 13376 3801 13379
rect 3436 13348 3801 13376
rect 3789 13345 3801 13348
rect 3835 13376 3847 13379
rect 4522 13376 4528 13388
rect 3835 13348 4528 13376
rect 3835 13345 3847 13348
rect 3789 13339 3847 13345
rect 4522 13336 4528 13348
rect 4580 13336 4586 13388
rect 4706 13336 4712 13388
rect 4764 13336 4770 13388
rect 4798 13336 4804 13388
rect 4856 13385 4862 13388
rect 4856 13379 4884 13385
rect 4872 13345 4884 13379
rect 4856 13339 4884 13345
rect 4856 13336 4862 13339
rect 4982 13336 4988 13388
rect 5040 13336 5046 13388
rect 6638 13336 6644 13388
rect 6696 13376 6702 13388
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 6696 13348 7481 13376
rect 6696 13336 6702 13348
rect 7469 13345 7481 13348
rect 7515 13345 7527 13379
rect 7469 13339 7527 13345
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 2038 13308 2044 13320
rect 1719 13280 2044 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 2038 13268 2044 13280
rect 2096 13268 2102 13320
rect 2499 13311 2557 13317
rect 2499 13277 2511 13311
rect 2545 13308 2557 13311
rect 3050 13308 3056 13320
rect 2545 13280 3056 13308
rect 2545 13277 2557 13280
rect 2499 13271 2557 13277
rect 3050 13268 3056 13280
rect 3108 13268 3114 13320
rect 3252 13308 3280 13336
rect 3694 13308 3700 13320
rect 3252 13280 3700 13308
rect 3694 13268 3700 13280
rect 3752 13308 3758 13320
rect 3973 13311 4031 13317
rect 3973 13308 3985 13311
rect 3752 13280 3985 13308
rect 3752 13268 3758 13280
rect 3973 13277 3985 13280
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13308 5871 13311
rect 7374 13308 7380 13320
rect 5859 13280 7380 13308
rect 5859 13277 5871 13280
rect 5813 13271 5871 13277
rect 7374 13268 7380 13280
rect 7432 13268 7438 13320
rect 7743 13311 7801 13317
rect 7743 13277 7755 13311
rect 7789 13308 7801 13311
rect 8404 13308 8432 13484
rect 8938 13472 8944 13484
rect 8996 13472 9002 13524
rect 9674 13472 9680 13524
rect 9732 13512 9738 13524
rect 10134 13512 10140 13524
rect 9732 13484 10140 13512
rect 9732 13472 9738 13484
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 10226 13472 10232 13524
rect 10284 13512 10290 13524
rect 10284 13484 10732 13512
rect 10284 13472 10290 13484
rect 8481 13447 8539 13453
rect 8481 13413 8493 13447
rect 8527 13444 8539 13447
rect 9585 13447 9643 13453
rect 9585 13444 9597 13447
rect 8527 13416 9597 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 9585 13413 9597 13416
rect 9631 13413 9643 13447
rect 9585 13407 9643 13413
rect 10704 13444 10732 13484
rect 10778 13472 10784 13524
rect 10836 13472 10842 13524
rect 12710 13512 12716 13524
rect 10980 13484 12716 13512
rect 10980 13444 11008 13484
rect 10704 13416 11008 13444
rect 8570 13336 8576 13388
rect 8628 13376 8634 13388
rect 9125 13379 9183 13385
rect 9125 13376 9137 13379
rect 8628 13348 9137 13376
rect 8628 13336 8634 13348
rect 9125 13345 9137 13348
rect 9171 13376 9183 13379
rect 9490 13376 9496 13388
rect 9171 13348 9496 13376
rect 9171 13345 9183 13348
rect 9125 13339 9183 13345
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 9978 13379 10036 13385
rect 9978 13376 9990 13379
rect 9732 13348 9990 13376
rect 9732 13336 9738 13348
rect 9978 13345 9990 13348
rect 10024 13345 10036 13379
rect 9978 13339 10036 13345
rect 10134 13336 10140 13388
rect 10192 13336 10198 13388
rect 10704 13376 10732 13416
rect 10778 13376 10784 13388
rect 10704 13348 10784 13376
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 10870 13336 10876 13388
rect 10928 13336 10934 13388
rect 12268 13385 12296 13484
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 15562 13512 15568 13524
rect 15344 13484 15568 13512
rect 15344 13472 15350 13484
rect 15562 13472 15568 13484
rect 15620 13512 15626 13524
rect 15620 13484 16436 13512
rect 15620 13472 15626 13484
rect 15470 13404 15476 13456
rect 15528 13404 15534 13456
rect 16206 13404 16212 13456
rect 16264 13444 16270 13456
rect 16301 13447 16359 13453
rect 16301 13444 16313 13447
rect 16264 13416 16313 13444
rect 16264 13404 16270 13416
rect 16301 13413 16313 13416
rect 16347 13413 16359 13447
rect 16301 13407 16359 13413
rect 12253 13379 12311 13385
rect 12253 13345 12265 13379
rect 12299 13345 12311 13379
rect 15488 13376 15516 13404
rect 15654 13376 15660 13388
rect 15488 13348 15660 13376
rect 12253 13339 12311 13345
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 16408 13376 16436 13484
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 16850 13512 16856 13524
rect 16632 13484 16856 13512
rect 16632 13472 16638 13484
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 17494 13472 17500 13524
rect 17552 13472 17558 13524
rect 17862 13472 17868 13524
rect 17920 13512 17926 13524
rect 18230 13512 18236 13524
rect 17920 13484 18236 13512
rect 17920 13472 17926 13484
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 19702 13472 19708 13524
rect 19760 13512 19766 13524
rect 19797 13515 19855 13521
rect 19797 13512 19809 13515
rect 19760 13484 19809 13512
rect 19760 13472 19766 13484
rect 19797 13481 19809 13484
rect 19843 13481 19855 13515
rect 19797 13475 19855 13481
rect 22278 13472 22284 13524
rect 22336 13472 22342 13524
rect 23017 13515 23075 13521
rect 23017 13512 23029 13515
rect 22480 13484 23029 13512
rect 19058 13444 19064 13456
rect 18064 13416 19064 13444
rect 16694 13379 16752 13385
rect 16694 13376 16706 13379
rect 16408 13348 16706 13376
rect 16694 13345 16706 13348
rect 16740 13345 16752 13379
rect 16694 13339 16752 13345
rect 16853 13379 16911 13385
rect 16853 13345 16865 13379
rect 16899 13376 16911 13379
rect 17678 13376 17684 13388
rect 16899 13348 17684 13376
rect 16899 13345 16911 13348
rect 16853 13339 16911 13345
rect 17678 13336 17684 13348
rect 17736 13336 17742 13388
rect 18064 13385 18092 13416
rect 19058 13404 19064 13416
rect 19116 13404 19122 13456
rect 18049 13379 18107 13385
rect 18049 13345 18061 13379
rect 18095 13345 18107 13379
rect 18693 13379 18751 13385
rect 18693 13376 18705 13379
rect 18049 13339 18107 13345
rect 18156 13348 18705 13376
rect 7789 13280 8432 13308
rect 8941 13311 8999 13317
rect 7789 13277 7801 13280
rect 7743 13271 7801 13277
rect 7944 13252 7972 13280
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 2606 13212 3372 13240
rect 1762 13132 1768 13184
rect 1820 13172 1826 13184
rect 2606 13172 2634 13212
rect 1820 13144 2634 13172
rect 1820 13132 1826 13144
rect 3234 13132 3240 13184
rect 3292 13132 3298 13184
rect 3344 13172 3372 13212
rect 7926 13200 7932 13252
rect 7984 13200 7990 13252
rect 5629 13175 5687 13181
rect 5629 13172 5641 13175
rect 3344 13144 5641 13172
rect 5629 13141 5641 13144
rect 5675 13141 5687 13175
rect 8956 13172 8984 13271
rect 9858 13268 9864 13320
rect 9916 13268 9922 13320
rect 11164 13307 11468 13308
rect 11147 13301 11468 13307
rect 11147 13267 11159 13301
rect 11193 13280 11468 13301
rect 11193 13267 11205 13280
rect 11147 13261 11205 13267
rect 11440 13240 11468 13280
rect 11514 13268 11520 13320
rect 11572 13308 11578 13320
rect 12526 13308 12532 13320
rect 11572 13280 12296 13308
rect 12487 13280 12532 13308
rect 11572 13268 11578 13280
rect 12268 13252 12296 13280
rect 12526 13268 12532 13280
rect 12584 13268 12590 13320
rect 15841 13311 15899 13317
rect 15841 13277 15853 13311
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 11440 13212 12002 13240
rect 9490 13172 9496 13184
rect 8956 13144 9496 13172
rect 5629 13135 5687 13141
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 9858 13132 9864 13184
rect 9916 13172 9922 13184
rect 11790 13172 11796 13184
rect 9916 13144 11796 13172
rect 9916 13132 9922 13144
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 11882 13132 11888 13184
rect 11940 13132 11946 13184
rect 11974 13172 12002 13212
rect 12250 13200 12256 13252
rect 12308 13240 12314 13252
rect 12308 13212 15424 13240
rect 12308 13200 12314 13212
rect 15396 13184 15424 13212
rect 12618 13172 12624 13184
rect 11974 13144 12624 13172
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 13262 13132 13268 13184
rect 13320 13132 13326 13184
rect 15378 13132 15384 13184
rect 15436 13132 15442 13184
rect 15856 13172 15884 13271
rect 16574 13268 16580 13320
rect 16632 13268 16638 13320
rect 18156 13317 18184 13348
rect 18693 13345 18705 13348
rect 18739 13345 18751 13379
rect 19076 13376 19104 13404
rect 22480 13385 22508 13484
rect 23017 13481 23029 13484
rect 23063 13481 23075 13515
rect 23017 13475 23075 13481
rect 23198 13472 23204 13524
rect 23256 13472 23262 13524
rect 22922 13444 22928 13456
rect 22572 13416 22928 13444
rect 18693 13339 18751 13345
rect 18892 13348 19104 13376
rect 19981 13379 20039 13385
rect 18141 13311 18199 13317
rect 18141 13277 18153 13311
rect 18187 13277 18199 13311
rect 18141 13271 18199 13277
rect 18598 13268 18604 13320
rect 18656 13268 18662 13320
rect 18892 13317 18920 13348
rect 19981 13345 19993 13379
rect 20027 13376 20039 13379
rect 20165 13379 20223 13385
rect 20165 13376 20177 13379
rect 20027 13348 20177 13376
rect 20027 13345 20039 13348
rect 19981 13339 20039 13345
rect 20165 13345 20177 13348
rect 20211 13345 20223 13379
rect 20165 13339 20223 13345
rect 22465 13379 22523 13385
rect 22465 13345 22477 13379
rect 22511 13345 22523 13379
rect 22465 13339 22523 13345
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13277 18935 13311
rect 18877 13271 18935 13277
rect 19061 13311 19119 13317
rect 19061 13277 19073 13311
rect 19107 13308 19119 13311
rect 19426 13308 19432 13320
rect 19107 13280 19432 13308
rect 19107 13277 19119 13280
rect 19061 13271 19119 13277
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 19705 13311 19763 13317
rect 19705 13277 19717 13311
rect 19751 13277 19763 13311
rect 20070 13308 20076 13320
rect 19705 13271 19763 13277
rect 19904 13280 20076 13308
rect 18414 13200 18420 13252
rect 18472 13200 18478 13252
rect 18509 13243 18567 13249
rect 18509 13209 18521 13243
rect 18555 13240 18567 13243
rect 18969 13243 19027 13249
rect 18969 13240 18981 13243
rect 18555 13212 18981 13240
rect 18555 13209 18567 13212
rect 18509 13203 18567 13209
rect 18969 13209 18981 13212
rect 19015 13209 19027 13243
rect 19720 13240 19748 13271
rect 19904 13240 19932 13280
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 20254 13268 20260 13320
rect 20312 13268 20318 13320
rect 22189 13311 22247 13317
rect 22189 13277 22201 13311
rect 22235 13308 22247 13311
rect 22572 13308 22600 13416
rect 22922 13404 22928 13416
rect 22980 13444 22986 13456
rect 22980 13416 23058 13444
rect 22980 13404 22986 13416
rect 22646 13336 22652 13388
rect 22704 13336 22710 13388
rect 22235 13280 22600 13308
rect 22235 13277 22247 13280
rect 22189 13271 22247 13277
rect 19720 13212 19932 13240
rect 19996 13212 22094 13240
rect 18969 13203 19027 13209
rect 16390 13172 16396 13184
rect 15856 13144 16396 13172
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 19996 13181 20024 13212
rect 19981 13175 20039 13181
rect 19981 13141 19993 13175
rect 20027 13141 20039 13175
rect 19981 13135 20039 13141
rect 20162 13132 20168 13184
rect 20220 13172 20226 13184
rect 20530 13172 20536 13184
rect 20220 13144 20536 13172
rect 20220 13132 20226 13144
rect 20530 13132 20536 13144
rect 20588 13132 20594 13184
rect 22066 13172 22094 13212
rect 22370 13172 22376 13184
rect 22066 13144 22376 13172
rect 22370 13132 22376 13144
rect 22428 13132 22434 13184
rect 22462 13132 22468 13184
rect 22520 13132 22526 13184
rect 22664 13181 22692 13336
rect 22931 13311 22989 13317
rect 22833 13287 22891 13293
rect 22833 13253 22845 13287
rect 22879 13253 22891 13287
rect 22931 13277 22943 13311
rect 22977 13308 22989 13311
rect 23030 13308 23058 13416
rect 23216 13376 23244 13472
rect 23385 13447 23443 13453
rect 23385 13413 23397 13447
rect 23431 13444 23443 13447
rect 24670 13444 24676 13456
rect 23431 13416 24676 13444
rect 23431 13413 23443 13416
rect 23385 13407 23443 13413
rect 24670 13404 24676 13416
rect 24728 13404 24734 13456
rect 23124 13348 23244 13376
rect 23124 13317 23152 13348
rect 22977 13280 23058 13308
rect 23109 13311 23167 13317
rect 22977 13277 22989 13280
rect 22931 13271 22989 13277
rect 23109 13277 23121 13311
rect 23155 13277 23167 13311
rect 23109 13271 23167 13277
rect 23201 13311 23259 13317
rect 23201 13277 23213 13311
rect 23247 13308 23259 13311
rect 23290 13308 23296 13320
rect 23247 13280 23296 13308
rect 23247 13277 23259 13280
rect 23201 13271 23259 13277
rect 23290 13268 23296 13280
rect 23348 13268 23354 13320
rect 23661 13311 23719 13317
rect 23661 13277 23673 13311
rect 23707 13308 23719 13311
rect 25682 13308 25688 13320
rect 23707 13280 25688 13308
rect 23707 13277 23719 13280
rect 23661 13271 23719 13277
rect 25682 13268 25688 13280
rect 25740 13268 25746 13320
rect 22833 13247 22891 13253
rect 22649 13175 22707 13181
rect 22649 13141 22661 13175
rect 22695 13141 22707 13175
rect 22848 13172 22876 13247
rect 24026 13200 24032 13252
rect 24084 13200 24090 13252
rect 23106 13172 23112 13184
rect 22848 13144 23112 13172
rect 22649 13135 22707 13141
rect 23106 13132 23112 13144
rect 23164 13132 23170 13184
rect 1104 13082 25000 13104
rect 1104 13030 6884 13082
rect 6936 13030 6948 13082
rect 7000 13030 7012 13082
rect 7064 13030 7076 13082
rect 7128 13030 7140 13082
rect 7192 13030 12818 13082
rect 12870 13030 12882 13082
rect 12934 13030 12946 13082
rect 12998 13030 13010 13082
rect 13062 13030 13074 13082
rect 13126 13030 18752 13082
rect 18804 13030 18816 13082
rect 18868 13030 18880 13082
rect 18932 13030 18944 13082
rect 18996 13030 19008 13082
rect 19060 13030 24686 13082
rect 24738 13030 24750 13082
rect 24802 13030 24814 13082
rect 24866 13030 24878 13082
rect 24930 13030 24942 13082
rect 24994 13030 25000 13082
rect 1104 13008 25000 13030
rect 1670 12928 1676 12980
rect 1728 12928 1734 12980
rect 2038 12928 2044 12980
rect 2096 12968 2102 12980
rect 2682 12968 2688 12980
rect 2096 12940 2688 12968
rect 2096 12928 2102 12940
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 3050 12928 3056 12980
rect 3108 12968 3114 12980
rect 3326 12968 3332 12980
rect 3108 12940 3332 12968
rect 3108 12928 3114 12940
rect 3326 12928 3332 12940
rect 3384 12928 3390 12980
rect 3510 12928 3516 12980
rect 3568 12968 3574 12980
rect 4157 12971 4215 12977
rect 4157 12968 4169 12971
rect 3568 12940 4169 12968
rect 3568 12928 3574 12940
rect 4157 12937 4169 12940
rect 4203 12937 4215 12971
rect 4157 12931 4215 12937
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 18414 12968 18420 12980
rect 4580 12940 18420 12968
rect 4580 12928 4586 12940
rect 18414 12928 18420 12940
rect 18472 12928 18478 12980
rect 18598 12928 18604 12980
rect 18656 12928 18662 12980
rect 19426 12928 19432 12980
rect 19484 12928 19490 12980
rect 19978 12928 19984 12980
rect 20036 12968 20042 12980
rect 20438 12968 20444 12980
rect 20036 12940 20444 12968
rect 20036 12928 20042 12940
rect 20438 12928 20444 12940
rect 20496 12928 20502 12980
rect 22462 12928 22468 12980
rect 22520 12928 22526 12980
rect 24397 12971 24455 12977
rect 24397 12937 24409 12971
rect 24443 12968 24455 12971
rect 24486 12968 24492 12980
rect 24443 12940 24492 12968
rect 24443 12937 24455 12940
rect 24397 12931 24455 12937
rect 24486 12928 24492 12940
rect 24544 12928 24550 12980
rect 3878 12860 3884 12912
rect 3936 12900 3942 12912
rect 3936 12872 4200 12900
rect 3936 12860 3942 12872
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12832 1639 12835
rect 1627 12804 2360 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 1946 12724 1952 12776
rect 2004 12724 2010 12776
rect 2041 12767 2099 12773
rect 2041 12733 2053 12767
rect 2087 12764 2099 12767
rect 2130 12764 2136 12776
rect 2087 12736 2136 12764
rect 2087 12733 2099 12736
rect 2041 12727 2099 12733
rect 2130 12724 2136 12736
rect 2188 12724 2194 12776
rect 2225 12767 2283 12773
rect 2225 12733 2237 12767
rect 2271 12733 2283 12767
rect 2332 12764 2360 12804
rect 3050 12792 3056 12844
rect 3108 12841 3114 12844
rect 3108 12835 3136 12841
rect 3124 12801 3136 12835
rect 3108 12795 3136 12801
rect 3108 12792 3114 12795
rect 3970 12792 3976 12844
rect 4028 12792 4034 12844
rect 4065 12835 4123 12841
rect 4065 12801 4077 12835
rect 4111 12801 4123 12835
rect 4065 12795 4123 12801
rect 2774 12764 2780 12776
rect 2332 12736 2780 12764
rect 2225 12727 2283 12733
rect 1964 12696 1992 12724
rect 2240 12696 2268 12727
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 2958 12724 2964 12776
rect 3016 12724 3022 12776
rect 3237 12767 3295 12773
rect 3237 12733 3249 12767
rect 3283 12764 3295 12767
rect 3988 12764 4016 12792
rect 3283 12736 4016 12764
rect 3283 12733 3295 12736
rect 3237 12727 3295 12733
rect 2406 12696 2412 12708
rect 1964 12668 2412 12696
rect 2406 12656 2412 12668
rect 2464 12656 2470 12708
rect 2682 12656 2688 12708
rect 2740 12656 2746 12708
rect 4080 12696 4108 12795
rect 4172 12764 4200 12872
rect 6546 12860 6552 12912
rect 6604 12860 6610 12912
rect 14458 12860 14464 12912
rect 14516 12860 14522 12912
rect 14642 12860 14648 12912
rect 14700 12860 14706 12912
rect 15378 12860 15384 12912
rect 15436 12900 15442 12912
rect 16574 12900 16580 12912
rect 15436 12872 16580 12900
rect 15436 12860 15442 12872
rect 16574 12860 16580 12872
rect 16632 12860 16638 12912
rect 18616 12900 18644 12928
rect 22480 12900 22508 12928
rect 24121 12903 24179 12909
rect 24121 12900 24133 12903
rect 17696 12872 18644 12900
rect 18892 12872 20576 12900
rect 22480 12872 24133 12900
rect 4614 12792 4620 12844
rect 4672 12832 4678 12844
rect 5135 12835 5193 12841
rect 5135 12832 5147 12835
rect 4672 12804 5147 12832
rect 4672 12792 4678 12804
rect 5135 12801 5147 12804
rect 5181 12801 5193 12835
rect 6564 12832 6592 12860
rect 6639 12835 6697 12841
rect 6639 12832 6651 12835
rect 6564 12804 6651 12832
rect 5135 12795 5193 12801
rect 6639 12801 6651 12804
rect 6685 12801 6697 12835
rect 6639 12795 6697 12801
rect 9582 12792 9588 12844
rect 9640 12792 9646 12844
rect 11241 12835 11299 12841
rect 11241 12801 11253 12835
rect 11287 12832 11299 12835
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 11287 12804 11529 12832
rect 11287 12801 11299 12804
rect 11241 12795 11299 12801
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 13538 12792 13544 12844
rect 13596 12792 13602 12844
rect 13630 12792 13636 12844
rect 13688 12841 13694 12844
rect 13688 12835 13716 12841
rect 13704 12801 13716 12835
rect 13688 12795 13716 12801
rect 13688 12792 13694 12795
rect 13814 12792 13820 12844
rect 13872 12792 13878 12844
rect 14550 12792 14556 12844
rect 14608 12792 14614 12844
rect 14660 12832 14688 12860
rect 14795 12835 14853 12841
rect 14795 12832 14807 12835
rect 14660 12804 14807 12832
rect 14795 12801 14807 12804
rect 14841 12801 14853 12835
rect 14795 12795 14853 12801
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 4172 12736 4905 12764
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 4893 12727 4951 12733
rect 6365 12767 6423 12773
rect 6365 12733 6377 12767
rect 6411 12733 6423 12767
rect 6365 12727 6423 12733
rect 9401 12767 9459 12773
rect 9401 12733 9413 12767
rect 9447 12764 9459 12767
rect 9490 12764 9496 12776
rect 9447 12736 9496 12764
rect 9447 12733 9459 12736
rect 9401 12727 9459 12733
rect 3620 12668 4108 12696
rect 1946 12588 1952 12640
rect 2004 12628 2010 12640
rect 3620 12628 3648 12668
rect 2004 12600 3648 12628
rect 2004 12588 2010 12600
rect 3694 12588 3700 12640
rect 3752 12628 3758 12640
rect 3881 12631 3939 12637
rect 3881 12628 3893 12631
rect 3752 12600 3893 12628
rect 3752 12588 3758 12600
rect 3881 12597 3893 12600
rect 3927 12597 3939 12631
rect 4908 12628 4936 12727
rect 6380 12696 6408 12727
rect 9490 12724 9496 12736
rect 9548 12724 9554 12776
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 10152 12736 10333 12764
rect 5552 12668 6408 12696
rect 5552 12628 5580 12668
rect 4908 12600 5580 12628
rect 3881 12591 3939 12597
rect 5902 12588 5908 12640
rect 5960 12588 5966 12640
rect 6380 12628 6408 12668
rect 10042 12656 10048 12708
rect 10100 12656 10106 12708
rect 6638 12628 6644 12640
rect 6380 12600 6644 12628
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 7377 12631 7435 12637
rect 7377 12628 7389 12631
rect 7156 12600 7389 12628
rect 7156 12588 7162 12600
rect 7377 12597 7389 12600
rect 7423 12597 7435 12631
rect 7377 12591 7435 12597
rect 9214 12588 9220 12640
rect 9272 12628 9278 12640
rect 9398 12628 9404 12640
rect 9272 12600 9404 12628
rect 9272 12588 9278 12600
rect 9398 12588 9404 12600
rect 9456 12588 9462 12640
rect 10152 12628 10180 12736
rect 10321 12733 10333 12736
rect 10367 12733 10379 12767
rect 10321 12727 10379 12733
rect 10410 12724 10416 12776
rect 10468 12773 10474 12776
rect 10468 12767 10496 12773
rect 10484 12733 10496 12767
rect 10468 12727 10496 12733
rect 10468 12724 10474 12727
rect 10594 12724 10600 12776
rect 10652 12724 10658 12776
rect 12621 12767 12679 12773
rect 12621 12733 12633 12767
rect 12667 12733 12679 12767
rect 12621 12727 12679 12733
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12764 12863 12767
rect 12851 12736 13216 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 11514 12656 11520 12708
rect 11572 12656 11578 12708
rect 12636 12696 12664 12727
rect 13078 12696 13084 12708
rect 12636 12668 13084 12696
rect 13078 12656 13084 12668
rect 13136 12656 13142 12708
rect 11532 12628 11560 12656
rect 10152 12600 11560 12628
rect 11606 12588 11612 12640
rect 11664 12628 11670 12640
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 11664 12600 11713 12628
rect 11664 12588 11670 12600
rect 11701 12597 11713 12600
rect 11747 12597 11759 12631
rect 13188 12628 13216 12736
rect 13262 12724 13268 12776
rect 13320 12724 13326 12776
rect 13998 12724 14004 12776
rect 14056 12764 14062 12776
rect 14568 12764 14596 12792
rect 14056 12736 14596 12764
rect 14056 12724 14062 12736
rect 17696 12705 17724 12872
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12832 17923 12835
rect 18224 12835 18282 12841
rect 18224 12832 18236 12835
rect 17911 12804 18236 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 18224 12801 18236 12804
rect 18270 12832 18282 12835
rect 18892 12832 18920 12872
rect 20548 12844 20576 12872
rect 24121 12869 24133 12872
rect 24167 12869 24179 12903
rect 24121 12863 24179 12869
rect 19613 12835 19671 12841
rect 19613 12832 19625 12835
rect 18270 12804 18920 12832
rect 19352 12804 19625 12832
rect 18270 12801 18282 12804
rect 18224 12795 18282 12801
rect 17954 12724 17960 12776
rect 18012 12724 18018 12776
rect 19352 12705 19380 12804
rect 19613 12801 19625 12804
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 20530 12792 20536 12844
rect 20588 12792 20594 12844
rect 20901 12835 20959 12841
rect 20901 12801 20913 12835
rect 20947 12801 20959 12835
rect 20901 12795 20959 12801
rect 20916 12764 20944 12795
rect 21174 12792 21180 12844
rect 21232 12792 21238 12844
rect 21358 12792 21364 12844
rect 21416 12792 21422 12844
rect 21450 12792 21456 12844
rect 21508 12832 21514 12844
rect 21637 12835 21695 12841
rect 21637 12832 21649 12835
rect 21508 12804 21649 12832
rect 21508 12792 21514 12804
rect 21637 12801 21649 12804
rect 21683 12801 21695 12835
rect 21637 12795 21695 12801
rect 22370 12792 22376 12844
rect 22428 12832 22434 12844
rect 23474 12832 23480 12844
rect 22428 12804 23480 12832
rect 22428 12792 22434 12804
rect 23474 12792 23480 12804
rect 23532 12792 23538 12844
rect 23569 12835 23627 12841
rect 23569 12801 23581 12835
rect 23615 12832 23627 12835
rect 25314 12832 25320 12844
rect 23615 12804 25320 12832
rect 23615 12801 23627 12804
rect 23569 12795 23627 12801
rect 25314 12792 25320 12804
rect 25372 12792 25378 12844
rect 20916 12736 21496 12764
rect 21468 12705 21496 12736
rect 17681 12699 17739 12705
rect 17681 12665 17693 12699
rect 17727 12665 17739 12699
rect 17681 12659 17739 12665
rect 19337 12699 19395 12705
rect 19337 12665 19349 12699
rect 19383 12665 19395 12699
rect 19337 12659 19395 12665
rect 21453 12699 21511 12705
rect 21453 12665 21465 12699
rect 21499 12665 21511 12699
rect 21453 12659 21511 12665
rect 25314 12656 25320 12708
rect 25372 12696 25378 12708
rect 25682 12696 25688 12708
rect 25372 12668 25688 12696
rect 25372 12656 25378 12668
rect 25682 12656 25688 12668
rect 25740 12656 25746 12708
rect 14550 12628 14556 12640
rect 13188 12600 14556 12628
rect 11701 12591 11759 12597
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 15562 12588 15568 12640
rect 15620 12588 15626 12640
rect 15654 12588 15660 12640
rect 15712 12628 15718 12640
rect 17494 12628 17500 12640
rect 15712 12600 17500 12628
rect 15712 12588 15718 12600
rect 17494 12588 17500 12600
rect 17552 12588 17558 12640
rect 20990 12588 20996 12640
rect 21048 12588 21054 12640
rect 21266 12588 21272 12640
rect 21324 12588 21330 12640
rect 23842 12588 23848 12640
rect 23900 12588 23906 12640
rect 1104 12538 24840 12560
rect 1104 12486 3917 12538
rect 3969 12486 3981 12538
rect 4033 12486 4045 12538
rect 4097 12486 4109 12538
rect 4161 12486 4173 12538
rect 4225 12486 9851 12538
rect 9903 12486 9915 12538
rect 9967 12486 9979 12538
rect 10031 12486 10043 12538
rect 10095 12486 10107 12538
rect 10159 12486 15785 12538
rect 15837 12486 15849 12538
rect 15901 12486 15913 12538
rect 15965 12486 15977 12538
rect 16029 12486 16041 12538
rect 16093 12486 21719 12538
rect 21771 12486 21783 12538
rect 21835 12486 21847 12538
rect 21899 12486 21911 12538
rect 21963 12486 21975 12538
rect 22027 12486 24840 12538
rect 1104 12464 24840 12486
rect 1394 12384 1400 12436
rect 1452 12384 1458 12436
rect 2682 12384 2688 12436
rect 2740 12384 2746 12436
rect 4522 12384 4528 12436
rect 4580 12424 4586 12436
rect 5166 12424 5172 12436
rect 4580 12396 5172 12424
rect 4580 12384 4586 12396
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 5534 12384 5540 12436
rect 5592 12384 5598 12436
rect 5902 12424 5908 12436
rect 5644 12396 5908 12424
rect 3602 12316 3608 12368
rect 3660 12356 3666 12368
rect 5350 12356 5356 12368
rect 3660 12328 5356 12356
rect 3660 12316 3666 12328
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 1486 12248 1492 12300
rect 1544 12288 1550 12300
rect 1673 12291 1731 12297
rect 1673 12288 1685 12291
rect 1544 12260 1685 12288
rect 1544 12248 1550 12260
rect 1673 12257 1685 12260
rect 1719 12257 1731 12291
rect 1673 12251 1731 12257
rect 2406 12248 2412 12300
rect 2464 12288 2470 12300
rect 5166 12288 5172 12300
rect 2464 12260 5172 12288
rect 2464 12248 2470 12260
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 5552 12288 5580 12384
rect 5644 12365 5672 12396
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 5994 12384 6000 12436
rect 6052 12424 6058 12436
rect 8757 12427 8815 12433
rect 8757 12424 8769 12427
rect 6052 12396 8769 12424
rect 6052 12384 6058 12396
rect 8757 12393 8769 12396
rect 8803 12393 8815 12427
rect 10870 12424 10876 12436
rect 8757 12387 8815 12393
rect 9784 12396 10876 12424
rect 5629 12359 5687 12365
rect 5629 12325 5641 12359
rect 5675 12325 5687 12359
rect 5629 12319 5687 12325
rect 6638 12316 6644 12368
rect 6696 12356 6702 12368
rect 6696 12328 7144 12356
rect 6696 12316 6702 12328
rect 6022 12291 6080 12297
rect 6022 12288 6034 12291
rect 5552 12260 6034 12288
rect 6022 12257 6034 12260
rect 6068 12257 6080 12291
rect 6022 12251 6080 12257
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12288 6239 12291
rect 7006 12288 7012 12300
rect 6227 12260 7012 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 7116 12297 7144 12328
rect 7558 12316 7564 12368
rect 7616 12316 7622 12368
rect 7101 12291 7159 12297
rect 7101 12257 7113 12291
rect 7147 12257 7159 12291
rect 7101 12251 7159 12257
rect 7466 12248 7472 12300
rect 7524 12288 7530 12300
rect 7524 12260 7972 12288
rect 7524 12248 7530 12260
rect 1581 12223 1639 12229
rect 1581 12189 1593 12223
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 1947 12223 2005 12229
rect 1947 12189 1959 12223
rect 1993 12220 2005 12223
rect 2314 12220 2320 12232
rect 1993 12192 2320 12220
rect 1993 12189 2005 12192
rect 1947 12183 2005 12189
rect 1302 12112 1308 12164
rect 1360 12152 1366 12164
rect 1596 12152 1624 12183
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 3881 12223 3939 12229
rect 2746 12192 3832 12220
rect 2746 12152 2774 12192
rect 1360 12124 1532 12152
rect 1596 12124 2774 12152
rect 1360 12112 1366 12124
rect 1504 12084 1532 12124
rect 3142 12112 3148 12164
rect 3200 12112 3206 12164
rect 3804 12152 3832 12192
rect 3881 12189 3893 12223
rect 3927 12220 3939 12223
rect 4614 12220 4620 12232
rect 3927 12192 4620 12220
rect 3927 12189 3939 12192
rect 3881 12183 3939 12189
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 4985 12223 5043 12229
rect 4985 12189 4997 12223
rect 5031 12220 5043 12223
rect 5074 12220 5080 12232
rect 5031 12192 5080 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 5902 12180 5908 12232
rect 5960 12180 5966 12232
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 4706 12152 4712 12164
rect 3804 12124 4712 12152
rect 4706 12112 4712 12124
rect 4764 12112 4770 12164
rect 3237 12087 3295 12093
rect 3237 12084 3249 12087
rect 1504 12056 3249 12084
rect 3237 12053 3249 12056
rect 3283 12053 3295 12087
rect 3237 12047 3295 12053
rect 3970 12044 3976 12096
rect 4028 12044 4034 12096
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 6825 12087 6883 12093
rect 6825 12084 6837 12087
rect 5224 12056 6837 12084
rect 5224 12044 5230 12056
rect 6825 12053 6837 12056
rect 6871 12053 6883 12087
rect 6932 12084 6960 12183
rect 7834 12180 7840 12232
rect 7892 12180 7898 12232
rect 7944 12229 7972 12260
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9490 12288 9496 12300
rect 9364 12260 9496 12288
rect 9364 12248 9370 12260
rect 9490 12248 9496 12260
rect 9548 12248 9554 12300
rect 9784 12297 9812 12396
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 12618 12384 12624 12436
rect 12676 12424 12682 12436
rect 13262 12424 13268 12436
rect 12676 12396 13268 12424
rect 12676 12384 12682 12396
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 15565 12427 15623 12433
rect 15565 12393 15577 12427
rect 15611 12424 15623 12427
rect 15654 12424 15660 12436
rect 15611 12396 15660 12424
rect 15611 12393 15623 12396
rect 15565 12387 15623 12393
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 16298 12384 16304 12436
rect 16356 12424 16362 12436
rect 16850 12424 16856 12436
rect 16356 12396 16856 12424
rect 16356 12384 16362 12396
rect 16850 12384 16856 12396
rect 16908 12424 16914 12436
rect 16908 12396 17172 12424
rect 16908 12384 16914 12396
rect 10781 12359 10839 12365
rect 10781 12325 10793 12359
rect 10827 12325 10839 12359
rect 10781 12319 10839 12325
rect 9769 12291 9827 12297
rect 9769 12257 9781 12291
rect 9815 12257 9827 12291
rect 10796 12288 10824 12319
rect 17034 12316 17040 12368
rect 17092 12316 17098 12368
rect 14280 12300 14332 12306
rect 10796 12260 11178 12288
rect 9769 12251 9827 12257
rect 13078 12248 13084 12300
rect 13136 12288 13142 12300
rect 13136 12260 13860 12288
rect 13136 12248 13142 12260
rect 7944 12223 8012 12229
rect 7944 12192 7966 12223
rect 7954 12189 7966 12192
rect 8000 12189 8012 12223
rect 7954 12183 8012 12189
rect 8110 12180 8116 12232
rect 8168 12180 8174 12232
rect 10042 12180 10048 12232
rect 10100 12180 10106 12232
rect 11698 12180 11704 12232
rect 11756 12180 11762 12232
rect 11974 12180 11980 12232
rect 12032 12180 12038 12232
rect 12069 12223 12127 12229
rect 12069 12189 12081 12223
rect 12115 12220 12127 12223
rect 12710 12220 12716 12232
rect 12115 12192 12716 12220
rect 12115 12189 12127 12192
rect 12069 12183 12127 12189
rect 12710 12180 12716 12192
rect 12768 12220 12774 12232
rect 13170 12220 13176 12232
rect 12768 12192 13176 12220
rect 12768 12180 12774 12192
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 11609 12155 11667 12161
rect 9732 12124 11468 12152
rect 9732 12112 9738 12124
rect 8202 12084 8208 12096
rect 6932 12056 8208 12084
rect 6825 12047 6883 12053
rect 8202 12044 8208 12056
rect 8260 12084 8266 12096
rect 8754 12084 8760 12096
rect 8260 12056 8760 12084
rect 8260 12044 8266 12056
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 11330 12044 11336 12096
rect 11388 12044 11394 12096
rect 11440 12084 11468 12124
rect 11609 12121 11621 12155
rect 11655 12152 11667 12155
rect 11992 12152 12020 12180
rect 13832 12152 13860 12260
rect 15378 12248 15384 12300
rect 15436 12288 15442 12300
rect 16298 12288 16304 12300
rect 15436 12260 16304 12288
rect 15436 12248 15442 12260
rect 16298 12248 16304 12260
rect 16356 12288 16362 12300
rect 16577 12291 16635 12297
rect 16577 12288 16589 12291
rect 16356 12260 16589 12288
rect 16356 12248 16362 12260
rect 16577 12257 16589 12260
rect 16623 12257 16635 12291
rect 17144 12288 17172 12396
rect 17310 12384 17316 12436
rect 17368 12424 17374 12436
rect 20441 12427 20499 12433
rect 17368 12396 20300 12424
rect 17368 12384 17374 12396
rect 18322 12316 18328 12368
rect 18380 12356 18386 12368
rect 19242 12356 19248 12368
rect 18380 12328 19248 12356
rect 18380 12316 18386 12328
rect 19242 12316 19248 12328
rect 19300 12316 19306 12368
rect 17313 12291 17371 12297
rect 17313 12288 17325 12291
rect 17144 12260 17325 12288
rect 16577 12251 16635 12257
rect 17313 12257 17325 12260
rect 17359 12257 17371 12291
rect 17313 12251 17371 12257
rect 17589 12291 17647 12297
rect 17589 12257 17601 12291
rect 17635 12288 17647 12291
rect 18138 12288 18144 12300
rect 17635 12260 18144 12288
rect 17635 12257 17647 12260
rect 17589 12251 17647 12257
rect 14280 12242 14332 12248
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12220 14703 12223
rect 15562 12220 15568 12232
rect 14691 12192 15568 12220
rect 14691 12189 14703 12192
rect 14645 12183 14703 12189
rect 15562 12180 15568 12192
rect 15620 12180 15626 12232
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 13906 12152 13912 12164
rect 11655 12124 12020 12152
rect 12082 12124 12664 12152
rect 13832 12124 13912 12152
rect 11655 12121 11667 12124
rect 11609 12115 11667 12121
rect 12082 12084 12110 12124
rect 11440 12056 12110 12084
rect 12434 12044 12440 12096
rect 12492 12044 12498 12096
rect 12636 12093 12664 12124
rect 13906 12112 13912 12124
rect 13964 12152 13970 12164
rect 14458 12152 14464 12164
rect 13964 12124 14464 12152
rect 13964 12112 13970 12124
rect 14458 12112 14464 12124
rect 14516 12152 14522 12164
rect 14553 12155 14611 12161
rect 14553 12152 14565 12155
rect 14516 12124 14565 12152
rect 14516 12112 14522 12124
rect 14553 12121 14565 12124
rect 14599 12121 14611 12155
rect 15013 12155 15071 12161
rect 15013 12152 15025 12155
rect 14553 12115 14611 12121
rect 14660 12124 15025 12152
rect 14660 12096 14688 12124
rect 15013 12121 15025 12124
rect 15059 12121 15071 12155
rect 15013 12115 15071 12121
rect 15194 12112 15200 12164
rect 15252 12152 15258 12164
rect 16408 12152 16436 12183
rect 15252 12124 16436 12152
rect 15252 12112 15258 12124
rect 12621 12087 12679 12093
rect 12621 12053 12633 12087
rect 12667 12053 12679 12087
rect 12621 12047 12679 12053
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 14090 12084 14096 12096
rect 13872 12056 14096 12084
rect 13872 12044 13878 12056
rect 14090 12044 14096 12056
rect 14148 12084 14154 12096
rect 14277 12087 14335 12093
rect 14277 12084 14289 12087
rect 14148 12056 14289 12084
rect 14148 12044 14154 12056
rect 14277 12053 14289 12056
rect 14323 12053 14335 12087
rect 14277 12047 14335 12053
rect 14642 12044 14648 12096
rect 14700 12044 14706 12096
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 14918 12084 14924 12096
rect 14792 12056 14924 12084
rect 14792 12044 14798 12056
rect 14918 12044 14924 12056
rect 14976 12084 14982 12096
rect 15381 12087 15439 12093
rect 15381 12084 15393 12087
rect 14976 12056 15393 12084
rect 14976 12044 14982 12056
rect 15381 12053 15393 12056
rect 15427 12053 15439 12087
rect 16592 12084 16620 12251
rect 18138 12248 18144 12260
rect 18196 12248 18202 12300
rect 17494 12229 17500 12232
rect 17451 12223 17500 12229
rect 17451 12189 17463 12223
rect 17497 12189 17500 12223
rect 17451 12183 17500 12189
rect 17494 12180 17500 12183
rect 17552 12180 17558 12232
rect 19426 12180 19432 12232
rect 19484 12180 19490 12232
rect 19703 12223 19761 12229
rect 19703 12189 19715 12223
rect 19749 12220 19761 12223
rect 20162 12220 20168 12232
rect 19749 12192 20168 12220
rect 19749 12189 19761 12192
rect 19703 12183 19761 12189
rect 20162 12180 20168 12192
rect 20220 12180 20226 12232
rect 20272 12220 20300 12396
rect 20441 12393 20453 12427
rect 20487 12424 20499 12427
rect 20714 12424 20720 12436
rect 20487 12396 20720 12424
rect 20487 12393 20499 12396
rect 20441 12387 20499 12393
rect 20714 12384 20720 12396
rect 20772 12424 20778 12436
rect 21174 12424 21180 12436
rect 20772 12396 21180 12424
rect 20772 12384 20778 12396
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 21542 12384 21548 12436
rect 21600 12424 21606 12436
rect 21600 12396 22094 12424
rect 21600 12384 21606 12396
rect 22066 12356 22094 12396
rect 22646 12384 22652 12436
rect 22704 12384 22710 12436
rect 22066 12328 22692 12356
rect 20806 12248 20812 12300
rect 20864 12248 20870 12300
rect 22002 12248 22008 12300
rect 22060 12248 22066 12300
rect 22020 12220 22048 12248
rect 22664 12232 22692 12328
rect 20272 12192 22048 12220
rect 22646 12180 22652 12232
rect 22704 12220 22710 12232
rect 22833 12223 22891 12229
rect 22833 12220 22845 12223
rect 22704 12192 22845 12220
rect 22704 12180 22710 12192
rect 22833 12189 22845 12192
rect 22879 12220 22891 12223
rect 22879 12192 22968 12220
rect 22879 12189 22891 12192
rect 22833 12183 22891 12189
rect 22940 12164 22968 12192
rect 23091 12193 23149 12199
rect 21082 12161 21088 12164
rect 21076 12152 21088 12161
rect 21043 12124 21088 12152
rect 21076 12115 21088 12124
rect 21140 12152 21146 12164
rect 21450 12152 21456 12164
rect 21140 12124 21456 12152
rect 21082 12112 21088 12115
rect 21140 12112 21146 12124
rect 21450 12112 21456 12124
rect 21508 12112 21514 12164
rect 21542 12112 21548 12164
rect 21600 12152 21606 12164
rect 22557 12155 22615 12161
rect 22557 12152 22569 12155
rect 21600 12124 22569 12152
rect 21600 12112 21606 12124
rect 22557 12121 22569 12124
rect 22603 12121 22615 12155
rect 22557 12115 22615 12121
rect 22922 12112 22928 12164
rect 22980 12112 22986 12164
rect 23091 12159 23103 12193
rect 23137 12190 23149 12193
rect 23137 12159 23152 12190
rect 23091 12153 23152 12159
rect 23124 12152 23152 12153
rect 23124 12124 25728 12152
rect 18046 12084 18052 12096
rect 16592 12056 18052 12084
rect 15381 12047 15439 12053
rect 18046 12044 18052 12056
rect 18104 12044 18110 12096
rect 18230 12044 18236 12096
rect 18288 12044 18294 12096
rect 22186 12044 22192 12096
rect 22244 12044 22250 12096
rect 22462 12044 22468 12096
rect 22520 12084 22526 12096
rect 23124 12084 23152 12124
rect 25700 12096 25728 12124
rect 22520 12056 23152 12084
rect 22520 12044 22526 12056
rect 23842 12044 23848 12096
rect 23900 12044 23906 12096
rect 25682 12044 25688 12096
rect 25740 12044 25746 12096
rect 1104 11994 25000 12016
rect 1104 11942 6884 11994
rect 6936 11942 6948 11994
rect 7000 11942 7012 11994
rect 7064 11942 7076 11994
rect 7128 11942 7140 11994
rect 7192 11942 12818 11994
rect 12870 11942 12882 11994
rect 12934 11942 12946 11994
rect 12998 11942 13010 11994
rect 13062 11942 13074 11994
rect 13126 11942 18752 11994
rect 18804 11942 18816 11994
rect 18868 11942 18880 11994
rect 18932 11942 18944 11994
rect 18996 11942 19008 11994
rect 19060 11942 24686 11994
rect 24738 11942 24750 11994
rect 24802 11942 24814 11994
rect 24866 11942 24878 11994
rect 24930 11942 24942 11994
rect 24994 11942 25000 11994
rect 1104 11920 25000 11942
rect 1486 11840 1492 11892
rect 1544 11880 1550 11892
rect 1544 11852 3096 11880
rect 1544 11840 1550 11852
rect 2130 11812 2136 11824
rect 1504 11784 2136 11812
rect 1504 11753 1532 11784
rect 2130 11772 2136 11784
rect 2188 11772 2194 11824
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11713 1547 11747
rect 2283 11747 2341 11753
rect 2283 11744 2295 11747
rect 1489 11707 1547 11713
rect 1688 11716 2295 11744
rect 106 11636 112 11688
rect 164 11676 170 11688
rect 1688 11676 1716 11716
rect 2283 11713 2295 11716
rect 2329 11744 2341 11747
rect 2866 11744 2872 11756
rect 2329 11716 2872 11744
rect 2329 11713 2341 11716
rect 2283 11707 2341 11713
rect 2866 11704 2872 11716
rect 2924 11704 2930 11756
rect 164 11648 1716 11676
rect 1765 11679 1823 11685
rect 164 11636 170 11648
rect 1765 11645 1777 11679
rect 1811 11676 1823 11679
rect 1854 11676 1860 11688
rect 1811 11648 1860 11676
rect 1811 11645 1823 11648
rect 1765 11639 1823 11645
rect 1854 11636 1860 11648
rect 1912 11636 1918 11688
rect 2041 11679 2099 11685
rect 2041 11645 2053 11679
rect 2087 11645 2099 11679
rect 3068 11676 3096 11852
rect 3142 11840 3148 11892
rect 3200 11880 3206 11892
rect 3421 11883 3479 11889
rect 3421 11880 3433 11883
rect 3200 11852 3433 11880
rect 3200 11840 3206 11852
rect 3421 11849 3433 11852
rect 3467 11849 3479 11883
rect 3421 11843 3479 11849
rect 5166 11840 5172 11892
rect 5224 11840 5230 11892
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 5994 11880 6000 11892
rect 5316 11852 6000 11880
rect 5316 11840 5322 11852
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 6546 11840 6552 11892
rect 6604 11880 6610 11892
rect 6604 11852 7512 11880
rect 6604 11840 6610 11852
rect 5184 11812 5212 11840
rect 7374 11812 7380 11824
rect 3620 11784 5212 11812
rect 7116 11784 7380 11812
rect 3620 11753 3648 11784
rect 7116 11783 7144 11784
rect 7083 11777 7144 11783
rect 3605 11747 3663 11753
rect 3605 11713 3617 11747
rect 3651 11713 3663 11747
rect 3605 11707 3663 11713
rect 3971 11747 4029 11753
rect 3971 11713 3983 11747
rect 4017 11744 4029 11747
rect 4062 11744 4068 11756
rect 4017 11716 4068 11744
rect 4017 11713 4029 11716
rect 3971 11707 4029 11713
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 4338 11704 4344 11756
rect 4396 11744 4402 11756
rect 5442 11744 5448 11756
rect 4396 11716 5448 11744
rect 4396 11704 4402 11716
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 7083 11743 7095 11777
rect 7129 11746 7144 11777
rect 7374 11772 7380 11784
rect 7432 11772 7438 11824
rect 7129 11743 7141 11746
rect 7083 11737 7141 11743
rect 7484 11744 7512 11852
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 7837 11883 7895 11889
rect 7837 11880 7849 11883
rect 7616 11852 7849 11880
rect 7616 11840 7622 11852
rect 7837 11849 7849 11852
rect 7883 11849 7895 11883
rect 7837 11843 7895 11849
rect 8110 11840 8116 11892
rect 8168 11880 8174 11892
rect 9217 11883 9275 11889
rect 9217 11880 9229 11883
rect 8168 11852 9229 11880
rect 8168 11840 8174 11852
rect 9217 11849 9229 11852
rect 9263 11849 9275 11883
rect 9217 11843 9275 11849
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 10318 11880 10324 11892
rect 10100 11852 10324 11880
rect 10100 11840 10106 11852
rect 10318 11840 10324 11852
rect 10376 11840 10382 11892
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 10652 11852 10701 11880
rect 10652 11840 10658 11852
rect 10689 11849 10701 11852
rect 10735 11849 10747 11883
rect 10689 11843 10747 11849
rect 10796 11852 14228 11880
rect 8754 11772 8760 11824
rect 8812 11812 8818 11824
rect 10796 11812 10824 11852
rect 8812 11784 10824 11812
rect 8812 11772 8818 11784
rect 12342 11772 12348 11824
rect 12400 11772 12406 11824
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 13170 11812 13176 11824
rect 12492 11784 13176 11812
rect 12492 11772 12498 11784
rect 13170 11772 13176 11784
rect 13228 11772 13234 11824
rect 13372 11784 14044 11812
rect 8447 11747 8505 11753
rect 8447 11744 8459 11747
rect 7484 11716 8459 11744
rect 8447 11713 8459 11716
rect 8493 11713 8505 11747
rect 9919 11747 9977 11753
rect 9919 11744 9931 11747
rect 8447 11707 8505 11713
rect 9600 11716 9931 11744
rect 9600 11688 9628 11716
rect 9919 11713 9931 11716
rect 9965 11744 9977 11747
rect 10962 11744 10968 11756
rect 9965 11716 10968 11744
rect 9965 11713 9977 11716
rect 9919 11707 9977 11713
rect 10962 11704 10968 11716
rect 11020 11744 11026 11756
rect 12360 11744 12388 11772
rect 13372 11753 13400 11784
rect 14016 11756 14044 11784
rect 11020 11716 12388 11744
rect 13357 11747 13415 11753
rect 11020 11704 11026 11716
rect 13357 11713 13369 11747
rect 13403 11713 13415 11747
rect 13630 11744 13636 11756
rect 13591 11716 13636 11744
rect 13357 11707 13415 11713
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 13998 11704 14004 11756
rect 14056 11704 14062 11756
rect 3697 11679 3755 11685
rect 3697 11676 3709 11679
rect 3068 11648 3709 11676
rect 2041 11639 2099 11645
rect 3697 11645 3709 11648
rect 3743 11645 3755 11679
rect 3697 11639 3755 11645
rect 2056 11540 2084 11639
rect 2406 11540 2412 11552
rect 2056 11512 2412 11540
rect 2406 11500 2412 11512
rect 2464 11500 2470 11552
rect 3050 11500 3056 11552
rect 3108 11500 3114 11552
rect 3712 11540 3740 11639
rect 4614 11636 4620 11688
rect 4672 11676 4678 11688
rect 5534 11676 5540 11688
rect 4672 11648 5540 11676
rect 4672 11636 4678 11648
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 8205 11679 8263 11685
rect 8205 11645 8217 11679
rect 8251 11645 8263 11679
rect 8205 11639 8263 11645
rect 4798 11568 4804 11620
rect 4856 11608 4862 11620
rect 5074 11608 5080 11620
rect 4856 11580 5080 11608
rect 4856 11568 4862 11580
rect 5074 11568 5080 11580
rect 5132 11568 5138 11620
rect 4154 11540 4160 11552
rect 3712 11512 4160 11540
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 4709 11543 4767 11549
rect 4709 11540 4721 11543
rect 4672 11512 4721 11540
rect 4672 11500 4678 11512
rect 4709 11509 4721 11512
rect 4755 11509 4767 11543
rect 6840 11540 6868 11639
rect 8220 11540 8248 11639
rect 9582 11636 9588 11688
rect 9640 11636 9646 11688
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11645 9735 11679
rect 9677 11639 9735 11645
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 9692 11608 9720 11639
rect 10778 11636 10784 11688
rect 10836 11636 10842 11688
rect 10796 11608 10824 11636
rect 13078 11608 13084 11620
rect 8996 11580 9720 11608
rect 10334 11580 13084 11608
rect 8996 11568 9002 11580
rect 9214 11540 9220 11552
rect 6840 11512 9220 11540
rect 4709 11503 4767 11509
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 9646 11540 9674 11580
rect 10334 11540 10362 11580
rect 13078 11568 13084 11580
rect 13136 11568 13142 11620
rect 9646 11512 10362 11540
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 13446 11540 13452 11552
rect 10836 11512 13452 11540
rect 10836 11500 10842 11512
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 14200 11540 14228 11852
rect 14274 11840 14280 11892
rect 14332 11880 14338 11892
rect 14369 11883 14427 11889
rect 14369 11880 14381 11883
rect 14332 11852 14381 11880
rect 14332 11840 14338 11852
rect 14369 11849 14381 11852
rect 14415 11849 14427 11883
rect 14369 11843 14427 11849
rect 16942 11840 16948 11892
rect 17000 11880 17006 11892
rect 17000 11852 17724 11880
rect 17000 11840 17006 11852
rect 14458 11772 14464 11824
rect 14516 11812 14522 11824
rect 17310 11812 17316 11824
rect 14516 11784 17316 11812
rect 14516 11772 14522 11784
rect 17310 11772 17316 11784
rect 17368 11772 17374 11824
rect 17696 11756 17724 11852
rect 18138 11840 18144 11892
rect 18196 11840 18202 11892
rect 18322 11840 18328 11892
rect 18380 11880 18386 11892
rect 18380 11852 19334 11880
rect 18380 11840 18386 11852
rect 18156 11812 18184 11840
rect 19306 11812 19334 11852
rect 21358 11840 21364 11892
rect 21416 11880 21422 11892
rect 21821 11883 21879 11889
rect 21821 11880 21833 11883
rect 21416 11852 21833 11880
rect 21416 11840 21422 11852
rect 21821 11849 21833 11852
rect 21867 11849 21879 11883
rect 21821 11843 21879 11849
rect 22186 11840 22192 11892
rect 22244 11840 22250 11892
rect 22373 11883 22431 11889
rect 22373 11849 22385 11883
rect 22419 11880 22431 11883
rect 23750 11880 23756 11892
rect 22419 11852 23756 11880
rect 22419 11849 22431 11852
rect 22373 11843 22431 11849
rect 23750 11840 23756 11852
rect 23808 11840 23814 11892
rect 23842 11840 23848 11892
rect 23900 11840 23906 11892
rect 24394 11840 24400 11892
rect 24452 11840 24458 11892
rect 21910 11812 21916 11824
rect 18156 11784 18460 11812
rect 19306 11784 21916 11812
rect 14274 11704 14280 11756
rect 14332 11744 14338 11756
rect 16482 11744 16488 11756
rect 14332 11716 16488 11744
rect 14332 11704 14338 11716
rect 16482 11704 16488 11716
rect 16540 11744 16546 11756
rect 16911 11747 16969 11753
rect 16911 11744 16923 11747
rect 16540 11716 16923 11744
rect 16540 11704 16546 11716
rect 16911 11713 16923 11716
rect 16957 11713 16969 11747
rect 16911 11707 16969 11713
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17092 11716 17356 11744
rect 17092 11704 17098 11716
rect 14642 11636 14648 11688
rect 14700 11676 14706 11688
rect 16666 11676 16672 11688
rect 14700 11648 16672 11676
rect 14700 11636 14706 11648
rect 16666 11636 16672 11648
rect 16724 11636 16730 11688
rect 17328 11608 17356 11716
rect 17678 11704 17684 11756
rect 17736 11744 17742 11756
rect 18323 11747 18381 11753
rect 18323 11744 18335 11747
rect 17736 11716 18335 11744
rect 17736 11704 17742 11716
rect 18323 11713 18335 11716
rect 18369 11713 18381 11747
rect 18432 11744 18460 11784
rect 21910 11772 21916 11784
rect 21968 11772 21974 11824
rect 18432 11716 19104 11744
rect 18323 11707 18381 11713
rect 17494 11636 17500 11688
rect 17552 11676 17558 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 17552 11648 18061 11676
rect 17552 11636 17558 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 19076 11617 19104 11716
rect 20714 11704 20720 11756
rect 20772 11704 20778 11756
rect 20990 11704 20996 11756
rect 21048 11704 21054 11756
rect 21358 11704 21364 11756
rect 21416 11704 21422 11756
rect 22005 11747 22063 11753
rect 22005 11713 22017 11747
rect 22051 11744 22063 11747
rect 22204 11744 22232 11840
rect 23860 11812 23888 11840
rect 22664 11784 23888 11812
rect 22051 11716 22232 11744
rect 22557 11747 22615 11753
rect 22051 11713 22063 11716
rect 22005 11707 22063 11713
rect 22557 11713 22569 11747
rect 22603 11744 22615 11747
rect 22664 11744 22692 11784
rect 22603 11716 22692 11744
rect 22603 11713 22615 11716
rect 22557 11707 22615 11713
rect 22830 11704 22836 11756
rect 22888 11744 22894 11756
rect 22923 11747 22981 11753
rect 22923 11744 22935 11747
rect 22888 11716 22935 11744
rect 22888 11704 22894 11716
rect 22923 11713 22935 11716
rect 22969 11713 22981 11747
rect 22923 11707 22981 11713
rect 23474 11704 23480 11756
rect 23532 11744 23538 11756
rect 24213 11747 24271 11753
rect 24213 11744 24225 11747
rect 23532 11716 24225 11744
rect 23532 11704 23538 11716
rect 24213 11713 24225 11716
rect 24259 11713 24271 11747
rect 24213 11707 24271 11713
rect 19242 11636 19248 11688
rect 19300 11676 19306 11688
rect 19300 11648 21496 11676
rect 19300 11636 19306 11648
rect 17681 11611 17739 11617
rect 17681 11608 17693 11611
rect 17328 11580 17693 11608
rect 17681 11577 17693 11580
rect 17727 11577 17739 11611
rect 17681 11571 17739 11577
rect 19061 11611 19119 11617
rect 19061 11577 19073 11611
rect 19107 11577 19119 11611
rect 19061 11571 19119 11577
rect 21361 11611 21419 11617
rect 21361 11577 21373 11611
rect 21407 11577 21419 11611
rect 21468 11608 21496 11648
rect 22462 11636 22468 11688
rect 22520 11636 22526 11688
rect 22646 11636 22652 11688
rect 22704 11636 22710 11688
rect 22480 11608 22508 11636
rect 21468 11580 22508 11608
rect 21361 11571 21419 11577
rect 21376 11540 21404 11571
rect 14200 11512 21404 11540
rect 22462 11500 22468 11552
rect 22520 11540 22526 11552
rect 23474 11540 23480 11552
rect 22520 11512 23480 11540
rect 22520 11500 22526 11512
rect 23474 11500 23480 11512
rect 23532 11500 23538 11552
rect 23658 11500 23664 11552
rect 23716 11500 23722 11552
rect 1104 11450 24840 11472
rect 1104 11398 3917 11450
rect 3969 11398 3981 11450
rect 4033 11398 4045 11450
rect 4097 11398 4109 11450
rect 4161 11398 4173 11450
rect 4225 11398 9851 11450
rect 9903 11398 9915 11450
rect 9967 11398 9979 11450
rect 10031 11398 10043 11450
rect 10095 11398 10107 11450
rect 10159 11398 15785 11450
rect 15837 11398 15849 11450
rect 15901 11398 15913 11450
rect 15965 11398 15977 11450
rect 16029 11398 16041 11450
rect 16093 11398 21719 11450
rect 21771 11398 21783 11450
rect 21835 11398 21847 11450
rect 21899 11398 21911 11450
rect 21963 11398 21975 11450
rect 22027 11398 24840 11450
rect 1104 11376 24840 11398
rect 1762 11296 1768 11348
rect 1820 11296 1826 11348
rect 1854 11296 1860 11348
rect 1912 11336 1918 11348
rect 2222 11336 2228 11348
rect 1912 11308 2228 11336
rect 1912 11296 1918 11308
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 3050 11336 3056 11348
rect 2424 11308 3056 11336
rect 750 11160 756 11212
rect 808 11160 814 11212
rect 1780 11200 1808 11296
rect 2424 11277 2452 11308
rect 3050 11296 3056 11308
rect 3108 11296 3114 11348
rect 4614 11296 4620 11348
rect 4672 11296 4678 11348
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 10137 11339 10195 11345
rect 5868 11308 10088 11336
rect 5868 11296 5874 11308
rect 2409 11271 2467 11277
rect 2409 11237 2421 11271
rect 2455 11237 2467 11271
rect 2409 11231 2467 11237
rect 4525 11271 4583 11277
rect 4525 11237 4537 11271
rect 4571 11268 4583 11271
rect 4632 11268 4660 11296
rect 4571 11240 4660 11268
rect 4571 11237 4583 11240
rect 4525 11231 4583 11237
rect 7374 11228 7380 11280
rect 7432 11268 7438 11280
rect 8294 11268 8300 11280
rect 7432 11240 8300 11268
rect 7432 11228 7438 11240
rect 8294 11228 8300 11240
rect 8352 11228 8358 11280
rect 10060 11268 10088 11308
rect 10137 11305 10149 11339
rect 10183 11336 10195 11339
rect 10226 11336 10232 11348
rect 10183 11308 10232 11336
rect 10183 11305 10195 11308
rect 10137 11299 10195 11305
rect 10226 11296 10232 11308
rect 10284 11296 10290 11348
rect 17037 11339 17095 11345
rect 17037 11336 17049 11339
rect 10336 11308 17049 11336
rect 10336 11268 10364 11308
rect 17037 11305 17049 11308
rect 17083 11305 17095 11339
rect 18141 11339 18199 11345
rect 18141 11336 18153 11339
rect 17037 11299 17095 11305
rect 17144 11308 18153 11336
rect 10060 11240 10364 11268
rect 12434 11228 12440 11280
rect 12492 11268 12498 11280
rect 14274 11268 14280 11280
rect 12492 11240 14280 11268
rect 12492 11228 12498 11240
rect 14274 11228 14280 11240
rect 14332 11228 14338 11280
rect 15304 11240 15976 11268
rect 15304 11212 15332 11240
rect 1596 11172 1808 11200
rect 2823 11203 2881 11209
rect 768 11064 796 11160
rect 1596 11141 1624 11172
rect 2823 11169 2835 11203
rect 2869 11200 2881 11203
rect 3326 11200 3332 11212
rect 2869 11172 3332 11200
rect 2869 11169 2881 11172
rect 2823 11163 2881 11169
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 3605 11203 3663 11209
rect 3605 11169 3617 11203
rect 3651 11200 3663 11203
rect 4246 11200 4252 11212
rect 3651 11172 4252 11200
rect 3651 11169 3663 11172
rect 3605 11163 3663 11169
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 4798 11160 4804 11212
rect 4856 11160 4862 11212
rect 4982 11209 4988 11212
rect 4939 11203 4988 11209
rect 4939 11169 4951 11203
rect 4985 11169 4988 11203
rect 4939 11163 4988 11169
rect 4982 11160 4988 11163
rect 5040 11160 5046 11212
rect 5626 11160 5632 11212
rect 5684 11200 5690 11212
rect 5994 11200 6000 11212
rect 5684 11172 6000 11200
rect 5684 11160 5690 11172
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 6638 11160 6644 11212
rect 6696 11200 6702 11212
rect 7466 11200 7472 11212
rect 6696 11172 7472 11200
rect 6696 11160 6702 11172
rect 7466 11160 7472 11172
rect 7524 11200 7530 11212
rect 8754 11200 8760 11212
rect 7524 11172 8760 11200
rect 7524 11160 7530 11172
rect 8754 11160 8760 11172
rect 8812 11160 8818 11212
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 11146 11200 11152 11212
rect 10192 11172 11152 11200
rect 10192 11160 10198 11172
rect 11146 11160 11152 11172
rect 11204 11200 11210 11212
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 11204 11172 11713 11200
rect 11204 11160 11210 11172
rect 11701 11169 11713 11172
rect 11747 11169 11759 11203
rect 11701 11163 11759 11169
rect 13078 11160 13084 11212
rect 13136 11200 13142 11212
rect 14642 11200 14648 11212
rect 13136 11172 14648 11200
rect 13136 11160 13142 11172
rect 14642 11160 14648 11172
rect 14700 11160 14706 11212
rect 15286 11160 15292 11212
rect 15344 11160 15350 11212
rect 15838 11160 15844 11212
rect 15896 11160 15902 11212
rect 15948 11200 15976 11240
rect 16393 11203 16451 11209
rect 15948 11172 16277 11200
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11101 1639 11135
rect 1581 11095 1639 11101
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11132 1823 11135
rect 1854 11132 1860 11144
rect 1811 11104 1860 11132
rect 1811 11101 1823 11104
rect 1765 11095 1823 11101
rect 1854 11092 1860 11104
rect 1912 11092 1918 11144
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11101 2007 11135
rect 1949 11095 2007 11101
rect 1964 11064 1992 11095
rect 2682 11092 2688 11144
rect 2740 11092 2746 11144
rect 2958 11092 2964 11144
rect 3016 11092 3022 11144
rect 3878 11092 3884 11144
rect 3936 11092 3942 11144
rect 3970 11092 3976 11144
rect 4028 11132 4034 11144
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 4028 11104 4077 11132
rect 4028 11092 4034 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 5074 11092 5080 11144
rect 5132 11092 5138 11144
rect 6362 11092 6368 11144
rect 6420 11132 6426 11144
rect 7650 11132 7656 11144
rect 6420 11104 7656 11132
rect 6420 11092 6426 11104
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 8018 11092 8024 11144
rect 8076 11132 8082 11144
rect 8938 11132 8944 11144
rect 8076 11104 8944 11132
rect 8076 11092 8082 11104
rect 8938 11092 8944 11104
rect 8996 11132 9002 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8996 11104 9137 11132
rect 8996 11092 9002 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 11975 11135 12033 11141
rect 9125 11095 9183 11101
rect 9383 11105 9441 11111
rect 3988 11064 4016 11092
rect 768 11036 1992 11064
rect 1394 10956 1400 11008
rect 1452 10956 1458 11008
rect 1964 10996 1992 11036
rect 3436 11036 4016 11064
rect 3436 10996 3464 11036
rect 5626 11024 5632 11076
rect 5684 11064 5690 11076
rect 5721 11067 5779 11073
rect 5721 11064 5733 11067
rect 5684 11036 5733 11064
rect 5684 11024 5690 11036
rect 5721 11033 5733 11036
rect 5767 11033 5779 11067
rect 5721 11027 5779 11033
rect 6546 11024 6552 11076
rect 6604 11064 6610 11076
rect 7558 11064 7564 11076
rect 6604 11036 7564 11064
rect 6604 11024 6610 11036
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 9383 11071 9395 11105
rect 9429 11102 9441 11105
rect 9429 11071 9444 11102
rect 11975 11101 11987 11135
rect 12021 11132 12033 11135
rect 15010 11132 15016 11144
rect 12021 11104 15016 11132
rect 12021 11101 12033 11104
rect 11975 11095 12033 11101
rect 15010 11092 15016 11104
rect 15068 11092 15074 11144
rect 15194 11092 15200 11144
rect 15252 11092 15258 11144
rect 15378 11092 15384 11144
rect 15436 11092 15442 11144
rect 16114 11092 16120 11144
rect 16172 11092 16178 11144
rect 16249 11141 16277 11172
rect 16393 11169 16405 11203
rect 16439 11200 16451 11203
rect 17144 11200 17172 11308
rect 18141 11305 18153 11308
rect 18187 11305 18199 11339
rect 18141 11299 18199 11305
rect 22189 11339 22247 11345
rect 22189 11305 22201 11339
rect 22235 11336 22247 11339
rect 22462 11336 22468 11348
rect 22235 11308 22468 11336
rect 22235 11305 22247 11308
rect 22189 11299 22247 11305
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 23658 11336 23664 11348
rect 22664 11308 23664 11336
rect 16439 11172 17172 11200
rect 16439 11169 16451 11172
rect 16393 11163 16451 11169
rect 16234 11135 16292 11141
rect 16234 11101 16246 11135
rect 16280 11101 16292 11135
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 16234 11095 16292 11101
rect 16960 11104 17141 11132
rect 16960 11076 16988 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17129 11095 17187 11101
rect 17371 11135 17429 11141
rect 17371 11101 17383 11135
rect 17417 11101 17429 11135
rect 17371 11095 17429 11101
rect 9383 11065 9444 11071
rect 9416 11064 9444 11065
rect 9490 11064 9496 11076
rect 9416 11036 9496 11064
rect 9490 11024 9496 11036
rect 9548 11064 9554 11076
rect 10502 11064 10508 11076
rect 9548 11036 10508 11064
rect 9548 11024 9554 11036
rect 10502 11024 10508 11036
rect 10560 11024 10566 11076
rect 11992 11036 12848 11064
rect 1964 10968 3464 10996
rect 4982 10956 4988 11008
rect 5040 10996 5046 11008
rect 11992 10996 12020 11036
rect 5040 10968 12020 10996
rect 5040 10956 5046 10968
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 12713 10999 12771 11005
rect 12713 10996 12725 10999
rect 12124 10968 12725 10996
rect 12124 10956 12130 10968
rect 12713 10965 12725 10968
rect 12759 10965 12771 10999
rect 12820 10996 12848 11036
rect 16942 11024 16948 11076
rect 17000 11024 17006 11076
rect 17218 11024 17224 11076
rect 17276 11064 17282 11076
rect 17386 11064 17414 11095
rect 17770 11092 17776 11144
rect 17828 11132 17834 11144
rect 17828 11104 19196 11132
rect 17828 11092 17834 11104
rect 17276 11036 17414 11064
rect 17276 11024 17282 11036
rect 18230 11024 18236 11076
rect 18288 11024 18294 11076
rect 19168 11064 19196 11104
rect 19242 11092 19248 11144
rect 19300 11092 19306 11144
rect 19519 11135 19577 11141
rect 19519 11132 19531 11135
rect 19343 11104 19531 11132
rect 19343 11064 19371 11104
rect 19519 11101 19531 11104
rect 19565 11132 19577 11135
rect 22094 11132 22100 11144
rect 19565 11104 22100 11132
rect 19565 11101 19577 11104
rect 19519 11095 19577 11101
rect 22094 11092 22100 11104
rect 22152 11092 22158 11144
rect 22664 11141 22692 11308
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 22373 11135 22431 11141
rect 22373 11101 22385 11135
rect 22419 11101 22431 11135
rect 22373 11095 22431 11101
rect 22649 11135 22707 11141
rect 22649 11101 22661 11135
rect 22695 11101 22707 11135
rect 22649 11095 22707 11101
rect 22741 11135 22799 11141
rect 22741 11101 22753 11135
rect 22787 11132 22799 11135
rect 22922 11132 22928 11144
rect 22787 11104 22928 11132
rect 22787 11101 22799 11104
rect 22741 11095 22799 11101
rect 19168 11036 19371 11064
rect 22388 11064 22416 11095
rect 22922 11092 22928 11104
rect 22980 11092 22986 11144
rect 23014 11092 23020 11144
rect 23072 11092 23078 11144
rect 22388 11036 23796 11064
rect 18248 10996 18276 11024
rect 12820 10968 18276 10996
rect 12713 10959 12771 10965
rect 19334 10956 19340 11008
rect 19392 10996 19398 11008
rect 20257 10999 20315 11005
rect 20257 10996 20269 10999
rect 19392 10968 20269 10996
rect 19392 10956 19398 10968
rect 20257 10965 20269 10968
rect 20303 10965 20315 10999
rect 20257 10959 20315 10965
rect 22465 10999 22523 11005
rect 22465 10965 22477 10999
rect 22511 10996 22523 10999
rect 23658 10996 23664 11008
rect 22511 10968 23664 10996
rect 22511 10965 22523 10968
rect 22465 10959 22523 10965
rect 23658 10956 23664 10968
rect 23716 10956 23722 11008
rect 23768 11005 23796 11036
rect 23753 10999 23811 11005
rect 23753 10965 23765 10999
rect 23799 10965 23811 10999
rect 23753 10959 23811 10965
rect 1104 10906 25000 10928
rect 1104 10854 6884 10906
rect 6936 10854 6948 10906
rect 7000 10854 7012 10906
rect 7064 10854 7076 10906
rect 7128 10854 7140 10906
rect 7192 10854 12818 10906
rect 12870 10854 12882 10906
rect 12934 10854 12946 10906
rect 12998 10854 13010 10906
rect 13062 10854 13074 10906
rect 13126 10854 18752 10906
rect 18804 10854 18816 10906
rect 18868 10854 18880 10906
rect 18932 10854 18944 10906
rect 18996 10854 19008 10906
rect 19060 10854 24686 10906
rect 24738 10854 24750 10906
rect 24802 10854 24814 10906
rect 24866 10854 24878 10906
rect 24930 10854 24942 10906
rect 24994 10854 25000 10906
rect 1104 10832 25000 10854
rect 1949 10795 2007 10801
rect 1949 10792 1961 10795
rect 1504 10764 1961 10792
rect 1504 10733 1532 10764
rect 1949 10761 1961 10764
rect 1995 10761 2007 10795
rect 1949 10755 2007 10761
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 3421 10795 3479 10801
rect 3421 10792 3433 10795
rect 3016 10764 3433 10792
rect 3016 10752 3022 10764
rect 3421 10761 3433 10764
rect 3467 10761 3479 10795
rect 4982 10792 4988 10804
rect 3421 10755 3479 10761
rect 3528 10764 4988 10792
rect 1489 10727 1547 10733
rect 1489 10693 1501 10727
rect 1535 10693 1547 10727
rect 3528 10724 3556 10764
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 5074 10752 5080 10804
rect 5132 10792 5138 10804
rect 5261 10795 5319 10801
rect 5261 10792 5273 10795
rect 5132 10764 5273 10792
rect 5132 10752 5138 10764
rect 5261 10761 5273 10764
rect 5307 10761 5319 10795
rect 5261 10755 5319 10761
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5592 10764 5641 10792
rect 5592 10752 5598 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 5629 10755 5687 10761
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 11790 10792 11796 10804
rect 5960 10764 11796 10792
rect 5960 10752 5966 10764
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 12250 10752 12256 10804
rect 12308 10792 12314 10804
rect 12989 10795 13047 10801
rect 12989 10792 13001 10795
rect 12308 10764 13001 10792
rect 12308 10752 12314 10764
rect 12989 10761 13001 10764
rect 13035 10792 13047 10795
rect 13538 10792 13544 10804
rect 13035 10764 13544 10792
rect 13035 10761 13047 10764
rect 12989 10755 13047 10761
rect 13538 10752 13544 10764
rect 13596 10752 13602 10804
rect 14182 10792 14188 10804
rect 13832 10764 14188 10792
rect 10134 10724 10140 10736
rect 1489 10687 1547 10693
rect 2148 10696 3556 10724
rect 3896 10696 4534 10724
rect 2148 10665 2176 10696
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10625 2191 10659
rect 2133 10619 2191 10625
rect 2590 10616 2596 10668
rect 2648 10656 2654 10668
rect 2683 10659 2741 10665
rect 2683 10656 2695 10659
rect 2648 10628 2695 10656
rect 2648 10616 2654 10628
rect 2683 10625 2695 10628
rect 2729 10656 2741 10659
rect 3896 10656 3924 10696
rect 4506 10695 4534 10696
rect 10060 10696 10140 10724
rect 4506 10689 4565 10695
rect 2729 10628 3924 10656
rect 2729 10625 2741 10628
rect 2683 10619 2741 10625
rect 3970 10616 3976 10668
rect 4028 10616 4034 10668
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4249 10659 4307 10665
rect 4249 10656 4261 10659
rect 4212 10628 4261 10656
rect 4212 10616 4218 10628
rect 4249 10625 4261 10628
rect 4295 10625 4307 10659
rect 4506 10658 4519 10689
rect 4507 10655 4519 10658
rect 4553 10655 4565 10689
rect 4507 10649 4565 10655
rect 4249 10619 4307 10625
rect 5810 10616 5816 10668
rect 5868 10616 5874 10668
rect 6365 10659 6423 10665
rect 6365 10625 6377 10659
rect 6411 10656 6423 10659
rect 6730 10656 6736 10668
rect 6411 10628 6736 10656
rect 6411 10625 6423 10628
rect 6365 10619 6423 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 7423 10659 7481 10665
rect 7423 10625 7435 10659
rect 7469 10625 7481 10659
rect 7423 10619 7481 10625
rect 2406 10548 2412 10600
rect 2464 10548 2470 10600
rect 3694 10548 3700 10600
rect 3752 10588 3758 10600
rect 4062 10588 4068 10600
rect 3752 10560 4068 10588
rect 3752 10548 3758 10560
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 6546 10548 6552 10600
rect 6604 10548 6610 10600
rect 7282 10548 7288 10600
rect 7340 10548 7346 10600
rect 7438 10588 7466 10619
rect 7558 10616 7564 10668
rect 7616 10616 7622 10668
rect 10060 10665 10088 10696
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 11606 10724 11612 10736
rect 11388 10696 11612 10724
rect 11388 10684 11394 10696
rect 11606 10684 11612 10696
rect 11664 10724 11670 10736
rect 11701 10727 11759 10733
rect 11701 10724 11713 10727
rect 11664 10696 11713 10724
rect 11664 10684 11670 10696
rect 11701 10693 11713 10696
rect 11747 10693 11759 10727
rect 11701 10687 11759 10693
rect 11974 10684 11980 10736
rect 12032 10684 12038 10736
rect 12066 10684 12072 10736
rect 12124 10684 12130 10736
rect 12437 10727 12495 10733
rect 12437 10693 12449 10727
rect 12483 10724 12495 10727
rect 12710 10724 12716 10736
rect 12483 10696 12716 10724
rect 12483 10693 12495 10696
rect 12437 10687 12495 10693
rect 12710 10684 12716 10696
rect 12768 10684 12774 10736
rect 12805 10727 12863 10733
rect 12805 10693 12817 10727
rect 12851 10724 12863 10727
rect 13170 10724 13176 10736
rect 12851 10696 13176 10724
rect 12851 10693 12863 10696
rect 12805 10687 12863 10693
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 13722 10684 13728 10736
rect 13780 10684 13786 10736
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10625 10103 10659
rect 10045 10619 10103 10625
rect 10319 10659 10377 10665
rect 10319 10625 10331 10659
rect 10365 10656 10377 10659
rect 13832 10656 13860 10764
rect 14182 10752 14188 10764
rect 14240 10792 14246 10804
rect 15013 10795 15071 10801
rect 14240 10764 14964 10792
rect 14240 10752 14246 10764
rect 13906 10684 13912 10736
rect 13964 10684 13970 10736
rect 14826 10684 14832 10736
rect 14884 10684 14890 10736
rect 14936 10724 14964 10764
rect 15013 10761 15025 10795
rect 15059 10792 15071 10795
rect 15286 10792 15292 10804
rect 15059 10764 15292 10792
rect 15059 10761 15071 10764
rect 15013 10755 15071 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16209 10795 16267 10801
rect 16209 10792 16221 10795
rect 15896 10764 16221 10792
rect 15896 10752 15902 10764
rect 16209 10761 16221 10764
rect 16255 10761 16267 10795
rect 16209 10755 16267 10761
rect 16666 10752 16672 10804
rect 16724 10792 16730 10804
rect 16942 10792 16948 10804
rect 16724 10764 16948 10792
rect 16724 10752 16730 10764
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 17034 10752 17040 10804
rect 17092 10792 17098 10804
rect 17092 10764 20024 10792
rect 17092 10752 17098 10764
rect 16960 10724 16988 10752
rect 17494 10724 17500 10736
rect 14936 10696 15498 10724
rect 16960 10696 17500 10724
rect 10365 10628 13860 10656
rect 13924 10656 13952 10684
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13924 10628 14013 10656
rect 10365 10625 10377 10628
rect 10319 10619 10377 10625
rect 14001 10625 14013 10628
rect 14047 10625 14059 10659
rect 14001 10619 14059 10625
rect 14090 10616 14096 10668
rect 14148 10616 14154 10668
rect 14458 10616 14464 10668
rect 14516 10616 14522 10668
rect 14642 10616 14648 10668
rect 14700 10656 14706 10668
rect 15470 10665 15498 10696
rect 17494 10684 17500 10696
rect 17552 10684 17558 10736
rect 18046 10684 18052 10736
rect 18104 10724 18110 10736
rect 19153 10727 19211 10733
rect 19153 10724 19165 10727
rect 18104 10696 19165 10724
rect 18104 10684 18110 10696
rect 19153 10693 19165 10696
rect 19199 10693 19211 10727
rect 19153 10687 19211 10693
rect 19245 10727 19303 10733
rect 19245 10693 19257 10727
rect 19291 10724 19303 10727
rect 19429 10727 19487 10733
rect 19429 10724 19441 10727
rect 19291 10696 19441 10724
rect 19291 10693 19303 10696
rect 19245 10687 19303 10693
rect 19429 10693 19441 10696
rect 19475 10693 19487 10727
rect 19429 10687 19487 10693
rect 19702 10684 19708 10736
rect 19760 10684 19766 10736
rect 19886 10695 19892 10736
rect 19871 10689 19892 10695
rect 15455 10659 15513 10665
rect 14700 10628 14854 10656
rect 14700 10616 14706 10628
rect 14826 10600 14854 10628
rect 15455 10625 15467 10659
rect 15501 10656 15513 10659
rect 15562 10656 15568 10668
rect 15501 10628 15568 10656
rect 15501 10625 15513 10628
rect 15455 10619 15513 10625
rect 15562 10616 15568 10628
rect 15620 10616 15626 10668
rect 18874 10616 18880 10668
rect 18932 10616 18938 10668
rect 19061 10659 19119 10665
rect 19061 10625 19073 10659
rect 19107 10656 19119 10659
rect 19334 10656 19340 10668
rect 19107 10628 19340 10656
rect 19107 10625 19119 10628
rect 19061 10619 19119 10625
rect 19334 10616 19340 10628
rect 19392 10616 19398 10668
rect 19518 10616 19524 10668
rect 19576 10616 19582 10668
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10656 19671 10659
rect 19720 10656 19748 10684
rect 19659 10628 19748 10656
rect 19871 10655 19883 10689
rect 19944 10684 19950 10736
rect 19996 10724 20024 10764
rect 20162 10752 20168 10804
rect 20220 10792 20226 10804
rect 20220 10764 23336 10792
rect 20220 10752 20226 10764
rect 19996 10696 23152 10724
rect 19917 10658 19932 10684
rect 19917 10655 19929 10658
rect 19871 10649 19929 10655
rect 19659 10625 19671 10628
rect 19613 10619 19671 10625
rect 22370 10616 22376 10668
rect 22428 10616 22434 10668
rect 22646 10616 22652 10668
rect 22704 10616 22710 10668
rect 8110 10588 8116 10600
rect 7438 10560 8116 10588
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 3418 10480 3424 10532
rect 3476 10520 3482 10532
rect 3476 10492 3924 10520
rect 3476 10480 3482 10492
rect 1578 10412 1584 10464
rect 1636 10412 1642 10464
rect 2866 10412 2872 10464
rect 2924 10452 2930 10464
rect 3789 10455 3847 10461
rect 3789 10452 3801 10455
rect 2924 10424 3801 10452
rect 2924 10412 2930 10424
rect 3789 10421 3801 10424
rect 3835 10421 3847 10455
rect 3896 10452 3924 10492
rect 5534 10480 5540 10532
rect 5592 10520 5598 10532
rect 7009 10523 7067 10529
rect 7009 10520 7021 10523
rect 5592 10492 7021 10520
rect 5592 10480 5598 10492
rect 7009 10489 7021 10492
rect 7055 10489 7067 10523
rect 7009 10483 7067 10489
rect 11057 10523 11115 10529
rect 11057 10489 11069 10523
rect 11103 10520 11115 10523
rect 11532 10520 11560 10574
rect 13630 10548 13636 10600
rect 13688 10548 13694 10600
rect 14826 10548 14832 10600
rect 14884 10588 14890 10600
rect 15197 10591 15255 10597
rect 15197 10588 15209 10591
rect 14884 10560 15209 10588
rect 14884 10548 14890 10560
rect 15197 10557 15209 10560
rect 15243 10557 15255 10591
rect 15197 10551 15255 10557
rect 22005 10591 22063 10597
rect 22005 10557 22017 10591
rect 22051 10588 22063 10591
rect 22094 10588 22100 10600
rect 22051 10560 22100 10588
rect 22051 10557 22063 10560
rect 22005 10551 22063 10557
rect 22094 10548 22100 10560
rect 22152 10548 22158 10600
rect 22649 10523 22707 10529
rect 22649 10520 22661 10523
rect 11103 10492 11560 10520
rect 20272 10492 22661 10520
rect 11103 10489 11115 10492
rect 11057 10483 11115 10489
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 3896 10424 8217 10452
rect 3789 10415 3847 10421
rect 8205 10421 8217 10424
rect 8251 10421 8263 10455
rect 8205 10415 8263 10421
rect 15286 10412 15292 10464
rect 15344 10452 15350 10464
rect 20272 10452 20300 10492
rect 22649 10489 22661 10492
rect 22695 10489 22707 10523
rect 23124 10520 23152 10696
rect 23198 10616 23204 10668
rect 23256 10616 23262 10668
rect 23308 10588 23336 10764
rect 23474 10684 23480 10736
rect 23532 10724 23538 10736
rect 23569 10727 23627 10733
rect 23569 10724 23581 10727
rect 23532 10696 23581 10724
rect 23532 10684 23538 10696
rect 23569 10693 23581 10696
rect 23615 10693 23627 10727
rect 23569 10687 23627 10693
rect 23658 10684 23664 10736
rect 23716 10724 23722 10736
rect 24121 10727 24179 10733
rect 24121 10724 24133 10727
rect 23716 10696 24133 10724
rect 23716 10684 23722 10696
rect 24121 10693 24133 10696
rect 24167 10693 24179 10727
rect 24121 10687 24179 10693
rect 24486 10616 24492 10668
rect 24544 10616 24550 10668
rect 25590 10588 25596 10600
rect 23308 10560 25596 10588
rect 25590 10548 25596 10560
rect 25648 10548 25654 10600
rect 25406 10520 25412 10532
rect 23124 10492 25412 10520
rect 22649 10483 22707 10489
rect 25406 10480 25412 10492
rect 25464 10480 25470 10532
rect 15344 10424 20300 10452
rect 20625 10455 20683 10461
rect 15344 10412 15350 10424
rect 20625 10421 20637 10455
rect 20671 10452 20683 10455
rect 20898 10452 20904 10464
rect 20671 10424 20904 10452
rect 20671 10421 20683 10424
rect 20625 10415 20683 10421
rect 20898 10412 20904 10424
rect 20956 10412 20962 10464
rect 22830 10412 22836 10464
rect 22888 10452 22894 10464
rect 23017 10455 23075 10461
rect 23017 10452 23029 10455
rect 22888 10424 23029 10452
rect 22888 10412 22894 10424
rect 23017 10421 23029 10424
rect 23063 10421 23075 10455
rect 23017 10415 23075 10421
rect 23842 10412 23848 10464
rect 23900 10412 23906 10464
rect 1104 10362 24840 10384
rect 1104 10310 3917 10362
rect 3969 10310 3981 10362
rect 4033 10310 4045 10362
rect 4097 10310 4109 10362
rect 4161 10310 4173 10362
rect 4225 10310 9851 10362
rect 9903 10310 9915 10362
rect 9967 10310 9979 10362
rect 10031 10310 10043 10362
rect 10095 10310 10107 10362
rect 10159 10310 15785 10362
rect 15837 10310 15849 10362
rect 15901 10310 15913 10362
rect 15965 10310 15977 10362
rect 16029 10310 16041 10362
rect 16093 10310 21719 10362
rect 21771 10310 21783 10362
rect 21835 10310 21847 10362
rect 21899 10310 21911 10362
rect 21963 10310 21975 10362
rect 22027 10310 24840 10362
rect 1104 10288 24840 10310
rect 3234 10208 3240 10260
rect 3292 10208 3298 10260
rect 3344 10220 5212 10248
rect 1670 10140 1676 10192
rect 1728 10140 1734 10192
rect 2317 10115 2375 10121
rect 2317 10081 2329 10115
rect 2363 10112 2375 10115
rect 2774 10112 2780 10124
rect 2363 10084 2780 10112
rect 2363 10081 2375 10084
rect 2317 10075 2375 10081
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 3344 10112 3372 10220
rect 5184 10180 5212 10220
rect 5534 10208 5540 10260
rect 5592 10208 5598 10260
rect 5902 10208 5908 10260
rect 5960 10208 5966 10260
rect 6822 10208 6828 10260
rect 6880 10208 6886 10260
rect 6914 10208 6920 10260
rect 6972 10208 6978 10260
rect 10781 10251 10839 10257
rect 10781 10248 10793 10251
rect 7024 10220 10793 10248
rect 5920 10180 5948 10208
rect 5184 10152 5948 10180
rect 6840 10180 6868 10208
rect 7024 10180 7052 10220
rect 10781 10217 10793 10220
rect 10827 10217 10839 10251
rect 12250 10248 12256 10260
rect 10781 10211 10839 10217
rect 10980 10220 12256 10248
rect 6840 10152 7052 10180
rect 7484 10152 9720 10180
rect 3068 10084 3372 10112
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 1489 10047 1547 10053
rect 1489 10013 1501 10047
rect 1535 10044 1547 10047
rect 3068 10044 3096 10084
rect 4338 10072 4344 10124
rect 4396 10112 4402 10124
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 4396 10084 4537 10112
rect 4396 10072 4402 10084
rect 4525 10081 4537 10084
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 1535 10016 3096 10044
rect 3145 10047 3203 10053
rect 1535 10013 1547 10016
rect 1489 10007 1547 10013
rect 3145 10013 3157 10047
rect 3191 10013 3203 10047
rect 3145 10007 3203 10013
rect 1412 9976 1440 10004
rect 2041 9979 2099 9985
rect 2041 9976 2053 9979
rect 1412 9948 2053 9976
rect 2041 9945 2053 9948
rect 2087 9945 2099 9979
rect 2041 9939 2099 9945
rect 2593 9979 2651 9985
rect 2593 9945 2605 9979
rect 2639 9976 2651 9979
rect 2682 9976 2688 9988
rect 2639 9948 2688 9976
rect 2639 9945 2651 9948
rect 2593 9939 2651 9945
rect 2682 9936 2688 9948
rect 2740 9936 2746 9988
rect 2958 9936 2964 9988
rect 3016 9976 3022 9988
rect 3160 9976 3188 10007
rect 3016 9948 3188 9976
rect 3016 9936 3022 9948
rect 3878 9936 3884 9988
rect 3936 9936 3942 9988
rect 4540 9976 4568 10075
rect 4798 10044 4804 10056
rect 4759 10016 4804 10044
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 6163 10017 6221 10023
rect 5810 9976 5816 9988
rect 4540 9948 5816 9976
rect 5810 9936 5816 9948
rect 5868 9976 5874 9988
rect 5920 9976 5948 10007
rect 6163 9983 6175 10017
rect 6209 10014 6221 10017
rect 6209 9983 6224 10014
rect 6163 9977 6224 9983
rect 5868 9948 5948 9976
rect 6196 9976 6224 9977
rect 6270 9976 6276 9988
rect 6196 9948 6276 9976
rect 5868 9936 5874 9948
rect 6270 9936 6276 9948
rect 6328 9936 6334 9988
rect 2866 9868 2872 9920
rect 2924 9868 2930 9920
rect 3326 9868 3332 9920
rect 3384 9908 3390 9920
rect 3973 9911 4031 9917
rect 3973 9908 3985 9911
rect 3384 9880 3985 9908
rect 3384 9868 3390 9880
rect 3973 9877 3985 9880
rect 4019 9877 4031 9911
rect 3973 9871 4031 9877
rect 5442 9868 5448 9920
rect 5500 9908 5506 9920
rect 7484 9908 7512 10152
rect 9122 10112 9128 10124
rect 8312 10084 9128 10112
rect 8312 10056 8340 10084
rect 9122 10072 9128 10084
rect 9180 10072 9186 10124
rect 9582 10072 9588 10124
rect 9640 10072 9646 10124
rect 9692 10112 9720 10152
rect 9858 10112 9864 10124
rect 9692 10084 9864 10112
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 9999 10115 10057 10121
rect 9999 10081 10011 10115
rect 10045 10112 10057 10115
rect 10980 10112 11008 10220
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 12492 10220 12572 10248
rect 12492 10208 12498 10220
rect 10045 10084 11008 10112
rect 10045 10081 10057 10084
rect 9999 10075 10057 10081
rect 8294 10004 8300 10056
rect 8352 10004 8358 10056
rect 8754 10004 8760 10056
rect 8812 10044 8818 10056
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8812 10016 8953 10044
rect 8812 10004 8818 10016
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 10134 10004 10140 10056
rect 10192 10004 10198 10056
rect 10870 10004 10876 10056
rect 10928 10044 10934 10056
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10928 10016 10977 10044
rect 10928 10004 10934 10016
rect 10965 10013 10977 10016
rect 11011 10013 11023 10047
rect 11239 10047 11297 10053
rect 11239 10044 11251 10047
rect 10965 10007 11023 10013
rect 11070 10016 11251 10044
rect 5500 9880 7512 9908
rect 5500 9868 5506 9880
rect 10410 9868 10416 9920
rect 10468 9908 10474 9920
rect 11070 9908 11098 10016
rect 11239 10013 11251 10016
rect 11285 10044 11297 10047
rect 12342 10044 12348 10056
rect 11285 10016 12348 10044
rect 11285 10013 11297 10016
rect 11239 10007 11297 10013
rect 12342 10004 12348 10016
rect 12400 10004 12406 10056
rect 12544 10044 12572 10220
rect 12694 10220 13308 10248
rect 12694 10180 12722 10220
rect 12636 10152 12722 10180
rect 13280 10180 13308 10220
rect 13630 10208 13636 10260
rect 13688 10208 13694 10260
rect 14090 10208 14096 10260
rect 14148 10248 14154 10260
rect 15105 10251 15163 10257
rect 15105 10248 15117 10251
rect 14148 10220 15117 10248
rect 14148 10208 14154 10220
rect 15105 10217 15117 10220
rect 15151 10217 15163 10251
rect 15105 10211 15163 10217
rect 18785 10251 18843 10257
rect 18785 10217 18797 10251
rect 18831 10248 18843 10251
rect 18874 10248 18880 10260
rect 18831 10220 18880 10248
rect 18831 10217 18843 10220
rect 18785 10211 18843 10217
rect 18874 10208 18880 10220
rect 18932 10208 18938 10260
rect 19518 10208 19524 10260
rect 19576 10208 19582 10260
rect 22370 10208 22376 10260
rect 22428 10208 22434 10260
rect 22646 10208 22652 10260
rect 22704 10208 22710 10260
rect 22830 10208 22836 10260
rect 22888 10208 22894 10260
rect 19245 10183 19303 10189
rect 13280 10152 14044 10180
rect 12636 10121 12664 10152
rect 14016 10124 14044 10152
rect 19245 10149 19257 10183
rect 19291 10149 19303 10183
rect 19245 10143 19303 10149
rect 21913 10183 21971 10189
rect 21913 10149 21925 10183
rect 21959 10180 21971 10183
rect 22094 10180 22100 10192
rect 21959 10152 22100 10180
rect 21959 10149 21971 10152
rect 21913 10143 21971 10149
rect 12621 10115 12679 10121
rect 12621 10081 12633 10115
rect 12667 10081 12679 10115
rect 12621 10075 12679 10081
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 14056 10084 14105 10112
rect 14056 10072 14062 10084
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 14366 10053 14372 10056
rect 12863 10047 12921 10053
rect 12863 10044 12875 10047
rect 12544 10016 12875 10044
rect 12863 10013 12875 10016
rect 12909 10013 12921 10047
rect 12863 10007 12921 10013
rect 14351 10047 14372 10053
rect 14351 10013 14363 10047
rect 14351 10007 14372 10013
rect 14366 10004 14372 10007
rect 14424 10004 14430 10056
rect 16850 10004 16856 10056
rect 16908 10044 16914 10056
rect 17402 10044 17408 10056
rect 16908 10016 17408 10044
rect 16908 10004 16914 10016
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10044 18751 10047
rect 19260 10044 19288 10143
rect 22094 10140 22100 10152
rect 22152 10180 22158 10192
rect 22152 10152 22600 10180
rect 22152 10140 22158 10152
rect 18739 10016 19288 10044
rect 19429 10047 19487 10053
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 19429 10013 19441 10047
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 11330 9936 11336 9988
rect 11388 9976 11394 9988
rect 14366 9976 14394 10004
rect 17678 9976 17684 9988
rect 11388 9948 14394 9976
rect 17236 9948 17684 9976
rect 11388 9936 11394 9948
rect 10468 9880 11098 9908
rect 10468 9868 10474 9880
rect 11882 9868 11888 9920
rect 11940 9908 11946 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 11940 9880 11989 9908
rect 11940 9868 11946 9880
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 11977 9871 12035 9877
rect 12066 9868 12072 9920
rect 12124 9908 12130 9920
rect 17236 9908 17264 9948
rect 17678 9936 17684 9948
rect 17736 9936 17742 9988
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 19444 9976 19472 10007
rect 19702 10004 19708 10056
rect 19760 10004 19766 10056
rect 21174 10053 21180 10056
rect 20901 10047 20959 10053
rect 20901 10013 20913 10047
rect 20947 10044 20959 10047
rect 21143 10047 21180 10053
rect 20947 10016 21036 10044
rect 20947 10013 20959 10016
rect 20901 10007 20959 10013
rect 21008 9988 21036 10016
rect 21143 10013 21155 10047
rect 21143 10007 21180 10013
rect 21174 10004 21180 10007
rect 21232 10004 21238 10056
rect 21726 10004 21732 10056
rect 21784 10044 21790 10056
rect 22572 10053 22600 10152
rect 22848 10112 22876 10208
rect 22756 10084 22876 10112
rect 22756 10053 22784 10084
rect 22281 10047 22339 10053
rect 22281 10044 22293 10047
rect 21784 10016 22293 10044
rect 21784 10004 21790 10016
rect 22281 10013 22293 10016
rect 22327 10013 22339 10047
rect 22281 10007 22339 10013
rect 22557 10047 22615 10053
rect 22557 10013 22569 10047
rect 22603 10013 22615 10047
rect 22557 10007 22615 10013
rect 22741 10047 22799 10053
rect 22741 10013 22753 10047
rect 22787 10013 22799 10047
rect 22741 10007 22799 10013
rect 22833 10047 22891 10053
rect 22833 10013 22845 10047
rect 22879 10044 22891 10047
rect 22879 10016 22968 10044
rect 22879 10013 22891 10016
rect 22833 10007 22891 10013
rect 22940 9988 22968 10016
rect 23091 10017 23149 10023
rect 19978 9976 19984 9988
rect 19392 9948 19984 9976
rect 19392 9936 19398 9948
rect 19978 9936 19984 9948
rect 20036 9936 20042 9988
rect 20990 9936 20996 9988
rect 21048 9976 21054 9988
rect 21542 9976 21548 9988
rect 21048 9948 21548 9976
rect 21048 9936 21054 9948
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 22922 9936 22928 9988
rect 22980 9936 22986 9988
rect 23091 9983 23103 10017
rect 23137 10014 23149 10017
rect 23137 9983 23152 10014
rect 23091 9977 23152 9983
rect 12124 9880 17264 9908
rect 12124 9868 12130 9880
rect 17310 9868 17316 9920
rect 17368 9908 17374 9920
rect 23124 9908 23152 9977
rect 17368 9880 23152 9908
rect 23845 9911 23903 9917
rect 17368 9868 17374 9880
rect 23845 9877 23857 9911
rect 23891 9908 23903 9911
rect 24118 9908 24124 9920
rect 23891 9880 24124 9908
rect 23891 9877 23903 9880
rect 23845 9871 23903 9877
rect 24118 9868 24124 9880
rect 24176 9868 24182 9920
rect 1104 9818 25000 9840
rect 1104 9766 6884 9818
rect 6936 9766 6948 9818
rect 7000 9766 7012 9818
rect 7064 9766 7076 9818
rect 7128 9766 7140 9818
rect 7192 9766 12818 9818
rect 12870 9766 12882 9818
rect 12934 9766 12946 9818
rect 12998 9766 13010 9818
rect 13062 9766 13074 9818
rect 13126 9766 18752 9818
rect 18804 9766 18816 9818
rect 18868 9766 18880 9818
rect 18932 9766 18944 9818
rect 18996 9766 19008 9818
rect 19060 9766 24686 9818
rect 24738 9766 24750 9818
rect 24802 9766 24814 9818
rect 24866 9766 24878 9818
rect 24930 9766 24942 9818
rect 24994 9766 25000 9818
rect 1104 9744 25000 9766
rect 1762 9664 1768 9716
rect 1820 9664 1826 9716
rect 2314 9664 2320 9716
rect 2372 9664 2378 9716
rect 3237 9707 3295 9713
rect 3237 9673 3249 9707
rect 3283 9704 3295 9707
rect 3878 9704 3884 9716
rect 3283 9676 3884 9704
rect 3283 9673 3295 9676
rect 3237 9667 3295 9673
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 6546 9704 6552 9716
rect 5776 9676 6552 9704
rect 5776 9664 5782 9676
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 8297 9707 8355 9713
rect 7116 9676 7586 9704
rect 2777 9639 2835 9645
rect 2777 9605 2789 9639
rect 2823 9636 2835 9639
rect 2823 9608 3096 9636
rect 2823 9605 2835 9608
rect 2777 9599 2835 9605
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 1688 9500 1716 9531
rect 2222 9528 2228 9580
rect 2280 9528 2286 9580
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 2958 9568 2964 9580
rect 2648 9540 2964 9568
rect 2648 9528 2654 9540
rect 2958 9528 2964 9540
rect 3016 9528 3022 9580
rect 3068 9568 3096 9608
rect 3142 9596 3148 9648
rect 3200 9596 3206 9648
rect 3344 9608 4660 9636
rect 3344 9568 3372 9608
rect 3068 9540 3372 9568
rect 3418 9528 3424 9580
rect 3476 9528 3482 9580
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 3787 9571 3845 9577
rect 3787 9537 3799 9571
rect 3833 9568 3845 9571
rect 4338 9568 4344 9580
rect 3833 9540 4344 9568
rect 3833 9537 3845 9540
rect 3787 9531 3845 9537
rect 3528 9500 3556 9531
rect 4338 9528 4344 9540
rect 4396 9568 4402 9580
rect 4522 9568 4528 9580
rect 4396 9540 4528 9568
rect 4396 9528 4402 9540
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 1688 9472 2774 9500
rect 2746 9364 2774 9472
rect 3436 9472 3556 9500
rect 4632 9500 4660 9608
rect 6086 9596 6092 9648
rect 6144 9596 6150 9648
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9568 5135 9571
rect 5166 9568 5172 9580
rect 5123 9540 5172 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 5350 9528 5356 9580
rect 5408 9528 5414 9580
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 5644 9500 5672 9531
rect 5902 9528 5908 9580
rect 5960 9528 5966 9580
rect 6104 9568 6132 9596
rect 7116 9568 7144 9676
rect 7558 9607 7586 9676
rect 8297 9673 8309 9707
rect 8343 9704 8355 9707
rect 9582 9704 9588 9716
rect 8343 9676 9588 9704
rect 8343 9673 8355 9676
rect 8297 9667 8355 9673
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 9677 9707 9735 9713
rect 9677 9673 9689 9707
rect 9723 9704 9735 9707
rect 10134 9704 10140 9716
rect 9723 9676 10140 9704
rect 9723 9673 9735 9676
rect 9677 9667 9735 9673
rect 10134 9664 10140 9676
rect 10192 9664 10198 9716
rect 12989 9707 13047 9713
rect 12989 9704 13001 9707
rect 10980 9676 13001 9704
rect 6104 9540 7144 9568
rect 7543 9601 7601 9607
rect 7543 9567 7555 9601
rect 7589 9567 7601 9601
rect 9030 9596 9036 9648
rect 9088 9636 9094 9648
rect 10980 9636 11008 9676
rect 12989 9673 13001 9676
rect 13035 9673 13047 9707
rect 19429 9707 19487 9713
rect 12989 9667 13047 9673
rect 16592 9676 17080 9704
rect 9088 9608 11008 9636
rect 9088 9596 9094 9608
rect 11054 9596 11060 9648
rect 11112 9636 11118 9648
rect 11606 9636 11612 9648
rect 11112 9608 11612 9636
rect 11112 9596 11118 9608
rect 11606 9596 11612 9608
rect 11664 9636 11670 9648
rect 11701 9639 11759 9645
rect 11701 9636 11713 9639
rect 11664 9608 11713 9636
rect 11664 9596 11670 9608
rect 11701 9605 11713 9608
rect 11747 9605 11759 9639
rect 11701 9599 11759 9605
rect 11974 9596 11980 9648
rect 12032 9596 12038 9648
rect 12360 9608 12756 9636
rect 12360 9580 12388 9608
rect 7543 9561 7601 9567
rect 8939 9571 8997 9577
rect 8939 9537 8951 9571
rect 8985 9568 8997 9571
rect 8985 9540 10916 9568
rect 8985 9537 8997 9540
rect 8939 9531 8997 9537
rect 7190 9500 7196 9512
rect 4632 9472 5488 9500
rect 5644 9472 7196 9500
rect 3436 9444 3464 9472
rect 3418 9392 3424 9444
rect 3476 9392 3482 9444
rect 5460 9441 5488 9472
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 4893 9435 4951 9441
rect 4893 9432 4905 9435
rect 4172 9404 4905 9432
rect 4172 9364 4200 9404
rect 4893 9401 4905 9404
rect 4939 9401 4951 9435
rect 4893 9395 4951 9401
rect 5445 9435 5503 9441
rect 5445 9401 5457 9435
rect 5491 9401 5503 9435
rect 5445 9395 5503 9401
rect 5810 9392 5816 9444
rect 5868 9432 5874 9444
rect 6730 9432 6736 9444
rect 5868 9404 6736 9432
rect 5868 9392 5874 9404
rect 6730 9392 6736 9404
rect 6788 9432 6794 9444
rect 7300 9432 7328 9463
rect 6788 9404 7420 9432
rect 6788 9392 6794 9404
rect 2746 9336 4200 9364
rect 4522 9324 4528 9376
rect 4580 9324 4586 9376
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 5169 9367 5227 9373
rect 5169 9364 5181 9367
rect 4672 9336 5181 9364
rect 4672 9324 4678 9336
rect 5169 9333 5181 9336
rect 5215 9333 5227 9367
rect 5169 9327 5227 9333
rect 5718 9324 5724 9376
rect 5776 9324 5782 9376
rect 7392 9364 7420 9404
rect 8680 9364 8708 9463
rect 7392 9336 8708 9364
rect 8938 9324 8944 9376
rect 8996 9364 9002 9376
rect 9600 9364 9628 9540
rect 10888 9500 10916 9540
rect 10962 9528 10968 9580
rect 11020 9568 11026 9580
rect 11790 9568 11796 9580
rect 11020 9540 11796 9568
rect 11020 9528 11026 9540
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9568 12127 9571
rect 12250 9568 12256 9580
rect 12115 9540 12256 9568
rect 12115 9537 12127 9540
rect 12069 9531 12127 9537
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 12342 9528 12348 9580
rect 12400 9528 12406 9580
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9568 12495 9571
rect 12526 9568 12532 9580
rect 12483 9540 12532 9568
rect 12483 9537 12495 9540
rect 12437 9531 12495 9537
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12728 9568 12756 9608
rect 12802 9596 12808 9648
rect 12860 9596 12866 9648
rect 16592 9568 16620 9676
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 17052 9636 17080 9676
rect 17880 9676 19380 9704
rect 17218 9636 17224 9648
rect 16724 9608 16804 9636
rect 17052 9608 17224 9636
rect 16724 9596 16730 9608
rect 16776 9568 16804 9608
rect 17218 9596 17224 9608
rect 17276 9636 17282 9648
rect 17880 9636 17908 9676
rect 17276 9608 17908 9636
rect 18316 9639 18374 9645
rect 17276 9596 17282 9608
rect 18316 9605 18328 9639
rect 18362 9636 18374 9639
rect 19242 9636 19248 9648
rect 18362 9608 19248 9636
rect 18362 9605 18374 9608
rect 18316 9599 18374 9605
rect 19242 9596 19248 9608
rect 19300 9596 19306 9648
rect 19352 9636 19380 9676
rect 19429 9673 19441 9707
rect 19475 9704 19487 9707
rect 19702 9704 19708 9716
rect 19475 9676 19708 9704
rect 19475 9673 19487 9676
rect 19429 9667 19487 9673
rect 19702 9664 19708 9676
rect 19760 9664 19766 9716
rect 21266 9704 21272 9716
rect 19812 9676 21272 9704
rect 19812 9636 19840 9676
rect 21266 9664 21272 9676
rect 21324 9664 21330 9716
rect 21453 9707 21511 9713
rect 21453 9673 21465 9707
rect 21499 9704 21511 9707
rect 21726 9704 21732 9716
rect 21499 9676 21732 9704
rect 21499 9673 21511 9676
rect 21453 9667 21511 9673
rect 21726 9664 21732 9676
rect 21784 9664 21790 9716
rect 22370 9664 22376 9716
rect 22428 9704 22434 9716
rect 23106 9704 23112 9716
rect 22428 9676 23112 9704
rect 22428 9664 22434 9676
rect 23106 9664 23112 9676
rect 23164 9664 23170 9716
rect 23198 9664 23204 9716
rect 23256 9664 23262 9716
rect 24210 9664 24216 9716
rect 24268 9704 24274 9716
rect 24946 9704 24952 9716
rect 24268 9676 24952 9704
rect 24268 9664 24274 9676
rect 24946 9664 24952 9676
rect 25004 9664 25010 9716
rect 19352 9608 19840 9636
rect 23750 9596 23756 9648
rect 23808 9636 23814 9648
rect 24121 9639 24179 9645
rect 24121 9636 24133 9639
rect 23808 9608 24133 9636
rect 23808 9596 23814 9608
rect 24121 9605 24133 9608
rect 24167 9605 24179 9639
rect 24121 9599 24179 9605
rect 24489 9639 24547 9645
rect 24489 9605 24501 9639
rect 24535 9636 24547 9639
rect 25038 9636 25044 9648
rect 24535 9608 25044 9636
rect 24535 9605 24547 9608
rect 24489 9599 24547 9605
rect 25038 9596 25044 9608
rect 25096 9596 25102 9648
rect 16943 9571 17001 9577
rect 16943 9568 16955 9571
rect 12728 9540 12940 9568
rect 16592 9540 16712 9568
rect 16776 9540 16955 9568
rect 11330 9500 11336 9512
rect 10888 9472 11336 9500
rect 11330 9460 11336 9472
rect 11388 9460 11394 9512
rect 11882 9460 11888 9512
rect 11940 9460 11946 9512
rect 8996 9336 9628 9364
rect 12912 9364 12940 9540
rect 16684 9512 16712 9540
rect 16943 9537 16955 9540
rect 16989 9568 17001 9571
rect 17034 9568 17040 9580
rect 16989 9540 17040 9568
rect 16989 9537 17001 9540
rect 16943 9531 17001 9537
rect 17034 9528 17040 9540
rect 17092 9568 17098 9580
rect 19763 9571 19821 9577
rect 19763 9568 19775 9571
rect 17092 9540 19775 9568
rect 17092 9528 17098 9540
rect 19763 9537 19775 9540
rect 19809 9537 19821 9571
rect 19763 9531 19821 9537
rect 21637 9571 21695 9577
rect 21637 9537 21649 9571
rect 21683 9568 21695 9571
rect 22088 9571 22146 9577
rect 22088 9568 22100 9571
rect 21683 9540 22100 9568
rect 21683 9537 21695 9540
rect 21637 9531 21695 9537
rect 22088 9537 22100 9540
rect 22134 9568 22146 9571
rect 22134 9540 22876 9568
rect 22134 9537 22146 9540
rect 22088 9531 22146 9537
rect 16666 9460 16672 9512
rect 16724 9460 16730 9512
rect 18046 9460 18052 9512
rect 18104 9460 18110 9512
rect 19521 9503 19579 9509
rect 19521 9469 19533 9503
rect 19567 9469 19579 9503
rect 19521 9463 19579 9469
rect 19426 9392 19432 9444
rect 19484 9432 19490 9444
rect 19536 9432 19564 9463
rect 20806 9460 20812 9512
rect 20864 9500 20870 9512
rect 21542 9500 21548 9512
rect 20864 9472 21548 9500
rect 20864 9460 20870 9472
rect 21542 9460 21548 9472
rect 21600 9500 21606 9512
rect 21821 9503 21879 9509
rect 21821 9500 21833 9503
rect 21600 9472 21833 9500
rect 21600 9460 21606 9472
rect 21821 9469 21833 9472
rect 21867 9469 21879 9503
rect 22848 9500 22876 9540
rect 23566 9528 23572 9580
rect 23624 9528 23630 9580
rect 23934 9528 23940 9580
rect 23992 9528 23998 9580
rect 24210 9528 24216 9580
rect 24268 9528 24274 9580
rect 24228 9500 24256 9528
rect 22848 9472 24256 9500
rect 21821 9463 21879 9469
rect 20990 9432 20996 9444
rect 19484 9404 19564 9432
rect 19484 9392 19490 9404
rect 17126 9364 17132 9376
rect 12912 9336 17132 9364
rect 8996 9324 9002 9336
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 17678 9324 17684 9376
rect 17736 9324 17742 9376
rect 19536 9364 19564 9404
rect 20180 9404 20996 9432
rect 20180 9364 20208 9404
rect 20990 9392 20996 9404
rect 21048 9392 21054 9444
rect 19536 9336 20208 9364
rect 20438 9324 20444 9376
rect 20496 9364 20502 9376
rect 20533 9367 20591 9373
rect 20533 9364 20545 9367
rect 20496 9336 20545 9364
rect 20496 9324 20502 9336
rect 20533 9333 20545 9336
rect 20579 9333 20591 9367
rect 20533 9327 20591 9333
rect 21358 9324 21364 9376
rect 21416 9364 21422 9376
rect 23106 9364 23112 9376
rect 21416 9336 23112 9364
rect 21416 9324 21422 9336
rect 23106 9324 23112 9336
rect 23164 9324 23170 9376
rect 1104 9274 24840 9296
rect 1104 9222 3917 9274
rect 3969 9222 3981 9274
rect 4033 9222 4045 9274
rect 4097 9222 4109 9274
rect 4161 9222 4173 9274
rect 4225 9222 9851 9274
rect 9903 9222 9915 9274
rect 9967 9222 9979 9274
rect 10031 9222 10043 9274
rect 10095 9222 10107 9274
rect 10159 9222 15785 9274
rect 15837 9222 15849 9274
rect 15901 9222 15913 9274
rect 15965 9222 15977 9274
rect 16029 9222 16041 9274
rect 16093 9222 21719 9274
rect 21771 9222 21783 9274
rect 21835 9222 21847 9274
rect 21899 9222 21911 9274
rect 21963 9222 21975 9274
rect 22027 9222 24840 9274
rect 1104 9200 24840 9222
rect 1302 9120 1308 9172
rect 1360 9120 1366 9172
rect 1489 9163 1547 9169
rect 1489 9129 1501 9163
rect 1535 9160 1547 9163
rect 2222 9160 2228 9172
rect 1535 9132 2228 9160
rect 1535 9129 1547 9132
rect 1489 9123 1547 9129
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 4338 9160 4344 9172
rect 3016 9132 4344 9160
rect 3016 9120 3022 9132
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 4522 9160 4528 9172
rect 4448 9132 4528 9160
rect 1320 9024 1348 9120
rect 2590 9092 2596 9104
rect 2516 9064 2596 9092
rect 1765 9027 1823 9033
rect 1765 9024 1777 9027
rect 1320 8996 1777 9024
rect 1765 8993 1777 8996
rect 1811 8993 1823 9027
rect 1765 8987 1823 8993
rect 1670 8916 1676 8968
rect 1728 8916 1734 8968
rect 2039 8959 2097 8965
rect 2039 8925 2051 8959
rect 2085 8956 2097 8959
rect 2516 8956 2544 9064
rect 2590 9052 2596 9064
rect 2648 9052 2654 9104
rect 3418 9052 3424 9104
rect 3476 9092 3482 9104
rect 4154 9092 4160 9104
rect 3476 9064 4160 9092
rect 3476 9052 3482 9064
rect 4154 9052 4160 9064
rect 4212 9052 4218 9104
rect 4448 9101 4476 9132
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 4764 9132 5641 9160
rect 4764 9120 4770 9132
rect 5629 9129 5641 9132
rect 5675 9129 5687 9163
rect 5629 9123 5687 9129
rect 7190 9120 7196 9172
rect 7248 9160 7254 9172
rect 12158 9160 12164 9172
rect 7248 9132 12164 9160
rect 7248 9120 7254 9132
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 12250 9120 12256 9172
rect 12308 9160 12314 9172
rect 12897 9163 12955 9169
rect 12897 9160 12909 9163
rect 12308 9132 12909 9160
rect 12308 9120 12314 9132
rect 12897 9129 12909 9132
rect 12943 9129 12955 9163
rect 12897 9123 12955 9129
rect 17126 9120 17132 9172
rect 17184 9160 17190 9172
rect 17184 9132 22094 9160
rect 17184 9120 17190 9132
rect 4433 9095 4491 9101
rect 4433 9061 4445 9095
rect 4479 9061 4491 9095
rect 4433 9055 4491 9061
rect 7356 9052 7362 9104
rect 7414 9101 7420 9104
rect 7414 9095 7435 9101
rect 7423 9061 7435 9095
rect 7414 9055 7435 9061
rect 7414 9052 7420 9055
rect 8386 9052 8392 9104
rect 8444 9092 8450 9104
rect 8444 9064 9674 9092
rect 8444 9052 8450 9064
rect 4522 9024 4528 9036
rect 3252 8996 4528 9024
rect 2085 8928 2544 8956
rect 2085 8925 2097 8928
rect 2039 8919 2097 8925
rect 2590 8916 2596 8968
rect 2648 8956 2654 8968
rect 3252 8965 3280 8996
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 4890 9033 4896 9036
rect 4847 9027 4896 9033
rect 4847 8993 4859 9027
rect 4893 8993 4896 9027
rect 4847 8987 4896 8993
rect 4890 8984 4896 8987
rect 4948 8984 4954 9036
rect 6914 8984 6920 9036
rect 6972 8984 6978 9036
rect 7650 9024 7656 9036
rect 7024 8996 7656 9024
rect 3237 8959 3295 8965
rect 2648 8928 3188 8956
rect 2648 8916 2654 8928
rect 1302 8848 1308 8900
rect 1360 8888 1366 8900
rect 3160 8888 3188 8928
rect 3237 8925 3249 8959
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3660 8928 3801 8956
rect 3660 8916 3666 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 3970 8916 3976 8968
rect 4028 8916 4034 8968
rect 4706 8916 4712 8968
rect 4764 8916 4770 8968
rect 4982 8916 4988 8968
rect 5040 8916 5046 8968
rect 6733 8959 6791 8965
rect 6733 8956 6745 8959
rect 5552 8928 6745 8956
rect 3620 8888 3648 8916
rect 5552 8900 5580 8928
rect 6733 8925 6745 8928
rect 6779 8925 6791 8959
rect 7024 8956 7052 8996
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 7791 9027 7849 9033
rect 7791 8993 7803 9027
rect 7837 9024 7849 9027
rect 8110 9024 8116 9036
rect 7837 8996 8116 9024
rect 7837 8993 7849 8996
rect 7791 8987 7849 8993
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 9309 9027 9367 9033
rect 9309 9024 9321 9027
rect 8536 8996 9321 9024
rect 8536 8984 8542 8996
rect 9309 8993 9321 8996
rect 9355 8993 9367 9027
rect 9646 9024 9674 9064
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 9953 9095 10011 9101
rect 9953 9092 9965 9095
rect 9824 9064 9965 9092
rect 9824 9052 9830 9064
rect 9953 9061 9965 9064
rect 9999 9061 10011 9095
rect 9953 9055 10011 9061
rect 16482 9052 16488 9104
rect 16540 9052 16546 9104
rect 18138 9052 18144 9104
rect 18196 9092 18202 9104
rect 20993 9095 21051 9101
rect 20993 9092 21005 9095
rect 18196 9064 21005 9092
rect 18196 9052 18202 9064
rect 20993 9061 21005 9064
rect 21039 9061 21051 9095
rect 22066 9092 22094 9132
rect 23937 9095 23995 9101
rect 23937 9092 23949 9095
rect 22066 9064 23949 9092
rect 20993 9055 21051 9061
rect 23937 9061 23949 9064
rect 23983 9061 23995 9095
rect 23937 9055 23995 9061
rect 10229 9027 10287 9033
rect 10229 9024 10241 9027
rect 9646 8996 10241 9024
rect 9309 8987 9367 8993
rect 10229 8993 10241 8996
rect 10275 8993 10287 9027
rect 16500 9024 16528 9052
rect 16669 9027 16727 9033
rect 16669 9024 16681 9027
rect 16500 8996 16681 9024
rect 10229 8987 10287 8993
rect 16669 8993 16681 8996
rect 16715 8993 16727 9027
rect 16669 8987 16727 8993
rect 17126 8984 17132 9036
rect 17184 8984 17190 9036
rect 18322 8984 18328 9036
rect 18380 8984 18386 9036
rect 19981 9027 20039 9033
rect 19981 8993 19993 9027
rect 20027 9024 20039 9027
rect 21453 9027 21511 9033
rect 21453 9024 21465 9027
rect 20027 8996 20576 9024
rect 20027 8993 20039 8996
rect 19981 8987 20039 8993
rect 6733 8919 6791 8925
rect 6840 8928 7052 8956
rect 1360 8860 3096 8888
rect 3160 8860 3648 8888
rect 1360 8848 1366 8860
rect 2774 8780 2780 8832
rect 2832 8780 2838 8832
rect 3068 8820 3096 8860
rect 5534 8848 5540 8900
rect 5592 8848 5598 8900
rect 6178 8848 6184 8900
rect 6236 8888 6242 8900
rect 6840 8888 6868 8928
rect 7926 8916 7932 8968
rect 7984 8916 7990 8968
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 10410 8965 10416 8968
rect 9493 8959 9551 8965
rect 9493 8956 9505 8959
rect 9180 8928 9505 8956
rect 9180 8916 9186 8928
rect 9493 8925 9505 8928
rect 9539 8925 9551 8959
rect 9493 8919 9551 8925
rect 10367 8959 10416 8965
rect 10367 8925 10379 8959
rect 10413 8925 10416 8959
rect 10367 8919 10416 8925
rect 10410 8916 10416 8919
rect 10468 8916 10474 8968
rect 10502 8916 10508 8968
rect 10560 8916 10566 8968
rect 11882 8916 11888 8968
rect 11940 8916 11946 8968
rect 12066 8916 12072 8968
rect 12124 8956 12130 8968
rect 12159 8959 12217 8965
rect 12159 8956 12171 8959
rect 12124 8928 12171 8956
rect 12124 8916 12130 8928
rect 12159 8925 12171 8928
rect 12205 8925 12217 8959
rect 12159 8919 12217 8925
rect 14826 8916 14832 8968
rect 14884 8956 14890 8968
rect 15105 8959 15163 8965
rect 15105 8956 15117 8959
rect 14884 8928 15117 8956
rect 14884 8916 14890 8928
rect 15105 8925 15117 8928
rect 15151 8925 15163 8959
rect 15363 8959 15421 8965
rect 15363 8956 15375 8959
rect 15105 8919 15163 8925
rect 15212 8928 15375 8956
rect 15212 8888 15240 8928
rect 15363 8925 15375 8928
rect 15409 8956 15421 8959
rect 15409 8925 15424 8956
rect 15363 8919 15424 8925
rect 6236 8860 6868 8888
rect 10980 8860 15240 8888
rect 15396 8888 15424 8919
rect 15470 8916 15476 8968
rect 15528 8956 15534 8968
rect 16485 8959 16543 8965
rect 16485 8956 16497 8959
rect 15528 8928 16497 8956
rect 15528 8916 15534 8928
rect 16485 8925 16497 8928
rect 16531 8925 16543 8959
rect 16485 8919 16543 8925
rect 17402 8916 17408 8968
rect 17460 8916 17466 8968
rect 17494 8916 17500 8968
rect 17552 8965 17558 8968
rect 17552 8959 17580 8965
rect 17568 8925 17580 8959
rect 17552 8919 17580 8925
rect 17552 8918 17565 8919
rect 17552 8916 17558 8918
rect 17678 8916 17684 8968
rect 17736 8916 17742 8968
rect 19889 8959 19947 8965
rect 19889 8925 19901 8959
rect 19935 8925 19947 8959
rect 19889 8919 19947 8925
rect 20349 8959 20407 8965
rect 20349 8925 20361 8959
rect 20395 8956 20407 8959
rect 20438 8956 20444 8968
rect 20395 8928 20444 8956
rect 20395 8925 20407 8928
rect 20349 8919 20407 8925
rect 15562 8888 15568 8900
rect 15396 8860 15568 8888
rect 6236 8848 6242 8860
rect 3329 8823 3387 8829
rect 3329 8820 3341 8823
rect 3068 8792 3341 8820
rect 3329 8789 3341 8792
rect 3375 8789 3387 8823
rect 3329 8783 3387 8789
rect 3418 8780 3424 8832
rect 3476 8820 3482 8832
rect 4706 8820 4712 8832
rect 3476 8792 4712 8820
rect 3476 8780 3482 8792
rect 4706 8780 4712 8792
rect 4764 8820 4770 8832
rect 5074 8820 5080 8832
rect 4764 8792 5080 8820
rect 4764 8780 4770 8792
rect 5074 8780 5080 8792
rect 5132 8820 5138 8832
rect 6454 8820 6460 8832
rect 5132 8792 6460 8820
rect 5132 8780 5138 8792
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 7466 8780 7472 8832
rect 7524 8820 7530 8832
rect 8573 8823 8631 8829
rect 8573 8820 8585 8823
rect 7524 8792 8585 8820
rect 7524 8780 7530 8792
rect 8573 8789 8585 8792
rect 8619 8789 8631 8823
rect 8573 8783 8631 8789
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 10980 8820 11008 8860
rect 15028 8832 15056 8860
rect 15562 8848 15568 8860
rect 15620 8848 15626 8900
rect 10284 8792 11008 8820
rect 10284 8780 10290 8792
rect 11146 8780 11152 8832
rect 11204 8780 11210 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 14090 8820 14096 8832
rect 12492 8792 14096 8820
rect 12492 8780 12498 8792
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 15010 8780 15016 8832
rect 15068 8780 15074 8832
rect 16114 8780 16120 8832
rect 16172 8780 16178 8832
rect 19904 8820 19932 8919
rect 20364 8888 20392 8919
rect 20438 8916 20444 8928
rect 20496 8916 20502 8968
rect 20548 8965 20576 8996
rect 21100 8996 21465 9024
rect 21100 8965 21128 8996
rect 21453 8993 21465 8996
rect 21499 8993 21511 9027
rect 21453 8987 21511 8993
rect 21634 8984 21640 9036
rect 21692 9024 21698 9036
rect 25498 9024 25504 9036
rect 21692 8996 25504 9024
rect 21692 8984 21698 8996
rect 25498 8984 25504 8996
rect 25556 8984 25562 9036
rect 20533 8959 20591 8965
rect 20533 8925 20545 8959
rect 20579 8925 20591 8959
rect 20533 8919 20591 8925
rect 21085 8959 21143 8965
rect 21085 8925 21097 8959
rect 21131 8925 21143 8959
rect 21361 8959 21419 8965
rect 21361 8956 21373 8959
rect 21085 8919 21143 8925
rect 21192 8928 21373 8956
rect 21192 8888 21220 8928
rect 21361 8925 21373 8928
rect 21407 8925 21419 8959
rect 21361 8919 21419 8925
rect 21545 8959 21603 8965
rect 21545 8925 21557 8959
rect 21591 8956 21603 8959
rect 21591 8928 21680 8956
rect 21591 8925 21603 8928
rect 21545 8919 21603 8925
rect 20364 8860 21220 8888
rect 20806 8820 20812 8832
rect 19904 8792 20812 8820
rect 20806 8780 20812 8792
rect 20864 8780 20870 8832
rect 21652 8829 21680 8928
rect 21818 8916 21824 8968
rect 21876 8916 21882 8968
rect 23017 8959 23075 8965
rect 23017 8925 23029 8959
rect 23063 8925 23075 8959
rect 23017 8919 23075 8925
rect 23032 8888 23060 8919
rect 23290 8916 23296 8968
rect 23348 8916 23354 8968
rect 23474 8916 23480 8968
rect 23532 8916 23538 8968
rect 24026 8916 24032 8968
rect 24084 8916 24090 8968
rect 23934 8888 23940 8900
rect 23032 8860 23940 8888
rect 23934 8848 23940 8860
rect 23992 8848 23998 8900
rect 21637 8823 21695 8829
rect 21637 8789 21649 8823
rect 21683 8789 21695 8823
rect 21637 8783 21695 8789
rect 22833 8823 22891 8829
rect 22833 8789 22845 8823
rect 22879 8820 22891 8823
rect 23198 8820 23204 8832
rect 22879 8792 23204 8820
rect 22879 8789 22891 8792
rect 22833 8783 22891 8789
rect 23198 8780 23204 8792
rect 23256 8780 23262 8832
rect 1104 8730 25000 8752
rect 1104 8678 6884 8730
rect 6936 8678 6948 8730
rect 7000 8678 7012 8730
rect 7064 8678 7076 8730
rect 7128 8678 7140 8730
rect 7192 8678 12818 8730
rect 12870 8678 12882 8730
rect 12934 8678 12946 8730
rect 12998 8678 13010 8730
rect 13062 8678 13074 8730
rect 13126 8678 18752 8730
rect 18804 8678 18816 8730
rect 18868 8678 18880 8730
rect 18932 8678 18944 8730
rect 18996 8678 19008 8730
rect 19060 8678 24686 8730
rect 24738 8678 24750 8730
rect 24802 8678 24814 8730
rect 24866 8678 24878 8730
rect 24930 8678 24942 8730
rect 24994 8678 25000 8730
rect 1104 8656 25000 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 1728 8588 3893 8616
rect 1728 8576 1734 8588
rect 3881 8585 3893 8588
rect 3927 8585 3939 8619
rect 3881 8579 3939 8585
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 5040 8588 5089 8616
rect 5040 8576 5046 8588
rect 5077 8585 5089 8588
rect 5123 8585 5135 8619
rect 5077 8579 5135 8585
rect 5258 8576 5264 8628
rect 5316 8616 5322 8628
rect 5534 8616 5540 8628
rect 5316 8588 5540 8616
rect 5316 8576 5322 8588
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 7190 8616 7196 8628
rect 6788 8588 7196 8616
rect 6788 8576 6794 8588
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 7282 8576 7288 8628
rect 7340 8616 7346 8628
rect 7558 8616 7564 8628
rect 7340 8588 7564 8616
rect 7340 8576 7346 8588
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 8113 8619 8171 8625
rect 8113 8616 8125 8619
rect 7984 8588 8125 8616
rect 7984 8576 7990 8588
rect 8113 8585 8125 8588
rect 8159 8585 8171 8619
rect 8113 8579 8171 8585
rect 10502 8576 10508 8628
rect 10560 8576 10566 8628
rect 10594 8576 10600 8628
rect 10652 8576 10658 8628
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 11882 8616 11888 8628
rect 10928 8588 11888 8616
rect 10928 8576 10934 8588
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 12161 8619 12219 8625
rect 12161 8585 12173 8619
rect 12207 8616 12219 8619
rect 14458 8616 14464 8628
rect 12207 8588 12848 8616
rect 12207 8585 12219 8588
rect 12161 8579 12219 8585
rect 1394 8508 1400 8560
rect 1452 8548 1458 8560
rect 1949 8551 2007 8557
rect 1949 8548 1961 8551
rect 1452 8520 1961 8548
rect 1452 8508 1458 8520
rect 1949 8517 1961 8520
rect 1995 8517 2007 8551
rect 5736 8548 5764 8576
rect 1949 8511 2007 8517
rect 3896 8520 5764 8548
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 2056 8452 2452 8480
rect 1596 8344 1624 8443
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 2056 8421 2084 8452
rect 2041 8415 2099 8421
rect 2041 8412 2053 8415
rect 1728 8384 2053 8412
rect 1728 8372 1734 8384
rect 2041 8381 2053 8384
rect 2087 8381 2099 8415
rect 2041 8375 2099 8381
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8412 2283 8415
rect 2314 8412 2320 8424
rect 2271 8384 2320 8412
rect 2271 8381 2283 8384
rect 2225 8375 2283 8381
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 2424 8412 2452 8452
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 2590 8412 2596 8424
rect 2424 8384 2596 8412
rect 2590 8372 2596 8384
rect 2648 8372 2654 8424
rect 2685 8415 2743 8421
rect 2685 8381 2697 8415
rect 2731 8412 2743 8415
rect 2774 8412 2780 8424
rect 2731 8384 2780 8412
rect 2731 8381 2743 8384
rect 2685 8375 2743 8381
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 2958 8372 2964 8424
rect 3016 8372 3022 8424
rect 3099 8415 3157 8421
rect 3099 8381 3111 8415
rect 3145 8412 3157 8415
rect 3418 8412 3424 8424
rect 3145 8384 3424 8412
rect 3145 8381 3157 8384
rect 3099 8375 3157 8381
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 3896 8344 3924 8520
rect 7300 8510 7328 8576
rect 7359 8513 7417 8519
rect 7359 8510 7371 8513
rect 4307 8483 4365 8489
rect 4307 8480 4319 8483
rect 3988 8452 4319 8480
rect 3988 8424 4016 8452
rect 4307 8449 4319 8452
rect 4353 8480 4365 8483
rect 6546 8480 6552 8492
rect 4353 8452 6552 8480
rect 4353 8449 4365 8452
rect 4307 8443 4365 8449
rect 6546 8440 6552 8452
rect 6604 8440 6610 8492
rect 7300 8482 7371 8510
rect 7359 8479 7371 8482
rect 7405 8479 7417 8513
rect 7650 8508 7656 8560
rect 7708 8548 7714 8560
rect 10612 8548 10640 8576
rect 12250 8548 12256 8560
rect 7708 8520 12256 8548
rect 7708 8508 7714 8520
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 12434 8508 12440 8560
rect 12492 8508 12498 8560
rect 7359 8473 7417 8479
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 9735 8483 9793 8489
rect 9735 8480 9747 8483
rect 7984 8452 9747 8480
rect 7984 8440 7990 8452
rect 9735 8449 9747 8452
rect 9781 8449 9793 8483
rect 9735 8443 9793 8449
rect 12342 8440 12348 8492
rect 12400 8480 12406 8492
rect 12529 8483 12587 8489
rect 12529 8480 12541 8483
rect 12400 8452 12541 8480
rect 12400 8440 12406 8452
rect 12529 8449 12541 8452
rect 12575 8449 12587 8483
rect 12820 8480 12848 8588
rect 13188 8588 14464 8616
rect 13188 8560 13216 8588
rect 14458 8576 14464 8588
rect 14516 8616 14522 8628
rect 14516 8588 14596 8616
rect 14516 8576 14522 8588
rect 12897 8551 12955 8557
rect 12897 8517 12909 8551
rect 12943 8548 12955 8551
rect 13170 8548 13176 8560
rect 12943 8520 13176 8548
rect 12943 8517 12955 8520
rect 12897 8511 12955 8517
rect 13170 8508 13176 8520
rect 13228 8508 13234 8560
rect 13265 8551 13323 8557
rect 13265 8517 13277 8551
rect 13311 8548 13323 8551
rect 13311 8520 13400 8548
rect 13311 8517 13323 8520
rect 13265 8511 13323 8517
rect 13372 8480 13400 8520
rect 13630 8508 13636 8560
rect 13688 8548 13694 8560
rect 14568 8557 14596 8588
rect 16574 8576 16580 8628
rect 16632 8576 16638 8628
rect 16758 8576 16764 8628
rect 16816 8616 16822 8628
rect 17034 8616 17040 8628
rect 16816 8588 17040 8616
rect 16816 8576 16822 8588
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17681 8619 17739 8625
rect 17681 8616 17693 8619
rect 17184 8588 17693 8616
rect 17184 8576 17190 8588
rect 17681 8585 17693 8588
rect 17727 8585 17739 8619
rect 17681 8579 17739 8585
rect 21453 8619 21511 8625
rect 21453 8585 21465 8619
rect 21499 8616 21511 8619
rect 21818 8616 21824 8628
rect 21499 8588 21824 8616
rect 21499 8585 21511 8588
rect 21453 8579 21511 8585
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 22925 8619 22983 8625
rect 22925 8585 22937 8619
rect 22971 8616 22983 8619
rect 23474 8616 23480 8628
rect 22971 8588 23480 8616
rect 22971 8585 22983 8588
rect 22925 8579 22983 8585
rect 23474 8576 23480 8588
rect 23532 8576 23538 8628
rect 13817 8551 13875 8557
rect 13817 8548 13829 8551
rect 13688 8520 13829 8548
rect 13688 8508 13694 8520
rect 13817 8517 13829 8520
rect 13863 8517 13875 8551
rect 14553 8551 14611 8557
rect 13817 8511 13875 8517
rect 14016 8520 14320 8548
rect 14016 8492 14044 8520
rect 13998 8480 14004 8492
rect 12820 8452 13308 8480
rect 13372 8452 14004 8480
rect 12529 8443 12587 8449
rect 3970 8372 3976 8424
rect 4028 8372 4034 8424
rect 4065 8415 4123 8421
rect 4065 8381 4077 8415
rect 4111 8381 4123 8415
rect 6638 8412 6644 8424
rect 4065 8375 4123 8381
rect 4724 8384 6644 8412
rect 1596 8316 2820 8344
rect 2792 8276 2820 8316
rect 3620 8316 3924 8344
rect 4080 8344 4108 8375
rect 4080 8316 4200 8344
rect 3620 8276 3648 8316
rect 4172 8288 4200 8316
rect 2792 8248 3648 8276
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4724 8276 4752 8384
rect 6638 8372 6644 8384
rect 6696 8412 6702 8424
rect 7101 8415 7159 8421
rect 7101 8412 7113 8415
rect 6696 8384 7113 8412
rect 6696 8372 6702 8384
rect 7101 8381 7113 8384
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 9493 8415 9551 8421
rect 9493 8412 9505 8415
rect 9364 8384 9505 8412
rect 9364 8372 9370 8384
rect 9493 8381 9505 8384
rect 9539 8381 9551 8415
rect 9493 8375 9551 8381
rect 12986 8372 12992 8424
rect 13044 8372 13050 8424
rect 13280 8412 13308 8452
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 14090 8440 14096 8492
rect 14148 8440 14154 8492
rect 14182 8440 14188 8492
rect 14240 8440 14246 8492
rect 14292 8480 14320 8520
rect 14553 8517 14565 8551
rect 14599 8517 14611 8551
rect 14553 8511 14611 8517
rect 14918 8508 14924 8560
rect 14976 8508 14982 8560
rect 16592 8548 16620 8576
rect 19426 8548 19432 8560
rect 16592 8520 16896 8548
rect 14936 8480 14964 8508
rect 14292 8452 14964 8480
rect 16666 8440 16672 8492
rect 16724 8440 16730 8492
rect 16868 8480 16896 8520
rect 17604 8520 19432 8548
rect 16927 8483 16985 8489
rect 16927 8480 16939 8483
rect 16868 8452 16939 8480
rect 16927 8449 16939 8452
rect 16973 8480 16985 8483
rect 17604 8480 17632 8520
rect 19426 8508 19432 8520
rect 19484 8508 19490 8560
rect 23658 8548 23664 8560
rect 20088 8520 21588 8548
rect 16973 8452 17632 8480
rect 16973 8449 16985 8452
rect 16927 8443 16985 8449
rect 18046 8440 18052 8492
rect 18104 8480 18110 8492
rect 19242 8480 19248 8492
rect 18104 8452 19248 8480
rect 18104 8440 18110 8452
rect 19242 8440 19248 8452
rect 19300 8480 19306 8492
rect 20088 8489 20116 8520
rect 20073 8483 20131 8489
rect 20073 8480 20085 8483
rect 19300 8452 20085 8480
rect 19300 8440 19306 8452
rect 20073 8449 20085 8452
rect 20119 8449 20131 8483
rect 20073 8443 20131 8449
rect 20340 8483 20398 8489
rect 20340 8449 20352 8483
rect 20386 8480 20398 8483
rect 21082 8480 21088 8492
rect 20386 8452 21088 8480
rect 20386 8449 20398 8452
rect 20340 8443 20398 8449
rect 21082 8440 21088 8452
rect 21140 8440 21146 8492
rect 21560 8424 21588 8520
rect 22848 8520 23664 8548
rect 22848 8489 22876 8520
rect 23658 8508 23664 8520
rect 23716 8508 23722 8560
rect 22833 8483 22891 8489
rect 22833 8449 22845 8483
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 23198 8440 23204 8492
rect 23256 8480 23262 8492
rect 23365 8483 23423 8489
rect 23365 8480 23377 8483
rect 23256 8452 23377 8480
rect 23256 8440 23262 8452
rect 23365 8449 23377 8452
rect 23411 8480 23423 8483
rect 23750 8480 23756 8492
rect 23411 8452 23756 8480
rect 23411 8449 23423 8452
rect 23365 8443 23423 8449
rect 23750 8440 23756 8452
rect 23808 8440 23814 8492
rect 13280 8384 13400 8412
rect 5166 8304 5172 8356
rect 5224 8344 5230 8356
rect 6086 8344 6092 8356
rect 5224 8316 6092 8344
rect 5224 8304 5230 8316
rect 6086 8304 6092 8316
rect 6144 8304 6150 8356
rect 4212 8248 4752 8276
rect 4212 8236 4218 8248
rect 6822 8236 6828 8288
rect 6880 8276 6886 8288
rect 9214 8276 9220 8288
rect 6880 8248 9220 8276
rect 6880 8236 6886 8248
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 9490 8236 9496 8288
rect 9548 8276 9554 8288
rect 11054 8276 11060 8288
rect 9548 8248 11060 8276
rect 9548 8236 9554 8248
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 13372 8276 13400 8384
rect 13446 8304 13452 8356
rect 13504 8304 13510 8356
rect 13832 8288 13860 8398
rect 21542 8372 21548 8424
rect 21600 8412 21606 8424
rect 23109 8415 23167 8421
rect 23109 8412 23121 8415
rect 21600 8384 23121 8412
rect 21600 8372 21606 8384
rect 23109 8381 23121 8384
rect 23155 8381 23167 8415
rect 23109 8375 23167 8381
rect 15105 8347 15163 8353
rect 15105 8313 15117 8347
rect 15151 8344 15163 8347
rect 16390 8344 16396 8356
rect 15151 8316 16396 8344
rect 15151 8313 15163 8316
rect 15105 8307 15163 8313
rect 16390 8304 16396 8316
rect 16448 8304 16454 8356
rect 21634 8344 21640 8356
rect 19306 8316 20116 8344
rect 13630 8276 13636 8288
rect 13372 8248 13636 8276
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 13814 8236 13820 8288
rect 13872 8236 13878 8288
rect 15010 8236 15016 8288
rect 15068 8276 15074 8288
rect 19306 8276 19334 8316
rect 15068 8248 19334 8276
rect 20088 8276 20116 8316
rect 21008 8316 21640 8344
rect 21008 8276 21036 8316
rect 21634 8304 21640 8316
rect 21692 8304 21698 8356
rect 20088 8248 21036 8276
rect 15068 8236 15074 8248
rect 22094 8236 22100 8288
rect 22152 8276 22158 8288
rect 24489 8279 24547 8285
rect 24489 8276 24501 8279
rect 22152 8248 24501 8276
rect 22152 8236 22158 8248
rect 24489 8245 24501 8248
rect 24535 8245 24547 8279
rect 24489 8239 24547 8245
rect 1104 8186 24840 8208
rect 1104 8134 3917 8186
rect 3969 8134 3981 8186
rect 4033 8134 4045 8186
rect 4097 8134 4109 8186
rect 4161 8134 4173 8186
rect 4225 8134 9851 8186
rect 9903 8134 9915 8186
rect 9967 8134 9979 8186
rect 10031 8134 10043 8186
rect 10095 8134 10107 8186
rect 10159 8134 15785 8186
rect 15837 8134 15849 8186
rect 15901 8134 15913 8186
rect 15965 8134 15977 8186
rect 16029 8134 16041 8186
rect 16093 8134 21719 8186
rect 21771 8134 21783 8186
rect 21835 8134 21847 8186
rect 21899 8134 21911 8186
rect 21963 8134 21975 8186
rect 22027 8134 24840 8186
rect 1104 8112 24840 8134
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 1544 8044 1593 8072
rect 1544 8032 1550 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 1581 8035 1639 8041
rect 1946 8032 1952 8084
rect 2004 8032 2010 8084
rect 2498 8032 2504 8084
rect 2556 8072 2562 8084
rect 2556 8044 3188 8072
rect 2556 8032 2562 8044
rect 3160 8004 3188 8044
rect 3234 8032 3240 8084
rect 3292 8032 3298 8084
rect 4338 8032 4344 8084
rect 4396 8072 4402 8084
rect 6822 8072 6828 8084
rect 4396 8044 6828 8072
rect 4396 8032 4402 8044
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 8389 8075 8447 8081
rect 8389 8072 8401 8075
rect 7392 8044 8401 8072
rect 3789 8007 3847 8013
rect 3789 8004 3801 8007
rect 3160 7976 3801 8004
rect 3789 7973 3801 7976
rect 3835 7973 3847 8007
rect 3789 7967 3847 7973
rect 5077 8007 5135 8013
rect 5077 7973 5089 8007
rect 5123 8004 5135 8007
rect 6089 8007 6147 8013
rect 6089 8004 6101 8007
rect 5123 7976 6101 8004
rect 5123 7973 5135 7976
rect 5077 7967 5135 7973
rect 6089 7973 6101 7976
rect 6135 7973 6147 8007
rect 6089 7967 6147 7973
rect 7282 7964 7288 8016
rect 7340 7964 7346 8016
rect 1210 7896 1216 7948
rect 1268 7936 1274 7948
rect 2225 7939 2283 7945
rect 2225 7936 2237 7939
rect 1268 7908 2237 7936
rect 1268 7896 1274 7908
rect 2225 7905 2237 7908
rect 2271 7905 2283 7939
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 2225 7899 2283 7905
rect 3436 7908 4077 7936
rect 2130 7828 2136 7880
rect 2188 7828 2194 7880
rect 1486 7760 1492 7812
rect 1544 7760 1550 7812
rect 2240 7800 2268 7899
rect 2499 7871 2557 7877
rect 2499 7837 2511 7871
rect 2545 7868 2557 7871
rect 3326 7868 3332 7880
rect 2545 7840 3332 7868
rect 2545 7837 2557 7840
rect 2499 7831 2557 7837
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 3436 7800 3464 7908
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 5994 7936 6000 7948
rect 4065 7899 4123 7905
rect 5368 7908 6000 7936
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4339 7871 4397 7877
rect 4339 7837 4351 7871
rect 4385 7868 4397 7871
rect 5368 7868 5396 7908
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6178 7896 6184 7948
rect 6236 7936 6242 7948
rect 6365 7939 6423 7945
rect 6365 7936 6377 7939
rect 6236 7908 6377 7936
rect 6236 7896 6242 7908
rect 6365 7905 6377 7908
rect 6411 7905 6423 7939
rect 6365 7899 6423 7905
rect 6454 7896 6460 7948
rect 6512 7945 6518 7948
rect 6512 7939 6540 7945
rect 6528 7905 6540 7939
rect 6512 7899 6540 7905
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7936 6699 7939
rect 7392 7936 7420 8044
rect 8389 8041 8401 8044
rect 8435 8041 8447 8075
rect 8389 8035 8447 8041
rect 9048 8044 9628 8072
rect 8662 8004 8668 8016
rect 8404 7976 8668 8004
rect 8404 7948 8432 7976
rect 8662 7964 8668 7976
rect 8720 8004 8726 8016
rect 9048 8004 9076 8044
rect 8720 7976 9076 8004
rect 9600 8004 9628 8044
rect 9766 8032 9772 8084
rect 9824 8072 9830 8084
rect 9953 8075 10011 8081
rect 9953 8072 9965 8075
rect 9824 8044 9965 8072
rect 9824 8032 9830 8044
rect 9953 8041 9965 8044
rect 9999 8041 10011 8075
rect 16482 8072 16488 8084
rect 9953 8035 10011 8041
rect 10888 8044 12434 8072
rect 10888 8004 10916 8044
rect 9600 7976 10916 8004
rect 12406 8004 12434 8044
rect 15948 8044 16488 8072
rect 13446 8004 13452 8016
rect 12406 7976 13452 8004
rect 8720 7964 8726 7976
rect 13446 7964 13452 7976
rect 13504 7964 13510 8016
rect 6687 7908 7420 7936
rect 6687 7905 6699 7908
rect 6641 7899 6699 7905
rect 6512 7896 6518 7899
rect 8386 7896 8392 7948
rect 8444 7896 8450 7948
rect 11790 7896 11796 7948
rect 11848 7936 11854 7948
rect 15565 7939 15623 7945
rect 15565 7936 15577 7939
rect 11848 7908 15577 7936
rect 11848 7896 11854 7908
rect 15565 7905 15577 7908
rect 15611 7936 15623 7939
rect 15948 7936 15976 8044
rect 16482 8032 16488 8044
rect 16540 8072 16546 8084
rect 16540 8044 20208 8072
rect 16540 8032 16546 8044
rect 16025 8007 16083 8013
rect 16025 7973 16037 8007
rect 16071 8004 16083 8007
rect 16114 8004 16120 8016
rect 16071 7976 16120 8004
rect 16071 7973 16083 7976
rect 16025 7967 16083 7973
rect 16114 7964 16120 7976
rect 16172 7964 16178 8016
rect 20180 8013 20208 8044
rect 20622 8032 20628 8084
rect 20680 8072 20686 8084
rect 20990 8072 20996 8084
rect 20680 8044 20852 8072
rect 20680 8032 20686 8044
rect 20165 8007 20223 8013
rect 20165 7973 20177 8007
rect 20211 7973 20223 8007
rect 20165 7967 20223 7973
rect 15611 7908 15976 7936
rect 15611 7905 15623 7908
rect 15565 7899 15623 7905
rect 16298 7896 16304 7948
rect 16356 7896 16362 7948
rect 16390 7896 16396 7948
rect 16448 7945 16454 7948
rect 16448 7939 16476 7945
rect 16464 7905 16476 7939
rect 20625 7939 20683 7945
rect 20625 7936 20637 7939
rect 16448 7899 16476 7905
rect 20272 7908 20637 7936
rect 16448 7896 16454 7899
rect 4385 7840 5396 7868
rect 5445 7871 5503 7877
rect 4385 7837 4397 7840
rect 4339 7831 4397 7837
rect 5445 7837 5457 7871
rect 5491 7868 5503 7871
rect 5534 7868 5540 7880
rect 5491 7840 5540 7868
rect 5491 7837 5503 7840
rect 5445 7831 5503 7837
rect 2240 7772 3464 7800
rect 3988 7732 4016 7831
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 5626 7828 5632 7880
rect 5684 7828 5690 7880
rect 7377 7871 7435 7877
rect 7377 7868 7389 7871
rect 7208 7840 7389 7868
rect 7208 7812 7236 7840
rect 7377 7837 7389 7840
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 7558 7828 7564 7880
rect 7616 7868 7622 7880
rect 7651 7871 7709 7877
rect 7651 7868 7663 7871
rect 7616 7840 7663 7868
rect 7616 7828 7622 7840
rect 7651 7837 7663 7840
rect 7697 7837 7709 7871
rect 7651 7831 7709 7837
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 7190 7760 7196 7812
rect 7248 7760 7254 7812
rect 8956 7800 8984 7831
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7837 10839 7871
rect 10781 7831 10839 7837
rect 11055 7871 11113 7877
rect 11055 7837 11067 7871
rect 11101 7868 11113 7871
rect 11698 7868 11704 7880
rect 11101 7840 11704 7868
rect 11101 7837 11113 7840
rect 11055 7831 11113 7837
rect 9306 7800 9312 7812
rect 8956 7772 9312 7800
rect 9306 7760 9312 7772
rect 9364 7800 9370 7812
rect 9858 7800 9864 7812
rect 9364 7772 9864 7800
rect 9364 7760 9370 7772
rect 9858 7760 9864 7772
rect 9916 7800 9922 7812
rect 10796 7800 10824 7831
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 15381 7871 15439 7877
rect 15381 7868 15393 7871
rect 15252 7840 15393 7868
rect 15252 7828 15258 7840
rect 15381 7837 15393 7840
rect 15427 7868 15439 7871
rect 15470 7868 15476 7880
rect 15427 7840 15476 7868
rect 15427 7837 15439 7840
rect 15381 7831 15439 7837
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 16574 7828 16580 7880
rect 16632 7828 16638 7880
rect 19521 7871 19579 7877
rect 19521 7837 19533 7871
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 9916 7772 10824 7800
rect 11624 7772 12434 7800
rect 9916 7760 9922 7772
rect 11624 7732 11652 7772
rect 3988 7704 11652 7732
rect 11698 7692 11704 7744
rect 11756 7732 11762 7744
rect 11793 7735 11851 7741
rect 11793 7732 11805 7735
rect 11756 7704 11805 7732
rect 11756 7692 11762 7704
rect 11793 7701 11805 7704
rect 11839 7701 11851 7735
rect 12406 7732 12434 7772
rect 12986 7760 12992 7812
rect 13044 7800 13050 7812
rect 13906 7800 13912 7812
rect 13044 7772 13912 7800
rect 13044 7760 13050 7772
rect 13906 7760 13912 7772
rect 13964 7760 13970 7812
rect 19536 7800 19564 7831
rect 19702 7828 19708 7880
rect 19760 7828 19766 7880
rect 20272 7877 20300 7908
rect 20625 7905 20637 7908
rect 20671 7905 20683 7939
rect 20625 7899 20683 7905
rect 20257 7871 20315 7877
rect 20257 7837 20269 7871
rect 20303 7837 20315 7871
rect 20533 7871 20591 7877
rect 20533 7868 20545 7871
rect 20257 7831 20315 7837
rect 20364 7840 20545 7868
rect 20162 7800 20168 7812
rect 19536 7772 20168 7800
rect 20162 7760 20168 7772
rect 20220 7800 20226 7812
rect 20364 7800 20392 7840
rect 20533 7837 20545 7840
rect 20579 7837 20591 7871
rect 20533 7831 20591 7837
rect 20714 7828 20720 7880
rect 20772 7828 20778 7880
rect 20824 7868 20852 8044
rect 20916 8044 20996 8072
rect 20916 7945 20944 8044
rect 20990 8032 20996 8044
rect 21048 8072 21054 8084
rect 21048 8044 22094 8072
rect 21048 8032 21054 8044
rect 20901 7939 20959 7945
rect 20901 7905 20913 7939
rect 20947 7905 20959 7939
rect 22066 7936 22094 8044
rect 23290 8032 23296 8084
rect 23348 8072 23354 8084
rect 23474 8072 23480 8084
rect 23348 8044 23480 8072
rect 23348 8032 23354 8044
rect 23474 8032 23480 8044
rect 23532 8032 23538 8084
rect 23566 8032 23572 8084
rect 23624 8072 23630 8084
rect 23937 8075 23995 8081
rect 23937 8072 23949 8075
rect 23624 8044 23949 8072
rect 23624 8032 23630 8044
rect 23937 8041 23949 8044
rect 23983 8041 23995 8075
rect 23937 8035 23995 8041
rect 23661 8007 23719 8013
rect 23661 7973 23673 8007
rect 23707 8004 23719 8007
rect 24210 8004 24216 8016
rect 23707 7976 24216 8004
rect 23707 7973 23719 7976
rect 23661 7967 23719 7973
rect 24210 7964 24216 7976
rect 24268 7964 24274 8016
rect 22281 7939 22339 7945
rect 22281 7936 22293 7939
rect 22066 7908 22293 7936
rect 20901 7899 20959 7905
rect 22204 7880 22232 7908
rect 22281 7905 22293 7908
rect 22327 7905 22339 7939
rect 22281 7899 22339 7905
rect 21143 7871 21201 7877
rect 21143 7868 21155 7871
rect 20824 7840 21155 7868
rect 21143 7837 21155 7840
rect 21189 7837 21201 7871
rect 21143 7831 21201 7837
rect 22186 7828 22192 7880
rect 22244 7828 22250 7880
rect 22554 7828 22560 7880
rect 22612 7828 22618 7880
rect 23842 7828 23848 7880
rect 23900 7828 23906 7880
rect 24118 7828 24124 7880
rect 24176 7828 24182 7880
rect 24210 7800 24216 7812
rect 20220 7772 20392 7800
rect 20548 7772 24216 7800
rect 20220 7760 20226 7772
rect 20548 7744 20576 7772
rect 24210 7760 24216 7772
rect 24268 7760 24274 7812
rect 17221 7735 17279 7741
rect 17221 7732 17233 7735
rect 12406 7704 17233 7732
rect 11793 7695 11851 7701
rect 17221 7701 17233 7704
rect 17267 7701 17279 7735
rect 17221 7695 17279 7701
rect 20530 7692 20536 7744
rect 20588 7692 20594 7744
rect 21913 7735 21971 7741
rect 21913 7701 21925 7735
rect 21959 7732 21971 7735
rect 22094 7732 22100 7744
rect 21959 7704 22100 7732
rect 21959 7701 21971 7704
rect 21913 7695 21971 7701
rect 22094 7692 22100 7704
rect 22152 7692 22158 7744
rect 22186 7692 22192 7744
rect 22244 7732 22250 7744
rect 22554 7732 22560 7744
rect 22244 7704 22560 7732
rect 22244 7692 22250 7704
rect 22554 7692 22560 7704
rect 22612 7692 22618 7744
rect 1104 7642 25000 7664
rect 1104 7590 6884 7642
rect 6936 7590 6948 7642
rect 7000 7590 7012 7642
rect 7064 7590 7076 7642
rect 7128 7590 7140 7642
rect 7192 7590 12818 7642
rect 12870 7590 12882 7642
rect 12934 7590 12946 7642
rect 12998 7590 13010 7642
rect 13062 7590 13074 7642
rect 13126 7590 18752 7642
rect 18804 7590 18816 7642
rect 18868 7590 18880 7642
rect 18932 7590 18944 7642
rect 18996 7590 19008 7642
rect 19060 7590 24686 7642
rect 24738 7590 24750 7642
rect 24802 7590 24814 7642
rect 24866 7590 24878 7642
rect 24930 7590 24942 7642
rect 24994 7590 25000 7642
rect 1104 7568 25000 7590
rect 1302 7488 1308 7540
rect 1360 7528 1366 7540
rect 3237 7531 3295 7537
rect 3237 7528 3249 7531
rect 1360 7500 3249 7528
rect 1360 7488 1366 7500
rect 3237 7497 3249 7500
rect 3283 7497 3295 7531
rect 3237 7491 3295 7497
rect 3789 7531 3847 7537
rect 3789 7497 3801 7531
rect 3835 7497 3847 7531
rect 3789 7491 3847 7497
rect 1854 7420 1860 7472
rect 1912 7420 1918 7472
rect 2409 7463 2467 7469
rect 2409 7429 2421 7463
rect 2455 7460 2467 7463
rect 2866 7460 2872 7472
rect 2455 7432 2872 7460
rect 2455 7429 2467 7432
rect 2409 7423 2467 7429
rect 2866 7420 2872 7432
rect 2924 7420 2930 7472
rect 3145 7463 3203 7469
rect 3145 7429 3157 7463
rect 3191 7460 3203 7463
rect 3804 7460 3832 7491
rect 4246 7488 4252 7540
rect 4304 7488 4310 7540
rect 7282 7488 7288 7540
rect 7340 7488 7346 7540
rect 7374 7488 7380 7540
rect 7432 7528 7438 7540
rect 7469 7531 7527 7537
rect 7469 7528 7481 7531
rect 7432 7500 7481 7528
rect 7432 7488 7438 7500
rect 7469 7497 7481 7500
rect 7515 7497 7527 7531
rect 7469 7491 7527 7497
rect 7650 7488 7656 7540
rect 7708 7488 7714 7540
rect 9398 7488 9404 7540
rect 9456 7488 9462 7540
rect 13725 7531 13783 7537
rect 9508 7500 13032 7528
rect 3191 7432 3832 7460
rect 3191 7429 3203 7432
rect 3145 7423 3203 7429
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7392 1547 7395
rect 1946 7392 1952 7404
rect 1535 7364 1952 7392
rect 1535 7361 1547 7364
rect 1489 7355 1547 7361
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 2056 7324 2084 7355
rect 2498 7352 2504 7404
rect 2556 7392 2562 7404
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2556 7364 2605 7392
rect 2556 7352 2562 7364
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 3694 7352 3700 7404
rect 3752 7392 3758 7404
rect 4264 7401 4292 7488
rect 7300 7460 7328 7488
rect 4540 7432 7328 7460
rect 7668 7460 7696 7488
rect 7926 7460 7932 7472
rect 7668 7432 7932 7460
rect 4540 7401 4568 7432
rect 7926 7420 7932 7432
rect 7984 7460 7990 7472
rect 9508 7460 9536 7500
rect 7984 7432 9536 7460
rect 7984 7420 7990 7432
rect 9858 7420 9864 7472
rect 9916 7420 9922 7472
rect 12526 7460 12532 7472
rect 11072 7432 12532 7460
rect 10027 7425 10085 7431
rect 3973 7395 4031 7401
rect 3973 7392 3985 7395
rect 3752 7364 3985 7392
rect 3752 7352 3758 7364
rect 3973 7361 3985 7364
rect 4019 7361 4031 7395
rect 3973 7355 4031 7361
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 6699 7395 6757 7401
rect 6699 7392 6711 7395
rect 6052 7364 6711 7392
rect 6052 7352 6058 7364
rect 6699 7361 6711 7364
rect 6745 7361 6757 7395
rect 6699 7355 6757 7361
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7282 7392 7288 7404
rect 6880 7364 7288 7392
rect 6880 7352 6886 7364
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7392 9275 7395
rect 9674 7392 9680 7404
rect 9263 7364 9680 7392
rect 9263 7361 9275 7364
rect 9217 7355 9275 7361
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7392 9827 7395
rect 9876 7392 9904 7420
rect 9815 7364 9904 7392
rect 10027 7391 10039 7425
rect 10073 7392 10085 7425
rect 10962 7392 10968 7404
rect 10073 7391 10968 7392
rect 10027 7385 10968 7391
rect 10042 7364 10968 7385
rect 9815 7361 9827 7364
rect 9769 7355 9827 7361
rect 2056 7296 4384 7324
rect 1302 7216 1308 7268
rect 1360 7256 1366 7268
rect 1360 7228 2728 7256
rect 1360 7216 1366 7228
rect 2700 7197 2728 7228
rect 2958 7216 2964 7268
rect 3016 7216 3022 7268
rect 3694 7216 3700 7268
rect 3752 7256 3758 7268
rect 4356 7265 4384 7296
rect 6086 7284 6092 7336
rect 6144 7324 6150 7336
rect 6457 7327 6515 7333
rect 6457 7324 6469 7327
rect 6144 7296 6469 7324
rect 6144 7284 6150 7296
rect 6457 7293 6469 7296
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 4065 7259 4123 7265
rect 4065 7256 4077 7259
rect 3752 7228 4077 7256
rect 3752 7216 3758 7228
rect 4065 7225 4077 7228
rect 4111 7225 4123 7259
rect 4065 7219 4123 7225
rect 4341 7259 4399 7265
rect 4341 7225 4353 7259
rect 4387 7225 4399 7259
rect 6178 7256 6184 7268
rect 4341 7219 4399 7225
rect 5000 7228 6184 7256
rect 2685 7191 2743 7197
rect 2685 7157 2697 7191
rect 2731 7157 2743 7191
rect 2976 7188 3004 7216
rect 5000 7188 5028 7228
rect 6178 7216 6184 7228
rect 6236 7216 6242 7268
rect 9214 7216 9220 7268
rect 9272 7256 9278 7268
rect 9784 7256 9812 7355
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11072 7256 11100 7432
rect 12526 7420 12532 7432
rect 12584 7420 12590 7472
rect 13004 7431 13032 7500
rect 13725 7497 13737 7531
rect 13771 7528 13783 7531
rect 13814 7528 13820 7540
rect 13771 7500 13820 7528
rect 13771 7497 13783 7500
rect 13725 7491 13783 7497
rect 13814 7488 13820 7500
rect 13872 7488 13878 7540
rect 14182 7488 14188 7540
rect 14240 7528 14246 7540
rect 15105 7531 15163 7537
rect 15105 7528 15117 7531
rect 14240 7500 15117 7528
rect 14240 7488 14246 7500
rect 15105 7497 15117 7500
rect 15151 7497 15163 7531
rect 15105 7491 15163 7497
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 17681 7531 17739 7537
rect 17681 7528 17693 7531
rect 16632 7500 17693 7528
rect 16632 7488 16638 7500
rect 17681 7497 17693 7500
rect 17727 7497 17739 7531
rect 17681 7491 17739 7497
rect 18693 7531 18751 7537
rect 18693 7497 18705 7531
rect 18739 7497 18751 7531
rect 18693 7491 18751 7497
rect 19061 7531 19119 7537
rect 19061 7497 19073 7531
rect 19107 7528 19119 7531
rect 19702 7528 19708 7540
rect 19107 7500 19708 7528
rect 19107 7497 19119 7500
rect 19061 7491 19119 7497
rect 12971 7425 13032 7431
rect 11882 7352 11888 7404
rect 11940 7392 11946 7404
rect 11940 7364 12756 7392
rect 12971 7391 12983 7425
rect 13017 7394 13032 7425
rect 13262 7420 13268 7472
rect 13320 7460 13326 7472
rect 18708 7460 18736 7491
rect 19702 7488 19708 7500
rect 19760 7488 19766 7540
rect 20530 7488 20536 7540
rect 20588 7488 20594 7540
rect 20625 7531 20683 7537
rect 20625 7497 20637 7531
rect 20671 7497 20683 7531
rect 20625 7491 20683 7497
rect 19512 7463 19570 7469
rect 19512 7460 19524 7463
rect 13320 7432 16436 7460
rect 18708 7432 19012 7460
rect 13320 7420 13326 7432
rect 16408 7404 16436 7432
rect 16927 7405 16985 7411
rect 13017 7391 13029 7394
rect 12971 7385 13029 7391
rect 11940 7352 11946 7364
rect 12728 7333 12756 7364
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 14335 7395 14393 7401
rect 14335 7392 14347 7395
rect 13504 7364 14347 7392
rect 13504 7352 13510 7364
rect 14335 7361 14347 7364
rect 14381 7361 14393 7395
rect 14335 7355 14393 7361
rect 16390 7352 16396 7404
rect 16448 7392 16454 7404
rect 16927 7392 16939 7405
rect 16448 7371 16939 7392
rect 16973 7371 16985 7405
rect 16448 7365 16985 7371
rect 16448 7364 16970 7365
rect 16448 7352 16454 7364
rect 18230 7352 18236 7404
rect 18288 7352 18294 7404
rect 18601 7395 18659 7401
rect 18601 7361 18613 7395
rect 18647 7392 18659 7395
rect 18782 7392 18788 7404
rect 18647 7364 18788 7392
rect 18647 7361 18659 7364
rect 18601 7355 18659 7361
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 18984 7401 19012 7432
rect 19168 7432 19524 7460
rect 18877 7395 18935 7401
rect 18877 7361 18889 7395
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 18969 7395 19027 7401
rect 18969 7361 18981 7395
rect 19015 7361 19027 7395
rect 18969 7355 19027 7361
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 14093 7327 14151 7333
rect 14093 7293 14105 7327
rect 14139 7293 14151 7327
rect 14093 7287 14151 7293
rect 9272 7228 9812 7256
rect 10428 7228 11100 7256
rect 9272 7216 9278 7228
rect 2976 7160 5028 7188
rect 2685 7151 2743 7157
rect 5074 7148 5080 7200
rect 5132 7188 5138 7200
rect 10428 7188 10456 7228
rect 5132 7160 10456 7188
rect 10781 7191 10839 7197
rect 5132 7148 5138 7160
rect 10781 7157 10793 7191
rect 10827 7188 10839 7191
rect 11054 7188 11060 7200
rect 10827 7160 11060 7188
rect 10827 7157 10839 7160
rect 10781 7151 10839 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 12728 7188 12756 7287
rect 14108 7256 14136 7287
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 16666 7324 16672 7336
rect 14884 7296 16672 7324
rect 14884 7284 14890 7296
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 18322 7284 18328 7336
rect 18380 7284 18386 7336
rect 18892 7324 18920 7355
rect 19168 7324 19196 7432
rect 19512 7429 19524 7432
rect 19558 7460 19570 7463
rect 20548 7460 20576 7488
rect 19558 7432 20576 7460
rect 20640 7460 20668 7491
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 20993 7531 21051 7537
rect 20993 7528 21005 7531
rect 20772 7500 21005 7528
rect 20772 7488 20778 7500
rect 20993 7497 21005 7500
rect 21039 7497 21051 7531
rect 20993 7491 21051 7497
rect 21450 7488 21456 7540
rect 21508 7528 21514 7540
rect 23293 7531 23351 7537
rect 23293 7528 23305 7531
rect 21508 7500 23305 7528
rect 21508 7488 21514 7500
rect 23293 7497 23305 7500
rect 23339 7497 23351 7531
rect 23293 7491 23351 7497
rect 23658 7488 23664 7540
rect 23716 7488 23722 7540
rect 24026 7488 24032 7540
rect 24084 7488 24090 7540
rect 24210 7488 24216 7540
rect 24268 7528 24274 7540
rect 24397 7531 24455 7537
rect 24397 7528 24409 7531
rect 24268 7500 24409 7528
rect 24268 7488 24274 7500
rect 24397 7497 24409 7500
rect 24443 7497 24455 7531
rect 24397 7491 24455 7497
rect 22002 7460 22008 7472
rect 20640 7432 21220 7460
rect 19558 7429 19570 7432
rect 19512 7423 19570 7429
rect 19242 7352 19248 7404
rect 19300 7352 19306 7404
rect 21192 7401 21220 7432
rect 21652 7432 22008 7460
rect 21652 7401 21680 7432
rect 22002 7420 22008 7432
rect 22060 7420 22066 7472
rect 22296 7432 24164 7460
rect 20901 7395 20959 7401
rect 20901 7361 20913 7395
rect 20947 7392 20959 7395
rect 21177 7395 21235 7401
rect 20947 7364 21128 7392
rect 20947 7361 20959 7364
rect 20901 7355 20959 7361
rect 21100 7336 21128 7364
rect 21177 7361 21189 7395
rect 21223 7361 21235 7395
rect 21177 7355 21235 7361
rect 21637 7395 21695 7401
rect 21637 7361 21649 7395
rect 21683 7361 21695 7395
rect 21637 7355 21695 7361
rect 21913 7395 21971 7401
rect 21913 7361 21925 7395
rect 21959 7361 21971 7395
rect 21913 7355 21971 7361
rect 18892 7296 19196 7324
rect 21082 7284 21088 7336
rect 21140 7284 21146 7336
rect 21266 7284 21272 7336
rect 21324 7324 21330 7336
rect 21928 7324 21956 7355
rect 22094 7352 22100 7404
rect 22152 7392 22158 7404
rect 22189 7395 22247 7401
rect 22189 7392 22201 7395
rect 22152 7364 22201 7392
rect 22152 7352 22158 7364
rect 22189 7361 22201 7364
rect 22235 7361 22247 7395
rect 22189 7355 22247 7361
rect 21324 7296 21956 7324
rect 21324 7284 21330 7296
rect 18233 7259 18291 7265
rect 14108 7228 14228 7256
rect 14200 7200 14228 7228
rect 18233 7225 18245 7259
rect 18279 7225 18291 7259
rect 21453 7259 21511 7265
rect 18233 7219 18291 7225
rect 20180 7228 21128 7256
rect 14182 7188 14188 7200
rect 12728 7160 14188 7188
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 15286 7148 15292 7200
rect 15344 7188 15350 7200
rect 15562 7188 15568 7200
rect 15344 7160 15568 7188
rect 15344 7148 15350 7160
rect 15562 7148 15568 7160
rect 15620 7188 15626 7200
rect 18248 7188 18276 7219
rect 15620 7160 18276 7188
rect 15620 7148 15626 7160
rect 18414 7148 18420 7200
rect 18472 7188 18478 7200
rect 20180 7188 20208 7228
rect 21100 7200 21128 7228
rect 21453 7225 21465 7259
rect 21499 7256 21511 7259
rect 22296 7256 22324 7432
rect 22373 7395 22431 7401
rect 22373 7361 22385 7395
rect 22419 7392 22431 7395
rect 22419 7364 22600 7392
rect 22419 7361 22431 7364
rect 22373 7355 22431 7361
rect 22572 7265 22600 7364
rect 22738 7352 22744 7404
rect 22796 7352 22802 7404
rect 23198 7352 23204 7404
rect 23256 7352 23262 7404
rect 23474 7352 23480 7404
rect 23532 7352 23538 7404
rect 23566 7352 23572 7404
rect 23624 7352 23630 7404
rect 23750 7352 23756 7404
rect 23808 7392 23814 7404
rect 24136 7401 24164 7432
rect 23845 7395 23903 7401
rect 23845 7392 23857 7395
rect 23808 7364 23857 7392
rect 23808 7352 23814 7364
rect 23845 7361 23857 7364
rect 23891 7361 23903 7395
rect 23845 7355 23903 7361
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 24121 7395 24179 7401
rect 24121 7361 24133 7395
rect 24167 7361 24179 7395
rect 24121 7355 24179 7361
rect 23584 7324 23612 7352
rect 23952 7324 23980 7355
rect 24210 7352 24216 7404
rect 24268 7352 24274 7404
rect 23584 7296 23980 7324
rect 21499 7228 22324 7256
rect 22557 7259 22615 7265
rect 21499 7225 21511 7228
rect 21453 7219 21511 7225
rect 22557 7225 22569 7259
rect 22603 7225 22615 7259
rect 22557 7219 22615 7225
rect 18472 7160 20208 7188
rect 20717 7191 20775 7197
rect 18472 7148 18478 7160
rect 20717 7157 20729 7191
rect 20763 7188 20775 7191
rect 20806 7188 20812 7200
rect 20763 7160 20812 7188
rect 20763 7157 20775 7160
rect 20717 7151 20775 7157
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 21082 7148 21088 7200
rect 21140 7148 21146 7200
rect 22005 7191 22063 7197
rect 22005 7157 22017 7191
rect 22051 7188 22063 7191
rect 22186 7188 22192 7200
rect 22051 7160 22192 7188
rect 22051 7157 22063 7160
rect 22005 7151 22063 7157
rect 22186 7148 22192 7160
rect 22244 7148 22250 7200
rect 22278 7148 22284 7200
rect 22336 7148 22342 7200
rect 23014 7148 23020 7200
rect 23072 7148 23078 7200
rect 1104 7098 24840 7120
rect 1104 7046 3917 7098
rect 3969 7046 3981 7098
rect 4033 7046 4045 7098
rect 4097 7046 4109 7098
rect 4161 7046 4173 7098
rect 4225 7046 9851 7098
rect 9903 7046 9915 7098
rect 9967 7046 9979 7098
rect 10031 7046 10043 7098
rect 10095 7046 10107 7098
rect 10159 7046 15785 7098
rect 15837 7046 15849 7098
rect 15901 7046 15913 7098
rect 15965 7046 15977 7098
rect 16029 7046 16041 7098
rect 16093 7046 21719 7098
rect 21771 7046 21783 7098
rect 21835 7046 21847 7098
rect 21899 7046 21911 7098
rect 21963 7046 21975 7098
rect 22027 7046 24840 7098
rect 1104 7024 24840 7046
rect 1762 6944 1768 6996
rect 1820 6944 1826 6996
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 4706 6984 4712 6996
rect 2004 6956 4712 6984
rect 2004 6944 2010 6956
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 11146 6984 11152 6996
rect 4816 6956 11152 6984
rect 2958 6876 2964 6928
rect 3016 6916 3022 6928
rect 4816 6916 4844 6956
rect 11146 6944 11152 6956
rect 11204 6944 11210 6996
rect 17236 6956 17908 6984
rect 3016 6888 4844 6916
rect 3016 6876 3022 6888
rect 6086 6876 6092 6928
rect 6144 6916 6150 6928
rect 6638 6916 6644 6928
rect 6144 6888 6644 6916
rect 6144 6876 6150 6888
rect 6638 6876 6644 6888
rect 6696 6916 6702 6928
rect 6696 6888 6960 6916
rect 6696 6876 6702 6888
rect 1210 6808 1216 6860
rect 1268 6848 1274 6860
rect 2501 6851 2559 6857
rect 2501 6848 2513 6851
rect 1268 6820 2513 6848
rect 1268 6808 1274 6820
rect 2501 6817 2513 6820
rect 2547 6817 2559 6851
rect 2501 6811 2559 6817
rect 3050 6808 3056 6860
rect 3108 6808 3114 6860
rect 3326 6808 3332 6860
rect 3384 6848 3390 6860
rect 4157 6851 4215 6857
rect 4157 6848 4169 6851
rect 3384 6820 4169 6848
rect 3384 6808 3390 6820
rect 4157 6817 4169 6820
rect 4203 6817 4215 6851
rect 4157 6811 4215 6817
rect 4540 6820 4936 6848
rect 2130 6740 2136 6792
rect 2188 6780 2194 6792
rect 3421 6783 3479 6789
rect 2188 6752 2544 6780
rect 2188 6740 2194 6752
rect 2516 6724 2544 6752
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 1946 6712 1952 6724
rect 1719 6684 1952 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 1946 6672 1952 6684
rect 2004 6672 2010 6724
rect 2222 6672 2228 6724
rect 2280 6672 2286 6724
rect 2498 6672 2504 6724
rect 2556 6672 2562 6724
rect 2774 6672 2780 6724
rect 2832 6672 2838 6724
rect 3436 6712 3464 6743
rect 3694 6740 3700 6792
rect 3752 6780 3758 6792
rect 4540 6789 4568 6820
rect 3881 6783 3939 6789
rect 3881 6780 3893 6783
rect 3752 6752 3893 6780
rect 3752 6740 3758 6752
rect 3881 6749 3893 6752
rect 3927 6749 3939 6783
rect 3881 6743 3939 6749
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6749 4859 6783
rect 4908 6780 4936 6820
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 6362 6848 6368 6860
rect 5040 6820 6368 6848
rect 5040 6808 5046 6820
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 6932 6848 6960 6888
rect 11054 6876 11060 6928
rect 11112 6876 11118 6928
rect 12526 6916 12532 6928
rect 12176 6888 12532 6916
rect 6932 6820 7236 6848
rect 6638 6780 6644 6792
rect 4908 6752 6644 6780
rect 4801 6743 4859 6749
rect 4816 6712 4844 6743
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 7208 6789 7236 6820
rect 8018 6808 8024 6860
rect 8076 6848 8082 6860
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 8076 6820 8953 6848
rect 8076 6808 8082 6820
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 10410 6808 10416 6860
rect 10468 6848 10474 6860
rect 10689 6851 10747 6857
rect 10689 6848 10701 6851
rect 10468 6820 10701 6848
rect 10468 6808 10474 6820
rect 10689 6817 10701 6820
rect 10735 6817 10747 6851
rect 11072 6848 11100 6876
rect 11149 6851 11207 6857
rect 11149 6848 11161 6851
rect 11072 6820 11161 6848
rect 10689 6811 10747 6817
rect 11149 6817 11161 6820
rect 11195 6817 11207 6851
rect 11149 6811 11207 6817
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6848 11483 6851
rect 12176 6848 12204 6888
rect 12526 6876 12532 6888
rect 12584 6876 12590 6928
rect 17236 6857 17264 6956
rect 17880 6916 17908 6956
rect 18230 6944 18236 6996
rect 18288 6984 18294 6996
rect 18693 6987 18751 6993
rect 18693 6984 18705 6987
rect 18288 6956 18705 6984
rect 18288 6944 18294 6956
rect 18693 6953 18705 6956
rect 18739 6953 18751 6987
rect 18693 6947 18751 6953
rect 18782 6944 18788 6996
rect 18840 6984 18846 6996
rect 18969 6987 19027 6993
rect 18969 6984 18981 6987
rect 18840 6956 18981 6984
rect 18840 6944 18846 6956
rect 18969 6953 18981 6956
rect 19015 6953 19027 6987
rect 19610 6984 19616 6996
rect 18969 6947 19027 6953
rect 19168 6956 19616 6984
rect 19168 6916 19196 6956
rect 19610 6944 19616 6956
rect 19668 6944 19674 6996
rect 20162 6944 20168 6996
rect 20220 6984 20226 6996
rect 20257 6987 20315 6993
rect 20257 6984 20269 6987
rect 20220 6956 20269 6984
rect 20220 6944 20226 6956
rect 20257 6953 20269 6956
rect 20303 6953 20315 6987
rect 20257 6947 20315 6953
rect 21266 6944 21272 6996
rect 21324 6944 21330 6996
rect 21450 6944 21456 6996
rect 21508 6944 21514 6996
rect 21910 6944 21916 6996
rect 21968 6984 21974 6996
rect 22462 6984 22468 6996
rect 21968 6956 22468 6984
rect 21968 6944 21974 6956
rect 22462 6944 22468 6956
rect 22520 6944 22526 6996
rect 22738 6944 22744 6996
rect 22796 6984 22802 6996
rect 22925 6987 22983 6993
rect 22925 6984 22937 6987
rect 22796 6956 22937 6984
rect 22796 6944 22802 6956
rect 22925 6953 22937 6956
rect 22971 6953 22983 6987
rect 22925 6947 22983 6953
rect 17880 6888 19196 6916
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 11471 6820 12204 6848
rect 12268 6820 12633 6848
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6780 7251 6783
rect 7374 6780 7380 6792
rect 7239 6752 7380 6780
rect 7239 6749 7251 6752
rect 7193 6743 7251 6749
rect 7374 6740 7380 6752
rect 7432 6740 7438 6792
rect 7467 6783 7525 6789
rect 7467 6749 7479 6783
rect 7513 6780 7525 6783
rect 7558 6780 7564 6792
rect 7513 6752 7564 6780
rect 7513 6749 7525 6752
rect 7467 6743 7525 6749
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 9214 6759 9444 6780
rect 9199 6753 9444 6759
rect 8570 6712 8576 6724
rect 3436 6684 4752 6712
rect 4816 6684 8576 6712
rect 2038 6604 2044 6656
rect 2096 6644 2102 6656
rect 3237 6647 3295 6653
rect 3237 6644 3249 6647
rect 2096 6616 3249 6644
rect 2096 6604 2102 6616
rect 3237 6613 3249 6616
rect 3283 6613 3295 6647
rect 3237 6607 3295 6613
rect 3326 6604 3332 6656
rect 3384 6644 3390 6656
rect 3694 6644 3700 6656
rect 3384 6616 3700 6644
rect 3384 6604 3390 6616
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 4338 6604 4344 6656
rect 4396 6604 4402 6656
rect 4614 6604 4620 6656
rect 4672 6604 4678 6656
rect 4724 6644 4752 6684
rect 8570 6672 8576 6684
rect 8628 6672 8634 6724
rect 9199 6719 9211 6753
rect 9245 6752 9444 6753
rect 9245 6719 9257 6752
rect 9416 6724 9444 6752
rect 10502 6740 10508 6792
rect 10560 6740 10566 6792
rect 11514 6740 11520 6792
rect 11572 6789 11578 6792
rect 11572 6783 11600 6789
rect 11588 6749 11600 6783
rect 11572 6743 11600 6749
rect 11572 6740 11578 6743
rect 11698 6740 11704 6792
rect 11756 6740 11762 6792
rect 9199 6713 9257 6719
rect 9398 6672 9404 6724
rect 9456 6672 9462 6724
rect 12268 6656 12296 6820
rect 12621 6817 12633 6820
rect 12667 6817 12679 6851
rect 12621 6811 12679 6817
rect 17221 6851 17279 6857
rect 17221 6817 17233 6851
rect 17267 6817 17279 6851
rect 17221 6811 17279 6817
rect 17880 6792 17908 6888
rect 12342 6740 12348 6792
rect 12400 6780 12406 6792
rect 12863 6783 12921 6789
rect 12863 6780 12875 6783
rect 12400 6752 12875 6780
rect 12400 6740 12406 6752
rect 12863 6749 12875 6752
rect 12909 6749 12921 6783
rect 12863 6743 12921 6749
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 15654 6780 15660 6792
rect 15344 6752 15660 6780
rect 15344 6740 15350 6752
rect 15654 6740 15660 6752
rect 15712 6780 15718 6792
rect 17463 6783 17521 6789
rect 17463 6780 17475 6783
rect 15712 6752 17475 6780
rect 15712 6740 15718 6752
rect 17463 6749 17475 6752
rect 17509 6749 17521 6783
rect 17463 6743 17521 6749
rect 17862 6740 17868 6792
rect 17920 6740 17926 6792
rect 18598 6740 18604 6792
rect 18656 6740 18662 6792
rect 18877 6783 18935 6789
rect 18877 6749 18889 6783
rect 18923 6749 18935 6783
rect 18877 6743 18935 6749
rect 19061 6783 19119 6789
rect 19061 6749 19073 6783
rect 19107 6780 19119 6783
rect 19150 6780 19156 6792
rect 19107 6752 19156 6780
rect 19107 6749 19119 6752
rect 19061 6743 19119 6749
rect 12526 6672 12532 6724
rect 12584 6712 12590 6724
rect 13446 6712 13452 6724
rect 12584 6684 13452 6712
rect 12584 6672 12590 6684
rect 13446 6672 13452 6684
rect 13504 6712 13510 6724
rect 18892 6712 18920 6743
rect 19150 6740 19156 6752
rect 19208 6740 19214 6792
rect 19245 6783 19303 6789
rect 19245 6749 19257 6783
rect 19291 6749 19303 6783
rect 19245 6743 19303 6749
rect 13504 6684 17540 6712
rect 13504 6672 13510 6684
rect 17512 6656 17540 6684
rect 18340 6684 18920 6712
rect 19260 6712 19288 6743
rect 19426 6740 19432 6792
rect 19484 6780 19490 6792
rect 19519 6783 19577 6789
rect 19519 6780 19531 6783
rect 19484 6752 19531 6780
rect 19484 6740 19490 6752
rect 19519 6749 19531 6752
rect 19565 6749 19577 6783
rect 19519 6743 19577 6749
rect 19978 6740 19984 6792
rect 20036 6780 20042 6792
rect 21468 6789 21496 6944
rect 24029 6919 24087 6925
rect 24029 6885 24041 6919
rect 24075 6916 24087 6919
rect 24486 6916 24492 6928
rect 24075 6888 24492 6916
rect 24075 6885 24087 6888
rect 24029 6879 24087 6885
rect 24486 6876 24492 6888
rect 24544 6876 24550 6928
rect 21542 6808 21548 6860
rect 21600 6808 21606 6860
rect 21453 6783 21511 6789
rect 20036 6752 21404 6780
rect 20036 6740 20042 6752
rect 20714 6712 20720 6724
rect 19260 6684 20720 6712
rect 18340 6656 18368 6684
rect 20714 6672 20720 6684
rect 20772 6672 20778 6724
rect 21376 6712 21404 6752
rect 21453 6749 21465 6783
rect 21499 6780 21511 6783
rect 21801 6783 21859 6789
rect 21801 6780 21813 6783
rect 21499 6752 21813 6780
rect 21499 6749 21511 6752
rect 21453 6743 21511 6749
rect 21801 6749 21813 6752
rect 21847 6749 21859 6783
rect 21801 6743 21859 6749
rect 22738 6740 22744 6792
rect 22796 6780 22802 6792
rect 23109 6783 23167 6789
rect 23109 6780 23121 6783
rect 22796 6752 23121 6780
rect 22796 6740 22802 6752
rect 23109 6749 23121 6752
rect 23155 6749 23167 6783
rect 23109 6743 23167 6749
rect 23477 6783 23535 6789
rect 23477 6749 23489 6783
rect 23523 6749 23535 6783
rect 23477 6743 23535 6749
rect 21634 6712 21640 6724
rect 21376 6684 21640 6712
rect 21634 6672 21640 6684
rect 21692 6672 21698 6724
rect 7374 6644 7380 6656
rect 4724 6616 7380 6644
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 8018 6644 8024 6656
rect 7524 6616 8024 6644
rect 7524 6604 7530 6616
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 8202 6604 8208 6656
rect 8260 6604 8266 6656
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 9953 6647 10011 6653
rect 9953 6644 9965 6647
rect 9088 6616 9965 6644
rect 9088 6604 9094 6616
rect 9953 6613 9965 6616
rect 9999 6613 10011 6647
rect 9953 6607 10011 6613
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 12250 6644 12256 6656
rect 11296 6616 12256 6644
rect 11296 6604 11302 6616
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12342 6604 12348 6656
rect 12400 6604 12406 6656
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 13633 6647 13691 6653
rect 13633 6644 13645 6647
rect 12492 6616 13645 6644
rect 12492 6604 12498 6616
rect 13633 6613 13645 6616
rect 13679 6613 13691 6647
rect 13633 6607 13691 6613
rect 17494 6604 17500 6656
rect 17552 6604 17558 6656
rect 18233 6647 18291 6653
rect 18233 6613 18245 6647
rect 18279 6644 18291 6647
rect 18322 6644 18328 6656
rect 18279 6616 18328 6644
rect 18279 6613 18291 6616
rect 18233 6607 18291 6613
rect 18322 6604 18328 6616
rect 18380 6604 18386 6656
rect 21358 6604 21364 6656
rect 21416 6644 21422 6656
rect 23492 6644 23520 6743
rect 23566 6740 23572 6792
rect 23624 6780 23630 6792
rect 23937 6783 23995 6789
rect 23937 6780 23949 6783
rect 23624 6752 23949 6780
rect 23624 6740 23630 6752
rect 23937 6749 23949 6752
rect 23983 6749 23995 6783
rect 23937 6743 23995 6749
rect 21416 6616 23520 6644
rect 21416 6604 21422 6616
rect 1104 6554 25000 6576
rect 1104 6502 6884 6554
rect 6936 6502 6948 6554
rect 7000 6502 7012 6554
rect 7064 6502 7076 6554
rect 7128 6502 7140 6554
rect 7192 6502 12818 6554
rect 12870 6502 12882 6554
rect 12934 6502 12946 6554
rect 12998 6502 13010 6554
rect 13062 6502 13074 6554
rect 13126 6502 18752 6554
rect 18804 6502 18816 6554
rect 18868 6502 18880 6554
rect 18932 6502 18944 6554
rect 18996 6502 19008 6554
rect 19060 6502 24686 6554
rect 24738 6502 24750 6554
rect 24802 6502 24814 6554
rect 24866 6502 24878 6554
rect 24930 6502 24942 6554
rect 24994 6502 25000 6554
rect 1104 6480 25000 6502
rect 1578 6400 1584 6452
rect 1636 6400 1642 6452
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 3421 6443 3479 6449
rect 3421 6440 3433 6443
rect 2832 6412 3433 6440
rect 2832 6400 2838 6412
rect 3421 6409 3433 6412
rect 3467 6409 3479 6443
rect 4338 6440 4344 6452
rect 3421 6403 3479 6409
rect 3528 6412 4344 6440
rect 1489 6375 1547 6381
rect 1489 6341 1501 6375
rect 1535 6372 1547 6375
rect 3528 6372 3556 6412
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 5350 6400 5356 6452
rect 5408 6440 5414 6452
rect 8938 6440 8944 6452
rect 5408 6412 8944 6440
rect 5408 6400 5414 6412
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9674 6400 9680 6452
rect 9732 6400 9738 6452
rect 10502 6400 10508 6452
rect 10560 6400 10566 6452
rect 15562 6440 15568 6452
rect 10980 6412 15568 6440
rect 1535 6344 3556 6372
rect 1535 6341 1547 6344
rect 1489 6335 1547 6341
rect 1302 6264 1308 6316
rect 1360 6264 1366 6316
rect 1854 6264 1860 6316
rect 1912 6304 1918 6316
rect 2315 6307 2373 6313
rect 2315 6304 2327 6307
rect 1912 6276 2327 6304
rect 1912 6264 1918 6276
rect 2315 6273 2327 6276
rect 2361 6273 2373 6307
rect 2315 6267 2373 6273
rect 3602 6264 3608 6316
rect 3660 6264 3666 6316
rect 3694 6264 3700 6316
rect 3752 6264 3758 6316
rect 4614 6264 4620 6316
rect 4672 6264 4678 6316
rect 4890 6264 4896 6316
rect 4948 6264 4954 6316
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6304 5595 6307
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5583 6276 5825 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 8202 6264 8208 6316
rect 8260 6264 8266 6316
rect 8846 6264 8852 6316
rect 8904 6313 8910 6316
rect 8904 6307 8953 6313
rect 8904 6273 8907 6307
rect 8941 6273 8953 6307
rect 8904 6267 8953 6273
rect 8904 6264 8910 6267
rect 9030 6264 9036 6316
rect 9088 6264 9094 6316
rect 10410 6264 10416 6316
rect 10468 6264 10474 6316
rect 10520 6304 10548 6400
rect 10980 6304 11008 6412
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 17313 6443 17371 6449
rect 17313 6409 17325 6443
rect 17359 6440 17371 6443
rect 18598 6440 18604 6452
rect 17359 6412 18604 6440
rect 17359 6409 17371 6412
rect 17313 6403 17371 6409
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 19061 6443 19119 6449
rect 19061 6409 19073 6443
rect 19107 6440 19119 6443
rect 19150 6440 19156 6452
rect 19107 6412 19156 6440
rect 19107 6409 19119 6412
rect 19061 6403 19119 6409
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 20622 6400 20628 6452
rect 20680 6400 20686 6452
rect 20717 6443 20775 6449
rect 20717 6409 20729 6443
rect 20763 6440 20775 6443
rect 21358 6440 21364 6452
rect 20763 6412 21364 6440
rect 20763 6409 20775 6412
rect 20717 6403 20775 6409
rect 21358 6400 21364 6412
rect 21416 6400 21422 6452
rect 21450 6400 21456 6452
rect 21508 6440 21514 6452
rect 23014 6440 23020 6452
rect 21508 6412 23020 6440
rect 21508 6400 21514 6412
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 24489 6443 24547 6449
rect 24489 6409 24501 6443
rect 24535 6409 24547 6443
rect 24489 6403 24547 6409
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 15286 6372 15292 6384
rect 11112 6344 11652 6372
rect 11112 6332 11118 6344
rect 11624 6316 11652 6344
rect 15028 6344 15292 6372
rect 15028 6343 15056 6344
rect 14995 6337 15056 6343
rect 11517 6307 11575 6313
rect 11517 6304 11529 6307
rect 10520 6276 11529 6304
rect 11517 6273 11529 6276
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 11606 6264 11612 6316
rect 11664 6304 11670 6316
rect 11664 6276 11910 6304
rect 11664 6264 11670 6276
rect 1320 6236 1348 6264
rect 2041 6239 2099 6245
rect 2041 6236 2053 6239
rect 1320 6208 2053 6236
rect 1872 6180 1900 6208
rect 2041 6205 2053 6208
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 3510 6196 3516 6248
rect 3568 6236 3574 6248
rect 3881 6239 3939 6245
rect 3881 6236 3893 6239
rect 3568 6208 3893 6236
rect 3568 6196 3574 6208
rect 3881 6205 3893 6208
rect 3927 6205 3939 6239
rect 3881 6199 3939 6205
rect 4430 6196 4436 6248
rect 4488 6236 4494 6248
rect 4755 6239 4813 6245
rect 4755 6236 4767 6239
rect 4488 6208 4767 6236
rect 4488 6196 4494 6208
rect 4755 6205 4767 6208
rect 4801 6236 4813 6239
rect 5442 6236 5448 6248
rect 4801 6208 5448 6236
rect 4801 6205 4813 6208
rect 4755 6199 4813 6205
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 7834 6196 7840 6248
rect 7892 6196 7898 6248
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6205 8079 6239
rect 8220 6236 8248 6264
rect 8481 6239 8539 6245
rect 8481 6236 8493 6239
rect 8220 6208 8493 6236
rect 8021 6199 8079 6205
rect 8481 6205 8493 6208
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 8757 6239 8815 6245
rect 8757 6205 8769 6239
rect 8803 6236 8815 6239
rect 10428 6236 10456 6264
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 8803 6208 9674 6236
rect 10428 6208 11713 6236
rect 8803 6205 8815 6208
rect 8757 6199 8815 6205
rect 1854 6128 1860 6180
rect 1912 6128 1918 6180
rect 2884 6140 4200 6168
rect 2406 6060 2412 6112
rect 2464 6100 2470 6112
rect 2884 6100 2912 6140
rect 2464 6072 2912 6100
rect 2464 6060 2470 6072
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 3053 6103 3111 6109
rect 3053 6100 3065 6103
rect 3016 6072 3065 6100
rect 3016 6060 3022 6072
rect 3053 6069 3065 6072
rect 3099 6069 3111 6103
rect 4172 6100 4200 6140
rect 4338 6128 4344 6180
rect 4396 6128 4402 6180
rect 8036 6168 8064 6199
rect 8294 6168 8300 6180
rect 6104 6140 8300 6168
rect 6104 6112 6132 6140
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 9646 6168 9674 6208
rect 11701 6205 11713 6208
rect 11747 6236 11759 6239
rect 11790 6236 11796 6248
rect 11747 6208 11796 6236
rect 11747 6205 11759 6208
rect 11701 6199 11759 6205
rect 11790 6196 11796 6208
rect 11848 6196 11854 6248
rect 11882 6236 11910 6276
rect 12434 6264 12440 6316
rect 12492 6264 12498 6316
rect 14995 6303 15007 6337
rect 15041 6306 15056 6337
rect 15286 6332 15292 6344
rect 15344 6332 15350 6384
rect 19334 6372 19340 6384
rect 17604 6344 19340 6372
rect 17604 6313 17632 6344
rect 19334 6332 19340 6344
rect 19392 6332 19398 6384
rect 20640 6372 20668 6400
rect 24504 6372 24532 6403
rect 20640 6344 21036 6372
rect 17497 6307 17555 6313
rect 15041 6303 15053 6306
rect 14995 6297 15053 6303
rect 17497 6273 17509 6307
rect 17543 6273 17555 6307
rect 17497 6267 17555 6273
rect 17589 6307 17647 6313
rect 17589 6273 17601 6307
rect 17635 6273 17647 6307
rect 17856 6307 17914 6313
rect 17856 6304 17868 6307
rect 17589 6267 17647 6273
rect 17696 6276 17868 6304
rect 12554 6239 12612 6245
rect 12554 6236 12566 6239
rect 11882 6208 12566 6236
rect 12554 6205 12566 6208
rect 12600 6205 12612 6239
rect 12554 6199 12612 6205
rect 12710 6196 12716 6248
rect 12768 6196 12774 6248
rect 14737 6239 14795 6245
rect 14737 6205 14749 6239
rect 14783 6205 14795 6239
rect 14737 6199 14795 6205
rect 11054 6168 11060 6180
rect 9646 6140 11060 6168
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 11146 6128 11152 6180
rect 11204 6168 11210 6180
rect 12161 6171 12219 6177
rect 12161 6168 12173 6171
rect 11204 6140 12173 6168
rect 11204 6128 11210 6140
rect 12161 6137 12173 6140
rect 12207 6137 12219 6171
rect 12161 6131 12219 6137
rect 5629 6103 5687 6109
rect 5629 6100 5641 6103
rect 4172 6072 5641 6100
rect 3053 6063 3111 6069
rect 5629 6069 5641 6072
rect 5675 6069 5687 6103
rect 5629 6063 5687 6069
rect 6086 6060 6092 6112
rect 6144 6060 6150 6112
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 6362 6100 6368 6112
rect 6236 6072 6368 6100
rect 6236 6060 6242 6072
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 13357 6103 13415 6109
rect 13357 6100 13369 6103
rect 6696 6072 13369 6100
rect 6696 6060 6702 6072
rect 13357 6069 13369 6072
rect 13403 6069 13415 6103
rect 13357 6063 13415 6069
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14752 6100 14780 6199
rect 17218 6196 17224 6248
rect 17276 6196 17282 6248
rect 17512 6236 17540 6267
rect 17696 6236 17724 6276
rect 17856 6273 17868 6276
rect 17902 6304 17914 6307
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 17902 6276 18920 6304
rect 17902 6273 17914 6276
rect 17856 6267 17914 6273
rect 17512 6208 17724 6236
rect 16114 6168 16120 6180
rect 15394 6140 16120 6168
rect 15394 6100 15422 6140
rect 16114 6128 16120 6140
rect 16172 6168 16178 6180
rect 17236 6168 17264 6196
rect 16172 6140 17264 6168
rect 16172 6128 16178 6140
rect 13872 6072 15422 6100
rect 13872 6060 13878 6072
rect 15654 6060 15660 6112
rect 15712 6100 15718 6112
rect 15749 6103 15807 6109
rect 15749 6100 15761 6103
rect 15712 6072 15761 6100
rect 15712 6060 15718 6072
rect 15749 6069 15761 6072
rect 15795 6069 15807 6103
rect 15749 6063 15807 6069
rect 16482 6060 16488 6112
rect 16540 6100 16546 6112
rect 17494 6100 17500 6112
rect 16540 6072 17500 6100
rect 16540 6060 16546 6072
rect 17494 6060 17500 6072
rect 17552 6060 17558 6112
rect 18892 6100 18920 6276
rect 18984 6276 19257 6304
rect 18984 6177 19012 6276
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 20622 6264 20628 6316
rect 20680 6264 20686 6316
rect 18969 6171 19027 6177
rect 18969 6137 18981 6171
rect 19015 6137 19027 6171
rect 18969 6131 19027 6137
rect 19058 6128 19064 6180
rect 19116 6168 19122 6180
rect 20901 6171 20959 6177
rect 20901 6168 20913 6171
rect 19116 6140 20913 6168
rect 19116 6128 19122 6140
rect 20901 6137 20913 6140
rect 20947 6137 20959 6171
rect 21008 6168 21036 6344
rect 21100 6344 24532 6372
rect 21100 6313 21128 6344
rect 21085 6307 21143 6313
rect 21085 6273 21097 6307
rect 21131 6273 21143 6307
rect 21085 6267 21143 6273
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6304 21235 6307
rect 21266 6304 21272 6316
rect 21223 6276 21272 6304
rect 21223 6273 21235 6276
rect 21177 6267 21235 6273
rect 21266 6264 21272 6276
rect 21324 6264 21330 6316
rect 21358 6264 21364 6316
rect 21416 6304 21422 6316
rect 21453 6307 21511 6313
rect 21453 6304 21465 6307
rect 21416 6276 21465 6304
rect 21416 6264 21422 6276
rect 21453 6273 21465 6276
rect 21499 6273 21511 6307
rect 21453 6267 21511 6273
rect 22005 6307 22063 6313
rect 22005 6273 22017 6307
rect 22051 6304 22063 6307
rect 22094 6304 22100 6316
rect 22051 6276 22100 6304
rect 22051 6273 22063 6276
rect 22005 6267 22063 6273
rect 22094 6264 22100 6276
rect 22152 6264 22158 6316
rect 22186 6264 22192 6316
rect 22244 6264 22250 6316
rect 22278 6264 22284 6316
rect 22336 6304 22342 6316
rect 22649 6307 22707 6313
rect 22649 6304 22661 6307
rect 22336 6276 22661 6304
rect 22336 6264 22342 6276
rect 22649 6273 22661 6276
rect 22695 6273 22707 6307
rect 22649 6267 22707 6273
rect 23014 6264 23020 6316
rect 23072 6304 23078 6316
rect 23365 6307 23423 6313
rect 23365 6304 23377 6307
rect 23072 6276 23377 6304
rect 23072 6264 23078 6276
rect 23365 6273 23377 6276
rect 23411 6273 23423 6307
rect 23365 6267 23423 6273
rect 21542 6196 21548 6248
rect 21600 6236 21606 6248
rect 23109 6239 23167 6245
rect 23109 6236 23121 6239
rect 21600 6208 23121 6236
rect 21600 6196 21606 6208
rect 23109 6205 23121 6208
rect 23155 6205 23167 6239
rect 23109 6199 23167 6205
rect 21637 6171 21695 6177
rect 21637 6168 21649 6171
rect 21008 6140 21649 6168
rect 20901 6131 20959 6137
rect 21637 6137 21649 6140
rect 21683 6137 21695 6171
rect 21637 6131 21695 6137
rect 21910 6128 21916 6180
rect 21968 6168 21974 6180
rect 22186 6168 22192 6180
rect 21968 6140 22192 6168
rect 21968 6128 21974 6140
rect 22186 6128 22192 6140
rect 22244 6128 22250 6180
rect 22646 6128 22652 6180
rect 22704 6128 22710 6180
rect 20714 6100 20720 6112
rect 18892 6072 20720 6100
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 21174 6060 21180 6112
rect 21232 6100 21238 6112
rect 21361 6103 21419 6109
rect 21361 6100 21373 6103
rect 21232 6072 21373 6100
rect 21232 6060 21238 6072
rect 21361 6069 21373 6072
rect 21407 6069 21419 6103
rect 21361 6063 21419 6069
rect 21542 6060 21548 6112
rect 21600 6100 21606 6112
rect 23750 6100 23756 6112
rect 21600 6072 23756 6100
rect 21600 6060 21606 6072
rect 23750 6060 23756 6072
rect 23808 6060 23814 6112
rect 1104 6010 24840 6032
rect 1104 5958 3917 6010
rect 3969 5958 3981 6010
rect 4033 5958 4045 6010
rect 4097 5958 4109 6010
rect 4161 5958 4173 6010
rect 4225 5958 9851 6010
rect 9903 5958 9915 6010
rect 9967 5958 9979 6010
rect 10031 5958 10043 6010
rect 10095 5958 10107 6010
rect 10159 5958 15785 6010
rect 15837 5958 15849 6010
rect 15901 5958 15913 6010
rect 15965 5958 15977 6010
rect 16029 5958 16041 6010
rect 16093 5958 21719 6010
rect 21771 5958 21783 6010
rect 21835 5958 21847 6010
rect 21899 5958 21911 6010
rect 21963 5958 21975 6010
rect 22027 5958 24840 6010
rect 1104 5936 24840 5958
rect 1489 5899 1547 5905
rect 1489 5865 1501 5899
rect 1535 5896 1547 5899
rect 2222 5896 2228 5908
rect 1535 5868 2228 5896
rect 1535 5865 1547 5868
rect 1489 5859 1547 5865
rect 2222 5856 2228 5868
rect 2280 5856 2286 5908
rect 2774 5896 2780 5908
rect 2516 5868 2780 5896
rect 1762 5720 1768 5772
rect 1820 5720 1826 5772
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5760 2007 5763
rect 2314 5760 2320 5772
rect 1995 5732 2320 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 2314 5720 2320 5732
rect 2372 5720 2378 5772
rect 2406 5720 2412 5772
rect 2464 5720 2470 5772
rect 2516 5760 2544 5868
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3418 5896 3424 5908
rect 2924 5868 3424 5896
rect 2924 5856 2930 5868
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 3602 5856 3608 5908
rect 3660 5856 3666 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5077 5899 5135 5905
rect 5077 5896 5089 5899
rect 4948 5868 5089 5896
rect 4948 5856 4954 5868
rect 5077 5865 5089 5868
rect 5123 5865 5135 5899
rect 6086 5896 6092 5908
rect 5077 5859 5135 5865
rect 5460 5868 6092 5896
rect 2866 5769 2872 5772
rect 2685 5763 2743 5769
rect 2685 5760 2697 5763
rect 2516 5732 2697 5760
rect 2685 5729 2697 5732
rect 2731 5729 2743 5763
rect 2685 5723 2743 5729
rect 2823 5763 2872 5769
rect 2823 5729 2835 5763
rect 2869 5729 2872 5763
rect 2823 5723 2872 5729
rect 2866 5720 2872 5723
rect 2924 5720 2930 5772
rect 2958 5720 2964 5772
rect 3016 5720 3022 5772
rect 1670 5652 1676 5704
rect 1728 5652 1734 5704
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3752 5664 3985 5692
rect 3752 5652 3758 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4062 5652 4068 5704
rect 4120 5652 4126 5704
rect 4339 5695 4397 5701
rect 4339 5661 4351 5695
rect 4385 5692 4397 5695
rect 5350 5692 5356 5704
rect 4385 5664 5356 5692
rect 4385 5661 4397 5664
rect 4339 5655 4397 5661
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 3510 5584 3516 5636
rect 3568 5624 3574 5636
rect 5460 5624 5488 5868
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6196 5868 7144 5896
rect 5626 5788 5632 5840
rect 5684 5828 5690 5840
rect 6196 5828 6224 5868
rect 5684 5800 6224 5828
rect 7116 5828 7144 5868
rect 7374 5856 7380 5908
rect 7432 5856 7438 5908
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 8846 5896 8852 5908
rect 7892 5868 8852 5896
rect 7892 5856 7898 5868
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 11238 5896 11244 5908
rect 8956 5868 11244 5896
rect 8956 5828 8984 5868
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 11885 5899 11943 5905
rect 11885 5865 11897 5899
rect 11931 5896 11943 5899
rect 12710 5896 12716 5908
rect 11931 5868 12716 5896
rect 11931 5865 11943 5868
rect 11885 5859 11943 5865
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 13265 5899 13323 5905
rect 13265 5865 13277 5899
rect 13311 5896 13323 5899
rect 13906 5896 13912 5908
rect 13311 5868 13912 5896
rect 13311 5865 13323 5868
rect 13265 5859 13323 5865
rect 13906 5856 13912 5868
rect 13964 5856 13970 5908
rect 15654 5856 15660 5908
rect 15712 5856 15718 5908
rect 15746 5856 15752 5908
rect 15804 5896 15810 5908
rect 16298 5896 16304 5908
rect 15804 5868 16304 5896
rect 15804 5856 15810 5868
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 18141 5899 18199 5905
rect 18141 5896 18153 5899
rect 17052 5868 18153 5896
rect 12066 5828 12072 5840
rect 7116 5800 8984 5828
rect 11532 5800 12072 5828
rect 5684 5788 5690 5800
rect 5736 5769 5764 5800
rect 5721 5763 5779 5769
rect 5721 5729 5733 5763
rect 5767 5729 5779 5763
rect 5721 5723 5779 5729
rect 6178 5720 6184 5772
rect 6236 5720 6242 5772
rect 6546 5720 6552 5772
rect 6604 5769 6610 5772
rect 6604 5763 6632 5769
rect 6620 5729 6632 5763
rect 6604 5723 6632 5729
rect 6733 5763 6791 5769
rect 6733 5729 6745 5763
rect 6779 5760 6791 5763
rect 7374 5760 7380 5772
rect 6779 5732 7380 5760
rect 6779 5729 6791 5732
rect 6733 5723 6791 5729
rect 6604 5720 6610 5723
rect 7374 5720 7380 5732
rect 7432 5720 7438 5772
rect 10870 5720 10876 5772
rect 10928 5720 10934 5772
rect 5534 5652 5540 5704
rect 5592 5652 5598 5704
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 8754 5692 8760 5704
rect 7300 5664 8760 5692
rect 3568 5596 5488 5624
rect 3568 5584 3574 5596
rect 2314 5516 2320 5568
rect 2372 5556 2378 5568
rect 3789 5559 3847 5565
rect 3789 5556 3801 5559
rect 2372 5528 3801 5556
rect 2372 5516 2378 5528
rect 3789 5525 3801 5528
rect 3835 5525 3847 5559
rect 3789 5519 3847 5525
rect 4522 5516 4528 5568
rect 4580 5556 4586 5568
rect 5166 5556 5172 5568
rect 4580 5528 5172 5556
rect 4580 5516 4586 5528
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 5552 5556 5580 5652
rect 7300 5556 7328 5664
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 9122 5652 9128 5704
rect 9180 5652 9186 5704
rect 9306 5652 9312 5704
rect 9364 5701 9370 5704
rect 9364 5695 9425 5701
rect 9364 5661 9379 5695
rect 9413 5692 9425 5695
rect 10226 5692 10232 5704
rect 9413 5664 10232 5692
rect 9413 5661 9425 5664
rect 9364 5655 9425 5661
rect 9364 5652 9370 5655
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 7558 5584 7564 5636
rect 7616 5624 7622 5636
rect 10502 5624 10508 5636
rect 7616 5596 9352 5624
rect 7616 5584 7622 5596
rect 5552 5528 7328 5556
rect 9324 5556 9352 5596
rect 9646 5596 10508 5624
rect 9646 5556 9674 5596
rect 10502 5584 10508 5596
rect 10560 5584 10566 5636
rect 9324 5528 9674 5556
rect 10134 5516 10140 5568
rect 10192 5516 10198 5568
rect 10226 5516 10232 5568
rect 10284 5556 10290 5568
rect 10888 5556 10916 5720
rect 11147 5695 11205 5701
rect 11147 5692 11159 5695
rect 11072 5664 11159 5692
rect 11072 5636 11100 5664
rect 11147 5661 11159 5664
rect 11193 5692 11205 5695
rect 11532 5692 11560 5800
rect 12066 5788 12072 5800
rect 12124 5788 12130 5840
rect 15672 5828 15700 5856
rect 15841 5831 15899 5837
rect 15841 5828 15853 5831
rect 15672 5800 15853 5828
rect 15841 5797 15853 5800
rect 15887 5797 15899 5831
rect 15841 5791 15899 5797
rect 12250 5760 12256 5772
rect 11624 5732 12256 5760
rect 11624 5704 11652 5732
rect 12250 5720 12256 5732
rect 12308 5720 12314 5772
rect 16298 5769 16304 5772
rect 16117 5763 16175 5769
rect 16117 5760 16129 5763
rect 15580 5732 16129 5760
rect 15580 5704 15608 5732
rect 16117 5729 16129 5732
rect 16163 5729 16175 5763
rect 16117 5723 16175 5729
rect 16255 5763 16304 5769
rect 16255 5729 16267 5763
rect 16301 5729 16304 5763
rect 16255 5723 16304 5729
rect 16298 5720 16304 5723
rect 16356 5720 16362 5772
rect 16393 5763 16451 5769
rect 16393 5729 16405 5763
rect 16439 5760 16451 5763
rect 17052 5760 17080 5868
rect 18141 5865 18153 5868
rect 18187 5865 18199 5899
rect 18141 5859 18199 5865
rect 20257 5899 20315 5905
rect 20257 5865 20269 5899
rect 20303 5896 20315 5899
rect 20622 5896 20628 5908
rect 20303 5868 20628 5896
rect 20303 5865 20315 5868
rect 20257 5859 20315 5865
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 21174 5856 21180 5908
rect 21232 5856 21238 5908
rect 21542 5856 21548 5908
rect 21600 5856 21606 5908
rect 21634 5856 21640 5908
rect 21692 5896 21698 5908
rect 22281 5899 22339 5905
rect 22281 5896 22293 5899
rect 21692 5868 22293 5896
rect 21692 5856 21698 5868
rect 22281 5865 22293 5868
rect 22327 5865 22339 5899
rect 23753 5899 23811 5905
rect 23753 5896 23765 5899
rect 22281 5859 22339 5865
rect 22388 5868 23765 5896
rect 20717 5831 20775 5837
rect 20717 5828 20729 5831
rect 19306 5800 20729 5828
rect 16439 5732 17080 5760
rect 16439 5729 16451 5732
rect 16393 5723 16451 5729
rect 17126 5720 17132 5772
rect 17184 5720 17190 5772
rect 11193 5664 11560 5692
rect 11193 5661 11205 5664
rect 11147 5655 11205 5661
rect 11606 5652 11612 5704
rect 11664 5652 11670 5704
rect 11882 5652 11888 5704
rect 11940 5692 11946 5704
rect 11940 5671 12554 5692
rect 11940 5665 12569 5671
rect 11940 5664 12523 5665
rect 11940 5652 11946 5664
rect 11054 5584 11060 5636
rect 11112 5584 11118 5636
rect 12511 5631 12523 5664
rect 12557 5631 12569 5665
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 13320 5664 14780 5692
rect 13320 5652 13326 5664
rect 12511 5625 12569 5631
rect 10284 5528 10916 5556
rect 14752 5556 14780 5664
rect 15194 5652 15200 5704
rect 15252 5652 15258 5704
rect 15286 5652 15292 5704
rect 15344 5692 15350 5704
rect 15381 5695 15439 5701
rect 15381 5692 15393 5695
rect 15344 5664 15393 5692
rect 15344 5652 15350 5664
rect 15381 5661 15393 5664
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 15562 5652 15568 5704
rect 15620 5652 15626 5704
rect 17402 5692 17408 5704
rect 17363 5664 17408 5692
rect 17402 5652 17408 5664
rect 17460 5652 17466 5704
rect 17494 5652 17500 5704
rect 17552 5652 17558 5704
rect 17512 5624 17540 5652
rect 19306 5624 19334 5800
rect 20717 5797 20729 5800
rect 20763 5797 20775 5831
rect 21450 5828 21456 5840
rect 20717 5791 20775 5797
rect 20824 5800 21456 5828
rect 20824 5760 20852 5800
rect 21450 5788 21456 5800
rect 21508 5788 21514 5840
rect 21726 5788 21732 5840
rect 21784 5828 21790 5840
rect 21821 5831 21879 5837
rect 21821 5828 21833 5831
rect 21784 5800 21833 5828
rect 21784 5788 21790 5800
rect 21821 5797 21833 5800
rect 21867 5797 21879 5831
rect 21821 5791 21879 5797
rect 20456 5732 20852 5760
rect 20456 5701 20484 5732
rect 20898 5720 20904 5772
rect 20956 5720 20962 5772
rect 20990 5720 20996 5772
rect 21048 5760 21054 5772
rect 22388 5760 22416 5868
rect 23753 5865 23765 5868
rect 23799 5865 23811 5899
rect 23753 5859 23811 5865
rect 24210 5856 24216 5908
rect 24268 5856 24274 5908
rect 25866 5760 25872 5772
rect 21048 5732 22416 5760
rect 23860 5732 25872 5760
rect 21048 5720 21054 5732
rect 20441 5695 20499 5701
rect 20441 5661 20453 5695
rect 20487 5661 20499 5695
rect 20441 5655 20499 5661
rect 20717 5695 20775 5701
rect 20717 5661 20729 5695
rect 20763 5692 20775 5695
rect 21266 5692 21272 5704
rect 20763 5688 20852 5692
rect 20916 5688 21272 5692
rect 20763 5664 21272 5688
rect 20763 5661 20775 5664
rect 20717 5655 20775 5661
rect 20824 5660 20944 5664
rect 21266 5652 21272 5664
rect 21324 5652 21330 5704
rect 21376 5701 21404 5732
rect 21361 5695 21419 5701
rect 21361 5661 21373 5695
rect 21407 5661 21419 5695
rect 21361 5655 21419 5661
rect 21453 5695 21511 5701
rect 21453 5661 21465 5695
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 17512 5596 19334 5624
rect 21085 5627 21143 5633
rect 21085 5593 21097 5627
rect 21131 5593 21143 5627
rect 21085 5587 21143 5593
rect 17037 5559 17095 5565
rect 17037 5556 17049 5559
rect 14752 5528 17049 5556
rect 10284 5516 10290 5528
rect 17037 5525 17049 5528
rect 17083 5525 17095 5559
rect 17037 5519 17095 5525
rect 18046 5516 18052 5568
rect 18104 5556 18110 5568
rect 19058 5556 19064 5568
rect 18104 5528 19064 5556
rect 18104 5516 18110 5528
rect 19058 5516 19064 5528
rect 19116 5516 19122 5568
rect 20806 5516 20812 5568
rect 20864 5556 20870 5568
rect 21100 5556 21128 5587
rect 20864 5528 21128 5556
rect 21468 5556 21496 5655
rect 21634 5652 21640 5704
rect 21692 5652 21698 5704
rect 21729 5695 21787 5701
rect 21729 5661 21741 5695
rect 21775 5692 21787 5695
rect 21910 5692 21916 5704
rect 21775 5664 21916 5692
rect 21775 5661 21787 5664
rect 21729 5655 21787 5661
rect 21910 5652 21916 5664
rect 21968 5652 21974 5704
rect 22094 5652 22100 5704
rect 22152 5652 22158 5704
rect 22373 5695 22431 5701
rect 22373 5661 22385 5695
rect 22419 5692 22431 5695
rect 22554 5692 22560 5704
rect 22419 5664 22560 5692
rect 22419 5661 22431 5664
rect 22373 5655 22431 5661
rect 22554 5652 22560 5664
rect 22612 5652 22618 5704
rect 22647 5695 22705 5701
rect 22647 5661 22659 5695
rect 22693 5692 22705 5695
rect 23860 5692 23888 5732
rect 25866 5720 25872 5732
rect 25924 5720 25930 5772
rect 22693 5664 23888 5692
rect 22693 5661 22705 5664
rect 22647 5655 22705 5661
rect 23934 5652 23940 5704
rect 23992 5652 23998 5704
rect 24029 5695 24087 5701
rect 24029 5661 24041 5695
rect 24075 5692 24087 5695
rect 25314 5692 25320 5704
rect 24075 5664 25320 5692
rect 24075 5661 24087 5664
rect 24029 5655 24087 5661
rect 25314 5652 25320 5664
rect 25372 5652 25378 5704
rect 22922 5624 22928 5636
rect 22664 5596 22928 5624
rect 22664 5556 22692 5596
rect 22922 5584 22928 5596
rect 22980 5584 22986 5636
rect 21468 5528 22692 5556
rect 20864 5516 20870 5528
rect 22738 5516 22744 5568
rect 22796 5556 22802 5568
rect 23385 5559 23443 5565
rect 23385 5556 23397 5559
rect 22796 5528 23397 5556
rect 22796 5516 22802 5528
rect 23385 5525 23397 5528
rect 23431 5525 23443 5559
rect 23385 5519 23443 5525
rect 1104 5466 25000 5488
rect 1104 5414 6884 5466
rect 6936 5414 6948 5466
rect 7000 5414 7012 5466
rect 7064 5414 7076 5466
rect 7128 5414 7140 5466
rect 7192 5414 12818 5466
rect 12870 5414 12882 5466
rect 12934 5414 12946 5466
rect 12998 5414 13010 5466
rect 13062 5414 13074 5466
rect 13126 5414 18752 5466
rect 18804 5414 18816 5466
rect 18868 5414 18880 5466
rect 18932 5414 18944 5466
rect 18996 5414 19008 5466
rect 19060 5414 24686 5466
rect 24738 5414 24750 5466
rect 24802 5414 24814 5466
rect 24866 5414 24878 5466
rect 24930 5414 24942 5466
rect 24994 5414 25000 5466
rect 1104 5392 25000 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1452 5324 1593 5352
rect 1452 5312 1458 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 1581 5315 1639 5321
rect 2130 5312 2136 5364
rect 2188 5312 2194 5364
rect 2590 5312 2596 5364
rect 2648 5312 2654 5364
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 2869 5355 2927 5361
rect 2869 5352 2881 5355
rect 2832 5324 2881 5352
rect 2832 5312 2838 5324
rect 2869 5321 2881 5324
rect 2915 5321 2927 5355
rect 4062 5352 4068 5364
rect 2869 5315 2927 5321
rect 3160 5324 4068 5352
rect 2038 5244 2044 5296
rect 2096 5244 2102 5296
rect 2608 5284 2636 5312
rect 3160 5284 3188 5324
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4338 5312 4344 5364
rect 4396 5312 4402 5364
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 6178 5352 6184 5364
rect 5951 5324 6184 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 7374 5312 7380 5364
rect 7432 5312 7438 5364
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 9582 5352 9588 5364
rect 7524 5324 9588 5352
rect 7524 5312 7530 5324
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 9692 5324 11468 5352
rect 9692 5284 9720 5324
rect 2608 5256 3188 5284
rect 1489 5219 1547 5225
rect 1489 5185 1501 5219
rect 1535 5216 1547 5219
rect 1535 5188 2544 5216
rect 1535 5185 1547 5188
rect 1489 5179 1547 5185
rect 2516 5080 2544 5188
rect 2590 5176 2596 5228
rect 2648 5176 2654 5228
rect 3160 5148 3188 5256
rect 3252 5256 9720 5284
rect 3252 5225 3280 5256
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 3603 5219 3661 5225
rect 3603 5185 3615 5219
rect 3649 5216 3661 5219
rect 4522 5216 4528 5228
rect 3649 5188 4528 5216
rect 3649 5185 3661 5188
rect 3603 5179 3661 5185
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 4798 5176 4804 5228
rect 4856 5216 4862 5228
rect 5135 5219 5193 5225
rect 5135 5216 5147 5219
rect 4856 5188 5147 5216
rect 4856 5176 4862 5188
rect 5135 5185 5147 5188
rect 5181 5185 5193 5219
rect 5135 5179 5193 5185
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 6607 5219 6665 5225
rect 6607 5216 6619 5219
rect 6328 5188 6619 5216
rect 6328 5176 6334 5188
rect 6607 5185 6619 5188
rect 6653 5185 6665 5219
rect 6607 5179 6665 5185
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 8478 5216 8484 5228
rect 7340 5188 8484 5216
rect 7340 5176 7346 5188
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 9122 5176 9128 5228
rect 9180 5176 9186 5228
rect 9490 5176 9496 5228
rect 9548 5176 9554 5228
rect 10594 5225 10600 5228
rect 10551 5219 10600 5225
rect 10551 5185 10563 5219
rect 10597 5185 10600 5219
rect 10551 5179 10600 5185
rect 10594 5176 10600 5179
rect 10652 5176 10658 5228
rect 3329 5151 3387 5157
rect 3329 5148 3341 5151
rect 3160 5120 3341 5148
rect 3329 5117 3341 5120
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 4893 5151 4951 5157
rect 4893 5148 4905 5151
rect 4120 5120 4905 5148
rect 4120 5108 4126 5120
rect 4893 5117 4905 5120
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 6365 5151 6423 5157
rect 6365 5117 6377 5151
rect 6411 5117 6423 5151
rect 9140 5148 9168 5176
rect 6365 5111 6423 5117
rect 7024 5120 9168 5148
rect 2516 5052 3372 5080
rect 3344 5024 3372 5052
rect 3050 4972 3056 5024
rect 3108 4972 3114 5024
rect 3326 4972 3332 5024
rect 3384 4972 3390 5024
rect 4908 5012 4936 5111
rect 6380 5012 6408 5111
rect 7024 5012 7052 5120
rect 9674 5108 9680 5160
rect 9732 5108 9738 5160
rect 10134 5108 10140 5160
rect 10192 5108 10198 5160
rect 10410 5148 10416 5160
rect 10244 5120 10416 5148
rect 8294 5040 8300 5092
rect 8352 5080 8358 5092
rect 8662 5080 8668 5092
rect 8352 5052 8668 5080
rect 8352 5040 8358 5052
rect 8662 5040 8668 5052
rect 8720 5080 8726 5092
rect 10244 5080 10272 5120
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5148 10747 5151
rect 11238 5148 11244 5160
rect 10735 5120 11244 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 8720 5052 10272 5080
rect 8720 5040 8726 5052
rect 4908 4984 7052 5012
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 11333 5015 11391 5021
rect 11333 5012 11345 5015
rect 7432 4984 11345 5012
rect 7432 4972 7438 4984
rect 11333 4981 11345 4984
rect 11379 4981 11391 5015
rect 11440 5012 11468 5324
rect 13538 5312 13544 5364
rect 13596 5312 13602 5364
rect 14550 5312 14556 5364
rect 14608 5352 14614 5364
rect 15286 5352 15292 5364
rect 14608 5324 15292 5352
rect 14608 5312 14614 5324
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 16574 5312 16580 5364
rect 16632 5352 16638 5364
rect 20714 5352 20720 5364
rect 16632 5324 20720 5352
rect 16632 5312 16638 5324
rect 20714 5312 20720 5324
rect 20772 5312 20778 5364
rect 20898 5312 20904 5364
rect 20956 5312 20962 5364
rect 21174 5312 21180 5364
rect 21232 5312 21238 5364
rect 21266 5312 21272 5364
rect 21324 5352 21330 5364
rect 21361 5355 21419 5361
rect 21361 5352 21373 5355
rect 21324 5324 21373 5352
rect 21324 5312 21330 5324
rect 21361 5321 21373 5324
rect 21407 5321 21419 5355
rect 21361 5315 21419 5321
rect 21821 5355 21879 5361
rect 21821 5321 21833 5355
rect 21867 5352 21879 5355
rect 21867 5324 21956 5352
rect 21867 5321 21879 5324
rect 21821 5315 21879 5321
rect 12526 5255 12532 5296
rect 12511 5249 12532 5255
rect 12584 5284 12590 5296
rect 13556 5284 13584 5312
rect 18138 5284 18144 5296
rect 12584 5256 13584 5284
rect 15394 5256 18144 5284
rect 12511 5215 12523 5249
rect 12584 5244 12590 5256
rect 12557 5218 12572 5244
rect 12557 5215 12569 5218
rect 12511 5209 12569 5215
rect 13630 5176 13636 5228
rect 13688 5176 13694 5228
rect 14826 5176 14832 5228
rect 14884 5176 14890 5228
rect 12250 5108 12256 5160
rect 12308 5108 12314 5160
rect 13817 5151 13875 5157
rect 13817 5117 13829 5151
rect 13863 5148 13875 5151
rect 13998 5148 14004 5160
rect 13863 5120 14004 5148
rect 13863 5117 13875 5120
rect 13817 5111 13875 5117
rect 13998 5108 14004 5120
rect 14056 5108 14062 5160
rect 14550 5108 14556 5160
rect 14608 5108 14614 5160
rect 14642 5108 14648 5160
rect 14700 5157 14706 5160
rect 14700 5151 14749 5157
rect 14700 5117 14703 5151
rect 14737 5148 14749 5151
rect 15394 5148 15422 5256
rect 18138 5244 18144 5256
rect 18196 5244 18202 5296
rect 18690 5244 18696 5296
rect 18748 5284 18754 5296
rect 18748 5256 20484 5284
rect 18748 5244 18754 5256
rect 17402 5176 17408 5228
rect 17460 5216 17466 5228
rect 19027 5219 19085 5225
rect 19027 5216 19039 5219
rect 17460 5188 19039 5216
rect 17460 5176 17466 5188
rect 19027 5185 19039 5188
rect 19073 5185 19085 5219
rect 19027 5179 19085 5185
rect 19794 5176 19800 5228
rect 19852 5216 19858 5228
rect 20349 5219 20407 5225
rect 20349 5216 20361 5219
rect 19852 5188 20361 5216
rect 19852 5176 19858 5188
rect 20349 5185 20361 5188
rect 20395 5185 20407 5219
rect 20349 5179 20407 5185
rect 14737 5120 15422 5148
rect 14737 5117 14749 5120
rect 14700 5111 14749 5117
rect 14700 5108 14706 5111
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 17862 5148 17868 5160
rect 17276 5120 17868 5148
rect 17276 5108 17282 5120
rect 17862 5108 17868 5120
rect 17920 5148 17926 5160
rect 18785 5151 18843 5157
rect 18785 5148 18797 5151
rect 17920 5120 18797 5148
rect 17920 5108 17926 5120
rect 18785 5117 18797 5120
rect 18831 5117 18843 5151
rect 18785 5111 18843 5117
rect 20165 5151 20223 5157
rect 20165 5117 20177 5151
rect 20211 5117 20223 5151
rect 20165 5111 20223 5117
rect 13265 5083 13323 5089
rect 13265 5049 13277 5083
rect 13311 5080 13323 5083
rect 14277 5083 14335 5089
rect 14277 5080 14289 5083
rect 13311 5052 14289 5080
rect 13311 5049 13323 5052
rect 13265 5043 13323 5049
rect 14277 5049 14289 5052
rect 14323 5049 14335 5083
rect 14277 5043 14335 5049
rect 19797 5083 19855 5089
rect 19797 5049 19809 5083
rect 19843 5080 19855 5083
rect 19978 5080 19984 5092
rect 19843 5052 19984 5080
rect 19843 5049 19855 5052
rect 19797 5043 19855 5049
rect 19978 5040 19984 5052
rect 20036 5080 20042 5092
rect 20180 5080 20208 5111
rect 20036 5052 20208 5080
rect 20349 5083 20407 5089
rect 20036 5040 20042 5052
rect 20349 5049 20361 5083
rect 20395 5049 20407 5083
rect 20349 5043 20407 5049
rect 15473 5015 15531 5021
rect 15473 5012 15485 5015
rect 11440 4984 15485 5012
rect 11333 4975 11391 4981
rect 15473 4981 15485 4984
rect 15519 4981 15531 5015
rect 15473 4975 15531 4981
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 20364 5012 20392 5043
rect 17000 4984 20392 5012
rect 20456 5012 20484 5256
rect 20714 5176 20720 5228
rect 20772 5176 20778 5228
rect 20916 5216 20944 5312
rect 21192 5284 21220 5312
rect 21192 5256 21312 5284
rect 21284 5225 21312 5256
rect 20993 5219 21051 5225
rect 20993 5216 21005 5219
rect 20916 5188 21005 5216
rect 20993 5185 21005 5188
rect 21039 5185 21051 5219
rect 20993 5179 21051 5185
rect 21177 5219 21235 5225
rect 21177 5185 21189 5219
rect 21223 5185 21235 5219
rect 21177 5179 21235 5185
rect 21269 5219 21327 5225
rect 21269 5185 21281 5219
rect 21315 5185 21327 5219
rect 21928 5216 21956 5324
rect 22278 5312 22284 5364
rect 22336 5312 22342 5364
rect 22554 5312 22560 5364
rect 22612 5312 22618 5364
rect 22649 5355 22707 5361
rect 22649 5321 22661 5355
rect 22695 5352 22707 5355
rect 23658 5352 23664 5364
rect 22695 5324 23664 5352
rect 22695 5321 22707 5324
rect 22649 5315 22707 5321
rect 23658 5312 23664 5324
rect 23716 5312 23722 5364
rect 24394 5312 24400 5364
rect 24452 5312 24458 5364
rect 22570 5256 23428 5284
rect 21269 5179 21327 5185
rect 21376 5188 21956 5216
rect 22005 5219 22063 5225
rect 20806 5108 20812 5160
rect 20864 5148 20870 5160
rect 21085 5151 21143 5157
rect 21085 5148 21097 5151
rect 20864 5120 21097 5148
rect 20864 5108 20870 5120
rect 21085 5117 21097 5120
rect 21131 5117 21143 5151
rect 21192 5148 21220 5179
rect 21376 5148 21404 5188
rect 22005 5185 22017 5219
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 22097 5219 22155 5225
rect 22097 5185 22109 5219
rect 22143 5216 22155 5219
rect 22278 5216 22284 5228
rect 22143 5188 22284 5216
rect 22143 5185 22155 5188
rect 22097 5179 22155 5185
rect 21192 5120 21404 5148
rect 21085 5111 21143 5117
rect 21542 5108 21548 5160
rect 21600 5148 21606 5160
rect 22020 5148 22048 5179
rect 22278 5176 22284 5188
rect 22336 5176 22342 5228
rect 22373 5219 22431 5225
rect 22373 5185 22385 5219
rect 22419 5216 22431 5219
rect 22462 5216 22468 5228
rect 22419 5188 22468 5216
rect 22419 5185 22431 5188
rect 22373 5179 22431 5185
rect 22462 5176 22468 5188
rect 22520 5176 22526 5228
rect 21600 5120 22048 5148
rect 21600 5108 21606 5120
rect 22570 5012 22598 5256
rect 22833 5219 22891 5225
rect 22833 5214 22845 5219
rect 22725 5186 22845 5214
rect 22725 5080 22753 5186
rect 22833 5185 22845 5186
rect 22879 5185 22891 5219
rect 22833 5179 22891 5185
rect 22922 5176 22928 5228
rect 22980 5176 22986 5228
rect 23106 5176 23112 5228
rect 23164 5176 23170 5228
rect 23400 5225 23428 5256
rect 23750 5244 23756 5296
rect 23808 5244 23814 5296
rect 23385 5219 23443 5225
rect 23385 5185 23397 5219
rect 23431 5185 23443 5219
rect 23385 5179 23443 5185
rect 24026 5176 24032 5228
rect 24084 5176 24090 5228
rect 24305 5219 24363 5225
rect 24305 5185 24317 5219
rect 24351 5216 24363 5219
rect 25038 5216 25044 5228
rect 24351 5188 25044 5216
rect 24351 5185 24363 5188
rect 24305 5179 24363 5185
rect 25038 5176 25044 5188
rect 25096 5176 25102 5228
rect 22940 5148 22968 5176
rect 23201 5151 23259 5157
rect 23201 5148 23213 5151
rect 22940 5120 23213 5148
rect 23201 5117 23213 5120
rect 23247 5148 23259 5151
rect 24210 5148 24216 5160
rect 23247 5120 24216 5148
rect 23247 5117 23259 5120
rect 23201 5111 23259 5117
rect 24210 5108 24216 5120
rect 24268 5108 24274 5160
rect 23382 5080 23388 5092
rect 22725 5052 23388 5080
rect 23382 5040 23388 5052
rect 23440 5040 23446 5092
rect 23474 5040 23480 5092
rect 23532 5040 23538 5092
rect 20456 4984 22598 5012
rect 17000 4972 17006 4984
rect 22922 4972 22928 5024
rect 22980 4972 22986 5024
rect 23845 5015 23903 5021
rect 23845 4981 23857 5015
rect 23891 5012 23903 5015
rect 24118 5012 24124 5024
rect 23891 4984 24124 5012
rect 23891 4981 23903 4984
rect 23845 4975 23903 4981
rect 24118 4972 24124 4984
rect 24176 4972 24182 5024
rect 1104 4922 24840 4944
rect 1104 4870 3917 4922
rect 3969 4870 3981 4922
rect 4033 4870 4045 4922
rect 4097 4870 4109 4922
rect 4161 4870 4173 4922
rect 4225 4870 9851 4922
rect 9903 4870 9915 4922
rect 9967 4870 9979 4922
rect 10031 4870 10043 4922
rect 10095 4870 10107 4922
rect 10159 4870 15785 4922
rect 15837 4870 15849 4922
rect 15901 4870 15913 4922
rect 15965 4870 15977 4922
rect 16029 4870 16041 4922
rect 16093 4870 21719 4922
rect 21771 4870 21783 4922
rect 21835 4870 21847 4922
rect 21899 4870 21911 4922
rect 21963 4870 21975 4922
rect 22027 4870 24840 4922
rect 1104 4848 24840 4870
rect 1578 4768 1584 4820
rect 1636 4768 1642 4820
rect 2501 4811 2559 4817
rect 2501 4777 2513 4811
rect 2547 4808 2559 4811
rect 2590 4808 2596 4820
rect 2547 4780 2596 4808
rect 2547 4777 2559 4780
rect 2501 4771 2559 4777
rect 2590 4768 2596 4780
rect 2648 4768 2654 4820
rect 2682 4768 2688 4820
rect 2740 4808 2746 4820
rect 2777 4811 2835 4817
rect 2777 4808 2789 4811
rect 2740 4780 2789 4808
rect 2740 4768 2746 4780
rect 2777 4777 2789 4780
rect 2823 4777 2835 4811
rect 2777 4771 2835 4777
rect 3050 4768 3056 4820
rect 3108 4768 3114 4820
rect 4706 4768 4712 4820
rect 4764 4768 4770 4820
rect 8294 4808 8300 4820
rect 7576 4780 8300 4808
rect 3068 4740 3096 4768
rect 7576 4740 7604 4780
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 9732 4780 11100 4808
rect 9732 4768 9738 4780
rect 1504 4712 3096 4740
rect 3436 4712 7604 4740
rect 1504 4613 1532 4712
rect 1946 4632 1952 4684
rect 2004 4632 2010 4684
rect 3436 4672 3464 4712
rect 9122 4700 9128 4752
rect 9180 4740 9186 4752
rect 10042 4740 10048 4752
rect 9180 4712 10048 4740
rect 9180 4700 9186 4712
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 11072 4740 11100 4780
rect 11146 4768 11152 4820
rect 11204 4768 11210 4820
rect 12710 4808 12716 4820
rect 11716 4780 12716 4808
rect 11716 4740 11744 4780
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 14108 4780 14780 4808
rect 11072 4712 11744 4740
rect 12342 4700 12348 4752
rect 12400 4740 12406 4752
rect 14108 4740 14136 4780
rect 12400 4712 14136 4740
rect 14752 4740 14780 4780
rect 14826 4768 14832 4820
rect 14884 4808 14890 4820
rect 15105 4811 15163 4817
rect 15105 4808 15117 4811
rect 14884 4780 15117 4808
rect 14884 4768 14890 4780
rect 15105 4777 15117 4780
rect 15151 4777 15163 4811
rect 15105 4771 15163 4777
rect 15212 4780 18359 4808
rect 15212 4740 15240 4780
rect 14752 4712 15240 4740
rect 12400 4700 12406 4712
rect 7374 4672 7380 4684
rect 2976 4644 3464 4672
rect 3528 4644 7380 4672
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4573 1547 4607
rect 1489 4567 1547 4573
rect 1964 4536 1992 4632
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4604 2099 4607
rect 2314 4604 2320 4616
rect 2087 4576 2320 4604
rect 2087 4573 2099 4576
rect 2041 4567 2099 4573
rect 2314 4564 2320 4576
rect 2372 4564 2378 4616
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 2866 4604 2872 4616
rect 2731 4576 2872 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 2976 4613 3004 4644
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4573 3019 4607
rect 2961 4567 3019 4573
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4604 3295 4607
rect 3418 4604 3424 4616
rect 3283 4576 3424 4604
rect 3283 4573 3295 4576
rect 3237 4567 3295 4573
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 3528 4613 3556 4644
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 10134 4672 10140 4684
rect 8536 4644 10140 4672
rect 8536 4632 8542 4644
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 11606 4632 11612 4684
rect 11664 4632 11670 4684
rect 14108 4681 14136 4712
rect 14844 4684 14872 4712
rect 16942 4700 16948 4752
rect 17000 4700 17006 4752
rect 14093 4675 14151 4681
rect 14093 4641 14105 4675
rect 14139 4641 14151 4675
rect 14093 4635 14151 4641
rect 14826 4632 14832 4684
rect 14884 4632 14890 4684
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4604 4951 4607
rect 5166 4604 5172 4616
rect 4939 4576 5172 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 7282 4564 7288 4616
rect 7340 4604 7346 4616
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 7340 4576 7481 4604
rect 7340 4564 7346 4576
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 7743 4607 7801 4613
rect 7743 4573 7755 4607
rect 7789 4573 7801 4607
rect 9766 4604 9772 4616
rect 7743 4567 7801 4573
rect 8404 4576 9772 4604
rect 7758 4536 7786 4567
rect 1964 4508 2268 4536
rect 1118 4428 1124 4480
rect 1176 4468 1182 4480
rect 2133 4471 2191 4477
rect 2133 4468 2145 4471
rect 1176 4440 2145 4468
rect 1176 4428 1182 4440
rect 2133 4437 2145 4440
rect 2179 4437 2191 4471
rect 2240 4468 2268 4508
rect 2746 4508 3096 4536
rect 7758 4508 8064 4536
rect 2746 4468 2774 4508
rect 3068 4477 3096 4508
rect 2240 4440 2774 4468
rect 3053 4471 3111 4477
rect 2133 4431 2191 4437
rect 3053 4437 3065 4471
rect 3099 4437 3111 4471
rect 3053 4431 3111 4437
rect 3326 4428 3332 4480
rect 3384 4428 3390 4480
rect 4062 4428 4068 4480
rect 4120 4468 4126 4480
rect 7466 4468 7472 4480
rect 4120 4440 7472 4468
rect 4120 4428 4126 4440
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 8036 4468 8064 4508
rect 8404 4468 8432 4576
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 10318 4564 10324 4616
rect 10376 4604 10382 4616
rect 10411 4607 10469 4613
rect 10411 4604 10423 4607
rect 10376 4576 10423 4604
rect 10376 4564 10382 4576
rect 10411 4573 10423 4576
rect 10457 4573 10469 4607
rect 10411 4567 10469 4573
rect 10502 4564 10508 4616
rect 10560 4604 10566 4616
rect 12526 4604 12532 4616
rect 10560 4577 12532 4604
rect 10560 4576 11879 4577
rect 10560 4564 10566 4576
rect 11867 4543 11879 4576
rect 11913 4576 12532 4577
rect 11913 4546 11928 4576
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 14366 4604 14372 4616
rect 14327 4576 14372 4604
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 11913 4543 11925 4546
rect 11867 4537 11925 4543
rect 16960 4536 16988 4700
rect 17218 4564 17224 4616
rect 17276 4564 17282 4616
rect 17479 4577 17537 4583
rect 17479 4543 17491 4577
rect 17525 4543 17537 4577
rect 17479 4537 17537 4543
rect 11992 4508 16988 4536
rect 8036 4440 8432 4468
rect 8481 4471 8539 4477
rect 8481 4437 8493 4471
rect 8527 4468 8539 4471
rect 8754 4468 8760 4480
rect 8527 4440 8760 4468
rect 8527 4437 8539 4440
rect 8481 4431 8539 4437
rect 8754 4428 8760 4440
rect 8812 4428 8818 4480
rect 8846 4428 8852 4480
rect 8904 4468 8910 4480
rect 11992 4468 12020 4508
rect 8904 4440 12020 4468
rect 8904 4428 8910 4440
rect 12342 4428 12348 4480
rect 12400 4468 12406 4480
rect 12621 4471 12679 4477
rect 12621 4468 12633 4471
rect 12400 4440 12633 4468
rect 12400 4428 12406 4440
rect 12621 4437 12633 4440
rect 12667 4437 12679 4471
rect 12621 4431 12679 4437
rect 12710 4428 12716 4480
rect 12768 4468 12774 4480
rect 17310 4468 17316 4480
rect 12768 4440 17316 4468
rect 12768 4428 12774 4440
rect 17310 4428 17316 4440
rect 17368 4468 17374 4480
rect 17494 4468 17522 4537
rect 17368 4440 17522 4468
rect 17368 4428 17374 4440
rect 18230 4428 18236 4480
rect 18288 4428 18294 4480
rect 18331 4468 18359 4780
rect 18690 4768 18696 4820
rect 18748 4768 18754 4820
rect 18877 4811 18935 4817
rect 18877 4777 18889 4811
rect 18923 4808 18935 4811
rect 19702 4808 19708 4820
rect 18923 4780 19708 4808
rect 18923 4777 18935 4780
rect 18877 4771 18935 4777
rect 19702 4768 19708 4780
rect 19760 4768 19766 4820
rect 19794 4768 19800 4820
rect 19852 4768 19858 4820
rect 20073 4811 20131 4817
rect 20073 4777 20085 4811
rect 20119 4808 20131 4811
rect 20714 4808 20720 4820
rect 20119 4780 20720 4808
rect 20119 4777 20131 4780
rect 20073 4771 20131 4777
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 21542 4768 21548 4820
rect 21600 4768 21606 4820
rect 22370 4768 22376 4820
rect 22428 4808 22434 4820
rect 22465 4811 22523 4817
rect 22465 4808 22477 4811
rect 22428 4780 22477 4808
rect 22428 4768 22434 4780
rect 22465 4777 22477 4780
rect 22511 4777 22523 4811
rect 22465 4771 22523 4777
rect 24029 4811 24087 4817
rect 24029 4777 24041 4811
rect 24075 4808 24087 4811
rect 25406 4808 25412 4820
rect 24075 4780 25412 4808
rect 24075 4777 24087 4780
rect 24029 4771 24087 4777
rect 25406 4768 25412 4780
rect 25464 4768 25470 4820
rect 19429 4743 19487 4749
rect 19429 4709 19441 4743
rect 19475 4740 19487 4743
rect 20162 4740 20168 4752
rect 19475 4712 20168 4740
rect 19475 4709 19487 4712
rect 19429 4703 19487 4709
rect 20162 4700 20168 4712
rect 20220 4700 20226 4752
rect 21560 4740 21588 4768
rect 21913 4743 21971 4749
rect 21913 4740 21925 4743
rect 21560 4712 21925 4740
rect 21913 4709 21925 4712
rect 21959 4709 21971 4743
rect 21913 4703 21971 4709
rect 20530 4672 20536 4684
rect 19352 4644 20536 4672
rect 19352 4616 19380 4644
rect 20530 4632 20536 4644
rect 20588 4632 20594 4684
rect 22922 4672 22928 4684
rect 21560 4644 22928 4672
rect 18601 4607 18659 4613
rect 18601 4573 18613 4607
rect 18647 4573 18659 4607
rect 18601 4567 18659 4573
rect 18616 4536 18644 4567
rect 18690 4564 18696 4616
rect 18748 4604 18754 4616
rect 19061 4607 19119 4613
rect 19061 4604 19073 4607
rect 18748 4576 19073 4604
rect 18748 4564 18754 4576
rect 19061 4573 19073 4576
rect 19107 4573 19119 4607
rect 19061 4567 19119 4573
rect 19334 4564 19340 4616
rect 19392 4564 19398 4616
rect 19610 4564 19616 4616
rect 19668 4564 19674 4616
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4573 19763 4607
rect 19705 4567 19763 4573
rect 19518 4536 19524 4548
rect 18616 4508 19524 4536
rect 19518 4496 19524 4508
rect 19576 4496 19582 4548
rect 19720 4536 19748 4567
rect 19978 4564 19984 4616
rect 20036 4564 20042 4616
rect 20162 4564 20168 4616
rect 20220 4564 20226 4616
rect 20438 4564 20444 4616
rect 20496 4604 20502 4616
rect 21560 4604 21588 4644
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 23198 4632 23204 4684
rect 23256 4632 23262 4684
rect 22189 4607 22247 4613
rect 22189 4604 22201 4607
rect 20496 4576 21588 4604
rect 21652 4576 22201 4604
rect 20496 4564 20502 4576
rect 20800 4539 20858 4545
rect 19720 4508 20300 4536
rect 20162 4468 20168 4480
rect 18331 4440 20168 4468
rect 20162 4428 20168 4440
rect 20220 4428 20226 4480
rect 20272 4477 20300 4508
rect 20800 4505 20812 4539
rect 20846 4536 20858 4539
rect 20990 4536 20996 4548
rect 20846 4508 20996 4536
rect 20846 4505 20858 4508
rect 20800 4499 20858 4505
rect 20990 4496 20996 4508
rect 21048 4496 21054 4548
rect 21082 4496 21088 4548
rect 21140 4536 21146 4548
rect 21652 4536 21680 4576
rect 22189 4573 22201 4576
rect 22235 4573 22247 4607
rect 22189 4567 22247 4573
rect 22281 4607 22339 4613
rect 22281 4573 22293 4607
rect 22327 4604 22339 4607
rect 22554 4604 22560 4616
rect 22327 4576 22560 4604
rect 22327 4573 22339 4576
rect 22281 4567 22339 4573
rect 22554 4564 22560 4576
rect 22612 4564 22618 4616
rect 22646 4564 22652 4616
rect 22704 4564 22710 4616
rect 21140 4508 21680 4536
rect 21140 4496 21146 4508
rect 23658 4496 23664 4548
rect 23716 4536 23722 4548
rect 23937 4539 23995 4545
rect 23937 4536 23949 4539
rect 23716 4508 23949 4536
rect 23716 4496 23722 4508
rect 23937 4505 23949 4508
rect 23983 4505 23995 4539
rect 23937 4499 23995 4505
rect 20257 4471 20315 4477
rect 20257 4437 20269 4471
rect 20303 4437 20315 4471
rect 20257 4431 20315 4437
rect 20530 4428 20536 4480
rect 20588 4468 20594 4480
rect 22005 4471 22063 4477
rect 22005 4468 22017 4471
rect 20588 4440 22017 4468
rect 20588 4428 20594 4440
rect 22005 4437 22017 4440
rect 22051 4437 22063 4471
rect 22005 4431 22063 4437
rect 1104 4378 25000 4400
rect 1104 4326 6884 4378
rect 6936 4326 6948 4378
rect 7000 4326 7012 4378
rect 7064 4326 7076 4378
rect 7128 4326 7140 4378
rect 7192 4326 12818 4378
rect 12870 4326 12882 4378
rect 12934 4326 12946 4378
rect 12998 4326 13010 4378
rect 13062 4326 13074 4378
rect 13126 4326 18752 4378
rect 18804 4326 18816 4378
rect 18868 4326 18880 4378
rect 18932 4326 18944 4378
rect 18996 4326 19008 4378
rect 19060 4326 24686 4378
rect 24738 4326 24750 4378
rect 24802 4326 24814 4378
rect 24866 4326 24878 4378
rect 24930 4326 24942 4378
rect 24994 4326 25000 4378
rect 1104 4304 25000 4326
rect 1578 4224 1584 4276
rect 1636 4224 1642 4276
rect 3326 4264 3332 4276
rect 2746 4236 3332 4264
rect 1489 4199 1547 4205
rect 1489 4165 1501 4199
rect 1535 4196 1547 4199
rect 2746 4196 2774 4236
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 3694 4224 3700 4276
rect 3752 4264 3758 4276
rect 3752 4236 5028 4264
rect 3752 4224 3758 4236
rect 1535 4168 2774 4196
rect 5000 4196 5028 4236
rect 5166 4224 5172 4276
rect 5224 4224 5230 4276
rect 5368 4236 9260 4264
rect 5368 4205 5396 4236
rect 5353 4199 5411 4205
rect 5353 4196 5365 4199
rect 5000 4168 5365 4196
rect 1535 4165 1547 4168
rect 1489 4159 1547 4165
rect 5353 4165 5365 4168
rect 5399 4165 5411 4199
rect 9232 4196 9260 4236
rect 9398 4224 9404 4276
rect 9456 4224 9462 4276
rect 9508 4236 9674 4264
rect 9508 4196 9536 4236
rect 9232 4168 9536 4196
rect 5353 4159 5411 4165
rect 1854 4088 1860 4140
rect 1912 4128 1918 4140
rect 1949 4131 2007 4137
rect 1949 4128 1961 4131
rect 1912 4100 1961 4128
rect 1912 4088 1918 4100
rect 1949 4097 1961 4100
rect 1995 4097 2007 4131
rect 1949 4091 2007 4097
rect 2223 4131 2281 4137
rect 2223 4097 2235 4131
rect 2269 4128 2281 4131
rect 2590 4128 2596 4140
rect 2269 4100 2596 4128
rect 2269 4097 2281 4100
rect 2223 4091 2281 4097
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3292 4100 3341 4128
rect 3292 4088 3298 4100
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3510 4088 3516 4140
rect 3568 4088 3574 4140
rect 4430 4137 4436 4140
rect 4387 4131 4436 4137
rect 4387 4097 4399 4131
rect 4433 4097 4436 4131
rect 4387 4091 4436 4097
rect 4430 4088 4436 4091
rect 4488 4088 4494 4140
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4128 7619 4131
rect 7607 4100 7880 4128
rect 7607 4097 7619 4100
rect 7561 4091 7619 4097
rect 7852 4072 7880 4100
rect 8754 4088 8760 4140
rect 8812 4088 8818 4140
rect 9646 4128 9674 4236
rect 12158 4224 12164 4276
rect 12216 4224 12222 4276
rect 13265 4267 13323 4273
rect 13265 4264 13277 4267
rect 12360 4236 13277 4264
rect 12360 4132 12388 4236
rect 13265 4233 13277 4236
rect 13311 4233 13323 4267
rect 13265 4227 13323 4233
rect 13446 4224 13452 4276
rect 13504 4224 13510 4276
rect 15194 4264 15200 4276
rect 14844 4236 15200 4264
rect 12437 4199 12495 4205
rect 12437 4165 12449 4199
rect 12483 4165 12495 4199
rect 12437 4159 12495 4165
rect 12084 4128 12388 4132
rect 9646 4104 12388 4128
rect 12452 4128 12480 4159
rect 12526 4156 12532 4208
rect 12584 4156 12590 4208
rect 12897 4199 12955 4205
rect 12897 4165 12909 4199
rect 12943 4196 12955 4199
rect 13630 4196 13636 4208
rect 12943 4168 13636 4196
rect 12943 4165 12955 4168
rect 12897 4159 12955 4165
rect 13630 4156 13636 4168
rect 13688 4156 13694 4208
rect 12618 4128 12624 4140
rect 9646 4100 12112 4104
rect 12452 4100 12624 4128
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 14645 4131 14703 4137
rect 14645 4097 14657 4131
rect 14691 4128 14703 4131
rect 14844 4128 14872 4236
rect 15194 4224 15200 4236
rect 15252 4264 15258 4276
rect 19334 4264 19340 4276
rect 15252 4236 16436 4264
rect 15252 4224 15258 4236
rect 14691 4100 14872 4128
rect 14691 4097 14703 4100
rect 14645 4091 14703 4097
rect 15010 4088 15016 4140
rect 15068 4088 15074 4140
rect 15654 4088 15660 4140
rect 15712 4137 15718 4140
rect 15712 4131 15740 4137
rect 15728 4097 15740 4131
rect 16408 4128 16436 4236
rect 19168 4236 19340 4264
rect 18230 4196 18236 4208
rect 17972 4168 18236 4196
rect 17681 4131 17739 4137
rect 16408 4100 17172 4128
rect 15712 4091 15740 4097
rect 15712 4088 15718 4091
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 4080 4032 4261 4060
rect 2961 3995 3019 4001
rect 2961 3961 2973 3995
rect 3007 3992 3019 3995
rect 3973 3995 4031 4001
rect 3973 3992 3985 3995
rect 3007 3964 3985 3992
rect 3007 3961 3019 3964
rect 2961 3955 3019 3961
rect 3973 3961 3985 3964
rect 4019 3961 4031 3995
rect 3973 3955 4031 3961
rect 4080 3924 4108 4032
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 4522 4020 4528 4072
rect 4580 4020 4586 4072
rect 7745 4063 7803 4069
rect 7745 4029 7757 4063
rect 7791 4029 7803 4063
rect 7745 4023 7803 4029
rect 5534 3952 5540 4004
rect 5592 3952 5598 4004
rect 7760 3992 7788 4023
rect 7834 4020 7840 4072
rect 7892 4020 7898 4072
rect 8662 4069 8668 4072
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 8312 4032 8493 4060
rect 8110 3992 8116 4004
rect 7760 3964 8116 3992
rect 8110 3952 8116 3964
rect 8168 3952 8174 4004
rect 8202 3952 8208 4004
rect 8260 3952 8266 4004
rect 5258 3924 5264 3936
rect 4080 3896 5264 3924
rect 5258 3884 5264 3896
rect 5316 3924 5322 3936
rect 6638 3924 6644 3936
rect 5316 3896 6644 3924
rect 5316 3884 5322 3896
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 8312 3924 8340 4032
rect 8481 4029 8493 4032
rect 8527 4029 8539 4063
rect 8481 4023 8539 4029
rect 8619 4063 8668 4069
rect 8619 4029 8631 4063
rect 8665 4029 8668 4063
rect 8619 4023 8668 4029
rect 8662 4020 8668 4023
rect 8720 4060 8726 4072
rect 10962 4060 10968 4072
rect 8720 4032 10968 4060
rect 8720 4020 8726 4032
rect 10962 4020 10968 4032
rect 11020 4020 11026 4072
rect 12342 4020 12348 4072
rect 12400 4020 12406 4072
rect 14550 4020 14556 4072
rect 14608 4060 14614 4072
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 14608 4032 14841 4060
rect 14608 4020 14614 4032
rect 14829 4029 14841 4032
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 9766 3952 9772 4004
rect 9824 3992 9830 4004
rect 11606 3992 11612 4004
rect 9824 3964 11612 3992
rect 9824 3952 9830 3964
rect 11606 3952 11612 3964
rect 11664 3952 11670 4004
rect 13906 3952 13912 4004
rect 13964 3992 13970 4004
rect 15028 3992 15056 4088
rect 15562 4020 15568 4072
rect 15620 4020 15626 4072
rect 15841 4063 15899 4069
rect 15841 4029 15853 4063
rect 15887 4060 15899 4063
rect 17034 4060 17040 4072
rect 15887 4032 17040 4060
rect 15887 4029 15899 4032
rect 15841 4023 15899 4029
rect 17034 4020 17040 4032
rect 17092 4020 17098 4072
rect 17144 4060 17172 4100
rect 17681 4097 17693 4131
rect 17727 4128 17739 4131
rect 17865 4131 17923 4137
rect 17727 4100 17816 4128
rect 17727 4097 17739 4100
rect 17681 4091 17739 4097
rect 17788 4060 17816 4100
rect 17865 4097 17877 4131
rect 17911 4128 17923 4131
rect 17972 4128 18000 4168
rect 18230 4156 18236 4168
rect 18288 4156 18294 4208
rect 17911 4100 18000 4128
rect 18049 4131 18107 4137
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 18049 4097 18061 4131
rect 18095 4128 18107 4131
rect 18095 4100 18368 4128
rect 18095 4097 18107 4100
rect 18049 4091 18107 4097
rect 18138 4060 18144 4072
rect 17144 4032 17724 4060
rect 17788 4032 18144 4060
rect 13964 3964 15056 3992
rect 15289 3995 15347 4001
rect 13964 3952 13970 3964
rect 15289 3961 15301 3995
rect 15335 3992 15347 3995
rect 15378 3992 15384 4004
rect 15335 3964 15384 3992
rect 15335 3961 15347 3964
rect 15289 3955 15347 3961
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 17696 4001 17724 4032
rect 18138 4020 18144 4032
rect 18196 4020 18202 4072
rect 17681 3995 17739 4001
rect 17681 3961 17693 3995
rect 17727 3961 17739 3995
rect 17681 3955 17739 3961
rect 18340 3936 18368 4100
rect 18506 4088 18512 4140
rect 18564 4128 18570 4140
rect 19168 4137 19196 4236
rect 19334 4224 19340 4236
rect 19392 4224 19398 4276
rect 19610 4224 19616 4276
rect 19668 4264 19674 4276
rect 20533 4267 20591 4273
rect 20533 4264 20545 4267
rect 19668 4236 20545 4264
rect 19668 4224 19674 4236
rect 20533 4233 20545 4236
rect 20579 4233 20591 4267
rect 24394 4264 24400 4276
rect 20533 4227 20591 4233
rect 21008 4236 24400 4264
rect 19420 4199 19478 4205
rect 19420 4165 19432 4199
rect 19466 4196 19478 4199
rect 20438 4196 20444 4208
rect 19466 4168 20444 4196
rect 19466 4165 19478 4168
rect 19420 4159 19478 4165
rect 20438 4156 20444 4168
rect 20496 4156 20502 4208
rect 21008 4205 21036 4236
rect 24394 4224 24400 4236
rect 24452 4224 24458 4276
rect 20993 4199 21051 4205
rect 20993 4165 21005 4199
rect 21039 4165 21051 4199
rect 20993 4159 21051 4165
rect 22020 4168 22232 4196
rect 19061 4131 19119 4137
rect 19061 4128 19073 4131
rect 18564 4100 19073 4128
rect 18564 4088 18570 4100
rect 19061 4097 19073 4100
rect 19107 4097 19119 4131
rect 19061 4091 19119 4097
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4097 19211 4131
rect 19153 4091 19211 4097
rect 19794 4088 19800 4140
rect 19852 4128 19858 4140
rect 20809 4131 20867 4137
rect 20809 4128 20821 4131
rect 19852 4100 20821 4128
rect 19852 4088 19858 4100
rect 20809 4097 20821 4100
rect 20855 4097 20867 4131
rect 20809 4091 20867 4097
rect 21453 4131 21511 4137
rect 21453 4097 21465 4131
rect 21499 4128 21511 4131
rect 21542 4128 21548 4140
rect 21499 4100 21548 4128
rect 21499 4097 21511 4100
rect 21453 4091 21511 4097
rect 21542 4088 21548 4100
rect 21600 4088 21606 4140
rect 22020 4128 22048 4168
rect 21836 4100 22048 4128
rect 20438 4020 20444 4072
rect 20496 4060 20502 4072
rect 21836 4069 21864 4100
rect 22094 4088 22100 4140
rect 22152 4088 22158 4140
rect 22204 4128 22232 4168
rect 23201 4131 23259 4137
rect 23201 4128 23213 4131
rect 22204 4100 23213 4128
rect 23201 4097 23213 4100
rect 23247 4097 23259 4131
rect 23201 4091 23259 4097
rect 23475 4131 23533 4137
rect 23475 4097 23487 4131
rect 23521 4128 23533 4131
rect 25682 4128 25688 4140
rect 23521 4100 25688 4128
rect 23521 4097 23533 4100
rect 23475 4091 23533 4097
rect 25682 4088 25688 4100
rect 25740 4088 25746 4140
rect 21821 4063 21879 4069
rect 21821 4060 21833 4063
rect 20496 4032 21833 4060
rect 20496 4020 20502 4032
rect 21821 4029 21833 4032
rect 21867 4029 21879 4063
rect 21821 4023 21879 4029
rect 24210 4020 24216 4072
rect 24268 4020 24274 4072
rect 20162 3952 20168 4004
rect 20220 3992 20226 4004
rect 20625 3995 20683 4001
rect 20625 3992 20637 3995
rect 20220 3964 20637 3992
rect 20220 3952 20226 3964
rect 20625 3961 20637 3964
rect 20671 3961 20683 3995
rect 20625 3955 20683 3961
rect 8570 3924 8576 3936
rect 8312 3896 8576 3924
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 12066 3924 12072 3936
rect 9548 3896 12072 3924
rect 9548 3884 9554 3896
rect 12066 3884 12072 3896
rect 12124 3884 12130 3936
rect 14458 3884 14464 3936
rect 14516 3924 14522 3936
rect 16485 3927 16543 3933
rect 16485 3924 16497 3927
rect 14516 3896 16497 3924
rect 14516 3884 14522 3896
rect 16485 3893 16497 3896
rect 16531 3893 16543 3927
rect 16485 3887 16543 3893
rect 18322 3884 18328 3936
rect 18380 3884 18386 3936
rect 18874 3884 18880 3936
rect 18932 3884 18938 3936
rect 19150 3884 19156 3936
rect 19208 3924 19214 3936
rect 20990 3924 20996 3936
rect 19208 3896 20996 3924
rect 19208 3884 19214 3896
rect 20990 3884 20996 3896
rect 21048 3884 21054 3936
rect 21085 3927 21143 3933
rect 21085 3893 21097 3927
rect 21131 3924 21143 3927
rect 21174 3924 21180 3936
rect 21131 3896 21180 3924
rect 21131 3893 21143 3896
rect 21085 3887 21143 3893
rect 21174 3884 21180 3896
rect 21232 3884 21238 3936
rect 21450 3884 21456 3936
rect 21508 3924 21514 3936
rect 21545 3927 21603 3933
rect 21545 3924 21557 3927
rect 21508 3896 21557 3924
rect 21508 3884 21514 3896
rect 21545 3893 21557 3896
rect 21591 3893 21603 3927
rect 21545 3887 21603 3893
rect 22278 3884 22284 3936
rect 22336 3924 22342 3936
rect 24228 3933 24256 4020
rect 22833 3927 22891 3933
rect 22833 3924 22845 3927
rect 22336 3896 22845 3924
rect 22336 3884 22342 3896
rect 22833 3893 22845 3896
rect 22879 3893 22891 3927
rect 22833 3887 22891 3893
rect 24213 3927 24271 3933
rect 24213 3893 24225 3927
rect 24259 3893 24271 3927
rect 24213 3887 24271 3893
rect 1104 3834 24840 3856
rect 1104 3782 3917 3834
rect 3969 3782 3981 3834
rect 4033 3782 4045 3834
rect 4097 3782 4109 3834
rect 4161 3782 4173 3834
rect 4225 3782 9851 3834
rect 9903 3782 9915 3834
rect 9967 3782 9979 3834
rect 10031 3782 10043 3834
rect 10095 3782 10107 3834
rect 10159 3782 15785 3834
rect 15837 3782 15849 3834
rect 15901 3782 15913 3834
rect 15965 3782 15977 3834
rect 16029 3782 16041 3834
rect 16093 3782 21719 3834
rect 21771 3782 21783 3834
rect 21835 3782 21847 3834
rect 21899 3782 21911 3834
rect 21963 3782 21975 3834
rect 22027 3782 24840 3834
rect 1104 3760 24840 3782
rect 1397 3723 1455 3729
rect 1397 3689 1409 3723
rect 1443 3720 1455 3723
rect 1486 3720 1492 3732
rect 1443 3692 1492 3720
rect 1443 3689 1455 3692
rect 1397 3683 1455 3689
rect 1486 3680 1492 3692
rect 1544 3680 1550 3732
rect 2406 3680 2412 3732
rect 2464 3720 2470 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2464 3692 2697 3720
rect 2464 3680 2470 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 4522 3680 4528 3732
rect 4580 3720 4586 3732
rect 4801 3723 4859 3729
rect 4801 3720 4813 3723
rect 4580 3692 4813 3720
rect 4580 3680 4586 3692
rect 4801 3689 4813 3692
rect 4847 3689 4859 3723
rect 4801 3683 4859 3689
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 5902 3720 5908 3732
rect 5224 3692 5908 3720
rect 5224 3680 5230 3692
rect 5902 3680 5908 3692
rect 5960 3680 5966 3732
rect 7101 3723 7159 3729
rect 6104 3692 6776 3720
rect 6104 3593 6132 3692
rect 6748 3652 6776 3692
rect 7101 3689 7113 3723
rect 7147 3720 7159 3723
rect 8202 3720 8208 3732
rect 7147 3692 8208 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 14458 3720 14464 3732
rect 8352 3692 14464 3720
rect 8352 3680 8358 3692
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 14660 3692 15332 3720
rect 13262 3652 13268 3664
rect 6748 3624 7328 3652
rect 7300 3596 7328 3624
rect 11716 3624 13268 3652
rect 6089 3587 6147 3593
rect 6089 3553 6101 3587
rect 6135 3553 6147 3587
rect 6089 3547 6147 3553
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 7469 3587 7527 3593
rect 7469 3584 7481 3587
rect 7340 3556 7481 3584
rect 7340 3544 7346 3556
rect 7469 3553 7481 3556
rect 7515 3553 7527 3587
rect 7469 3547 7527 3553
rect 8864 3556 9536 3584
rect 1578 3476 1584 3528
rect 1636 3476 1642 3528
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 1854 3516 1860 3528
rect 1719 3488 1860 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 1854 3476 1860 3488
rect 1912 3476 1918 3528
rect 1947 3519 2005 3525
rect 1947 3485 1959 3519
rect 1993 3516 2005 3519
rect 2958 3516 2964 3528
rect 1993 3488 2964 3516
rect 1993 3485 2005 3488
rect 1947 3479 2005 3485
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 4063 3519 4121 3525
rect 4063 3485 4075 3519
rect 4109 3516 4121 3519
rect 6363 3519 6421 3525
rect 4109 3488 6040 3516
rect 4109 3485 4121 3488
rect 4063 3479 4121 3485
rect 1872 3448 1900 3476
rect 3804 3448 3832 3479
rect 1872 3420 3832 3448
rect 6012 3448 6040 3488
rect 6363 3485 6375 3519
rect 6409 3516 6421 3519
rect 6730 3516 6736 3528
rect 6409 3488 6736 3516
rect 6409 3485 6421 3488
rect 6363 3479 6421 3485
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 7743 3519 7801 3525
rect 7743 3485 7755 3519
rect 7789 3516 7801 3519
rect 8864 3516 8892 3556
rect 9508 3528 9536 3556
rect 9766 3544 9772 3596
rect 9824 3544 9830 3596
rect 7789 3488 8892 3516
rect 7789 3485 7801 3488
rect 7743 3479 7801 3485
rect 9122 3476 9128 3528
rect 9180 3476 9186 3528
rect 9490 3476 9496 3528
rect 9548 3476 9554 3528
rect 10043 3519 10101 3525
rect 10043 3485 10055 3519
rect 10089 3516 10101 3519
rect 11054 3516 11060 3528
rect 10089 3488 11060 3516
rect 10089 3485 10101 3488
rect 10043 3479 10101 3485
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 11716 3525 11744 3624
rect 13262 3612 13268 3624
rect 13320 3612 13326 3664
rect 13906 3612 13912 3664
rect 13964 3612 13970 3664
rect 12437 3587 12495 3593
rect 12437 3553 12449 3587
rect 12483 3584 12495 3587
rect 12710 3584 12716 3596
rect 12483 3556 12716 3584
rect 12483 3553 12495 3556
rect 12437 3547 12495 3553
rect 12710 3544 12716 3556
rect 12768 3544 12774 3596
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11204 3488 11713 3516
rect 11204 3476 11210 3488
rect 11701 3485 11713 3488
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 11974 3476 11980 3528
rect 12032 3516 12038 3528
rect 13357 3519 13415 3525
rect 13357 3516 13369 3519
rect 12032 3488 13369 3516
rect 12032 3476 12038 3488
rect 13357 3485 13369 3488
rect 13403 3516 13415 3519
rect 13817 3519 13875 3525
rect 13817 3516 13829 3519
rect 13403 3488 13829 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 13817 3485 13829 3488
rect 13863 3516 13875 3519
rect 13924 3516 13952 3612
rect 14660 3593 14688 3692
rect 15304 3652 15332 3692
rect 15378 3680 15384 3732
rect 15436 3720 15442 3732
rect 15657 3723 15715 3729
rect 15657 3720 15669 3723
rect 15436 3692 15669 3720
rect 15436 3680 15442 3692
rect 15657 3689 15669 3692
rect 15703 3689 15715 3723
rect 15657 3683 15715 3689
rect 16114 3680 16120 3732
rect 16172 3680 16178 3732
rect 17034 3680 17040 3732
rect 17092 3680 17098 3732
rect 18322 3680 18328 3732
rect 18380 3680 18386 3732
rect 19306 3692 20668 3720
rect 16132 3652 16160 3680
rect 19306 3652 19334 3692
rect 15304 3624 16160 3652
rect 17788 3624 19334 3652
rect 19435 3624 20300 3652
rect 16040 3593 16068 3624
rect 14645 3587 14703 3593
rect 14645 3553 14657 3587
rect 14691 3553 14703 3587
rect 14645 3547 14703 3553
rect 16025 3587 16083 3593
rect 16025 3553 16037 3587
rect 16071 3553 16083 3587
rect 16025 3547 16083 3553
rect 13863 3488 13952 3516
rect 13863 3485 13875 3488
rect 13817 3479 13875 3485
rect 14918 3476 14924 3528
rect 14976 3476 14982 3528
rect 16390 3516 16396 3528
rect 15672 3489 16396 3516
rect 15672 3488 16295 3489
rect 8386 3448 8392 3460
rect 6012 3420 8392 3448
rect 8386 3408 8392 3420
rect 8444 3408 8450 3460
rect 8570 3408 8576 3460
rect 8628 3448 8634 3460
rect 8628 3420 11744 3448
rect 8628 3408 8634 3420
rect 8481 3383 8539 3389
rect 8481 3349 8493 3383
rect 8527 3380 8539 3383
rect 8754 3380 8760 3392
rect 8527 3352 8760 3380
rect 8527 3349 8539 3352
rect 8481 3343 8539 3349
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 8938 3340 8944 3392
rect 8996 3340 9002 3392
rect 10226 3340 10232 3392
rect 10284 3380 10290 3392
rect 10781 3383 10839 3389
rect 10781 3380 10793 3383
rect 10284 3352 10793 3380
rect 10284 3340 10290 3352
rect 10781 3349 10793 3352
rect 10827 3349 10839 3383
rect 10781 3343 10839 3349
rect 11514 3340 11520 3392
rect 11572 3340 11578 3392
rect 11716 3380 11744 3420
rect 11790 3408 11796 3460
rect 11848 3448 11854 3460
rect 15562 3448 15568 3460
rect 11848 3420 15568 3448
rect 11848 3408 11854 3420
rect 15562 3408 15568 3420
rect 15620 3408 15626 3460
rect 13446 3380 13452 3392
rect 11716 3352 13452 3380
rect 13446 3340 13452 3352
rect 13504 3340 13510 3392
rect 13633 3383 13691 3389
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 13814 3380 13820 3392
rect 13679 3352 13820 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 13906 3340 13912 3392
rect 13964 3380 13970 3392
rect 15672 3380 15700 3488
rect 16283 3455 16295 3488
rect 16329 3488 16396 3489
rect 16329 3458 16342 3488
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 17586 3476 17592 3528
rect 17644 3516 17650 3528
rect 17788 3525 17816 3624
rect 18138 3544 18144 3596
rect 18196 3584 18202 3596
rect 18601 3587 18659 3593
rect 18601 3584 18613 3587
rect 18196 3556 18613 3584
rect 18196 3544 18202 3556
rect 18601 3553 18613 3556
rect 18647 3553 18659 3587
rect 18601 3547 18659 3553
rect 18874 3544 18880 3596
rect 18932 3584 18938 3596
rect 19435 3584 19463 3624
rect 19886 3584 19892 3596
rect 18932 3556 19463 3584
rect 19536 3556 19892 3584
rect 18932 3544 18938 3556
rect 17681 3519 17739 3525
rect 17681 3516 17693 3519
rect 17644 3488 17693 3516
rect 17644 3476 17650 3488
rect 17681 3485 17693 3488
rect 17727 3485 17739 3519
rect 17681 3479 17739 3485
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3485 17831 3519
rect 17773 3479 17831 3485
rect 17957 3519 18015 3525
rect 17957 3485 17969 3519
rect 18003 3485 18015 3519
rect 17957 3479 18015 3485
rect 16329 3455 16341 3458
rect 16283 3449 16341 3455
rect 17126 3408 17132 3460
rect 17184 3448 17190 3460
rect 17184 3420 17632 3448
rect 17184 3408 17190 3420
rect 13964 3352 15700 3380
rect 13964 3340 13970 3352
rect 17494 3340 17500 3392
rect 17552 3340 17558 3392
rect 17604 3380 17632 3420
rect 17862 3408 17868 3460
rect 17920 3408 17926 3460
rect 17972 3380 18000 3479
rect 18230 3476 18236 3528
rect 18288 3476 18294 3528
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 18432 3448 18460 3479
rect 18506 3476 18512 3528
rect 18564 3476 18570 3528
rect 18969 3519 19027 3525
rect 18969 3485 18981 3519
rect 19015 3516 19027 3519
rect 19242 3516 19248 3528
rect 19015 3488 19248 3516
rect 19015 3485 19027 3488
rect 18969 3479 19027 3485
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3516 19487 3519
rect 19536 3516 19564 3556
rect 19886 3544 19892 3556
rect 19944 3544 19950 3596
rect 20162 3544 20168 3596
rect 20220 3544 20226 3596
rect 20180 3516 20208 3544
rect 20272 3525 20300 3624
rect 19475 3488 19564 3516
rect 19628 3488 20208 3516
rect 20257 3519 20315 3525
rect 19475 3485 19487 3488
rect 19429 3479 19487 3485
rect 19628 3448 19656 3488
rect 20257 3485 20269 3519
rect 20303 3485 20315 3519
rect 20640 3516 20668 3692
rect 22462 3680 22468 3732
rect 22520 3720 22526 3732
rect 25590 3720 25596 3732
rect 22520 3692 25596 3720
rect 22520 3680 22526 3692
rect 25590 3680 25596 3692
rect 25648 3680 25654 3732
rect 21358 3612 21364 3664
rect 21416 3652 21422 3664
rect 22646 3652 22652 3664
rect 21416 3624 22652 3652
rect 21416 3612 21422 3624
rect 22646 3612 22652 3624
rect 22704 3612 22710 3664
rect 23566 3612 23572 3664
rect 23624 3652 23630 3664
rect 23937 3655 23995 3661
rect 23937 3652 23949 3655
rect 23624 3624 23949 3652
rect 23624 3612 23630 3624
rect 23937 3621 23949 3624
rect 23983 3621 23995 3655
rect 23937 3615 23995 3621
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 22189 3587 22247 3593
rect 22189 3584 22201 3587
rect 20772 3556 22201 3584
rect 20772 3544 20778 3556
rect 22189 3553 22201 3556
rect 22235 3553 22247 3587
rect 22189 3547 22247 3553
rect 22278 3544 22284 3596
rect 22336 3544 22342 3596
rect 23014 3544 23020 3596
rect 23072 3544 23078 3596
rect 21453 3519 21511 3525
rect 21453 3516 21465 3519
rect 20640 3488 21465 3516
rect 20257 3479 20315 3485
rect 21453 3485 21465 3488
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 18432 3420 19656 3448
rect 19702 3408 19708 3460
rect 19760 3408 19766 3460
rect 19886 3408 19892 3460
rect 19944 3448 19950 3460
rect 20809 3451 20867 3457
rect 19944 3420 20484 3448
rect 19944 3408 19950 3420
rect 17604 3352 18000 3380
rect 18598 3340 18604 3392
rect 18656 3380 18662 3392
rect 18785 3383 18843 3389
rect 18785 3380 18797 3383
rect 18656 3352 18797 3380
rect 18656 3340 18662 3352
rect 18785 3349 18797 3352
rect 18831 3349 18843 3383
rect 18785 3343 18843 3349
rect 19242 3340 19248 3392
rect 19300 3340 19306 3392
rect 19518 3340 19524 3392
rect 19576 3380 19582 3392
rect 19797 3383 19855 3389
rect 19797 3380 19809 3383
rect 19576 3352 19809 3380
rect 19576 3340 19582 3352
rect 19797 3349 19809 3352
rect 19843 3349 19855 3383
rect 19797 3343 19855 3349
rect 20162 3340 20168 3392
rect 20220 3380 20226 3392
rect 20349 3383 20407 3389
rect 20349 3380 20361 3383
rect 20220 3352 20361 3380
rect 20220 3340 20226 3352
rect 20349 3349 20361 3352
rect 20395 3349 20407 3383
rect 20456 3380 20484 3420
rect 20809 3417 20821 3451
rect 20855 3448 20867 3451
rect 20990 3448 20996 3460
rect 20855 3420 20996 3448
rect 20855 3417 20867 3420
rect 20809 3411 20867 3417
rect 20990 3408 20996 3420
rect 21048 3408 21054 3460
rect 21468 3448 21496 3479
rect 21634 3476 21640 3528
rect 21692 3476 21698 3528
rect 22094 3476 22100 3528
rect 22152 3476 22158 3528
rect 22296 3448 22324 3544
rect 22646 3476 22652 3528
rect 22704 3476 22710 3528
rect 23106 3476 23112 3528
rect 23164 3516 23170 3528
rect 23753 3519 23811 3525
rect 23753 3516 23765 3519
rect 23164 3488 23765 3516
rect 23164 3476 23170 3488
rect 23753 3485 23765 3488
rect 23799 3485 23811 3519
rect 23753 3479 23811 3485
rect 21468 3420 22324 3448
rect 20901 3383 20959 3389
rect 20901 3380 20913 3383
rect 20456 3352 20913 3380
rect 20349 3343 20407 3349
rect 20901 3349 20913 3352
rect 20947 3349 20959 3383
rect 20901 3343 20959 3349
rect 1104 3290 25000 3312
rect 1104 3238 6884 3290
rect 6936 3238 6948 3290
rect 7000 3238 7012 3290
rect 7064 3238 7076 3290
rect 7128 3238 7140 3290
rect 7192 3238 12818 3290
rect 12870 3238 12882 3290
rect 12934 3238 12946 3290
rect 12998 3238 13010 3290
rect 13062 3238 13074 3290
rect 13126 3238 18752 3290
rect 18804 3238 18816 3290
rect 18868 3238 18880 3290
rect 18932 3238 18944 3290
rect 18996 3238 19008 3290
rect 19060 3238 24686 3290
rect 24738 3238 24750 3290
rect 24802 3238 24814 3290
rect 24866 3238 24878 3290
rect 24930 3238 24942 3290
rect 24994 3238 25000 3290
rect 1104 3216 25000 3238
rect 1578 3136 1584 3188
rect 1636 3176 1642 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 1636 3148 9413 3176
rect 1636 3136 1642 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9401 3139 9459 3145
rect 9861 3179 9919 3185
rect 9861 3145 9873 3179
rect 9907 3176 9919 3179
rect 11146 3176 11152 3188
rect 9907 3148 11152 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 11514 3136 11520 3188
rect 11572 3136 11578 3188
rect 12526 3136 12532 3188
rect 12584 3176 12590 3188
rect 13265 3179 13323 3185
rect 13265 3176 13277 3179
rect 12584 3148 13277 3176
rect 12584 3136 12590 3148
rect 13265 3145 13277 3148
rect 13311 3145 13323 3179
rect 13265 3139 13323 3145
rect 14366 3136 14372 3188
rect 14424 3136 14430 3188
rect 17773 3179 17831 3185
rect 16500 3148 17540 3176
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 2961 3111 3019 3117
rect 2961 3108 2973 3111
rect 2004 3080 2973 3108
rect 2004 3068 2010 3080
rect 2961 3077 2973 3080
rect 3007 3108 3019 3111
rect 4338 3108 4344 3120
rect 3007 3080 4344 3108
rect 3007 3077 3019 3080
rect 2961 3071 3019 3077
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 4430 3068 4436 3120
rect 4488 3068 4494 3120
rect 5151 3073 5209 3079
rect 5151 3039 5163 3073
rect 5197 3040 5209 3073
rect 6178 3068 6184 3120
rect 6236 3108 6242 3120
rect 6236 3080 6960 3108
rect 6236 3068 6242 3080
rect 5197 3039 6592 3040
rect 5151 3033 6592 3039
rect 5166 3012 6592 3033
rect 566 2932 572 2984
rect 624 2972 630 2984
rect 3145 2975 3203 2981
rect 3145 2972 3157 2975
rect 624 2944 3157 2972
rect 624 2932 630 2944
rect 3145 2941 3157 2944
rect 3191 2941 3203 2975
rect 3145 2935 3203 2941
rect 4614 2932 4620 2984
rect 4672 2932 4678 2984
rect 4890 2932 4896 2984
rect 4948 2932 4954 2984
rect 6564 2972 6592 3012
rect 6638 3000 6644 3052
rect 6696 3000 6702 3052
rect 6932 3049 6960 3080
rect 10134 3068 10140 3120
rect 10192 3068 10198 3120
rect 10226 3068 10232 3120
rect 10284 3068 10290 3120
rect 10410 3068 10416 3120
rect 10468 3108 10474 3120
rect 10597 3111 10655 3117
rect 10597 3108 10609 3111
rect 10468 3080 10609 3108
rect 10468 3068 10474 3080
rect 10597 3077 10609 3080
rect 10643 3077 10655 3111
rect 10597 3071 10655 3077
rect 10965 3111 11023 3117
rect 10965 3077 10977 3111
rect 11011 3077 11023 3111
rect 10965 3071 11023 3077
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7190 3000 7196 3052
rect 7248 3000 7254 3052
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 7607 3012 7880 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 7484 2972 7512 3003
rect 7852 2984 7880 3012
rect 8478 3000 8484 3052
rect 8536 3000 8542 3052
rect 8662 3049 8668 3052
rect 8619 3043 8668 3049
rect 8619 3009 8631 3043
rect 8665 3009 8668 3043
rect 8619 3003 8668 3009
rect 8662 3000 8668 3003
rect 8720 3000 8726 3052
rect 8754 3000 8760 3052
rect 8812 3000 8818 3052
rect 9398 3000 9404 3052
rect 9456 3040 9462 3052
rect 10980 3040 11008 3071
rect 9456 3012 11008 3040
rect 11532 3040 11560 3136
rect 11606 3068 11612 3120
rect 11664 3108 11670 3120
rect 11664 3080 12020 3108
rect 11664 3068 11670 3080
rect 11885 3043 11943 3049
rect 11885 3040 11897 3043
rect 11532 3012 11897 3040
rect 9456 3000 9462 3012
rect 11885 3009 11897 3012
rect 11931 3009 11943 3043
rect 11885 3003 11943 3009
rect 7650 2972 7656 2984
rect 6564 2944 7420 2972
rect 7484 2944 7656 2972
rect 6546 2864 6552 2916
rect 6604 2904 6610 2916
rect 6604 2876 7052 2904
rect 6604 2864 6610 2876
rect 5350 2796 5356 2848
rect 5408 2836 5414 2848
rect 5905 2839 5963 2845
rect 5905 2836 5917 2839
rect 5408 2808 5917 2836
rect 5408 2796 5414 2808
rect 5905 2805 5917 2808
rect 5951 2805 5963 2839
rect 5905 2799 5963 2805
rect 6454 2796 6460 2848
rect 6512 2796 6518 2848
rect 6730 2796 6736 2848
rect 6788 2796 6794 2848
rect 7024 2845 7052 2876
rect 7009 2839 7067 2845
rect 7009 2805 7021 2839
rect 7055 2805 7067 2839
rect 7009 2799 7067 2805
rect 7282 2796 7288 2848
rect 7340 2796 7346 2848
rect 7392 2836 7420 2944
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 7745 2975 7803 2981
rect 7745 2941 7757 2975
rect 7791 2941 7803 2975
rect 7745 2935 7803 2941
rect 7760 2904 7788 2935
rect 7834 2932 7840 2984
rect 7892 2932 7898 2984
rect 8110 2932 8116 2984
rect 8168 2932 8174 2984
rect 10226 2932 10232 2984
rect 10284 2932 10290 2984
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11992 2972 12020 3080
rect 12066 3068 12072 3120
rect 12124 3108 12130 3120
rect 14384 3108 14412 3136
rect 12124 3080 12388 3108
rect 12124 3068 12130 3080
rect 12158 3000 12164 3052
rect 12216 3000 12222 3052
rect 12360 3040 12388 3080
rect 12820 3080 14412 3108
rect 12527 3043 12585 3049
rect 12527 3040 12539 3043
rect 12360 3012 12539 3040
rect 12527 3009 12539 3012
rect 12573 3040 12585 3043
rect 12820 3040 12848 3080
rect 12573 3012 12848 3040
rect 12573 3009 12585 3012
rect 12527 3003 12585 3009
rect 12894 3000 12900 3052
rect 12952 3040 12958 3052
rect 13722 3040 13728 3052
rect 12952 3012 13728 3040
rect 12952 3000 12958 3012
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 16298 3000 16304 3052
rect 16356 3000 16362 3052
rect 16500 3049 16528 3148
rect 17034 3068 17040 3120
rect 17092 3108 17098 3120
rect 17512 3108 17540 3148
rect 17773 3145 17785 3179
rect 17819 3176 17831 3179
rect 18506 3176 18512 3188
rect 17819 3148 18512 3176
rect 17819 3145 17831 3148
rect 17773 3139 17831 3145
rect 18506 3136 18512 3148
rect 18564 3136 18570 3188
rect 19334 3136 19340 3188
rect 19392 3136 19398 3188
rect 19426 3136 19432 3188
rect 19484 3136 19490 3188
rect 19705 3179 19763 3185
rect 19705 3176 19717 3179
rect 19527 3148 19717 3176
rect 17092 3080 17448 3108
rect 17512 3080 17908 3108
rect 17092 3068 17098 3080
rect 16485 3043 16543 3049
rect 16485 3009 16497 3043
rect 16531 3009 16543 3043
rect 16485 3003 16543 3009
rect 16850 3000 16856 3052
rect 16908 3000 16914 3052
rect 17420 3049 17448 3080
rect 17880 3052 17908 3080
rect 18230 3068 18236 3120
rect 18288 3108 18294 3120
rect 19352 3108 19380 3136
rect 19527 3108 19555 3148
rect 19705 3145 19717 3148
rect 19751 3145 19763 3179
rect 19705 3139 19763 3145
rect 18288 3080 19380 3108
rect 19435 3080 19555 3108
rect 18288 3068 18294 3080
rect 17129 3043 17187 3049
rect 17129 3009 17141 3043
rect 17175 3009 17187 3043
rect 17129 3003 17187 3009
rect 17405 3043 17463 3049
rect 17405 3009 17417 3043
rect 17451 3009 17463 3043
rect 17405 3003 17463 3009
rect 12253 2975 12311 2981
rect 12253 2972 12265 2975
rect 11020 2944 11744 2972
rect 11992 2944 12265 2972
rect 11020 2932 11026 2944
rect 8128 2904 8156 2932
rect 7760 2876 8156 2904
rect 8202 2864 8208 2916
rect 8260 2864 8266 2916
rect 9306 2864 9312 2916
rect 9364 2864 9370 2916
rect 11054 2864 11060 2916
rect 11112 2904 11118 2916
rect 11149 2907 11207 2913
rect 11149 2904 11161 2907
rect 11112 2876 11161 2904
rect 11112 2864 11118 2876
rect 11149 2873 11161 2876
rect 11195 2873 11207 2907
rect 11149 2867 11207 2873
rect 9324 2836 9352 2864
rect 11716 2845 11744 2944
rect 12253 2941 12265 2944
rect 12299 2941 12311 2975
rect 17144 2972 17172 3003
rect 17678 3000 17684 3052
rect 17736 3000 17742 3052
rect 17862 3000 17868 3052
rect 17920 3000 17926 3052
rect 17957 3043 18015 3049
rect 17957 3009 17969 3043
rect 18003 3038 18015 3043
rect 18316 3043 18374 3049
rect 18316 3040 18328 3043
rect 18156 3038 18328 3040
rect 18003 3012 18328 3038
rect 18003 3010 18184 3012
rect 18003 3009 18015 3010
rect 17957 3003 18015 3009
rect 18316 3009 18328 3012
rect 18362 3040 18374 3043
rect 19334 3040 19340 3052
rect 18362 3012 19340 3040
rect 18362 3009 18374 3012
rect 19306 3010 19340 3012
rect 18316 3003 18374 3009
rect 19334 3000 19340 3010
rect 19392 3000 19398 3052
rect 18049 2975 18107 2981
rect 17144 2944 18000 2972
rect 12253 2935 12311 2941
rect 7392 2808 9352 2836
rect 11701 2839 11759 2845
rect 11701 2805 11713 2839
rect 11747 2805 11759 2839
rect 11701 2799 11759 2805
rect 11790 2796 11796 2848
rect 11848 2836 11854 2848
rect 11977 2839 12035 2845
rect 11977 2836 11989 2839
rect 11848 2808 11989 2836
rect 11848 2796 11854 2808
rect 11977 2805 11989 2808
rect 12023 2805 12035 2839
rect 12268 2836 12296 2935
rect 17972 2916 18000 2944
rect 18049 2941 18061 2975
rect 18095 2941 18107 2975
rect 19435 2972 19463 3080
rect 19610 3068 19616 3120
rect 19668 3068 19674 3120
rect 20165 3111 20223 3117
rect 20165 3077 20177 3111
rect 20211 3108 20223 3111
rect 22738 3108 22744 3120
rect 20211 3080 22744 3108
rect 20211 3077 20223 3080
rect 20165 3071 20223 3077
rect 22738 3068 22744 3080
rect 22796 3068 22802 3120
rect 22830 3068 22836 3120
rect 22888 3068 22894 3120
rect 23014 3068 23020 3120
rect 23072 3108 23078 3120
rect 23376 3111 23434 3117
rect 23376 3108 23388 3111
rect 23072 3080 23388 3108
rect 23072 3068 23078 3080
rect 23376 3077 23388 3080
rect 23422 3108 23434 3111
rect 24118 3108 24124 3120
rect 23422 3080 24124 3108
rect 23422 3077 23434 3080
rect 23376 3071 23434 3077
rect 24118 3068 24124 3080
rect 24176 3068 24182 3120
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 21634 3040 21640 3052
rect 20855 3012 21640 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 21634 3000 21640 3012
rect 21692 3000 21698 3052
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3040 22247 3043
rect 22278 3040 22284 3052
rect 22235 3012 22284 3040
rect 22235 3009 22247 3012
rect 22189 3003 22247 3009
rect 22278 3000 22284 3012
rect 22336 3000 22342 3052
rect 18049 2935 18107 2941
rect 19306 2944 19463 2972
rect 17310 2904 17316 2916
rect 16960 2876 17316 2904
rect 14366 2836 14372 2848
rect 12268 2808 14372 2836
rect 11977 2799 12035 2805
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 16393 2839 16451 2845
rect 16393 2805 16405 2839
rect 16439 2836 16451 2839
rect 16574 2836 16580 2848
rect 16439 2808 16580 2836
rect 16439 2805 16451 2808
rect 16393 2799 16451 2805
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 16669 2839 16727 2845
rect 16669 2805 16681 2839
rect 16715 2836 16727 2839
rect 16850 2836 16856 2848
rect 16715 2808 16856 2836
rect 16715 2805 16727 2808
rect 16669 2799 16727 2805
rect 16850 2796 16856 2808
rect 16908 2796 16914 2848
rect 16960 2845 16988 2876
rect 17310 2864 17316 2876
rect 17368 2864 17374 2916
rect 17954 2864 17960 2916
rect 18012 2864 18018 2916
rect 16945 2839 17003 2845
rect 16945 2805 16957 2839
rect 16991 2805 17003 2839
rect 16945 2799 17003 2805
rect 17218 2796 17224 2848
rect 17276 2796 17282 2848
rect 17497 2839 17555 2845
rect 17497 2805 17509 2839
rect 17543 2836 17555 2839
rect 17678 2836 17684 2848
rect 17543 2808 17684 2836
rect 17543 2805 17555 2808
rect 17497 2799 17555 2805
rect 17678 2796 17684 2808
rect 17736 2796 17742 2848
rect 18064 2836 18092 2935
rect 19150 2864 19156 2916
rect 19208 2904 19214 2916
rect 19306 2904 19334 2944
rect 19702 2932 19708 2984
rect 19760 2972 19766 2984
rect 20898 2972 20904 2984
rect 19760 2944 20904 2972
rect 19760 2932 19766 2944
rect 20898 2932 20904 2944
rect 20956 2932 20962 2984
rect 20993 2975 21051 2981
rect 20993 2941 21005 2975
rect 21039 2941 21051 2975
rect 20993 2935 21051 2941
rect 19208 2876 19334 2904
rect 19208 2864 19214 2876
rect 19978 2864 19984 2916
rect 20036 2904 20042 2916
rect 20036 2876 20383 2904
rect 20036 2864 20042 2876
rect 18230 2836 18236 2848
rect 18064 2808 18236 2836
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 18414 2796 18420 2848
rect 18472 2836 18478 2848
rect 19518 2836 19524 2848
rect 18472 2808 19524 2836
rect 18472 2796 18478 2808
rect 19518 2796 19524 2808
rect 19576 2796 19582 2848
rect 19794 2796 19800 2848
rect 19852 2836 19858 2848
rect 20257 2839 20315 2845
rect 20257 2836 20269 2839
rect 19852 2808 20269 2836
rect 19852 2796 19858 2808
rect 20257 2805 20269 2808
rect 20303 2805 20315 2839
rect 20355 2836 20383 2876
rect 20714 2864 20720 2916
rect 20772 2904 20778 2916
rect 21008 2904 21036 2935
rect 22462 2932 22468 2984
rect 22520 2972 22526 2984
rect 23109 2975 23167 2981
rect 23109 2972 23121 2975
rect 22520 2944 23121 2972
rect 22520 2932 22526 2944
rect 23109 2941 23121 2944
rect 23155 2941 23167 2975
rect 23109 2935 23167 2941
rect 20772 2876 21036 2904
rect 20772 2864 20778 2876
rect 21266 2836 21272 2848
rect 20355 2808 21272 2836
rect 20257 2799 20315 2805
rect 21266 2796 21272 2808
rect 21324 2796 21330 2848
rect 21542 2796 21548 2848
rect 21600 2836 21606 2848
rect 24210 2836 24216 2848
rect 21600 2808 24216 2836
rect 21600 2796 21606 2808
rect 24210 2796 24216 2808
rect 24268 2796 24274 2848
rect 24486 2796 24492 2848
rect 24544 2796 24550 2848
rect 1104 2746 24840 2768
rect 1104 2694 3917 2746
rect 3969 2694 3981 2746
rect 4033 2694 4045 2746
rect 4097 2694 4109 2746
rect 4161 2694 4173 2746
rect 4225 2694 9851 2746
rect 9903 2694 9915 2746
rect 9967 2694 9979 2746
rect 10031 2694 10043 2746
rect 10095 2694 10107 2746
rect 10159 2694 15785 2746
rect 15837 2694 15849 2746
rect 15901 2694 15913 2746
rect 15965 2694 15977 2746
rect 16029 2694 16041 2746
rect 16093 2694 21719 2746
rect 21771 2694 21783 2746
rect 21835 2694 21847 2746
rect 21899 2694 21911 2746
rect 21963 2694 21975 2746
rect 22027 2694 24840 2746
rect 1104 2672 24840 2694
rect 1946 2592 1952 2644
rect 2004 2592 2010 2644
rect 2685 2635 2743 2641
rect 2685 2601 2697 2635
rect 2731 2632 2743 2635
rect 4430 2632 4436 2644
rect 2731 2604 4436 2632
rect 2731 2601 2743 2604
rect 2685 2595 2743 2601
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 4982 2632 4988 2644
rect 4939 2604 4988 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 4982 2592 4988 2604
rect 5040 2592 5046 2644
rect 5166 2592 5172 2644
rect 5224 2592 5230 2644
rect 6733 2635 6791 2641
rect 6733 2601 6745 2635
rect 6779 2632 6791 2635
rect 6822 2632 6828 2644
rect 6779 2604 6828 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 6822 2592 6828 2604
rect 6880 2632 6886 2644
rect 7929 2635 7987 2641
rect 6880 2604 7604 2632
rect 6880 2592 6886 2604
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2564 1639 2567
rect 7576 2564 7604 2604
rect 7929 2601 7941 2635
rect 7975 2632 7987 2635
rect 8202 2632 8208 2644
rect 7975 2604 8208 2632
rect 7975 2601 7987 2604
rect 7929 2595 7987 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 8386 2592 8392 2644
rect 8444 2592 8450 2644
rect 9398 2592 9404 2644
rect 9456 2592 9462 2644
rect 10244 2604 10916 2632
rect 8404 2564 8432 2592
rect 1627 2536 4568 2564
rect 7576 2536 8432 2564
rect 8941 2567 8999 2573
rect 1627 2533 1639 2536
rect 1581 2527 1639 2533
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 992 2400 1409 2428
rect 992 2388 998 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1486 2388 1492 2440
rect 1544 2428 1550 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 1544 2400 1777 2428
rect 1544 2388 1550 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2498 2388 2504 2440
rect 2556 2388 2562 2440
rect 4540 2372 4568 2536
rect 8941 2533 8953 2567
rect 8987 2564 8999 2567
rect 9674 2564 9680 2576
rect 8987 2536 9680 2564
rect 8987 2533 8999 2536
rect 8941 2527 8999 2533
rect 9674 2524 9680 2536
rect 9732 2524 9738 2576
rect 5350 2456 5356 2508
rect 5408 2456 5414 2508
rect 10244 2505 10272 2604
rect 10229 2499 10287 2505
rect 7852 2468 10180 2496
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 4706 2388 4712 2440
rect 4764 2388 4770 2440
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 750 2320 756 2372
rect 808 2360 814 2372
rect 808 2332 4108 2360
rect 808 2320 814 2332
rect 4080 2304 4108 2332
rect 4522 2320 4528 2372
rect 4580 2320 4586 2372
rect 5000 2360 5028 2391
rect 5718 2388 5724 2440
rect 5776 2388 5782 2440
rect 5902 2388 5908 2440
rect 5960 2428 5966 2440
rect 6917 2431 6975 2437
rect 5960 2400 6592 2428
rect 5960 2388 5966 2400
rect 5258 2360 5264 2372
rect 5000 2332 5264 2360
rect 5258 2320 5264 2332
rect 5316 2320 5322 2372
rect 5368 2332 5672 2360
rect 4062 2252 4068 2304
rect 4120 2252 4126 2304
rect 4433 2295 4491 2301
rect 4433 2261 4445 2295
rect 4479 2292 4491 2295
rect 5368 2292 5396 2332
rect 4479 2264 5396 2292
rect 5445 2295 5503 2301
rect 4479 2261 4491 2264
rect 4433 2255 4491 2261
rect 5445 2261 5457 2295
rect 5491 2292 5503 2295
rect 5534 2292 5540 2304
rect 5491 2264 5540 2292
rect 5491 2261 5503 2264
rect 5445 2255 5503 2261
rect 5534 2252 5540 2264
rect 5592 2252 5598 2304
rect 5644 2292 5672 2332
rect 5810 2320 5816 2372
rect 5868 2320 5874 2372
rect 6564 2369 6592 2400
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 7098 2428 7104 2440
rect 6963 2400 7104 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7191 2431 7249 2437
rect 7191 2397 7203 2431
rect 7237 2428 7249 2431
rect 7558 2428 7564 2440
rect 7237 2400 7564 2428
rect 7237 2397 7249 2400
rect 7191 2391 7249 2397
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 6181 2363 6239 2369
rect 6181 2329 6193 2363
rect 6227 2329 6239 2363
rect 6181 2323 6239 2329
rect 6549 2363 6607 2369
rect 6549 2329 6561 2363
rect 6595 2329 6607 2363
rect 6549 2323 6607 2329
rect 6196 2292 6224 2323
rect 5644 2264 6224 2292
rect 6362 2252 6368 2304
rect 6420 2292 6426 2304
rect 7852 2292 7880 2468
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 8754 2388 8760 2440
rect 8812 2388 8818 2440
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2397 9919 2431
rect 10152 2428 10180 2468
rect 10229 2465 10241 2499
rect 10275 2465 10287 2499
rect 10888 2496 10916 2604
rect 11054 2592 11060 2644
rect 11112 2592 11118 2644
rect 11238 2592 11244 2644
rect 11296 2592 11302 2644
rect 13998 2632 14004 2644
rect 11557 2604 14004 2632
rect 11072 2564 11100 2592
rect 11557 2564 11585 2604
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 16758 2592 16764 2644
rect 16816 2632 16822 2644
rect 17129 2635 17187 2641
rect 17129 2632 17141 2635
rect 16816 2604 17141 2632
rect 16816 2592 16822 2604
rect 17129 2601 17141 2604
rect 17175 2601 17187 2635
rect 17129 2595 17187 2601
rect 17402 2592 17408 2644
rect 17460 2632 17466 2644
rect 18325 2635 18383 2641
rect 18325 2632 18337 2635
rect 17460 2604 18337 2632
rect 17460 2592 17466 2604
rect 18325 2601 18337 2604
rect 18371 2601 18383 2635
rect 18325 2595 18383 2601
rect 19058 2592 19064 2644
rect 19116 2632 19122 2644
rect 19245 2635 19303 2641
rect 19245 2632 19257 2635
rect 19116 2604 19257 2632
rect 19116 2592 19122 2604
rect 19245 2601 19257 2604
rect 19291 2601 19303 2635
rect 19935 2635 19993 2641
rect 19245 2595 19303 2601
rect 19628 2604 19806 2632
rect 13906 2564 13912 2576
rect 11072 2536 11585 2564
rect 11624 2536 13912 2564
rect 11330 2496 11336 2508
rect 10888 2468 11336 2496
rect 10229 2459 10287 2465
rect 11330 2456 11336 2468
rect 11388 2456 11394 2508
rect 10471 2431 10529 2437
rect 10471 2428 10483 2431
rect 10152 2400 10483 2428
rect 9861 2391 9919 2397
rect 10471 2397 10483 2400
rect 10517 2428 10529 2431
rect 11624 2428 11652 2536
rect 13906 2524 13912 2536
rect 13964 2524 13970 2576
rect 15289 2567 15347 2573
rect 15289 2533 15301 2567
rect 15335 2533 15347 2567
rect 19628 2564 19656 2604
rect 15289 2527 15347 2533
rect 15764 2536 19656 2564
rect 19778 2564 19806 2604
rect 19935 2601 19947 2635
rect 19981 2632 19993 2635
rect 20070 2632 20076 2644
rect 19981 2604 20076 2632
rect 19981 2601 19993 2604
rect 19935 2595 19993 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 21910 2592 21916 2644
rect 21968 2592 21974 2644
rect 24121 2635 24179 2641
rect 22020 2604 23888 2632
rect 22020 2564 22048 2604
rect 23860 2573 23888 2604
rect 24121 2601 24133 2635
rect 24167 2632 24179 2635
rect 24578 2632 24584 2644
rect 24167 2604 24584 2632
rect 24167 2601 24179 2604
rect 24121 2595 24179 2601
rect 24578 2592 24584 2604
rect 24636 2592 24642 2644
rect 19778 2536 22048 2564
rect 23845 2567 23903 2573
rect 15304 2496 15332 2527
rect 10517 2400 11652 2428
rect 11716 2468 15332 2496
rect 10517 2397 10529 2400
rect 10471 2391 10529 2397
rect 8662 2320 8668 2372
rect 8720 2360 8726 2372
rect 9309 2363 9367 2369
rect 9309 2360 9321 2363
rect 8720 2332 9321 2360
rect 8720 2320 8726 2332
rect 9309 2329 9321 2332
rect 9355 2329 9367 2363
rect 9876 2360 9904 2391
rect 11514 2360 11520 2372
rect 9876 2332 11520 2360
rect 9309 2323 9367 2329
rect 11514 2320 11520 2332
rect 11572 2320 11578 2372
rect 11716 2304 11744 2468
rect 11974 2388 11980 2440
rect 12032 2388 12038 2440
rect 12253 2431 12311 2437
rect 12253 2397 12265 2431
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 6420 2264 7880 2292
rect 6420 2252 6426 2264
rect 7926 2252 7932 2304
rect 7984 2292 7990 2304
rect 8297 2295 8355 2301
rect 8297 2292 8309 2295
rect 7984 2264 8309 2292
rect 7984 2252 7990 2264
rect 8297 2261 8309 2264
rect 8343 2261 8355 2295
rect 8297 2255 8355 2261
rect 8570 2252 8576 2304
rect 8628 2252 8634 2304
rect 9582 2252 9588 2304
rect 9640 2252 9646 2304
rect 10045 2295 10103 2301
rect 10045 2261 10057 2295
rect 10091 2292 10103 2295
rect 10778 2292 10784 2304
rect 10091 2264 10784 2292
rect 10091 2261 10103 2264
rect 10045 2255 10103 2261
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 11698 2252 11704 2304
rect 11756 2252 11762 2304
rect 11790 2252 11796 2304
rect 11848 2252 11854 2304
rect 12066 2252 12072 2304
rect 12124 2252 12130 2304
rect 12268 2292 12296 2391
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 12492 2400 12541 2428
rect 12492 2388 12498 2400
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 12894 2388 12900 2440
rect 12952 2388 12958 2440
rect 13262 2388 13268 2440
rect 13320 2388 13326 2440
rect 13538 2388 13544 2440
rect 13596 2388 13602 2440
rect 13817 2431 13875 2437
rect 13817 2397 13829 2431
rect 13863 2428 13875 2431
rect 14734 2428 14740 2440
rect 13863 2400 14740 2428
rect 13863 2397 13875 2400
rect 13817 2391 13875 2397
rect 14734 2388 14740 2400
rect 14792 2388 14798 2440
rect 14826 2388 14832 2440
rect 14884 2388 14890 2440
rect 15102 2388 15108 2440
rect 15160 2388 15166 2440
rect 15470 2388 15476 2440
rect 15528 2388 15534 2440
rect 15764 2437 15792 2536
rect 23845 2533 23857 2567
rect 23891 2533 23903 2567
rect 23845 2527 23903 2533
rect 16942 2456 16948 2508
rect 17000 2456 17006 2508
rect 18322 2496 18328 2508
rect 17052 2468 18328 2496
rect 15749 2431 15807 2437
rect 15749 2397 15761 2431
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 16022 2388 16028 2440
rect 16080 2388 16086 2440
rect 16393 2431 16451 2437
rect 16393 2397 16405 2431
rect 16439 2428 16451 2431
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16439 2400 16865 2428
rect 16439 2397 16451 2400
rect 16393 2391 16451 2397
rect 16853 2397 16865 2400
rect 16899 2428 16911 2431
rect 16960 2428 16988 2456
rect 16899 2400 16988 2428
rect 16899 2397 16911 2400
rect 16853 2391 16911 2397
rect 17052 2369 17080 2468
rect 18322 2456 18328 2468
rect 18380 2456 18386 2508
rect 18598 2456 18604 2508
rect 18656 2496 18662 2508
rect 19751 2499 19809 2505
rect 18656 2468 19656 2496
rect 18656 2456 18662 2468
rect 17310 2388 17316 2440
rect 17368 2388 17374 2440
rect 17494 2388 17500 2440
rect 17552 2388 17558 2440
rect 18874 2388 18880 2440
rect 18932 2388 18938 2440
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 17037 2363 17095 2369
rect 15580 2332 16804 2360
rect 12345 2295 12403 2301
rect 12345 2292 12357 2295
rect 12268 2264 12357 2292
rect 12345 2261 12357 2264
rect 12391 2261 12403 2295
rect 12345 2255 12403 2261
rect 12434 2252 12440 2304
rect 12492 2292 12498 2304
rect 12713 2295 12771 2301
rect 12713 2292 12725 2295
rect 12492 2264 12725 2292
rect 12492 2252 12498 2264
rect 12713 2261 12725 2264
rect 12759 2261 12771 2295
rect 12713 2255 12771 2261
rect 13081 2295 13139 2301
rect 13081 2261 13093 2295
rect 13127 2292 13139 2295
rect 13170 2292 13176 2304
rect 13127 2264 13176 2292
rect 13127 2261 13139 2264
rect 13081 2255 13139 2261
rect 13170 2252 13176 2264
rect 13228 2252 13234 2304
rect 13354 2252 13360 2304
rect 13412 2252 13418 2304
rect 13630 2252 13636 2304
rect 13688 2252 13694 2304
rect 14550 2252 14556 2304
rect 14608 2292 14614 2304
rect 14645 2295 14703 2301
rect 14645 2292 14657 2295
rect 14608 2264 14657 2292
rect 14608 2252 14614 2264
rect 14645 2261 14657 2264
rect 14691 2261 14703 2295
rect 14645 2255 14703 2261
rect 14918 2252 14924 2304
rect 14976 2252 14982 2304
rect 15580 2301 15608 2332
rect 15565 2295 15623 2301
rect 15565 2261 15577 2295
rect 15611 2261 15623 2295
rect 15565 2255 15623 2261
rect 15838 2252 15844 2304
rect 15896 2252 15902 2304
rect 16666 2252 16672 2304
rect 16724 2252 16730 2304
rect 16776 2292 16804 2332
rect 17037 2329 17049 2363
rect 17083 2329 17095 2363
rect 17328 2360 17356 2388
rect 17681 2363 17739 2369
rect 17681 2360 17693 2363
rect 17328 2332 17693 2360
rect 17037 2323 17095 2329
rect 17681 2329 17693 2332
rect 17727 2329 17739 2363
rect 17681 2323 17739 2329
rect 18233 2363 18291 2369
rect 18233 2329 18245 2363
rect 18279 2360 18291 2363
rect 19334 2360 19340 2372
rect 18279 2332 19340 2360
rect 18279 2329 18291 2332
rect 18233 2323 18291 2329
rect 19334 2320 19340 2332
rect 19392 2320 19398 2372
rect 17126 2292 17132 2304
rect 16776 2264 17132 2292
rect 17126 2252 17132 2264
rect 17184 2252 17190 2304
rect 17310 2252 17316 2304
rect 17368 2252 17374 2304
rect 17770 2252 17776 2304
rect 17828 2252 17834 2304
rect 18598 2252 18604 2304
rect 18656 2292 18662 2304
rect 18693 2295 18751 2301
rect 18693 2292 18705 2295
rect 18656 2264 18705 2292
rect 18656 2252 18662 2264
rect 18693 2261 18705 2264
rect 18739 2261 18751 2295
rect 19444 2292 19472 2391
rect 19628 2360 19656 2468
rect 19751 2465 19763 2499
rect 19797 2496 19809 2499
rect 19797 2468 20668 2496
rect 19797 2465 19809 2468
rect 19751 2459 19809 2465
rect 20640 2428 20668 2468
rect 20806 2456 20812 2508
rect 20864 2496 20870 2508
rect 22462 2496 22468 2508
rect 20864 2468 22468 2496
rect 20864 2456 20870 2468
rect 22462 2456 22468 2468
rect 22520 2456 22526 2508
rect 23750 2428 23756 2440
rect 20640 2400 23756 2428
rect 23750 2388 23756 2400
rect 23808 2388 23814 2440
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24029 2431 24087 2437
rect 24029 2428 24041 2431
rect 23900 2400 24041 2428
rect 23900 2388 23906 2400
rect 24029 2397 24041 2400
rect 24075 2397 24087 2431
rect 24029 2391 24087 2397
rect 19628 2332 20024 2360
rect 19794 2292 19800 2304
rect 19444 2264 19800 2292
rect 18693 2255 18751 2261
rect 19794 2252 19800 2264
rect 19852 2252 19858 2304
rect 19996 2292 20024 2332
rect 20622 2320 20628 2372
rect 20680 2320 20686 2372
rect 21450 2320 21456 2372
rect 21508 2360 21514 2372
rect 21726 2360 21732 2372
rect 21508 2332 21732 2360
rect 21508 2320 21514 2332
rect 21726 2320 21732 2332
rect 21784 2320 21790 2372
rect 22710 2363 22768 2369
rect 22710 2329 22722 2363
rect 22756 2329 22768 2363
rect 22710 2323 22768 2329
rect 22725 2292 22753 2323
rect 23474 2320 23480 2372
rect 23532 2360 23538 2372
rect 25130 2360 25136 2372
rect 23532 2332 25136 2360
rect 23532 2320 23538 2332
rect 25130 2320 25136 2332
rect 25188 2320 25194 2372
rect 19996 2264 22753 2292
rect 1104 2202 25000 2224
rect 1104 2150 6884 2202
rect 6936 2150 6948 2202
rect 7000 2150 7012 2202
rect 7064 2150 7076 2202
rect 7128 2150 7140 2202
rect 7192 2150 12818 2202
rect 12870 2150 12882 2202
rect 12934 2150 12946 2202
rect 12998 2150 13010 2202
rect 13062 2150 13074 2202
rect 13126 2150 18752 2202
rect 18804 2150 18816 2202
rect 18868 2150 18880 2202
rect 18932 2150 18944 2202
rect 18996 2150 19008 2202
rect 19060 2150 24686 2202
rect 24738 2150 24750 2202
rect 24802 2150 24814 2202
rect 24866 2150 24878 2202
rect 24930 2150 24942 2202
rect 24994 2150 25000 2202
rect 1104 2128 25000 2150
rect 2133 2091 2191 2097
rect 2133 2057 2145 2091
rect 2179 2088 2191 2091
rect 3050 2088 3056 2100
rect 2179 2060 3056 2088
rect 2179 2057 2191 2060
rect 2133 2051 2191 2057
rect 3050 2048 3056 2060
rect 3108 2048 3114 2100
rect 3237 2091 3295 2097
rect 3237 2057 3249 2091
rect 3283 2088 3295 2091
rect 3602 2088 3608 2100
rect 3283 2060 3608 2088
rect 3283 2057 3295 2060
rect 3237 2051 3295 2057
rect 3602 2048 3608 2060
rect 3660 2048 3666 2100
rect 3789 2091 3847 2097
rect 3789 2057 3801 2091
rect 3835 2088 3847 2091
rect 3970 2088 3976 2100
rect 3835 2060 3976 2088
rect 3835 2057 3847 2060
rect 3789 2051 3847 2057
rect 3970 2048 3976 2060
rect 4028 2048 4034 2100
rect 4062 2048 4068 2100
rect 4120 2048 4126 2100
rect 4246 2048 4252 2100
rect 4304 2048 4310 2100
rect 4430 2048 4436 2100
rect 4488 2048 4494 2100
rect 4709 2091 4767 2097
rect 4709 2057 4721 2091
rect 4755 2088 4767 2091
rect 5074 2088 5080 2100
rect 4755 2060 5080 2088
rect 4755 2057 4767 2060
rect 4709 2051 4767 2057
rect 5074 2048 5080 2060
rect 5132 2048 5138 2100
rect 5166 2048 5172 2100
rect 5224 2088 5230 2100
rect 5224 2060 5764 2088
rect 5224 2048 5230 2060
rect 1673 2023 1731 2029
rect 1673 1989 1685 2023
rect 1719 2020 1731 2023
rect 2866 2020 2872 2032
rect 1719 1992 2872 2020
rect 1719 1989 1731 1992
rect 1673 1983 1731 1989
rect 2866 1980 2872 1992
rect 2924 1980 2930 2032
rect 4264 2020 4292 2048
rect 5626 2020 5632 2032
rect 2976 1992 4292 2020
rect 4632 1992 5632 2020
rect 198 1912 204 1964
rect 256 1952 262 1964
rect 1489 1955 1547 1961
rect 1489 1952 1501 1955
rect 256 1924 1501 1952
rect 256 1912 262 1924
rect 1489 1921 1501 1924
rect 1535 1921 1547 1955
rect 1489 1915 1547 1921
rect 1857 1955 1915 1961
rect 1857 1921 1869 1955
rect 1903 1921 1915 1955
rect 1857 1915 1915 1921
rect 2409 1955 2467 1961
rect 2409 1921 2421 1955
rect 2455 1921 2467 1955
rect 2409 1915 2467 1921
rect 842 1844 848 1896
rect 900 1884 906 1896
rect 1872 1884 1900 1915
rect 900 1856 1900 1884
rect 900 1844 906 1856
rect 1026 1776 1032 1828
rect 1084 1816 1090 1828
rect 2424 1816 2452 1915
rect 2774 1912 2780 1964
rect 2832 1912 2838 1964
rect 2976 1825 3004 1992
rect 3050 1912 3056 1964
rect 3108 1912 3114 1964
rect 3510 1912 3516 1964
rect 3568 1912 3574 1964
rect 3605 1955 3663 1961
rect 3605 1921 3617 1955
rect 3651 1921 3663 1955
rect 3605 1915 3663 1921
rect 3620 1884 3648 1915
rect 3694 1912 3700 1964
rect 3752 1952 3758 1964
rect 4632 1961 4660 1992
rect 5626 1980 5632 1992
rect 5684 1980 5690 2032
rect 5736 2020 5764 2060
rect 5810 2048 5816 2100
rect 5868 2088 5874 2100
rect 5905 2091 5963 2097
rect 5905 2088 5917 2091
rect 5868 2060 5917 2088
rect 5868 2048 5874 2060
rect 5905 2057 5917 2060
rect 5951 2057 5963 2091
rect 5905 2051 5963 2057
rect 5994 2048 6000 2100
rect 6052 2088 6058 2100
rect 6641 2091 6699 2097
rect 6641 2088 6653 2091
rect 6052 2060 6653 2088
rect 6052 2048 6058 2060
rect 6641 2057 6653 2060
rect 6687 2057 6699 2091
rect 6641 2051 6699 2057
rect 7006 2048 7012 2100
rect 7064 2048 7070 2100
rect 7742 2048 7748 2100
rect 7800 2048 7806 2100
rect 7926 2048 7932 2100
rect 7984 2048 7990 2100
rect 8110 2048 8116 2100
rect 8168 2048 8174 2100
rect 8478 2048 8484 2100
rect 8536 2048 8542 2100
rect 8570 2048 8576 2100
rect 8628 2048 8634 2100
rect 8846 2048 8852 2100
rect 8904 2048 8910 2100
rect 9858 2088 9864 2100
rect 9048 2060 9864 2088
rect 5736 1992 6500 2020
rect 3973 1955 4031 1961
rect 3973 1952 3985 1955
rect 3752 1924 3985 1952
rect 3752 1912 3758 1924
rect 3973 1921 3985 1924
rect 4019 1921 4031 1955
rect 3973 1915 4031 1921
rect 4249 1955 4307 1961
rect 4249 1921 4261 1955
rect 4295 1921 4307 1955
rect 4249 1915 4307 1921
rect 4617 1955 4675 1961
rect 4617 1921 4629 1955
rect 4663 1921 4675 1955
rect 4617 1915 4675 1921
rect 4893 1955 4951 1961
rect 4893 1921 4905 1955
rect 4939 1952 4951 1955
rect 5074 1952 5080 1964
rect 4939 1924 5080 1952
rect 4939 1921 4951 1924
rect 4893 1915 4951 1921
rect 4062 1884 4068 1896
rect 3620 1856 4068 1884
rect 4062 1844 4068 1856
rect 4120 1844 4126 1896
rect 1084 1788 2452 1816
rect 2593 1819 2651 1825
rect 1084 1776 1090 1788
rect 2593 1785 2605 1819
rect 2639 1816 2651 1819
rect 2961 1819 3019 1825
rect 2639 1788 2774 1816
rect 2639 1785 2651 1788
rect 2593 1779 2651 1785
rect 2746 1748 2774 1788
rect 2961 1785 2973 1819
rect 3007 1785 3019 1819
rect 4264 1816 4292 1915
rect 5074 1912 5080 1924
rect 5132 1912 5138 1964
rect 5167 1955 5225 1961
rect 5167 1921 5179 1955
rect 5213 1952 5225 1955
rect 6362 1952 6368 1964
rect 5213 1924 6368 1952
rect 5213 1921 5225 1924
rect 5167 1915 5225 1921
rect 6362 1912 6368 1924
rect 6420 1912 6426 1964
rect 5718 1844 5724 1896
rect 5776 1844 5782 1896
rect 6472 1884 6500 1992
rect 6546 1980 6552 2032
rect 6604 1980 6610 2032
rect 6917 2023 6975 2029
rect 6917 1989 6929 2023
rect 6963 2020 6975 2023
rect 7282 2020 7288 2032
rect 6963 1992 7288 2020
rect 6963 1989 6975 1992
rect 6917 1983 6975 1989
rect 7282 1980 7288 1992
rect 7340 1980 7346 2032
rect 7653 2023 7711 2029
rect 7653 1989 7665 2023
rect 7699 2020 7711 2023
rect 7944 2020 7972 2048
rect 7699 1992 7972 2020
rect 8021 2023 8079 2029
rect 7699 1989 7711 1992
rect 7653 1983 7711 1989
rect 8021 1989 8033 2023
rect 8067 2020 8079 2023
rect 8588 2020 8616 2048
rect 8067 1992 8616 2020
rect 8757 2023 8815 2029
rect 8067 1989 8079 1992
rect 8021 1983 8079 1989
rect 8757 1989 8769 2023
rect 8803 2020 8815 2023
rect 8938 2020 8944 2032
rect 8803 1992 8944 2020
rect 8803 1989 8815 1992
rect 8757 1983 8815 1989
rect 8938 1980 8944 1992
rect 8996 1980 9002 2032
rect 7193 1955 7251 1961
rect 7193 1921 7205 1955
rect 7239 1952 7251 1955
rect 7466 1952 7472 1964
rect 7239 1924 7472 1952
rect 7239 1921 7251 1924
rect 7193 1915 7251 1921
rect 7466 1912 7472 1924
rect 7524 1912 7530 1964
rect 7576 1924 8156 1952
rect 7576 1884 7604 1924
rect 6472 1856 7604 1884
rect 8018 1844 8024 1896
rect 8076 1844 8082 1896
rect 8128 1884 8156 1924
rect 8294 1912 8300 1964
rect 8352 1952 8358 1964
rect 9048 1961 9076 2060
rect 9858 2048 9864 2060
rect 9916 2048 9922 2100
rect 10045 2091 10103 2097
rect 10045 2057 10057 2091
rect 10091 2088 10103 2091
rect 10226 2088 10232 2100
rect 10091 2060 10232 2088
rect 10091 2057 10103 2060
rect 10045 2051 10103 2057
rect 10226 2048 10232 2060
rect 10284 2048 10290 2100
rect 13354 2088 13360 2100
rect 10520 2060 13360 2088
rect 10318 2020 10324 2032
rect 9324 1992 10324 2020
rect 9324 1991 9352 1992
rect 9291 1985 9352 1991
rect 8389 1955 8447 1961
rect 8389 1952 8401 1955
rect 8352 1924 8401 1952
rect 8352 1912 8358 1924
rect 8389 1921 8401 1924
rect 8435 1921 8447 1955
rect 8389 1915 8447 1921
rect 9033 1955 9091 1961
rect 9033 1921 9045 1955
rect 9079 1921 9091 1955
rect 9291 1951 9303 1985
rect 9337 1954 9352 1985
rect 10318 1980 10324 1992
rect 10376 1980 10382 2032
rect 9337 1951 9349 1954
rect 9291 1945 9349 1951
rect 9033 1915 9091 1921
rect 9048 1884 9076 1915
rect 9398 1912 9404 1964
rect 9456 1952 9462 1964
rect 10410 1952 10416 1964
rect 9456 1924 10416 1952
rect 9456 1912 9462 1924
rect 10410 1912 10416 1924
rect 10468 1912 10474 1964
rect 10520 1961 10548 2060
rect 13354 2048 13360 2060
rect 13412 2048 13418 2100
rect 13630 2048 13636 2100
rect 13688 2048 13694 2100
rect 14918 2048 14924 2100
rect 14976 2048 14982 2100
rect 15838 2048 15844 2100
rect 15896 2048 15902 2100
rect 17310 2048 17316 2100
rect 17368 2048 17374 2100
rect 18598 2048 18604 2100
rect 18656 2048 18662 2100
rect 19334 2048 19340 2100
rect 19392 2088 19398 2100
rect 19429 2091 19487 2097
rect 19429 2088 19441 2091
rect 19392 2060 19441 2088
rect 19392 2048 19398 2060
rect 19429 2057 19441 2060
rect 19475 2057 19487 2091
rect 19429 2051 19487 2057
rect 19794 2048 19800 2100
rect 19852 2088 19858 2100
rect 20346 2088 20352 2100
rect 19852 2060 20352 2088
rect 19852 2048 19858 2060
rect 20346 2048 20352 2060
rect 20404 2048 20410 2100
rect 21726 2048 21732 2100
rect 21784 2088 21790 2100
rect 23109 2091 23167 2097
rect 23109 2088 23121 2091
rect 21784 2060 23121 2088
rect 21784 2048 21790 2060
rect 23109 2057 23121 2060
rect 23155 2057 23167 2091
rect 23109 2051 23167 2057
rect 23474 2048 23480 2100
rect 23532 2048 23538 2100
rect 23845 2091 23903 2097
rect 23845 2057 23857 2091
rect 23891 2088 23903 2091
rect 23934 2088 23940 2100
rect 23891 2060 23940 2088
rect 23891 2057 23903 2060
rect 23845 2051 23903 2057
rect 23934 2048 23940 2060
rect 23992 2048 23998 2100
rect 24486 2048 24492 2100
rect 24544 2048 24550 2100
rect 10965 2023 11023 2029
rect 10965 1989 10977 2023
rect 11011 2020 11023 2023
rect 11698 2020 11704 2032
rect 11011 1992 11704 2020
rect 11011 1989 11023 1992
rect 10965 1983 11023 1989
rect 11698 1980 11704 1992
rect 11756 1980 11762 2032
rect 11793 2023 11851 2029
rect 11793 1989 11805 2023
rect 11839 2020 11851 2023
rect 13648 2020 13676 2048
rect 11839 1992 13676 2020
rect 11839 1989 11851 1992
rect 11793 1983 11851 1989
rect 10505 1955 10563 1961
rect 10505 1921 10517 1955
rect 10551 1921 10563 1955
rect 10505 1915 10563 1921
rect 12342 1912 12348 1964
rect 12400 1912 12406 1964
rect 13081 1955 13139 1961
rect 13081 1921 13093 1955
rect 13127 1952 13139 1955
rect 13541 1955 13599 1961
rect 13541 1952 13553 1955
rect 13127 1924 13553 1952
rect 13127 1921 13139 1924
rect 13081 1915 13139 1921
rect 13541 1921 13553 1924
rect 13587 1952 13599 1955
rect 13722 1952 13728 1964
rect 13587 1924 13728 1952
rect 13587 1921 13599 1924
rect 13541 1915 13599 1921
rect 13722 1912 13728 1924
rect 13780 1912 13786 1964
rect 13814 1912 13820 1964
rect 13872 1912 13878 1964
rect 14274 1912 14280 1964
rect 14332 1912 14338 1964
rect 14461 1955 14519 1961
rect 14461 1921 14473 1955
rect 14507 1921 14519 1955
rect 14461 1915 14519 1921
rect 14829 1955 14887 1961
rect 14829 1921 14841 1955
rect 14875 1952 14887 1955
rect 14936 1952 14964 2048
rect 15657 2023 15715 2029
rect 15657 1989 15669 2023
rect 15703 2020 15715 2023
rect 15856 2020 15884 2048
rect 15703 1992 15884 2020
rect 16761 2023 16819 2029
rect 15703 1989 15715 1992
rect 15657 1983 15715 1989
rect 16761 1989 16773 2023
rect 16807 2020 16819 2023
rect 17328 2020 17356 2048
rect 16807 1992 17356 2020
rect 16807 1989 16819 1992
rect 16761 1983 16819 1989
rect 17586 1980 17592 2032
rect 17644 2020 17650 2032
rect 17865 2023 17923 2029
rect 17865 2020 17877 2023
rect 17644 1992 17877 2020
rect 17644 1980 17650 1992
rect 17865 1989 17877 1992
rect 17911 1989 17923 2023
rect 17865 1983 17923 1989
rect 18417 2023 18475 2029
rect 18417 1989 18429 2023
rect 18463 2020 18475 2023
rect 18506 2020 18512 2032
rect 18463 1992 18512 2020
rect 18463 1989 18475 1992
rect 18417 1983 18475 1989
rect 18506 1980 18512 1992
rect 18564 1980 18570 2032
rect 18616 2020 18644 2048
rect 18969 2023 19027 2029
rect 18969 2020 18981 2023
rect 18616 1992 18981 2020
rect 18969 1989 18981 1992
rect 19015 1989 19027 2023
rect 23492 2020 23520 2048
rect 24504 2020 24532 2048
rect 18969 1983 19027 1989
rect 19076 1992 23520 2020
rect 24044 1992 24532 2020
rect 14875 1924 14964 1952
rect 15381 1955 15439 1961
rect 14875 1921 14887 1924
rect 14829 1915 14887 1921
rect 15381 1921 15393 1955
rect 15427 1921 15439 1955
rect 15381 1915 15439 1921
rect 11698 1884 11704 1896
rect 8128 1856 9076 1884
rect 10704 1856 11704 1884
rect 2961 1779 3019 1785
rect 3068 1788 4200 1816
rect 4264 1788 5028 1816
rect 3068 1748 3096 1788
rect 2746 1720 3096 1748
rect 3326 1708 3332 1760
rect 3384 1708 3390 1760
rect 4172 1748 4200 1788
rect 4798 1748 4804 1760
rect 4172 1720 4804 1748
rect 4798 1708 4804 1720
rect 4856 1708 4862 1760
rect 5000 1748 5028 1788
rect 5350 1748 5356 1760
rect 5000 1720 5356 1748
rect 5350 1708 5356 1720
rect 5408 1708 5414 1760
rect 5736 1748 5764 1844
rect 7377 1819 7435 1825
rect 7377 1785 7389 1819
rect 7423 1816 7435 1819
rect 8036 1816 8064 1844
rect 10704 1825 10732 1856
rect 11698 1844 11704 1856
rect 11756 1844 11762 1896
rect 14476 1884 14504 1915
rect 15396 1884 15424 1915
rect 16114 1912 16120 1964
rect 16172 1912 16178 1964
rect 16850 1912 16856 1964
rect 16908 1952 16914 1964
rect 17313 1955 17371 1961
rect 17313 1952 17325 1955
rect 16908 1924 17325 1952
rect 16908 1912 16914 1924
rect 17313 1921 17325 1924
rect 17359 1921 17371 1955
rect 17313 1915 17371 1921
rect 17681 1955 17739 1961
rect 17681 1921 17693 1955
rect 17727 1952 17739 1955
rect 18598 1952 18604 1964
rect 17727 1924 18604 1952
rect 17727 1921 17739 1924
rect 17681 1915 17739 1921
rect 18598 1912 18604 1924
rect 18656 1912 18662 1964
rect 19076 1884 19104 1992
rect 19518 1912 19524 1964
rect 19576 1952 19582 1964
rect 19613 1955 19671 1961
rect 19613 1952 19625 1955
rect 19576 1924 19625 1952
rect 19576 1912 19582 1924
rect 19613 1921 19625 1924
rect 19659 1921 19671 1955
rect 19613 1915 19671 1921
rect 19981 1955 20039 1961
rect 19981 1921 19993 1955
rect 20027 1952 20039 1955
rect 20254 1952 20260 1964
rect 20027 1924 20260 1952
rect 20027 1921 20039 1924
rect 19981 1915 20039 1921
rect 20254 1912 20260 1924
rect 20312 1912 20318 1964
rect 20714 1912 20720 1964
rect 20772 1912 20778 1964
rect 21358 1912 21364 1964
rect 21416 1952 21422 1964
rect 24044 1961 24072 1992
rect 21821 1955 21879 1961
rect 21821 1952 21833 1955
rect 21416 1924 21833 1952
rect 21416 1912 21422 1924
rect 21821 1921 21833 1924
rect 21867 1921 21879 1955
rect 21821 1915 21879 1921
rect 24029 1955 24087 1961
rect 24029 1921 24041 1955
rect 24075 1921 24087 1955
rect 24029 1915 24087 1921
rect 24302 1912 24308 1964
rect 24360 1912 24366 1964
rect 14476 1856 15240 1884
rect 15396 1856 19104 1884
rect 19705 1887 19763 1893
rect 7423 1788 8064 1816
rect 10689 1819 10747 1825
rect 7423 1785 7435 1788
rect 7377 1779 7435 1785
rect 10689 1785 10701 1819
rect 10735 1785 10747 1819
rect 10689 1779 10747 1785
rect 11146 1776 11152 1828
rect 11204 1776 11210 1828
rect 11882 1776 11888 1828
rect 11940 1816 11946 1828
rect 15212 1825 15240 1856
rect 19705 1853 19717 1887
rect 19751 1853 19763 1887
rect 19705 1847 19763 1853
rect 11977 1819 12035 1825
rect 11977 1816 11989 1819
rect 11940 1788 11989 1816
rect 11940 1776 11946 1788
rect 11977 1785 11989 1788
rect 12023 1785 12035 1819
rect 11977 1779 12035 1785
rect 15197 1819 15255 1825
rect 15197 1785 15209 1819
rect 15243 1785 15255 1819
rect 15197 1779 15255 1785
rect 15378 1776 15384 1828
rect 15436 1816 15442 1828
rect 15436 1788 16344 1816
rect 15436 1776 15442 1788
rect 12250 1748 12256 1760
rect 5736 1720 12256 1748
rect 12250 1708 12256 1720
rect 12308 1708 12314 1760
rect 12618 1708 12624 1760
rect 12676 1708 12682 1760
rect 13354 1708 13360 1760
rect 13412 1708 13418 1760
rect 13630 1708 13636 1760
rect 13688 1708 13694 1760
rect 14090 1708 14096 1760
rect 14148 1708 14154 1760
rect 14274 1708 14280 1760
rect 14332 1748 14338 1760
rect 14645 1751 14703 1757
rect 14645 1748 14657 1751
rect 14332 1720 14657 1748
rect 14332 1708 14338 1720
rect 14645 1717 14657 1720
rect 14691 1717 14703 1751
rect 14645 1711 14703 1717
rect 14734 1708 14740 1760
rect 14792 1748 14798 1760
rect 15013 1751 15071 1757
rect 15013 1748 15025 1751
rect 14792 1720 15025 1748
rect 14792 1708 14798 1720
rect 15013 1717 15025 1720
rect 15059 1717 15071 1751
rect 15013 1711 15071 1717
rect 15746 1708 15752 1760
rect 15804 1708 15810 1760
rect 16316 1757 16344 1788
rect 17126 1776 17132 1828
rect 17184 1816 17190 1828
rect 19720 1816 19748 1847
rect 19794 1844 19800 1896
rect 19852 1884 19858 1896
rect 20993 1887 21051 1893
rect 20993 1884 21005 1887
rect 19852 1856 21005 1884
rect 19852 1844 19858 1856
rect 20993 1853 21005 1856
rect 21039 1853 21051 1887
rect 25314 1884 25320 1896
rect 20993 1847 21051 1853
rect 22066 1856 25320 1884
rect 22066 1816 22094 1856
rect 25314 1844 25320 1856
rect 25372 1844 25378 1896
rect 17184 1788 19104 1816
rect 19720 1788 22094 1816
rect 17184 1776 17190 1788
rect 16301 1751 16359 1757
rect 16301 1717 16313 1751
rect 16347 1717 16359 1751
rect 16301 1711 16359 1717
rect 16850 1708 16856 1760
rect 16908 1708 16914 1760
rect 17954 1708 17960 1760
rect 18012 1708 18018 1760
rect 18138 1708 18144 1760
rect 18196 1748 18202 1760
rect 19076 1757 19104 1788
rect 22738 1776 22744 1828
rect 22796 1816 22802 1828
rect 24121 1819 24179 1825
rect 24121 1816 24133 1819
rect 22796 1788 24133 1816
rect 22796 1776 22802 1788
rect 24121 1785 24133 1788
rect 24167 1785 24179 1819
rect 24121 1779 24179 1785
rect 18509 1751 18567 1757
rect 18509 1748 18521 1751
rect 18196 1720 18521 1748
rect 18196 1708 18202 1720
rect 18509 1717 18521 1720
rect 18555 1717 18567 1751
rect 18509 1711 18567 1717
rect 19061 1751 19119 1757
rect 19061 1717 19073 1751
rect 19107 1717 19119 1751
rect 19061 1711 19119 1717
rect 19518 1708 19524 1760
rect 19576 1748 19582 1760
rect 20162 1748 20168 1760
rect 19576 1720 20168 1748
rect 19576 1708 19582 1720
rect 20162 1708 20168 1720
rect 20220 1708 20226 1760
rect 1104 1658 24840 1680
rect 1104 1606 3917 1658
rect 3969 1606 3981 1658
rect 4033 1606 4045 1658
rect 4097 1606 4109 1658
rect 4161 1606 4173 1658
rect 4225 1606 9851 1658
rect 9903 1606 9915 1658
rect 9967 1606 9979 1658
rect 10031 1606 10043 1658
rect 10095 1606 10107 1658
rect 10159 1606 15785 1658
rect 15837 1606 15849 1658
rect 15901 1606 15913 1658
rect 15965 1606 15977 1658
rect 16029 1606 16041 1658
rect 16093 1606 21719 1658
rect 21771 1606 21783 1658
rect 21835 1606 21847 1658
rect 21899 1606 21911 1658
rect 21963 1606 21975 1658
rect 22027 1606 24840 1658
rect 1104 1584 24840 1606
rect 3326 1504 3332 1556
rect 3384 1544 3390 1556
rect 4430 1544 4436 1556
rect 3384 1516 4436 1544
rect 3384 1504 3390 1516
rect 4430 1504 4436 1516
rect 4488 1504 4494 1556
rect 4522 1504 4528 1556
rect 4580 1544 4586 1556
rect 9030 1544 9036 1556
rect 4580 1516 9036 1544
rect 4580 1504 4586 1516
rect 9030 1504 9036 1516
rect 9088 1504 9094 1556
rect 10410 1504 10416 1556
rect 10468 1544 10474 1556
rect 10689 1547 10747 1553
rect 10689 1544 10701 1547
rect 10468 1516 10701 1544
rect 10468 1504 10474 1516
rect 10689 1513 10701 1516
rect 10735 1513 10747 1547
rect 10689 1507 10747 1513
rect 10962 1504 10968 1556
rect 11020 1504 11026 1556
rect 12434 1544 12440 1556
rect 11072 1516 12440 1544
rect 7742 1476 7748 1488
rect 4080 1448 7748 1476
rect 1670 1300 1676 1352
rect 1728 1340 1734 1352
rect 1765 1343 1823 1349
rect 1765 1340 1777 1343
rect 1728 1312 1777 1340
rect 1728 1300 1734 1312
rect 1765 1309 1777 1312
rect 1811 1309 1823 1343
rect 1765 1303 1823 1309
rect 2038 1300 2044 1352
rect 2096 1340 2102 1352
rect 2133 1343 2191 1349
rect 2133 1340 2145 1343
rect 2096 1312 2145 1340
rect 2096 1300 2102 1312
rect 2133 1309 2145 1312
rect 2179 1309 2191 1343
rect 2133 1303 2191 1309
rect 2222 1300 2228 1352
rect 2280 1300 2286 1352
rect 2501 1343 2559 1349
rect 2501 1309 2513 1343
rect 2547 1340 2559 1343
rect 2590 1340 2596 1352
rect 2547 1312 2596 1340
rect 2547 1309 2559 1312
rect 2501 1303 2559 1309
rect 2590 1300 2596 1312
rect 2648 1300 2654 1352
rect 3421 1343 3479 1349
rect 3421 1309 3433 1343
rect 3467 1340 3479 1343
rect 3786 1340 3792 1352
rect 3467 1312 3792 1340
rect 3467 1309 3479 1312
rect 3421 1303 3479 1309
rect 3786 1300 3792 1312
rect 3844 1300 3850 1352
rect 4080 1349 4108 1448
rect 7742 1436 7748 1448
rect 7800 1436 7806 1488
rect 10980 1476 11008 1504
rect 7852 1448 11008 1476
rect 6454 1368 6460 1420
rect 6512 1408 6518 1420
rect 6512 1380 6868 1408
rect 6512 1368 6518 1380
rect 4065 1343 4123 1349
rect 4065 1309 4077 1343
rect 4111 1309 4123 1343
rect 4065 1303 4123 1309
rect 4157 1343 4215 1349
rect 4157 1309 4169 1343
rect 4203 1309 4215 1343
rect 4157 1303 4215 1309
rect 1578 1232 1584 1284
rect 1636 1232 1642 1284
rect 1946 1232 1952 1284
rect 2004 1232 2010 1284
rect 2958 1232 2964 1284
rect 3016 1272 3022 1284
rect 3237 1275 3295 1281
rect 3237 1272 3249 1275
rect 3016 1244 3249 1272
rect 3016 1232 3022 1244
rect 3237 1241 3249 1244
rect 3283 1241 3295 1275
rect 3237 1235 3295 1241
rect 3878 1164 3884 1216
rect 3936 1164 3942 1216
rect 4062 1164 4068 1216
rect 4120 1204 4126 1216
rect 4172 1204 4200 1303
rect 4430 1300 4436 1352
rect 4488 1300 4494 1352
rect 5261 1343 5319 1349
rect 5261 1309 5273 1343
rect 5307 1340 5319 1343
rect 5810 1340 5816 1352
rect 5307 1312 5816 1340
rect 5307 1309 5319 1312
rect 5261 1303 5319 1309
rect 5810 1300 5816 1312
rect 5868 1300 5874 1352
rect 5905 1343 5963 1349
rect 5905 1309 5917 1343
rect 5951 1340 5963 1343
rect 6270 1340 6276 1352
rect 5951 1312 6276 1340
rect 5951 1309 5963 1312
rect 5905 1303 5963 1309
rect 6270 1300 6276 1312
rect 6328 1300 6334 1352
rect 6362 1300 6368 1352
rect 6420 1340 6426 1352
rect 6549 1343 6607 1349
rect 6549 1340 6561 1343
rect 6420 1312 6561 1340
rect 6420 1300 6426 1312
rect 6549 1309 6561 1312
rect 6595 1309 6607 1343
rect 6549 1303 6607 1309
rect 6730 1300 6736 1352
rect 6788 1300 6794 1352
rect 6840 1340 6868 1380
rect 6914 1368 6920 1420
rect 6972 1408 6978 1420
rect 7852 1408 7880 1448
rect 10226 1408 10232 1420
rect 6972 1380 7880 1408
rect 9508 1380 10232 1408
rect 6972 1368 6978 1380
rect 7009 1343 7067 1349
rect 7009 1340 7021 1343
rect 6840 1312 7021 1340
rect 7009 1309 7021 1312
rect 7055 1309 7067 1343
rect 7009 1303 7067 1309
rect 8202 1300 8208 1352
rect 8260 1340 8266 1352
rect 8481 1343 8539 1349
rect 8481 1340 8493 1343
rect 8260 1312 8493 1340
rect 8260 1300 8266 1312
rect 8481 1309 8493 1312
rect 8527 1309 8539 1343
rect 8481 1303 8539 1309
rect 8757 1343 8815 1349
rect 8757 1309 8769 1343
rect 8803 1340 8815 1343
rect 9030 1340 9036 1352
rect 8803 1312 9036 1340
rect 8803 1309 8815 1312
rect 8757 1303 8815 1309
rect 9030 1300 9036 1312
rect 9088 1300 9094 1352
rect 9125 1343 9183 1349
rect 9125 1309 9137 1343
rect 9171 1340 9183 1343
rect 9508 1340 9536 1380
rect 10226 1368 10232 1380
rect 10284 1368 10290 1420
rect 10321 1411 10379 1417
rect 10321 1377 10333 1411
rect 10367 1408 10379 1411
rect 10367 1380 11008 1408
rect 10367 1377 10379 1380
rect 10321 1371 10379 1377
rect 9171 1312 9536 1340
rect 9171 1309 9183 1312
rect 9125 1303 9183 1309
rect 9582 1300 9588 1352
rect 9640 1300 9646 1352
rect 9674 1300 9680 1352
rect 9732 1340 9738 1352
rect 10597 1343 10655 1349
rect 10597 1340 10609 1343
rect 9732 1312 10609 1340
rect 9732 1300 9738 1312
rect 10597 1309 10609 1312
rect 10643 1309 10655 1343
rect 10597 1303 10655 1309
rect 5445 1275 5503 1281
rect 5445 1241 5457 1275
rect 5491 1272 5503 1275
rect 5994 1272 6000 1284
rect 5491 1244 6000 1272
rect 5491 1241 5503 1244
rect 5445 1235 5503 1241
rect 5994 1232 6000 1244
rect 6052 1232 6058 1284
rect 7469 1275 7527 1281
rect 7469 1272 7481 1275
rect 6564 1244 7481 1272
rect 6564 1216 6592 1244
rect 7469 1241 7481 1244
rect 7515 1241 7527 1275
rect 7469 1235 7527 1241
rect 7837 1275 7895 1281
rect 7837 1241 7849 1275
rect 7883 1272 7895 1275
rect 9309 1275 9367 1281
rect 9309 1272 9321 1275
rect 7883 1244 8340 1272
rect 7883 1241 7895 1244
rect 7837 1235 7895 1241
rect 4120 1176 4200 1204
rect 4120 1164 4126 1176
rect 5074 1164 5080 1216
rect 5132 1164 5138 1216
rect 5534 1164 5540 1216
rect 5592 1164 5598 1216
rect 6086 1164 6092 1216
rect 6144 1164 6150 1216
rect 6365 1207 6423 1213
rect 6365 1173 6377 1207
rect 6411 1204 6423 1207
rect 6454 1204 6460 1216
rect 6411 1176 6460 1204
rect 6411 1173 6423 1176
rect 6365 1167 6423 1173
rect 6454 1164 6460 1176
rect 6512 1164 6518 1216
rect 6546 1164 6552 1216
rect 6604 1164 6610 1216
rect 6730 1164 6736 1216
rect 6788 1204 6794 1216
rect 6825 1207 6883 1213
rect 6825 1204 6837 1207
rect 6788 1176 6837 1204
rect 6788 1164 6794 1176
rect 6825 1173 6837 1176
rect 6871 1173 6883 1207
rect 6825 1167 6883 1173
rect 6914 1164 6920 1216
rect 6972 1204 6978 1216
rect 7193 1207 7251 1213
rect 7193 1204 7205 1207
rect 6972 1176 7205 1204
rect 6972 1164 6978 1176
rect 7193 1173 7205 1176
rect 7239 1173 7251 1207
rect 7193 1167 7251 1173
rect 7558 1164 7564 1216
rect 7616 1164 7622 1216
rect 7926 1164 7932 1216
rect 7984 1164 7990 1216
rect 8312 1213 8340 1244
rect 8588 1244 9321 1272
rect 8588 1213 8616 1244
rect 9309 1241 9321 1244
rect 9355 1241 9367 1275
rect 9309 1235 9367 1241
rect 9493 1275 9551 1281
rect 9493 1241 9505 1275
rect 9539 1272 9551 1275
rect 10045 1275 10103 1281
rect 9539 1244 9996 1272
rect 9539 1241 9551 1244
rect 9493 1235 9551 1241
rect 8297 1207 8355 1213
rect 8297 1173 8309 1207
rect 8343 1173 8355 1207
rect 8297 1167 8355 1173
rect 8573 1207 8631 1213
rect 8573 1173 8585 1207
rect 8619 1173 8631 1207
rect 8573 1167 8631 1173
rect 8938 1164 8944 1216
rect 8996 1164 9002 1216
rect 9766 1164 9772 1216
rect 9824 1164 9830 1216
rect 9968 1204 9996 1244
rect 10045 1241 10057 1275
rect 10091 1272 10103 1275
rect 10778 1272 10784 1284
rect 10091 1244 10784 1272
rect 10091 1241 10103 1244
rect 10045 1235 10103 1241
rect 10778 1232 10784 1244
rect 10836 1232 10842 1284
rect 10980 1272 11008 1380
rect 11072 1349 11100 1516
rect 12434 1504 12440 1516
rect 12492 1504 12498 1556
rect 12526 1504 12532 1556
rect 12584 1544 12590 1556
rect 12713 1547 12771 1553
rect 12713 1544 12725 1547
rect 12584 1516 12725 1544
rect 12584 1504 12590 1516
rect 12713 1513 12725 1516
rect 12759 1513 12771 1547
rect 12713 1507 12771 1513
rect 13354 1504 13360 1556
rect 13412 1504 13418 1556
rect 13722 1504 13728 1556
rect 13780 1544 13786 1556
rect 14277 1547 14335 1553
rect 14277 1544 14289 1547
rect 13780 1516 14289 1544
rect 13780 1504 13786 1516
rect 14277 1513 14289 1516
rect 14323 1513 14335 1547
rect 14277 1507 14335 1513
rect 14918 1504 14924 1556
rect 14976 1544 14982 1556
rect 15381 1547 15439 1553
rect 15381 1544 15393 1547
rect 14976 1516 15393 1544
rect 14976 1504 14982 1516
rect 15381 1513 15393 1516
rect 15427 1513 15439 1547
rect 15381 1507 15439 1513
rect 15933 1547 15991 1553
rect 15933 1513 15945 1547
rect 15979 1513 15991 1547
rect 15933 1507 15991 1513
rect 11698 1436 11704 1488
rect 11756 1476 11762 1488
rect 11974 1476 11980 1488
rect 11756 1448 11980 1476
rect 11756 1436 11762 1448
rect 11974 1436 11980 1448
rect 12032 1436 12038 1488
rect 12066 1436 12072 1488
rect 12124 1476 12130 1488
rect 12124 1448 12664 1476
rect 12124 1436 12130 1448
rect 11330 1368 11336 1420
rect 11388 1408 11394 1420
rect 12250 1408 12256 1420
rect 11388 1380 12256 1408
rect 11388 1368 11394 1380
rect 12250 1368 12256 1380
rect 12308 1368 12314 1420
rect 11057 1343 11115 1349
rect 11057 1309 11069 1343
rect 11103 1309 11115 1343
rect 11057 1303 11115 1309
rect 11517 1343 11575 1349
rect 11517 1309 11529 1343
rect 11563 1340 11575 1343
rect 11790 1340 11796 1352
rect 11563 1312 11796 1340
rect 11563 1309 11575 1312
rect 11517 1303 11575 1309
rect 11790 1300 11796 1312
rect 11848 1300 11854 1352
rect 12636 1349 12664 1448
rect 13372 1408 13400 1504
rect 14090 1436 14096 1488
rect 14148 1436 14154 1488
rect 14182 1436 14188 1488
rect 14240 1476 14246 1488
rect 14240 1448 15148 1476
rect 14240 1436 14246 1448
rect 14108 1408 14136 1436
rect 15120 1408 15148 1448
rect 15194 1436 15200 1488
rect 15252 1476 15258 1488
rect 15948 1476 15976 1507
rect 16114 1504 16120 1556
rect 16172 1544 16178 1556
rect 16301 1547 16359 1553
rect 16301 1544 16313 1547
rect 16172 1516 16313 1544
rect 16172 1504 16178 1516
rect 16301 1513 16313 1516
rect 16347 1513 16359 1547
rect 16301 1507 16359 1513
rect 16853 1547 16911 1553
rect 16853 1513 16865 1547
rect 16899 1513 16911 1547
rect 16853 1507 16911 1513
rect 17405 1547 17463 1553
rect 17405 1513 17417 1547
rect 17451 1513 17463 1547
rect 17405 1507 17463 1513
rect 15252 1448 15976 1476
rect 15252 1436 15258 1448
rect 16022 1436 16028 1488
rect 16080 1476 16086 1488
rect 16868 1476 16896 1507
rect 16080 1448 16896 1476
rect 16080 1436 16086 1448
rect 13372 1380 13768 1408
rect 14108 1380 14780 1408
rect 15120 1380 16160 1408
rect 12069 1343 12127 1349
rect 12069 1309 12081 1343
rect 12115 1340 12127 1343
rect 12345 1343 12403 1349
rect 12345 1340 12357 1343
rect 12115 1312 12357 1340
rect 12115 1309 12127 1312
rect 12069 1303 12127 1309
rect 12345 1309 12357 1312
rect 12391 1309 12403 1343
rect 12345 1303 12403 1309
rect 12621 1343 12679 1349
rect 12621 1309 12633 1343
rect 12667 1309 12679 1343
rect 12621 1303 12679 1309
rect 11146 1272 11152 1284
rect 10980 1244 11152 1272
rect 11146 1232 11152 1244
rect 11204 1232 11210 1284
rect 12084 1272 12112 1303
rect 13170 1300 13176 1352
rect 13228 1340 13234 1352
rect 13265 1343 13323 1349
rect 13265 1340 13277 1343
rect 13228 1312 13277 1340
rect 13228 1300 13234 1312
rect 13265 1309 13277 1312
rect 13311 1309 13323 1343
rect 13265 1303 13323 1309
rect 13630 1300 13636 1352
rect 13688 1300 13694 1352
rect 13740 1340 13768 1380
rect 14645 1343 14703 1349
rect 14645 1340 14657 1343
rect 13740 1312 14657 1340
rect 14645 1309 14657 1312
rect 14691 1309 14703 1343
rect 14752 1340 14780 1380
rect 15289 1343 15347 1349
rect 15289 1340 15301 1343
rect 14752 1312 15301 1340
rect 14645 1303 14703 1309
rect 15289 1309 15301 1312
rect 15335 1309 15347 1343
rect 15289 1303 15347 1309
rect 14185 1275 14243 1281
rect 14185 1272 14197 1275
rect 11532 1244 12112 1272
rect 13096 1244 14197 1272
rect 11532 1216 11560 1244
rect 10594 1204 10600 1216
rect 9968 1176 10600 1204
rect 10594 1164 10600 1176
rect 10652 1164 10658 1216
rect 11238 1164 11244 1216
rect 11296 1164 11302 1216
rect 11514 1164 11520 1216
rect 11572 1164 11578 1216
rect 11698 1164 11704 1216
rect 11756 1164 11762 1216
rect 11885 1207 11943 1213
rect 11885 1173 11897 1207
rect 11931 1204 11943 1207
rect 13096 1204 13124 1244
rect 14185 1241 14197 1244
rect 14231 1241 14243 1275
rect 14185 1235 14243 1241
rect 14550 1232 14556 1284
rect 14608 1272 14614 1284
rect 15841 1275 15899 1281
rect 15841 1272 15853 1275
rect 14608 1244 15853 1272
rect 14608 1232 14614 1244
rect 15841 1241 15853 1244
rect 15887 1241 15899 1275
rect 16132 1272 16160 1380
rect 16206 1368 16212 1420
rect 16264 1408 16270 1420
rect 17420 1408 17448 1507
rect 18322 1504 18328 1556
rect 18380 1544 18386 1556
rect 24486 1544 24492 1556
rect 18380 1516 24492 1544
rect 18380 1504 18386 1516
rect 24486 1504 24492 1516
rect 24544 1504 24550 1556
rect 21266 1436 21272 1488
rect 21324 1476 21330 1488
rect 23753 1479 23811 1485
rect 23753 1476 23765 1479
rect 21324 1448 23765 1476
rect 21324 1436 21330 1448
rect 23753 1445 23765 1448
rect 23799 1445 23811 1479
rect 23753 1439 23811 1445
rect 19794 1408 19800 1420
rect 16264 1380 17448 1408
rect 17512 1380 19800 1408
rect 16264 1368 16270 1380
rect 16482 1300 16488 1352
rect 16540 1300 16546 1352
rect 16666 1300 16672 1352
rect 16724 1340 16730 1352
rect 16761 1343 16819 1349
rect 16761 1340 16773 1343
rect 16724 1312 16773 1340
rect 16724 1300 16730 1312
rect 16761 1309 16773 1312
rect 16807 1309 16819 1343
rect 16761 1303 16819 1309
rect 17218 1300 17224 1352
rect 17276 1340 17282 1352
rect 17313 1343 17371 1349
rect 17313 1340 17325 1343
rect 17276 1312 17325 1340
rect 17276 1300 17282 1312
rect 17313 1309 17325 1312
rect 17359 1309 17371 1343
rect 17512 1340 17540 1380
rect 19794 1368 19800 1380
rect 19852 1368 19858 1420
rect 17313 1303 17371 1309
rect 17420 1312 17540 1340
rect 17420 1272 17448 1312
rect 17678 1300 17684 1352
rect 17736 1340 17742 1352
rect 17865 1343 17923 1349
rect 17865 1340 17877 1343
rect 17736 1312 17877 1340
rect 17736 1300 17742 1312
rect 17865 1309 17877 1312
rect 17911 1309 17923 1343
rect 17865 1303 17923 1309
rect 18506 1300 18512 1352
rect 18564 1340 18570 1352
rect 19061 1343 19119 1349
rect 19061 1340 19073 1343
rect 18564 1312 19073 1340
rect 18564 1300 18570 1312
rect 19061 1309 19073 1312
rect 19107 1309 19119 1343
rect 19061 1303 19119 1309
rect 19426 1300 19432 1352
rect 19484 1300 19490 1352
rect 20165 1343 20223 1349
rect 20165 1309 20177 1343
rect 20211 1340 20223 1343
rect 20346 1340 20352 1352
rect 20211 1312 20352 1340
rect 20211 1309 20223 1312
rect 20165 1303 20223 1309
rect 20346 1300 20352 1312
rect 20404 1300 20410 1352
rect 20438 1300 20444 1352
rect 20496 1300 20502 1352
rect 20990 1300 20996 1352
rect 21048 1340 21054 1352
rect 22005 1343 22063 1349
rect 22005 1340 22017 1343
rect 21048 1312 22017 1340
rect 21048 1300 21054 1312
rect 22005 1309 22017 1312
rect 22051 1309 22063 1343
rect 22005 1303 22063 1309
rect 22097 1343 22155 1349
rect 22097 1309 22109 1343
rect 22143 1340 22155 1343
rect 23014 1340 23020 1352
rect 22143 1312 23020 1340
rect 22143 1309 22155 1312
rect 22097 1303 22155 1309
rect 23014 1300 23020 1312
rect 23072 1300 23078 1352
rect 19610 1272 19616 1284
rect 16132 1244 17448 1272
rect 18892 1244 19616 1272
rect 15841 1235 15899 1241
rect 11931 1176 13124 1204
rect 11931 1173 11943 1176
rect 11885 1167 11943 1173
rect 13446 1164 13452 1216
rect 13504 1164 13510 1216
rect 13630 1164 13636 1216
rect 13688 1204 13694 1216
rect 13817 1207 13875 1213
rect 13817 1204 13829 1207
rect 13688 1176 13829 1204
rect 13688 1164 13694 1176
rect 13817 1173 13829 1176
rect 13863 1173 13875 1207
rect 13817 1167 13875 1173
rect 13998 1164 14004 1216
rect 14056 1204 14062 1216
rect 14829 1207 14887 1213
rect 14829 1204 14841 1207
rect 14056 1176 14841 1204
rect 14056 1164 14062 1176
rect 14829 1173 14841 1176
rect 14875 1173 14887 1207
rect 14829 1167 14887 1173
rect 16482 1164 16488 1216
rect 16540 1204 16546 1216
rect 18892 1213 18920 1244
rect 19610 1232 19616 1244
rect 19668 1232 19674 1284
rect 21266 1232 21272 1284
rect 21324 1232 21330 1284
rect 22186 1232 22192 1284
rect 22244 1232 22250 1284
rect 22462 1232 22468 1284
rect 22520 1232 22526 1284
rect 17957 1207 18015 1213
rect 17957 1204 17969 1207
rect 16540 1176 17969 1204
rect 16540 1164 16546 1176
rect 17957 1173 17969 1176
rect 18003 1173 18015 1207
rect 17957 1167 18015 1173
rect 18877 1207 18935 1213
rect 18877 1173 18889 1207
rect 18923 1173 18935 1207
rect 18877 1167 18935 1173
rect 20898 1164 20904 1216
rect 20956 1204 20962 1216
rect 21821 1207 21879 1213
rect 21821 1204 21833 1207
rect 20956 1176 21833 1204
rect 20956 1164 20962 1176
rect 21821 1173 21833 1176
rect 21867 1173 21879 1207
rect 22204 1204 22232 1232
rect 22281 1207 22339 1213
rect 22281 1204 22293 1207
rect 22204 1176 22293 1204
rect 21821 1167 21879 1173
rect 22281 1173 22293 1176
rect 22327 1173 22339 1207
rect 22281 1167 22339 1173
rect 1104 1114 25000 1136
rect 1104 1062 6884 1114
rect 6936 1062 6948 1114
rect 7000 1062 7012 1114
rect 7064 1062 7076 1114
rect 7128 1062 7140 1114
rect 7192 1062 12818 1114
rect 12870 1062 12882 1114
rect 12934 1062 12946 1114
rect 12998 1062 13010 1114
rect 13062 1062 13074 1114
rect 13126 1062 18752 1114
rect 18804 1062 18816 1114
rect 18868 1062 18880 1114
rect 18932 1062 18944 1114
rect 18996 1062 19008 1114
rect 19060 1062 24686 1114
rect 24738 1062 24750 1114
rect 24802 1062 24814 1114
rect 24866 1062 24878 1114
rect 24930 1062 24942 1114
rect 24994 1062 25000 1114
rect 1104 1040 25000 1062
rect 5074 960 5080 1012
rect 5132 1000 5138 1012
rect 8294 1000 8300 1012
rect 5132 972 8300 1000
rect 5132 960 5138 972
rect 8294 960 8300 972
rect 8352 960 8358 1012
rect 8662 960 8668 1012
rect 8720 960 8726 1012
rect 11238 960 11244 1012
rect 11296 1000 11302 1012
rect 12894 1000 12900 1012
rect 11296 972 12900 1000
rect 11296 960 11302 972
rect 12894 960 12900 972
rect 12952 960 12958 1012
rect 14366 960 14372 1012
rect 14424 1000 14430 1012
rect 21266 1000 21272 1012
rect 14424 972 21272 1000
rect 14424 960 14430 972
rect 21266 960 21272 972
rect 21324 960 21330 1012
rect 3878 892 3884 944
rect 3936 932 3942 944
rect 7466 932 7472 944
rect 3936 904 7472 932
rect 3936 892 3942 904
rect 7466 892 7472 904
rect 7524 892 7530 944
rect 6454 824 6460 876
rect 6512 864 6518 876
rect 8680 864 8708 960
rect 8938 892 8944 944
rect 8996 932 9002 944
rect 11330 932 11336 944
rect 8996 904 11336 932
rect 8996 892 9002 904
rect 11330 892 11336 904
rect 11388 892 11394 944
rect 19426 892 19432 944
rect 19484 932 19490 944
rect 22830 932 22836 944
rect 19484 904 22836 932
rect 19484 892 19490 904
rect 22830 892 22836 904
rect 22888 892 22894 944
rect 6512 836 8708 864
rect 6512 824 6518 836
rect 566 756 572 808
rect 624 796 630 808
rect 11514 796 11520 808
rect 624 768 11520 796
rect 624 756 630 768
rect 11514 756 11520 768
rect 11572 756 11578 808
rect 6178 688 6184 740
rect 6236 728 6242 740
rect 7098 728 7104 740
rect 6236 700 7104 728
rect 6236 688 6242 700
rect 7098 688 7104 700
rect 7156 688 7162 740
rect 7558 688 7564 740
rect 7616 688 7622 740
rect 9030 688 9036 740
rect 9088 728 9094 740
rect 9674 728 9680 740
rect 9088 700 9680 728
rect 9088 688 9094 700
rect 9674 688 9680 700
rect 9732 688 9738 740
rect 7576 660 7604 688
rect 12710 660 12716 672
rect 7576 632 12716 660
rect 12710 620 12716 632
rect 12768 620 12774 672
rect 21266 620 21272 672
rect 21324 660 21330 672
rect 22462 660 22468 672
rect 21324 632 22468 660
rect 21324 620 21330 632
rect 22462 620 22468 632
rect 22520 620 22526 672
rect 6362 552 6368 604
rect 6420 592 6426 604
rect 9582 592 9588 604
rect 6420 564 9588 592
rect 6420 552 6426 564
rect 9582 552 9588 564
rect 9640 552 9646 604
rect 5810 484 5816 536
rect 5868 524 5874 536
rect 9030 524 9036 536
rect 5868 496 9036 524
rect 5868 484 5874 496
rect 9030 484 9036 496
rect 9088 484 9094 536
rect 6730 348 6736 400
rect 6788 388 6794 400
rect 11422 388 11428 400
rect 6788 360 11428 388
rect 6788 348 6794 360
rect 11422 348 11428 360
rect 11480 348 11486 400
<< via1 >>
rect 17224 44888 17276 44940
rect 18512 44888 18564 44940
rect 8944 44752 8996 44804
rect 9588 44752 9640 44804
rect 3516 44004 3568 44056
rect 4620 44004 4672 44056
rect 3608 43800 3660 43852
rect 6368 43800 6420 43852
rect 4804 43732 4856 43784
rect 17040 43732 17092 43784
rect 18052 43732 18104 43784
rect 3424 43664 3476 43716
rect 10508 43664 10560 43716
rect 17592 43664 17644 43716
rect 18604 43664 18656 43716
rect 1768 43596 1820 43648
rect 3976 43596 4028 43648
rect 5264 43596 5316 43648
rect 9128 43596 9180 43648
rect 16856 43596 16908 43648
rect 17316 43596 17368 43648
rect 18328 43596 18380 43648
rect 19984 43596 20036 43648
rect 22652 43596 22704 43648
rect 6884 43494 6936 43546
rect 6948 43494 7000 43546
rect 7012 43494 7064 43546
rect 7076 43494 7128 43546
rect 7140 43494 7192 43546
rect 12818 43494 12870 43546
rect 12882 43494 12934 43546
rect 12946 43494 12998 43546
rect 13010 43494 13062 43546
rect 13074 43494 13126 43546
rect 18752 43494 18804 43546
rect 18816 43494 18868 43546
rect 18880 43494 18932 43546
rect 18944 43494 18996 43546
rect 19008 43494 19060 43546
rect 24686 43494 24738 43546
rect 24750 43494 24802 43546
rect 24814 43494 24866 43546
rect 24878 43494 24930 43546
rect 24942 43494 24994 43546
rect 2136 43392 2188 43444
rect 2412 43435 2464 43444
rect 2412 43401 2421 43435
rect 2421 43401 2455 43435
rect 2455 43401 2464 43435
rect 2412 43392 2464 43401
rect 2964 43435 3016 43444
rect 2964 43401 2973 43435
rect 2973 43401 3007 43435
rect 3007 43401 3016 43435
rect 2964 43392 3016 43401
rect 3516 43435 3568 43444
rect 3516 43401 3525 43435
rect 3525 43401 3559 43435
rect 3559 43401 3568 43435
rect 3516 43392 3568 43401
rect 3976 43392 4028 43444
rect 5172 43392 5224 43444
rect 5448 43392 5500 43444
rect 5724 43435 5776 43444
rect 5724 43401 5733 43435
rect 5733 43401 5767 43435
rect 5767 43401 5776 43435
rect 5724 43392 5776 43401
rect 6828 43392 6880 43444
rect 7932 43392 7984 43444
rect 8208 43392 8260 43444
rect 8944 43392 8996 43444
rect 9036 43392 9088 43444
rect 9864 43392 9916 43444
rect 10508 43435 10560 43444
rect 10508 43401 10517 43435
rect 10517 43401 10551 43435
rect 10551 43401 10560 43435
rect 10508 43392 10560 43401
rect 13176 43392 13228 43444
rect 1676 43256 1728 43308
rect 1768 43299 1820 43308
rect 1768 43265 1777 43299
rect 1777 43265 1811 43299
rect 1811 43265 1820 43299
rect 1768 43256 1820 43265
rect 2872 43299 2924 43308
rect 2872 43265 2881 43299
rect 2881 43265 2915 43299
rect 2915 43265 2924 43299
rect 2872 43256 2924 43265
rect 3608 43256 3660 43308
rect 4160 43299 4212 43308
rect 4160 43265 4169 43299
rect 4169 43265 4203 43299
rect 4203 43265 4212 43299
rect 4160 43256 4212 43265
rect 4528 43299 4580 43308
rect 4528 43265 4537 43299
rect 4537 43265 4571 43299
rect 4571 43265 4580 43299
rect 4528 43256 4580 43265
rect 4620 43299 4672 43308
rect 4620 43265 4629 43299
rect 4629 43265 4663 43299
rect 4663 43265 4672 43299
rect 4620 43256 4672 43265
rect 5448 43256 5500 43308
rect 11244 43324 11296 43376
rect 12440 43367 12492 43376
rect 12440 43333 12449 43367
rect 12449 43333 12483 43367
rect 12483 43333 12492 43367
rect 12440 43324 12492 43333
rect 12624 43324 12676 43376
rect 13452 43324 13504 43376
rect 16856 43435 16908 43444
rect 16856 43401 16865 43435
rect 16865 43401 16899 43435
rect 16899 43401 16908 43435
rect 16856 43392 16908 43401
rect 14740 43367 14792 43376
rect 14740 43333 14749 43367
rect 14749 43333 14783 43367
rect 14783 43333 14792 43367
rect 14740 43324 14792 43333
rect 14832 43324 14884 43376
rect 15568 43367 15620 43376
rect 15568 43333 15577 43367
rect 15577 43333 15611 43367
rect 15611 43333 15620 43367
rect 15568 43324 15620 43333
rect 15660 43324 15712 43376
rect 16120 43324 16172 43376
rect 16396 43324 16448 43376
rect 17684 43392 17736 43444
rect 17868 43392 17920 43444
rect 20444 43435 20496 43444
rect 20444 43401 20453 43435
rect 20453 43401 20487 43435
rect 20487 43401 20496 43435
rect 20444 43392 20496 43401
rect 20628 43392 20680 43444
rect 21364 43392 21416 43444
rect 6552 43299 6604 43308
rect 6552 43265 6561 43299
rect 6561 43265 6595 43299
rect 6595 43265 6604 43299
rect 6552 43256 6604 43265
rect 7472 43256 7524 43308
rect 8300 43256 8352 43308
rect 6368 43188 6420 43240
rect 5540 43052 5592 43104
rect 9956 43299 10008 43308
rect 9956 43265 9965 43299
rect 9965 43265 9999 43299
rect 9999 43265 10008 43299
rect 9956 43256 10008 43265
rect 10324 43299 10376 43308
rect 10324 43265 10333 43299
rect 10333 43265 10367 43299
rect 10367 43265 10376 43299
rect 10324 43256 10376 43265
rect 10692 43299 10744 43308
rect 10692 43265 10701 43299
rect 10701 43265 10735 43299
rect 10735 43265 10744 43299
rect 10692 43256 10744 43265
rect 11060 43299 11112 43308
rect 11060 43265 11069 43299
rect 11069 43265 11103 43299
rect 11103 43265 11112 43299
rect 11060 43256 11112 43265
rect 12072 43299 12124 43308
rect 12072 43265 12081 43299
rect 12081 43265 12115 43299
rect 12115 43265 12124 43299
rect 12072 43256 12124 43265
rect 12164 43256 12216 43308
rect 17224 43299 17276 43308
rect 17224 43265 17233 43299
rect 17233 43265 17267 43299
rect 17267 43265 17276 43299
rect 17224 43256 17276 43265
rect 17316 43256 17368 43308
rect 18236 43324 18288 43376
rect 13636 43188 13688 43240
rect 16764 43188 16816 43240
rect 18052 43299 18104 43308
rect 18052 43265 18061 43299
rect 18061 43265 18095 43299
rect 18095 43265 18104 43299
rect 18052 43256 18104 43265
rect 18328 43299 18380 43308
rect 18328 43265 18337 43299
rect 18337 43265 18371 43299
rect 18371 43265 18380 43299
rect 18328 43256 18380 43265
rect 17960 43188 18012 43240
rect 18604 43299 18656 43308
rect 18604 43265 18613 43299
rect 18613 43265 18647 43299
rect 18647 43265 18656 43299
rect 18604 43256 18656 43265
rect 19432 43299 19484 43308
rect 19432 43265 19441 43299
rect 19441 43265 19475 43299
rect 19475 43265 19484 43299
rect 19432 43256 19484 43265
rect 21272 43324 21324 43376
rect 21456 43324 21508 43376
rect 22652 43392 22704 43444
rect 23388 43392 23440 43444
rect 18512 43188 18564 43240
rect 19248 43188 19300 43240
rect 20352 43299 20404 43308
rect 20352 43265 20361 43299
rect 20361 43265 20395 43299
rect 20395 43265 20404 43299
rect 20352 43256 20404 43265
rect 20904 43299 20956 43308
rect 20904 43265 20913 43299
rect 20913 43265 20947 43299
rect 20947 43265 20956 43299
rect 20904 43256 20956 43265
rect 21088 43256 21140 43308
rect 21548 43256 21600 43308
rect 22100 43256 22152 43308
rect 22560 43256 22612 43308
rect 23388 43256 23440 43308
rect 23112 43188 23164 43240
rect 10324 43120 10376 43172
rect 11796 43163 11848 43172
rect 11796 43129 11805 43163
rect 11805 43129 11839 43163
rect 11839 43129 11848 43163
rect 11796 43120 11848 43129
rect 13084 43120 13136 43172
rect 14924 43163 14976 43172
rect 14924 43129 14933 43163
rect 14933 43129 14967 43163
rect 14967 43129 14976 43163
rect 14924 43120 14976 43129
rect 15292 43163 15344 43172
rect 15292 43129 15301 43163
rect 15301 43129 15335 43163
rect 15335 43129 15344 43163
rect 15292 43120 15344 43129
rect 16120 43163 16172 43172
rect 16120 43129 16129 43163
rect 16129 43129 16163 43163
rect 16163 43129 16172 43163
rect 16120 43120 16172 43129
rect 17408 43120 17460 43172
rect 17500 43120 17552 43172
rect 20076 43120 20128 43172
rect 9772 43052 9824 43104
rect 10416 43052 10468 43104
rect 10876 43095 10928 43104
rect 10876 43061 10885 43095
rect 10885 43061 10919 43095
rect 10919 43061 10928 43095
rect 10876 43052 10928 43061
rect 11244 43095 11296 43104
rect 11244 43061 11253 43095
rect 11253 43061 11287 43095
rect 11287 43061 11296 43095
rect 11244 43052 11296 43061
rect 12256 43095 12308 43104
rect 12256 43061 12265 43095
rect 12265 43061 12299 43095
rect 12299 43061 12308 43095
rect 12256 43052 12308 43061
rect 12900 43095 12952 43104
rect 12900 43061 12909 43095
rect 12909 43061 12943 43095
rect 12943 43061 12952 43095
rect 12900 43052 12952 43061
rect 13820 43095 13872 43104
rect 13820 43061 13829 43095
rect 13829 43061 13863 43095
rect 13863 43061 13872 43095
rect 13820 43052 13872 43061
rect 14280 43095 14332 43104
rect 14280 43061 14289 43095
rect 14289 43061 14323 43095
rect 14323 43061 14332 43095
rect 14280 43052 14332 43061
rect 15660 43095 15712 43104
rect 15660 43061 15669 43095
rect 15669 43061 15703 43095
rect 15703 43061 15712 43095
rect 15660 43052 15712 43061
rect 17592 43052 17644 43104
rect 18052 43052 18104 43104
rect 19340 43052 19392 43104
rect 20996 43052 21048 43104
rect 21916 43052 21968 43104
rect 3917 42950 3969 43002
rect 3981 42950 4033 43002
rect 4045 42950 4097 43002
rect 4109 42950 4161 43002
rect 4173 42950 4225 43002
rect 9851 42950 9903 43002
rect 9915 42950 9967 43002
rect 9979 42950 10031 43002
rect 10043 42950 10095 43002
rect 10107 42950 10159 43002
rect 15785 42950 15837 43002
rect 15849 42950 15901 43002
rect 15913 42950 15965 43002
rect 15977 42950 16029 43002
rect 16041 42950 16093 43002
rect 21719 42950 21771 43002
rect 21783 42950 21835 43002
rect 21847 42950 21899 43002
rect 21911 42950 21963 43002
rect 21975 42950 22027 43002
rect 3332 42891 3384 42900
rect 3332 42857 3341 42891
rect 3341 42857 3375 42891
rect 3375 42857 3384 42891
rect 3332 42848 3384 42857
rect 4344 42891 4396 42900
rect 4344 42857 4353 42891
rect 4353 42857 4387 42891
rect 4387 42857 4396 42891
rect 4344 42848 4396 42857
rect 6092 42891 6144 42900
rect 6092 42857 6101 42891
rect 6101 42857 6135 42891
rect 6135 42857 6144 42891
rect 6092 42848 6144 42857
rect 6644 42891 6696 42900
rect 6644 42857 6653 42891
rect 6653 42857 6687 42891
rect 6687 42857 6696 42891
rect 6644 42848 6696 42857
rect 7196 42891 7248 42900
rect 7196 42857 7205 42891
rect 7205 42857 7239 42891
rect 7239 42857 7248 42891
rect 7196 42848 7248 42857
rect 8300 42848 8352 42900
rect 2688 42712 2740 42764
rect 4528 42644 4580 42696
rect 1400 42619 1452 42628
rect 1400 42585 1409 42619
rect 1409 42585 1443 42619
rect 1443 42585 1452 42619
rect 1400 42576 1452 42585
rect 2044 42576 2096 42628
rect 3056 42576 3108 42628
rect 3240 42619 3292 42628
rect 3240 42585 3249 42619
rect 3249 42585 3283 42619
rect 3283 42585 3292 42619
rect 3240 42576 3292 42585
rect 4988 42712 5040 42764
rect 8760 42712 8812 42764
rect 13636 42848 13688 42900
rect 9772 42780 9824 42832
rect 4712 42644 4764 42696
rect 5540 42687 5592 42696
rect 5540 42653 5549 42687
rect 5549 42653 5583 42687
rect 5583 42653 5592 42687
rect 5540 42644 5592 42653
rect 7564 42687 7616 42696
rect 7564 42653 7573 42687
rect 7573 42653 7607 42687
rect 7607 42653 7616 42687
rect 7564 42644 7616 42653
rect 8116 42687 8168 42696
rect 8116 42653 8125 42687
rect 8125 42653 8159 42687
rect 8159 42653 8168 42687
rect 8116 42644 8168 42653
rect 9312 42712 9364 42764
rect 3792 42508 3844 42560
rect 6000 42619 6052 42628
rect 6000 42585 6009 42619
rect 6009 42585 6043 42619
rect 6043 42585 6052 42619
rect 6000 42576 6052 42585
rect 6736 42576 6788 42628
rect 7288 42576 7340 42628
rect 7656 42576 7708 42628
rect 7840 42576 7892 42628
rect 9128 42687 9180 42696
rect 9128 42653 9137 42687
rect 9137 42653 9171 42687
rect 9171 42653 9180 42687
rect 9128 42644 9180 42653
rect 9496 42619 9548 42628
rect 9496 42585 9505 42619
rect 9505 42585 9539 42619
rect 9539 42585 9548 42619
rect 9496 42576 9548 42585
rect 9680 42576 9732 42628
rect 5540 42508 5592 42560
rect 6276 42508 6328 42560
rect 7932 42551 7984 42560
rect 7932 42517 7941 42551
rect 7941 42517 7975 42551
rect 7975 42517 7984 42551
rect 7932 42508 7984 42517
rect 8300 42508 8352 42560
rect 9588 42508 9640 42560
rect 10324 42644 10376 42696
rect 10508 42687 10560 42696
rect 10508 42653 10517 42687
rect 10517 42653 10551 42687
rect 10551 42653 10560 42687
rect 10508 42644 10560 42653
rect 10876 42687 10928 42696
rect 10876 42653 10885 42687
rect 10885 42653 10919 42687
rect 10919 42653 10928 42687
rect 10876 42644 10928 42653
rect 13544 42712 13596 42764
rect 13820 42712 13872 42764
rect 17316 42848 17368 42900
rect 17408 42848 17460 42900
rect 18604 42823 18656 42832
rect 18604 42789 18613 42823
rect 18613 42789 18647 42823
rect 18647 42789 18656 42823
rect 18604 42780 18656 42789
rect 11612 42687 11664 42696
rect 11612 42653 11621 42687
rect 11621 42653 11655 42687
rect 11655 42653 11664 42687
rect 11612 42644 11664 42653
rect 11888 42687 11940 42696
rect 11888 42653 11897 42687
rect 11897 42653 11931 42687
rect 11931 42653 11940 42687
rect 11888 42644 11940 42653
rect 12348 42687 12400 42696
rect 12348 42653 12357 42687
rect 12357 42653 12391 42687
rect 12391 42653 12400 42687
rect 12348 42644 12400 42653
rect 12716 42644 12768 42696
rect 14096 42687 14148 42696
rect 14096 42653 14105 42687
rect 14105 42653 14139 42687
rect 14139 42653 14148 42687
rect 14096 42644 14148 42653
rect 14372 42687 14424 42696
rect 14372 42653 14381 42687
rect 14381 42653 14415 42687
rect 14415 42653 14424 42687
rect 14372 42644 14424 42653
rect 15108 42687 15160 42696
rect 15108 42653 15117 42687
rect 15117 42653 15151 42687
rect 15151 42653 15160 42687
rect 15108 42644 15160 42653
rect 15384 42687 15436 42696
rect 15384 42653 15393 42687
rect 15393 42653 15427 42687
rect 15427 42653 15436 42687
rect 15384 42644 15436 42653
rect 16488 42644 16540 42696
rect 10784 42576 10836 42628
rect 11152 42551 11204 42560
rect 11152 42517 11161 42551
rect 11161 42517 11195 42551
rect 11195 42517 11204 42551
rect 11152 42508 11204 42517
rect 11336 42508 11388 42560
rect 12532 42551 12584 42560
rect 12532 42517 12541 42551
rect 12541 42517 12575 42551
rect 12575 42517 12584 42551
rect 12532 42508 12584 42517
rect 13360 42576 13412 42628
rect 13268 42508 13320 42560
rect 14832 42551 14884 42560
rect 14832 42517 14841 42551
rect 14841 42517 14875 42551
rect 14875 42517 14884 42551
rect 14832 42508 14884 42517
rect 15108 42508 15160 42560
rect 15292 42551 15344 42560
rect 15292 42517 15301 42551
rect 15301 42517 15335 42551
rect 15335 42517 15344 42551
rect 15292 42508 15344 42517
rect 16396 42576 16448 42628
rect 17500 42644 17552 42696
rect 17868 42644 17920 42696
rect 18052 42644 18104 42696
rect 20260 42848 20312 42900
rect 21548 42848 21600 42900
rect 22928 42848 22980 42900
rect 19708 42780 19760 42832
rect 20076 42712 20128 42764
rect 20168 42712 20220 42764
rect 19616 42644 19668 42696
rect 21364 42687 21416 42696
rect 21364 42653 21373 42687
rect 21373 42653 21407 42687
rect 21407 42653 21416 42687
rect 21364 42644 21416 42653
rect 22284 42712 22336 42764
rect 23572 42712 23624 42764
rect 24124 42644 24176 42696
rect 19248 42619 19300 42628
rect 19248 42585 19257 42619
rect 19257 42585 19291 42619
rect 19291 42585 19300 42619
rect 19248 42576 19300 42585
rect 20996 42619 21048 42628
rect 20996 42585 21005 42619
rect 21005 42585 21039 42619
rect 21039 42585 21048 42619
rect 20996 42576 21048 42585
rect 16764 42551 16816 42560
rect 16764 42517 16773 42551
rect 16773 42517 16807 42551
rect 16807 42517 16816 42551
rect 16764 42508 16816 42517
rect 17224 42551 17276 42560
rect 17224 42517 17233 42551
rect 17233 42517 17267 42551
rect 17267 42517 17276 42551
rect 17224 42508 17276 42517
rect 17316 42508 17368 42560
rect 17776 42551 17828 42560
rect 17776 42517 17785 42551
rect 17785 42517 17819 42551
rect 17819 42517 17828 42551
rect 17776 42508 17828 42517
rect 18052 42551 18104 42560
rect 18052 42517 18061 42551
rect 18061 42517 18095 42551
rect 18095 42517 18104 42551
rect 18052 42508 18104 42517
rect 18328 42551 18380 42560
rect 18328 42517 18337 42551
rect 18337 42517 18371 42551
rect 18371 42517 18380 42551
rect 18328 42508 18380 42517
rect 18420 42508 18472 42560
rect 20720 42508 20772 42560
rect 22376 42576 22428 42628
rect 22836 42576 22888 42628
rect 23848 42576 23900 42628
rect 25044 42508 25096 42560
rect 6884 42406 6936 42458
rect 6948 42406 7000 42458
rect 7012 42406 7064 42458
rect 7076 42406 7128 42458
rect 7140 42406 7192 42458
rect 12818 42406 12870 42458
rect 12882 42406 12934 42458
rect 12946 42406 12998 42458
rect 13010 42406 13062 42458
rect 13074 42406 13126 42458
rect 18752 42406 18804 42458
rect 18816 42406 18868 42458
rect 18880 42406 18932 42458
rect 18944 42406 18996 42458
rect 19008 42406 19060 42458
rect 24686 42406 24738 42458
rect 24750 42406 24802 42458
rect 24814 42406 24866 42458
rect 24878 42406 24930 42458
rect 24942 42406 24994 42458
rect 1032 42304 1084 42356
rect 1584 42236 1636 42288
rect 3240 42304 3292 42356
rect 5632 42304 5684 42356
rect 6552 42304 6604 42356
rect 7380 42304 7432 42356
rect 8208 42304 8260 42356
rect 8852 42304 8904 42356
rect 10784 42304 10836 42356
rect 11152 42304 11204 42356
rect 1400 42211 1452 42220
rect 1400 42177 1409 42211
rect 1409 42177 1443 42211
rect 1443 42177 1452 42211
rect 1400 42168 1452 42177
rect 2504 42211 2556 42220
rect 2504 42177 2513 42211
rect 2513 42177 2547 42211
rect 2547 42177 2556 42211
rect 2504 42168 2556 42177
rect 3608 42211 3660 42220
rect 3608 42177 3617 42211
rect 3617 42177 3651 42211
rect 3651 42177 3660 42211
rect 3608 42168 3660 42177
rect 3792 42168 3844 42220
rect 4436 42168 4488 42220
rect 2228 42143 2280 42152
rect 2228 42109 2237 42143
rect 2237 42109 2271 42143
rect 2271 42109 2280 42143
rect 2228 42100 2280 42109
rect 5816 42236 5868 42288
rect 6092 42168 6144 42220
rect 6184 42211 6236 42220
rect 6184 42177 6193 42211
rect 6193 42177 6227 42211
rect 6227 42177 6236 42211
rect 6184 42168 6236 42177
rect 6644 42211 6696 42220
rect 6644 42177 6653 42211
rect 6653 42177 6687 42211
rect 6687 42177 6696 42211
rect 6644 42168 6696 42177
rect 7196 42168 7248 42220
rect 8300 42236 8352 42288
rect 9404 42236 9456 42288
rect 9588 42236 9640 42288
rect 7748 42168 7800 42220
rect 8024 42168 8076 42220
rect 8392 42211 8444 42220
rect 8392 42177 8401 42211
rect 8401 42177 8435 42211
rect 8435 42177 8444 42211
rect 8392 42168 8444 42177
rect 8668 42168 8720 42220
rect 12532 42304 12584 42356
rect 17224 42304 17276 42356
rect 17316 42304 17368 42356
rect 16212 42211 16264 42220
rect 16212 42177 16221 42211
rect 16221 42177 16255 42211
rect 16255 42177 16264 42211
rect 16212 42168 16264 42177
rect 17684 42304 17736 42356
rect 17776 42304 17828 42356
rect 18052 42304 18104 42356
rect 18328 42304 18380 42356
rect 18420 42236 18472 42288
rect 18604 42211 18656 42220
rect 18604 42177 18613 42211
rect 18613 42177 18647 42211
rect 18647 42177 18656 42211
rect 18604 42168 18656 42177
rect 18880 42168 18932 42220
rect 19340 42279 19392 42288
rect 19340 42245 19349 42279
rect 19349 42245 19383 42279
rect 19383 42245 19392 42279
rect 19340 42236 19392 42245
rect 19616 42347 19668 42356
rect 19616 42313 19625 42347
rect 19625 42313 19659 42347
rect 19659 42313 19668 42347
rect 19616 42304 19668 42313
rect 19984 42304 20036 42356
rect 20352 42304 20404 42356
rect 20904 42304 20956 42356
rect 23020 42304 23072 42356
rect 24216 42304 24268 42356
rect 20260 42236 20312 42288
rect 22100 42236 22152 42288
rect 23756 42236 23808 42288
rect 19156 42168 19208 42220
rect 19984 42168 20036 42220
rect 20444 42211 20496 42220
rect 20444 42177 20453 42211
rect 20453 42177 20487 42211
rect 20487 42177 20496 42211
rect 20444 42168 20496 42177
rect 480 42032 532 42084
rect 7840 42100 7892 42152
rect 9772 42100 9824 42152
rect 1308 41964 1360 42016
rect 4528 42032 4580 42084
rect 5908 42032 5960 42084
rect 8208 42032 8260 42084
rect 16396 42032 16448 42084
rect 16948 42075 17000 42084
rect 16948 42041 16957 42075
rect 16957 42041 16991 42075
rect 16991 42041 17000 42075
rect 16948 42032 17000 42041
rect 17316 42075 17368 42084
rect 17316 42041 17325 42075
rect 17325 42041 17359 42075
rect 17359 42041 17368 42075
rect 17316 42032 17368 42041
rect 18420 42075 18472 42084
rect 18420 42041 18429 42075
rect 18429 42041 18463 42075
rect 18463 42041 18472 42075
rect 18420 42032 18472 42041
rect 4804 42007 4856 42016
rect 4804 41973 4813 42007
rect 4813 41973 4847 42007
rect 4847 41973 4856 42007
rect 4804 41964 4856 41973
rect 5724 42007 5776 42016
rect 5724 41973 5733 42007
rect 5733 41973 5767 42007
rect 5767 41973 5776 42007
rect 5724 41964 5776 41973
rect 6276 41964 6328 42016
rect 6736 42007 6788 42016
rect 6736 41973 6745 42007
rect 6745 41973 6779 42007
rect 6779 41973 6788 42007
rect 6736 41964 6788 41973
rect 7196 41964 7248 42016
rect 7380 41964 7432 42016
rect 8300 41964 8352 42016
rect 9036 41964 9088 42016
rect 16304 42007 16356 42016
rect 16304 41973 16313 42007
rect 16313 41973 16347 42007
rect 16347 41973 16356 42007
rect 16304 41964 16356 41973
rect 17592 42007 17644 42016
rect 17592 41973 17601 42007
rect 17601 41973 17635 42007
rect 17635 41973 17644 42007
rect 17592 41964 17644 41973
rect 17960 42007 18012 42016
rect 17960 41973 17969 42007
rect 17969 41973 18003 42007
rect 18003 41973 18012 42007
rect 17960 41964 18012 41973
rect 18696 42007 18748 42016
rect 18696 41973 18705 42007
rect 18705 41973 18739 42007
rect 18739 41973 18748 42007
rect 18696 41964 18748 41973
rect 19064 42007 19116 42016
rect 19064 41973 19073 42007
rect 19073 41973 19107 42007
rect 19107 41973 19116 42007
rect 19064 41964 19116 41973
rect 19340 41964 19392 42016
rect 19892 41964 19944 42016
rect 22468 42211 22520 42220
rect 22468 42177 22477 42211
rect 22477 42177 22511 42211
rect 22511 42177 22520 42211
rect 22468 42168 22520 42177
rect 22560 42168 22612 42220
rect 23572 42211 23624 42220
rect 23572 42177 23581 42211
rect 23581 42177 23615 42211
rect 23615 42177 23624 42211
rect 23572 42168 23624 42177
rect 24032 42168 24084 42220
rect 24124 42211 24176 42220
rect 24124 42177 24133 42211
rect 24133 42177 24167 42211
rect 24167 42177 24176 42211
rect 24124 42168 24176 42177
rect 25044 42168 25096 42220
rect 23756 42100 23808 42152
rect 25596 42100 25648 42152
rect 25688 41964 25740 42016
rect 3917 41862 3969 41914
rect 3981 41862 4033 41914
rect 4045 41862 4097 41914
rect 4109 41862 4161 41914
rect 4173 41862 4225 41914
rect 9851 41862 9903 41914
rect 9915 41862 9967 41914
rect 9979 41862 10031 41914
rect 10043 41862 10095 41914
rect 10107 41862 10159 41914
rect 15785 41862 15837 41914
rect 15849 41862 15901 41914
rect 15913 41862 15965 41914
rect 15977 41862 16029 41914
rect 16041 41862 16093 41914
rect 21719 41862 21771 41914
rect 21783 41862 21835 41914
rect 21847 41862 21899 41914
rect 21911 41862 21963 41914
rect 21975 41862 22027 41914
rect 3792 41760 3844 41812
rect 3884 41760 3936 41812
rect 4620 41760 4672 41812
rect 5448 41803 5500 41812
rect 5448 41769 5457 41803
rect 5457 41769 5491 41803
rect 5491 41769 5500 41803
rect 5448 41760 5500 41769
rect 5724 41760 5776 41812
rect 5816 41803 5868 41812
rect 5816 41769 5825 41803
rect 5825 41769 5859 41803
rect 5859 41769 5868 41803
rect 5816 41760 5868 41769
rect 6000 41760 6052 41812
rect 6368 41760 6420 41812
rect 6736 41760 6788 41812
rect 6828 41803 6880 41812
rect 6828 41769 6837 41803
rect 6837 41769 6871 41803
rect 6871 41769 6880 41803
rect 6828 41760 6880 41769
rect 7288 41803 7340 41812
rect 7288 41769 7297 41803
rect 7297 41769 7331 41803
rect 7331 41769 7340 41803
rect 7288 41760 7340 41769
rect 7564 41760 7616 41812
rect 7932 41760 7984 41812
rect 8208 41760 8260 41812
rect 8300 41760 8352 41812
rect 8392 41803 8444 41812
rect 8392 41769 8401 41803
rect 8401 41769 8435 41803
rect 8435 41769 8444 41803
rect 8392 41760 8444 41769
rect 9128 41760 9180 41812
rect 756 41556 808 41608
rect 2412 41531 2464 41540
rect 2412 41497 2421 41531
rect 2421 41497 2455 41531
rect 2455 41497 2464 41531
rect 2412 41488 2464 41497
rect 2780 41420 2832 41472
rect 3700 41556 3752 41608
rect 3884 41599 3936 41608
rect 3884 41565 3893 41599
rect 3893 41565 3927 41599
rect 3927 41565 3936 41599
rect 3884 41556 3936 41565
rect 4528 41624 4580 41676
rect 4344 41599 4396 41608
rect 4344 41565 4353 41599
rect 4353 41565 4387 41599
rect 4387 41565 4396 41599
rect 4344 41556 4396 41565
rect 4620 41556 4672 41608
rect 5172 41599 5224 41608
rect 5172 41565 5181 41599
rect 5181 41565 5215 41599
rect 5215 41565 5224 41599
rect 5172 41556 5224 41565
rect 6000 41599 6052 41608
rect 6000 41565 6009 41599
rect 6009 41565 6043 41599
rect 6043 41565 6052 41599
rect 6000 41556 6052 41565
rect 6276 41556 6328 41608
rect 6736 41599 6788 41608
rect 6736 41565 6745 41599
rect 6745 41565 6779 41599
rect 6779 41565 6788 41599
rect 6736 41556 6788 41565
rect 8576 41692 8628 41744
rect 11336 41760 11388 41812
rect 16304 41760 16356 41812
rect 16396 41760 16448 41812
rect 16672 41760 16724 41812
rect 4160 41488 4212 41540
rect 4804 41488 4856 41540
rect 5908 41488 5960 41540
rect 6184 41488 6236 41540
rect 7472 41420 7524 41472
rect 9404 41463 9456 41472
rect 9404 41429 9413 41463
rect 9413 41429 9447 41463
rect 9447 41429 9456 41463
rect 9404 41420 9456 41429
rect 9772 41599 9824 41608
rect 9772 41565 9781 41599
rect 9781 41565 9815 41599
rect 9815 41565 9824 41599
rect 9772 41556 9824 41565
rect 18880 41803 18932 41812
rect 18880 41769 18889 41803
rect 18889 41769 18923 41803
rect 18923 41769 18932 41803
rect 18880 41760 18932 41769
rect 19340 41760 19392 41812
rect 19708 41760 19760 41812
rect 19984 41760 20036 41812
rect 20444 41760 20496 41812
rect 20996 41760 21048 41812
rect 18696 41556 18748 41608
rect 10048 41535 10073 41540
rect 10073 41535 10100 41540
rect 10048 41488 10100 41535
rect 10784 41463 10836 41472
rect 10784 41429 10793 41463
rect 10793 41429 10827 41463
rect 10827 41429 10836 41463
rect 10784 41420 10836 41429
rect 15108 41488 15160 41540
rect 19340 41556 19392 41608
rect 19524 41556 19576 41608
rect 19800 41624 19852 41676
rect 21456 41760 21508 41812
rect 21732 41803 21784 41812
rect 21732 41769 21741 41803
rect 21741 41769 21775 41803
rect 21775 41769 21784 41803
rect 21732 41760 21784 41769
rect 22284 41803 22336 41812
rect 22284 41769 22293 41803
rect 22293 41769 22327 41803
rect 22327 41769 22336 41803
rect 22284 41760 22336 41769
rect 23664 41760 23716 41812
rect 23940 41803 23992 41812
rect 23940 41769 23949 41803
rect 23949 41769 23983 41803
rect 23983 41769 23992 41803
rect 23940 41760 23992 41769
rect 24584 41760 24636 41812
rect 21548 41692 21600 41744
rect 19892 41556 19944 41608
rect 20628 41556 20680 41608
rect 21180 41599 21232 41608
rect 21180 41565 21189 41599
rect 21189 41565 21223 41599
rect 21223 41565 21232 41599
rect 21180 41556 21232 41565
rect 22008 41599 22060 41608
rect 22008 41565 22017 41599
rect 22017 41565 22051 41599
rect 22051 41565 22060 41599
rect 22008 41556 22060 41565
rect 15200 41420 15252 41472
rect 16212 41463 16264 41472
rect 16212 41429 16221 41463
rect 16221 41429 16255 41463
rect 16255 41429 16264 41463
rect 16212 41420 16264 41429
rect 18328 41463 18380 41472
rect 18328 41429 18337 41463
rect 18337 41429 18371 41463
rect 18371 41429 18380 41463
rect 18328 41420 18380 41429
rect 19156 41420 19208 41472
rect 20260 41420 20312 41472
rect 20352 41463 20404 41472
rect 20352 41429 20361 41463
rect 20361 41429 20395 41463
rect 20395 41429 20404 41463
rect 20352 41420 20404 41429
rect 20444 41420 20496 41472
rect 21640 41488 21692 41540
rect 22284 41420 22336 41472
rect 23296 41531 23348 41540
rect 23296 41497 23305 41531
rect 23305 41497 23339 41531
rect 23339 41497 23348 41531
rect 23296 41488 23348 41497
rect 23848 41531 23900 41540
rect 23848 41497 23857 41531
rect 23857 41497 23891 41531
rect 23891 41497 23900 41531
rect 23848 41488 23900 41497
rect 24492 41420 24544 41472
rect 6884 41318 6936 41370
rect 6948 41318 7000 41370
rect 7012 41318 7064 41370
rect 7076 41318 7128 41370
rect 7140 41318 7192 41370
rect 12818 41318 12870 41370
rect 12882 41318 12934 41370
rect 12946 41318 12998 41370
rect 13010 41318 13062 41370
rect 13074 41318 13126 41370
rect 18752 41318 18804 41370
rect 18816 41318 18868 41370
rect 18880 41318 18932 41370
rect 18944 41318 18996 41370
rect 19008 41318 19060 41370
rect 24686 41318 24738 41370
rect 24750 41318 24802 41370
rect 24814 41318 24866 41370
rect 24878 41318 24930 41370
rect 24942 41318 24994 41370
rect 204 41216 256 41268
rect 4160 41216 4212 41268
rect 4804 41216 4856 41268
rect 5264 41259 5316 41268
rect 5264 41225 5273 41259
rect 5273 41225 5307 41259
rect 5307 41225 5316 41259
rect 5264 41216 5316 41225
rect 5540 41259 5592 41268
rect 5540 41225 5549 41259
rect 5549 41225 5583 41259
rect 5583 41225 5592 41259
rect 5540 41216 5592 41225
rect 5816 41259 5868 41268
rect 5816 41225 5825 41259
rect 5825 41225 5859 41259
rect 5859 41225 5868 41259
rect 5816 41216 5868 41225
rect 6552 41216 6604 41268
rect 7840 41216 7892 41268
rect 8208 41216 8260 41268
rect 9220 41216 9272 41268
rect 9772 41216 9824 41268
rect 2136 41080 2188 41132
rect 2320 41123 2372 41132
rect 2320 41089 2329 41123
rect 2329 41089 2363 41123
rect 2363 41089 2372 41123
rect 2320 41080 2372 41089
rect 2688 41080 2740 41132
rect 3516 41080 3568 41132
rect 5080 41080 5132 41132
rect 2964 41012 3016 41064
rect 4436 41012 4488 41064
rect 4712 41012 4764 41064
rect 5448 41123 5500 41132
rect 5448 41089 5457 41123
rect 5457 41089 5491 41123
rect 5491 41089 5500 41123
rect 5448 41080 5500 41089
rect 5540 41080 5592 41132
rect 6552 41123 6604 41132
rect 6552 41089 6561 41123
rect 6561 41089 6595 41123
rect 6595 41089 6604 41123
rect 6552 41080 6604 41089
rect 6276 41012 6328 41064
rect 6368 41012 6420 41064
rect 7380 41080 7432 41132
rect 8116 41080 8168 41132
rect 8208 41123 8260 41132
rect 8208 41089 8217 41123
rect 8217 41089 8251 41123
rect 8251 41089 8260 41123
rect 8208 41080 8260 41089
rect 9588 41080 9640 41132
rect 9680 41123 9732 41132
rect 9680 41089 9689 41123
rect 9689 41089 9723 41123
rect 9723 41089 9732 41123
rect 9680 41080 9732 41089
rect 9864 41080 9916 41132
rect 10324 41123 10376 41132
rect 10324 41089 10331 41123
rect 10331 41089 10365 41123
rect 10365 41089 10376 41123
rect 10324 41080 10376 41089
rect 1676 40987 1728 40996
rect 1676 40953 1685 40987
rect 1685 40953 1719 40987
rect 1719 40953 1728 40987
rect 1676 40944 1728 40953
rect 3240 40944 3292 40996
rect 3792 40876 3844 40928
rect 6000 40944 6052 40996
rect 9128 40876 9180 40928
rect 10876 40944 10928 40996
rect 19616 41216 19668 41268
rect 19156 41148 19208 41200
rect 18512 41080 18564 41132
rect 20352 41216 20404 41268
rect 20628 41216 20680 41268
rect 21272 41216 21324 41268
rect 22192 41216 22244 41268
rect 22284 41216 22336 41268
rect 23204 41216 23256 41268
rect 24308 41216 24360 41268
rect 20352 41123 20404 41132
rect 20352 41089 20361 41123
rect 20361 41089 20395 41123
rect 20395 41089 20404 41123
rect 20352 41080 20404 41089
rect 20812 41080 20864 41132
rect 21456 41080 21508 41132
rect 22008 41123 22060 41132
rect 22008 41089 22017 41123
rect 22017 41089 22051 41123
rect 22051 41089 22060 41123
rect 22008 41080 22060 41089
rect 22100 41080 22152 41132
rect 22284 41123 22336 41132
rect 22284 41089 22293 41123
rect 22293 41089 22327 41123
rect 22327 41089 22336 41123
rect 22284 41080 22336 41089
rect 22652 41123 22704 41132
rect 22652 41089 22661 41123
rect 22661 41089 22695 41123
rect 22695 41089 22704 41123
rect 22652 41080 22704 41089
rect 23112 41080 23164 41132
rect 22192 41012 22244 41064
rect 17316 40944 17368 40996
rect 19156 40987 19208 40996
rect 19156 40953 19165 40987
rect 19165 40953 19199 40987
rect 19199 40953 19208 40987
rect 19156 40944 19208 40953
rect 21364 40944 21416 40996
rect 23388 40944 23440 40996
rect 11060 40919 11112 40928
rect 11060 40885 11069 40919
rect 11069 40885 11103 40919
rect 11103 40885 11112 40919
rect 11060 40876 11112 40885
rect 19432 40919 19484 40928
rect 19432 40885 19441 40919
rect 19441 40885 19475 40919
rect 19475 40885 19484 40919
rect 19432 40876 19484 40885
rect 20536 40876 20588 40928
rect 21180 40876 21232 40928
rect 21456 40919 21508 40928
rect 21456 40885 21465 40919
rect 21465 40885 21499 40919
rect 21499 40885 21508 40919
rect 21456 40876 21508 40885
rect 23664 40919 23716 40928
rect 23664 40885 23673 40919
rect 23673 40885 23707 40919
rect 23707 40885 23716 40919
rect 23664 40876 23716 40885
rect 3917 40774 3969 40826
rect 3981 40774 4033 40826
rect 4045 40774 4097 40826
rect 4109 40774 4161 40826
rect 4173 40774 4225 40826
rect 9851 40774 9903 40826
rect 9915 40774 9967 40826
rect 9979 40774 10031 40826
rect 10043 40774 10095 40826
rect 10107 40774 10159 40826
rect 15785 40774 15837 40826
rect 15849 40774 15901 40826
rect 15913 40774 15965 40826
rect 15977 40774 16029 40826
rect 16041 40774 16093 40826
rect 21719 40774 21771 40826
rect 21783 40774 21835 40826
rect 21847 40774 21899 40826
rect 21911 40774 21963 40826
rect 21975 40774 22027 40826
rect 3608 40672 3660 40724
rect 4252 40672 4304 40724
rect 6000 40672 6052 40724
rect 3240 40536 3292 40588
rect 1676 40511 1728 40520
rect 1676 40477 1685 40511
rect 1685 40477 1719 40511
rect 1719 40477 1728 40511
rect 1676 40468 1728 40477
rect 2596 40511 2648 40520
rect 2596 40477 2603 40511
rect 2603 40477 2637 40511
rect 2637 40477 2648 40511
rect 2596 40468 2648 40477
rect 3976 40511 4028 40520
rect 3976 40477 3985 40511
rect 3985 40477 4019 40511
rect 4019 40477 4028 40511
rect 3976 40468 4028 40477
rect 7932 40672 7984 40724
rect 8576 40672 8628 40724
rect 10324 40672 10376 40724
rect 4252 40511 4304 40520
rect 4252 40477 4261 40511
rect 4261 40477 4295 40511
rect 4295 40477 4304 40511
rect 4252 40468 4304 40477
rect 4160 40400 4212 40452
rect 5264 40468 5316 40520
rect 4804 40400 4856 40452
rect 6828 40468 6880 40520
rect 6920 40468 6972 40520
rect 7472 40511 7524 40520
rect 7472 40477 7481 40511
rect 7481 40477 7515 40511
rect 7515 40477 7524 40511
rect 7472 40468 7524 40477
rect 8300 40468 8352 40520
rect 9772 40604 9824 40656
rect 10784 40672 10836 40724
rect 20168 40672 20220 40724
rect 21088 40672 21140 40724
rect 22376 40672 22428 40724
rect 22560 40715 22612 40724
rect 22560 40681 22569 40715
rect 22569 40681 22603 40715
rect 22603 40681 22612 40715
rect 22560 40672 22612 40681
rect 23296 40672 23348 40724
rect 25320 40672 25372 40724
rect 20904 40604 20956 40656
rect 20996 40647 21048 40656
rect 20996 40613 21005 40647
rect 21005 40613 21039 40647
rect 21039 40613 21048 40647
rect 20996 40604 21048 40613
rect 21272 40647 21324 40656
rect 21272 40613 21281 40647
rect 21281 40613 21315 40647
rect 21315 40613 21324 40647
rect 21272 40604 21324 40613
rect 10784 40579 10836 40588
rect 10784 40545 10793 40579
rect 10793 40545 10827 40579
rect 10827 40545 10836 40579
rect 10784 40536 10836 40545
rect 11060 40579 11112 40588
rect 11060 40545 11069 40579
rect 11069 40545 11103 40579
rect 11103 40545 11112 40579
rect 11060 40536 11112 40545
rect 16580 40536 16632 40588
rect 9772 40468 9824 40520
rect 3240 40332 3292 40384
rect 5356 40375 5408 40384
rect 5356 40341 5365 40375
rect 5365 40341 5399 40375
rect 5399 40341 5408 40375
rect 5356 40332 5408 40341
rect 6460 40332 6512 40384
rect 6736 40375 6788 40384
rect 6736 40341 6745 40375
rect 6745 40341 6779 40375
rect 6779 40341 6788 40375
rect 6736 40332 6788 40341
rect 8484 40375 8536 40384
rect 8484 40341 8493 40375
rect 8493 40341 8527 40375
rect 8527 40341 8536 40375
rect 8484 40332 8536 40341
rect 10876 40511 10928 40520
rect 10876 40477 10910 40511
rect 10910 40477 10928 40511
rect 10876 40468 10928 40477
rect 19432 40468 19484 40520
rect 20536 40536 20588 40588
rect 22008 40604 22060 40656
rect 23940 40604 23992 40656
rect 24124 40604 24176 40656
rect 20076 40511 20128 40520
rect 20076 40477 20085 40511
rect 20085 40477 20119 40511
rect 20119 40477 20128 40511
rect 20076 40468 20128 40477
rect 20812 40468 20864 40520
rect 20904 40511 20956 40520
rect 20904 40477 20913 40511
rect 20913 40477 20947 40511
rect 20947 40477 20956 40511
rect 20904 40468 20956 40477
rect 11152 40332 11204 40384
rect 11336 40332 11388 40384
rect 20720 40400 20772 40452
rect 12440 40332 12492 40384
rect 19432 40375 19484 40384
rect 19432 40341 19441 40375
rect 19441 40341 19475 40375
rect 19475 40341 19484 40375
rect 19432 40332 19484 40341
rect 19892 40375 19944 40384
rect 19892 40341 19901 40375
rect 19901 40341 19935 40375
rect 19935 40341 19944 40375
rect 19892 40332 19944 40341
rect 21364 40468 21416 40520
rect 21456 40511 21508 40520
rect 21456 40477 21465 40511
rect 21465 40477 21499 40511
rect 21499 40477 21508 40511
rect 21456 40468 21508 40477
rect 21732 40511 21784 40520
rect 21732 40477 21741 40511
rect 21741 40477 21775 40511
rect 21775 40477 21784 40511
rect 21732 40468 21784 40477
rect 22284 40511 22336 40520
rect 22284 40477 22293 40511
rect 22293 40477 22327 40511
rect 22327 40477 22336 40511
rect 22284 40468 22336 40477
rect 21916 40400 21968 40452
rect 22928 40468 22980 40520
rect 23020 40400 23072 40452
rect 23204 40400 23256 40452
rect 23848 40443 23900 40452
rect 23848 40409 23857 40443
rect 23857 40409 23891 40443
rect 23891 40409 23900 40443
rect 23848 40400 23900 40409
rect 24216 40443 24268 40452
rect 24216 40409 24225 40443
rect 24225 40409 24259 40443
rect 24259 40409 24268 40443
rect 24216 40400 24268 40409
rect 6884 40230 6936 40282
rect 6948 40230 7000 40282
rect 7012 40230 7064 40282
rect 7076 40230 7128 40282
rect 7140 40230 7192 40282
rect 12818 40230 12870 40282
rect 12882 40230 12934 40282
rect 12946 40230 12998 40282
rect 13010 40230 13062 40282
rect 13074 40230 13126 40282
rect 18752 40230 18804 40282
rect 18816 40230 18868 40282
rect 18880 40230 18932 40282
rect 18944 40230 18996 40282
rect 19008 40230 19060 40282
rect 24686 40230 24738 40282
rect 24750 40230 24802 40282
rect 24814 40230 24866 40282
rect 24878 40230 24930 40282
rect 24942 40230 24994 40282
rect 2872 40128 2924 40180
rect 2964 40128 3016 40180
rect 3148 40128 3200 40180
rect 3792 40128 3844 40180
rect 3884 40128 3936 40180
rect 4160 40128 4212 40180
rect 5264 40128 5316 40180
rect 8392 40128 8444 40180
rect 3424 40060 3476 40112
rect 2504 39992 2556 40044
rect 2964 40035 3016 40044
rect 2964 40001 2973 40035
rect 2973 40001 3007 40035
rect 3007 40001 3016 40035
rect 2964 39992 3016 40001
rect 3332 39992 3384 40044
rect 3792 39992 3844 40044
rect 4528 40060 4580 40112
rect 4988 40060 5040 40112
rect 6828 40035 6880 40044
rect 6828 40001 6835 40035
rect 6835 40001 6869 40035
rect 6869 40001 6880 40035
rect 6828 39992 6880 40001
rect 8300 40060 8352 40112
rect 10876 40128 10928 40180
rect 9036 40103 9088 40112
rect 9036 40069 9045 40103
rect 9045 40069 9079 40103
rect 9079 40069 9088 40103
rect 9036 40060 9088 40069
rect 9312 40060 9364 40112
rect 11336 40060 11388 40112
rect 15200 40060 15252 40112
rect 16856 40060 16908 40112
rect 20260 40171 20312 40180
rect 20260 40137 20269 40171
rect 20269 40137 20303 40171
rect 20303 40137 20312 40171
rect 20260 40128 20312 40137
rect 20904 40128 20956 40180
rect 22008 40128 22060 40180
rect 20628 40060 20680 40112
rect 20812 40060 20864 40112
rect 21732 40060 21784 40112
rect 22192 40128 22244 40180
rect 23112 40128 23164 40180
rect 23664 40128 23716 40180
rect 23756 40171 23808 40180
rect 23756 40137 23765 40171
rect 23765 40137 23799 40171
rect 23799 40137 23808 40171
rect 23756 40128 23808 40137
rect 8576 39992 8628 40044
rect 8760 39992 8812 40044
rect 8944 40035 8996 40044
rect 8944 40001 8953 40035
rect 8953 40001 8987 40035
rect 8987 40001 8996 40035
rect 8944 39992 8996 40001
rect 9220 39992 9272 40044
rect 9772 40035 9824 40044
rect 9772 40001 9795 40035
rect 9795 40001 9824 40035
rect 9772 39992 9824 40001
rect 20168 40035 20220 40044
rect 20168 40001 20177 40035
rect 20177 40001 20211 40035
rect 20211 40001 20220 40035
rect 20168 39992 20220 40001
rect 20444 40035 20496 40044
rect 20444 40001 20453 40035
rect 20453 40001 20487 40035
rect 20487 40001 20496 40035
rect 20444 39992 20496 40001
rect 20720 40035 20772 40044
rect 20720 40001 20729 40035
rect 20729 40001 20763 40035
rect 20763 40001 20772 40035
rect 20720 39992 20772 40001
rect 3240 39924 3292 39976
rect 4804 39924 4856 39976
rect 6460 39924 6512 39976
rect 8484 39924 8536 39976
rect 21088 40035 21140 40044
rect 21088 40001 21097 40035
rect 21097 40001 21131 40035
rect 21131 40001 21140 40035
rect 21088 39992 21140 40001
rect 21548 39992 21600 40044
rect 22100 39992 22152 40044
rect 22560 40035 22612 40044
rect 22560 40001 22569 40035
rect 22569 40001 22603 40035
rect 22603 40001 22612 40035
rect 22560 39992 22612 40001
rect 23480 40060 23532 40112
rect 23296 40035 23348 40044
rect 23296 40001 23305 40035
rect 23305 40001 23339 40035
rect 23339 40001 23348 40035
rect 23296 39992 23348 40001
rect 23664 39992 23716 40044
rect 24032 39992 24084 40044
rect 20904 39899 20956 39908
rect 20904 39865 20913 39899
rect 20913 39865 20947 39899
rect 20947 39865 20956 39899
rect 20904 39856 20956 39865
rect 21272 39856 21324 39908
rect 1860 39788 1912 39840
rect 2596 39788 2648 39840
rect 5172 39788 5224 39840
rect 5908 39831 5960 39840
rect 5908 39797 5917 39831
rect 5917 39797 5951 39831
rect 5951 39797 5960 39831
rect 5908 39788 5960 39797
rect 7472 39788 7524 39840
rect 10232 39788 10284 39840
rect 10416 39788 10468 39840
rect 12532 39788 12584 39840
rect 16948 39788 17000 39840
rect 21364 39788 21416 39840
rect 22468 39924 22520 39976
rect 23388 39856 23440 39908
rect 24400 39831 24452 39840
rect 24400 39797 24409 39831
rect 24409 39797 24443 39831
rect 24443 39797 24452 39831
rect 24400 39788 24452 39797
rect 3917 39686 3969 39738
rect 3981 39686 4033 39738
rect 4045 39686 4097 39738
rect 4109 39686 4161 39738
rect 4173 39686 4225 39738
rect 9851 39686 9903 39738
rect 9915 39686 9967 39738
rect 9979 39686 10031 39738
rect 10043 39686 10095 39738
rect 10107 39686 10159 39738
rect 15785 39686 15837 39738
rect 15849 39686 15901 39738
rect 15913 39686 15965 39738
rect 15977 39686 16029 39738
rect 16041 39686 16093 39738
rect 21719 39686 21771 39738
rect 21783 39686 21835 39738
rect 21847 39686 21899 39738
rect 21911 39686 21963 39738
rect 21975 39686 22027 39738
rect 572 39584 624 39636
rect 1860 39516 1912 39568
rect 4344 39584 4396 39636
rect 3056 39516 3108 39568
rect 4436 39516 4488 39568
rect 5356 39584 5408 39636
rect 5908 39584 5960 39636
rect 6000 39584 6052 39636
rect 8392 39584 8444 39636
rect 12164 39584 12216 39636
rect 1584 39380 1636 39432
rect 1952 39380 2004 39432
rect 4528 39448 4580 39500
rect 6736 39559 6788 39568
rect 6736 39525 6745 39559
rect 6745 39525 6779 39559
rect 6779 39525 6788 39559
rect 6736 39516 6788 39525
rect 9128 39516 9180 39568
rect 6644 39448 6696 39500
rect 7472 39448 7524 39500
rect 8208 39448 8260 39500
rect 12532 39584 12584 39636
rect 21456 39584 21508 39636
rect 21640 39627 21692 39636
rect 21640 39593 21649 39627
rect 21649 39593 21683 39627
rect 21683 39593 21692 39627
rect 21640 39584 21692 39593
rect 20812 39559 20864 39568
rect 20812 39525 20821 39559
rect 20821 39525 20855 39559
rect 20855 39525 20864 39559
rect 20812 39516 20864 39525
rect 21916 39448 21968 39500
rect 2044 39312 2096 39364
rect 940 39244 992 39296
rect 4252 39380 4304 39432
rect 5172 39423 5224 39432
rect 5172 39389 5206 39423
rect 5206 39389 5224 39423
rect 5172 39380 5224 39389
rect 3148 39312 3200 39364
rect 3056 39287 3108 39296
rect 3056 39253 3065 39287
rect 3065 39253 3099 39287
rect 3099 39253 3108 39287
rect 3056 39244 3108 39253
rect 6092 39244 6144 39296
rect 7012 39423 7064 39432
rect 7012 39389 7021 39423
rect 7021 39389 7055 39423
rect 7055 39389 7064 39423
rect 7012 39380 7064 39389
rect 7196 39380 7248 39432
rect 9496 39423 9548 39432
rect 9496 39389 9503 39423
rect 9503 39389 9537 39423
rect 9537 39389 9548 39423
rect 9496 39380 9548 39389
rect 7932 39312 7984 39364
rect 11612 39380 11664 39432
rect 7196 39244 7248 39296
rect 10140 39244 10192 39296
rect 10232 39287 10284 39296
rect 10232 39253 10241 39287
rect 10241 39253 10275 39287
rect 10275 39253 10284 39287
rect 10232 39244 10284 39253
rect 11336 39312 11388 39364
rect 20168 39380 20220 39432
rect 21272 39423 21324 39432
rect 21272 39389 21281 39423
rect 21281 39389 21315 39423
rect 21315 39389 21324 39423
rect 21272 39380 21324 39389
rect 22468 39627 22520 39636
rect 22468 39593 22477 39627
rect 22477 39593 22511 39627
rect 22511 39593 22520 39627
rect 22468 39584 22520 39593
rect 22560 39584 22612 39636
rect 23572 39584 23624 39636
rect 22560 39448 22612 39500
rect 19340 39312 19392 39364
rect 22008 39312 22060 39364
rect 12716 39244 12768 39296
rect 13268 39287 13320 39296
rect 13268 39253 13277 39287
rect 13277 39253 13311 39287
rect 13311 39253 13320 39287
rect 13268 39244 13320 39253
rect 17960 39244 18012 39296
rect 21640 39244 21692 39296
rect 22100 39244 22152 39296
rect 22468 39380 22520 39432
rect 22744 39380 22796 39432
rect 22284 39312 22336 39364
rect 23020 39287 23072 39296
rect 23020 39253 23029 39287
rect 23029 39253 23063 39287
rect 23063 39253 23072 39287
rect 23020 39244 23072 39253
rect 24124 39287 24176 39296
rect 24124 39253 24133 39287
rect 24133 39253 24167 39287
rect 24167 39253 24176 39287
rect 24124 39244 24176 39253
rect 6884 39142 6936 39194
rect 6948 39142 7000 39194
rect 7012 39142 7064 39194
rect 7076 39142 7128 39194
rect 7140 39142 7192 39194
rect 12818 39142 12870 39194
rect 12882 39142 12934 39194
rect 12946 39142 12998 39194
rect 13010 39142 13062 39194
rect 13074 39142 13126 39194
rect 18752 39142 18804 39194
rect 18816 39142 18868 39194
rect 18880 39142 18932 39194
rect 18944 39142 18996 39194
rect 19008 39142 19060 39194
rect 24686 39142 24738 39194
rect 24750 39142 24802 39194
rect 24814 39142 24866 39194
rect 24878 39142 24930 39194
rect 24942 39142 24994 39194
rect 1860 39040 1912 39092
rect 3148 39083 3200 39092
rect 3148 39049 3157 39083
rect 3157 39049 3191 39083
rect 3191 39049 3200 39083
rect 3148 39040 3200 39049
rect 3424 39040 3476 39092
rect 3792 39040 3844 39092
rect 6092 39040 6144 39092
rect 6276 39040 6328 39092
rect 6460 39040 6512 39092
rect 6644 39040 6696 39092
rect 8392 39040 8444 39092
rect 1400 38947 1452 38956
rect 1400 38913 1409 38947
rect 1409 38913 1443 38947
rect 1443 38913 1452 38947
rect 1400 38904 1452 38913
rect 1860 38904 1912 38956
rect 2044 38904 2096 38956
rect 2780 38904 2832 38956
rect 3240 38904 3292 38956
rect 3424 38947 3476 38956
rect 3424 38913 3433 38947
rect 3433 38913 3467 38947
rect 3467 38913 3476 38947
rect 3424 38904 3476 38913
rect 3792 38904 3844 38956
rect 4344 38972 4396 39024
rect 4528 38972 4580 39024
rect 4804 38904 4856 38956
rect 5356 38904 5408 38956
rect 7196 38904 7248 38956
rect 7932 38904 7984 38956
rect 8300 38972 8352 39024
rect 8668 38904 8720 38956
rect 10232 39040 10284 39092
rect 12256 39040 12308 39092
rect 20168 39083 20220 39092
rect 20168 39049 20177 39083
rect 20177 39049 20211 39083
rect 20211 39049 20220 39083
rect 20168 39040 20220 39049
rect 20720 39040 20772 39092
rect 9404 38972 9456 39024
rect 9220 38904 9272 38956
rect 9680 38947 9732 38956
rect 9680 38913 9703 38947
rect 9703 38913 9732 38947
rect 9680 38904 9732 38913
rect 2228 38879 2280 38888
rect 2228 38845 2237 38879
rect 2237 38845 2271 38879
rect 2271 38845 2280 38879
rect 2228 38836 2280 38845
rect 2044 38768 2096 38820
rect 3056 38836 3108 38888
rect 4252 38836 4304 38888
rect 4528 38700 4580 38752
rect 18328 38972 18380 39024
rect 10232 38904 10284 38956
rect 11336 38904 11388 38956
rect 12440 38947 12492 38956
rect 12440 38913 12449 38947
rect 12449 38913 12483 38947
rect 12483 38913 12492 38947
rect 12440 38904 12492 38913
rect 12716 38947 12768 38956
rect 12716 38913 12725 38947
rect 12725 38913 12759 38947
rect 12759 38913 12768 38947
rect 12716 38904 12768 38913
rect 19432 38947 19484 38956
rect 19432 38913 19441 38947
rect 19441 38913 19475 38947
rect 19475 38913 19484 38947
rect 19432 38904 19484 38913
rect 20352 38947 20404 38956
rect 20352 38913 20361 38947
rect 20361 38913 20395 38947
rect 20395 38913 20404 38947
rect 20352 38904 20404 38913
rect 11520 38879 11572 38888
rect 11520 38845 11529 38879
rect 11529 38845 11563 38879
rect 11563 38845 11572 38879
rect 11520 38836 11572 38845
rect 11704 38879 11756 38888
rect 11704 38845 11713 38879
rect 11713 38845 11747 38879
rect 11747 38845 11756 38879
rect 11704 38836 11756 38845
rect 8392 38700 8444 38752
rect 11796 38700 11848 38752
rect 12624 38700 12676 38752
rect 21364 38836 21416 38888
rect 22652 38972 22704 39024
rect 22928 39083 22980 39092
rect 22928 39049 22937 39083
rect 22937 39049 22971 39083
rect 22971 39049 22980 39083
rect 22928 39040 22980 39049
rect 23020 39040 23072 39092
rect 23112 39040 23164 39092
rect 23296 39040 23348 39092
rect 22468 38947 22520 38956
rect 22468 38913 22477 38947
rect 22477 38913 22511 38947
rect 22511 38913 22520 38947
rect 22468 38904 22520 38913
rect 23388 38947 23440 38956
rect 23388 38913 23397 38947
rect 23397 38913 23431 38947
rect 23431 38913 23440 38947
rect 23388 38904 23440 38913
rect 25228 38972 25280 39024
rect 22928 38836 22980 38888
rect 23572 38836 23624 38888
rect 24032 38904 24084 38956
rect 13636 38743 13688 38752
rect 13636 38709 13645 38743
rect 13645 38709 13679 38743
rect 13679 38709 13688 38743
rect 13636 38700 13688 38709
rect 14280 38700 14332 38752
rect 16120 38700 16172 38752
rect 22376 38700 22428 38752
rect 22652 38743 22704 38752
rect 22652 38709 22661 38743
rect 22661 38709 22695 38743
rect 22695 38709 22704 38743
rect 22652 38700 22704 38709
rect 23480 38811 23532 38820
rect 23480 38777 23489 38811
rect 23489 38777 23523 38811
rect 23523 38777 23532 38811
rect 23480 38768 23532 38777
rect 23940 38768 23992 38820
rect 24400 38743 24452 38752
rect 24400 38709 24409 38743
rect 24409 38709 24443 38743
rect 24443 38709 24452 38743
rect 24400 38700 24452 38709
rect 3917 38598 3969 38650
rect 3981 38598 4033 38650
rect 4045 38598 4097 38650
rect 4109 38598 4161 38650
rect 4173 38598 4225 38650
rect 9851 38598 9903 38650
rect 9915 38598 9967 38650
rect 9979 38598 10031 38650
rect 10043 38598 10095 38650
rect 10107 38598 10159 38650
rect 15785 38598 15837 38650
rect 15849 38598 15901 38650
rect 15913 38598 15965 38650
rect 15977 38598 16029 38650
rect 16041 38598 16093 38650
rect 21719 38598 21771 38650
rect 21783 38598 21835 38650
rect 21847 38598 21899 38650
rect 21911 38598 21963 38650
rect 21975 38598 22027 38650
rect 2504 38360 2556 38412
rect 1400 38335 1452 38344
rect 1400 38301 1409 38335
rect 1409 38301 1443 38335
rect 1443 38301 1452 38335
rect 1400 38292 1452 38301
rect 3056 38360 3108 38412
rect 2688 38267 2740 38276
rect 2688 38233 2697 38267
rect 2697 38233 2731 38267
rect 2731 38233 2740 38267
rect 2688 38224 2740 38233
rect 1216 38156 1268 38208
rect 3240 38292 3292 38344
rect 3516 38292 3568 38344
rect 4804 38539 4856 38548
rect 4804 38505 4813 38539
rect 4813 38505 4847 38539
rect 4847 38505 4856 38539
rect 4804 38496 4856 38505
rect 6736 38496 6788 38548
rect 5356 38428 5408 38480
rect 8392 38496 8444 38548
rect 9220 38496 9272 38548
rect 8944 38428 8996 38480
rect 9312 38428 9364 38480
rect 4068 38335 4120 38344
rect 4068 38301 4075 38335
rect 4075 38301 4109 38335
rect 4109 38301 4120 38335
rect 4068 38292 4120 38301
rect 7288 38292 7340 38344
rect 10140 38292 10192 38344
rect 12624 38496 12676 38548
rect 13268 38496 13320 38548
rect 19432 38496 19484 38548
rect 22468 38496 22520 38548
rect 24032 38496 24084 38548
rect 11704 38360 11756 38412
rect 12348 38360 12400 38412
rect 13636 38360 13688 38412
rect 19248 38360 19300 38412
rect 19708 38360 19760 38412
rect 6000 38156 6052 38208
rect 8208 38224 8260 38276
rect 8484 38199 8536 38208
rect 8484 38165 8493 38199
rect 8493 38165 8527 38199
rect 8527 38165 8536 38199
rect 8484 38156 8536 38165
rect 9772 38156 9824 38208
rect 11152 38292 11204 38344
rect 13084 38335 13136 38344
rect 13084 38301 13118 38335
rect 13118 38301 13136 38335
rect 13084 38292 13136 38301
rect 13268 38335 13320 38344
rect 13268 38301 13277 38335
rect 13277 38301 13311 38335
rect 13311 38301 13320 38335
rect 13268 38292 13320 38301
rect 18144 38292 18196 38344
rect 19616 38335 19668 38344
rect 19616 38301 19625 38335
rect 19625 38301 19659 38335
rect 19659 38301 19668 38335
rect 19616 38292 19668 38301
rect 22100 38335 22152 38344
rect 22100 38301 22109 38335
rect 22109 38301 22143 38335
rect 22143 38301 22152 38335
rect 22100 38292 22152 38301
rect 22376 38335 22428 38344
rect 22376 38301 22385 38335
rect 22385 38301 22428 38335
rect 22376 38292 22428 38301
rect 22468 38292 22520 38344
rect 10600 38224 10652 38276
rect 10324 38156 10376 38208
rect 11244 38199 11296 38208
rect 11244 38165 11253 38199
rect 11253 38165 11287 38199
rect 11287 38165 11296 38199
rect 11244 38156 11296 38165
rect 21364 38224 21416 38276
rect 12440 38156 12492 38208
rect 12532 38156 12584 38208
rect 13084 38156 13136 38208
rect 20352 38156 20404 38208
rect 21456 38156 21508 38208
rect 22284 38156 22336 38208
rect 22928 38156 22980 38208
rect 24124 38199 24176 38208
rect 24124 38165 24133 38199
rect 24133 38165 24167 38199
rect 24167 38165 24176 38199
rect 24124 38156 24176 38165
rect 6884 38054 6936 38106
rect 6948 38054 7000 38106
rect 7012 38054 7064 38106
rect 7076 38054 7128 38106
rect 7140 38054 7192 38106
rect 12818 38054 12870 38106
rect 12882 38054 12934 38106
rect 12946 38054 12998 38106
rect 13010 38054 13062 38106
rect 13074 38054 13126 38106
rect 18752 38054 18804 38106
rect 18816 38054 18868 38106
rect 18880 38054 18932 38106
rect 18944 38054 18996 38106
rect 19008 38054 19060 38106
rect 24686 38054 24738 38106
rect 24750 38054 24802 38106
rect 24814 38054 24866 38106
rect 24878 38054 24930 38106
rect 24942 38054 24994 38106
rect 1308 37952 1360 38004
rect 2596 37859 2648 37868
rect 2596 37825 2605 37859
rect 2605 37825 2639 37859
rect 2639 37825 2648 37859
rect 2596 37816 2648 37825
rect 3332 37859 3384 37868
rect 3332 37825 3341 37859
rect 3341 37825 3375 37859
rect 3375 37825 3384 37859
rect 3332 37816 3384 37825
rect 6736 37952 6788 38004
rect 9496 37952 9548 38004
rect 10600 37952 10652 38004
rect 13268 37952 13320 38004
rect 18144 37995 18196 38004
rect 18144 37961 18153 37995
rect 18153 37961 18187 37995
rect 18187 37961 18196 37995
rect 18144 37952 18196 37961
rect 21456 37952 21508 38004
rect 23020 37952 23072 38004
rect 23388 37995 23440 38004
rect 23388 37961 23397 37995
rect 23397 37961 23431 37995
rect 23431 37961 23440 37995
rect 23388 37952 23440 37961
rect 8300 37884 8352 37936
rect 8668 37884 8720 37936
rect 4068 37816 4120 37868
rect 1768 37748 1820 37800
rect 2320 37791 2372 37800
rect 2320 37757 2329 37791
rect 2329 37757 2363 37791
rect 2363 37757 2372 37791
rect 2320 37748 2372 37757
rect 3148 37748 3200 37800
rect 3424 37748 3476 37800
rect 1860 37680 1912 37732
rect 2136 37680 2188 37732
rect 4160 37791 4212 37800
rect 4160 37757 4169 37791
rect 4169 37757 4203 37791
rect 4203 37757 4212 37791
rect 4160 37748 4212 37757
rect 4528 37748 4580 37800
rect 7564 37859 7616 37868
rect 7564 37825 7573 37859
rect 7573 37825 7607 37859
rect 7607 37825 7616 37859
rect 7564 37816 7616 37825
rect 9220 37859 9272 37868
rect 9220 37825 9229 37859
rect 9229 37825 9263 37859
rect 9263 37825 9272 37859
rect 9220 37816 9272 37825
rect 9588 37927 9640 37936
rect 9588 37893 9597 37927
rect 9597 37893 9631 37927
rect 9631 37893 9640 37927
rect 9588 37884 9640 37893
rect 9772 37884 9824 37936
rect 15200 37884 15252 37936
rect 9680 37816 9732 37868
rect 12440 37816 12492 37868
rect 22652 37884 22704 37936
rect 2504 37612 2556 37664
rect 3148 37612 3200 37664
rect 4436 37612 4488 37664
rect 7656 37748 7708 37800
rect 8484 37748 8536 37800
rect 5816 37680 5868 37732
rect 6460 37680 6512 37732
rect 6644 37680 6696 37732
rect 7932 37680 7984 37732
rect 21088 37859 21140 37868
rect 21088 37825 21097 37859
rect 21097 37825 21131 37859
rect 21131 37825 21140 37859
rect 21088 37816 21140 37825
rect 12716 37791 12768 37800
rect 12716 37757 12725 37791
rect 12725 37757 12759 37791
rect 12759 37757 12768 37791
rect 12716 37748 12768 37757
rect 15660 37748 15712 37800
rect 20260 37748 20312 37800
rect 20536 37748 20588 37800
rect 22192 37816 22244 37868
rect 23020 37816 23072 37868
rect 23296 37816 23348 37868
rect 23848 37859 23900 37868
rect 23848 37825 23857 37859
rect 23857 37825 23891 37859
rect 23891 37825 23900 37859
rect 23848 37816 23900 37825
rect 22284 37791 22336 37800
rect 22284 37757 22293 37791
rect 22293 37757 22327 37791
rect 22327 37757 22336 37791
rect 22284 37748 22336 37757
rect 20904 37680 20956 37732
rect 22560 37680 22612 37732
rect 5632 37655 5684 37664
rect 5632 37621 5641 37655
rect 5641 37621 5675 37655
rect 5675 37621 5684 37655
rect 5632 37612 5684 37621
rect 8208 37612 8260 37664
rect 11060 37612 11112 37664
rect 12716 37612 12768 37664
rect 23388 37612 23440 37664
rect 24032 37612 24084 37664
rect 24400 37655 24452 37664
rect 24400 37621 24409 37655
rect 24409 37621 24443 37655
rect 24443 37621 24452 37655
rect 24400 37612 24452 37621
rect 3917 37510 3969 37562
rect 3981 37510 4033 37562
rect 4045 37510 4097 37562
rect 4109 37510 4161 37562
rect 4173 37510 4225 37562
rect 9851 37510 9903 37562
rect 9915 37510 9967 37562
rect 9979 37510 10031 37562
rect 10043 37510 10095 37562
rect 10107 37510 10159 37562
rect 15785 37510 15837 37562
rect 15849 37510 15901 37562
rect 15913 37510 15965 37562
rect 15977 37510 16029 37562
rect 16041 37510 16093 37562
rect 21719 37510 21771 37562
rect 21783 37510 21835 37562
rect 21847 37510 21899 37562
rect 21911 37510 21963 37562
rect 21975 37510 22027 37562
rect 1768 37408 1820 37460
rect 2136 37408 2188 37460
rect 7656 37408 7708 37460
rect 4344 37340 4396 37392
rect 4988 37340 5040 37392
rect 7472 37340 7524 37392
rect 9680 37408 9732 37460
rect 19616 37408 19668 37460
rect 22468 37451 22520 37460
rect 22468 37417 22477 37451
rect 22477 37417 22511 37451
rect 22511 37417 22520 37451
rect 22468 37408 22520 37417
rect 23296 37408 23348 37460
rect 23848 37408 23900 37460
rect 19156 37340 19208 37392
rect 23756 37340 23808 37392
rect 2136 37204 2188 37256
rect 2780 37247 2832 37256
rect 2780 37213 2789 37247
rect 2789 37213 2823 37247
rect 2823 37213 2832 37247
rect 2780 37204 2832 37213
rect 3516 37272 3568 37324
rect 4528 37272 4580 37324
rect 6460 37272 6512 37324
rect 1308 37068 1360 37120
rect 3884 37204 3936 37256
rect 8208 37315 8260 37324
rect 8208 37281 8217 37315
rect 8217 37281 8251 37315
rect 8251 37281 8260 37315
rect 8208 37272 8260 37281
rect 13820 37272 13872 37324
rect 19340 37272 19392 37324
rect 4528 37136 4580 37188
rect 5172 37136 5224 37188
rect 7656 37204 7708 37256
rect 8024 37247 8076 37256
rect 8024 37213 8033 37247
rect 8033 37213 8067 37247
rect 8067 37213 8076 37247
rect 8024 37204 8076 37213
rect 8116 37204 8168 37256
rect 6644 37136 6696 37188
rect 5264 37068 5316 37120
rect 6184 37068 6236 37120
rect 6736 37068 6788 37120
rect 9128 37204 9180 37256
rect 9312 37204 9364 37256
rect 12624 37204 12676 37256
rect 16488 37204 16540 37256
rect 19432 37247 19484 37256
rect 19432 37213 19441 37247
rect 19441 37213 19475 37247
rect 19475 37213 19484 37247
rect 19432 37204 19484 37213
rect 7288 37068 7340 37120
rect 7748 37068 7800 37120
rect 9404 37136 9456 37188
rect 20352 37247 20404 37256
rect 20352 37213 20361 37247
rect 20361 37213 20395 37247
rect 20395 37213 20404 37247
rect 20352 37204 20404 37213
rect 20904 37204 20956 37256
rect 21088 37204 21140 37256
rect 21456 37204 21508 37256
rect 23296 37272 23348 37324
rect 8392 37068 8444 37120
rect 9312 37068 9364 37120
rect 11612 37068 11664 37120
rect 13636 37068 13688 37120
rect 21272 37068 21324 37120
rect 23480 37204 23532 37256
rect 23664 37204 23716 37256
rect 23848 37247 23900 37256
rect 23848 37213 23857 37247
rect 23857 37213 23891 37247
rect 23891 37213 23900 37247
rect 23848 37204 23900 37213
rect 23940 37247 23992 37256
rect 23940 37213 23949 37247
rect 23949 37213 23983 37247
rect 23983 37213 23992 37247
rect 23940 37204 23992 37213
rect 24124 37111 24176 37120
rect 24124 37077 24133 37111
rect 24133 37077 24167 37111
rect 24167 37077 24176 37111
rect 24124 37068 24176 37077
rect 6884 36966 6936 37018
rect 6948 36966 7000 37018
rect 7012 36966 7064 37018
rect 7076 36966 7128 37018
rect 7140 36966 7192 37018
rect 12818 36966 12870 37018
rect 12882 36966 12934 37018
rect 12946 36966 12998 37018
rect 13010 36966 13062 37018
rect 13074 36966 13126 37018
rect 18752 36966 18804 37018
rect 18816 36966 18868 37018
rect 18880 36966 18932 37018
rect 18944 36966 18996 37018
rect 19008 36966 19060 37018
rect 24686 36966 24738 37018
rect 24750 36966 24802 37018
rect 24814 36966 24866 37018
rect 24878 36966 24930 37018
rect 24942 36966 24994 37018
rect 3424 36864 3476 36916
rect 5724 36864 5776 36916
rect 7196 36864 7248 36916
rect 7564 36864 7616 36916
rect 8024 36864 8076 36916
rect 9128 36864 9180 36916
rect 9404 36864 9456 36916
rect 3608 36796 3660 36848
rect 4160 36796 4212 36848
rect 4344 36796 4396 36848
rect 4988 36796 5040 36848
rect 5172 36796 5224 36848
rect 5448 36796 5500 36848
rect 1216 36728 1268 36780
rect 2872 36728 2924 36780
rect 3792 36728 3844 36780
rect 4436 36728 4488 36780
rect 20 36660 72 36712
rect 1768 36660 1820 36712
rect 2320 36660 2372 36712
rect 3332 36660 3384 36712
rect 4344 36592 4396 36644
rect 4436 36567 4488 36576
rect 4436 36533 4445 36567
rect 4445 36533 4479 36567
rect 4479 36533 4488 36567
rect 4436 36524 4488 36533
rect 5724 36660 5776 36712
rect 10140 36864 10192 36916
rect 19432 36864 19484 36916
rect 20352 36864 20404 36916
rect 23572 36864 23624 36916
rect 23940 36864 23992 36916
rect 7196 36771 7248 36780
rect 7196 36737 7205 36771
rect 7205 36737 7239 36771
rect 7239 36737 7248 36771
rect 7196 36728 7248 36737
rect 7656 36771 7708 36780
rect 7656 36737 7665 36771
rect 7665 36737 7699 36771
rect 7699 36737 7708 36771
rect 7656 36728 7708 36737
rect 7564 36660 7616 36712
rect 10140 36771 10192 36780
rect 10140 36737 10147 36771
rect 10147 36737 10181 36771
rect 10181 36737 10192 36771
rect 10140 36728 10192 36737
rect 10784 36660 10836 36712
rect 22284 36728 22336 36780
rect 24032 36796 24084 36848
rect 16764 36592 16816 36644
rect 17776 36592 17828 36644
rect 18144 36592 18196 36644
rect 10876 36567 10928 36576
rect 10876 36533 10885 36567
rect 10885 36533 10919 36567
rect 10919 36533 10928 36567
rect 10876 36524 10928 36533
rect 12072 36524 12124 36576
rect 12532 36524 12584 36576
rect 13452 36524 13504 36576
rect 13728 36524 13780 36576
rect 22928 36524 22980 36576
rect 23020 36567 23072 36576
rect 23020 36533 23029 36567
rect 23029 36533 23063 36567
rect 23063 36533 23072 36567
rect 23020 36524 23072 36533
rect 24400 36567 24452 36576
rect 24400 36533 24409 36567
rect 24409 36533 24443 36567
rect 24443 36533 24452 36567
rect 24400 36524 24452 36533
rect 3917 36422 3969 36474
rect 3981 36422 4033 36474
rect 4045 36422 4097 36474
rect 4109 36422 4161 36474
rect 4173 36422 4225 36474
rect 9851 36422 9903 36474
rect 9915 36422 9967 36474
rect 9979 36422 10031 36474
rect 10043 36422 10095 36474
rect 10107 36422 10159 36474
rect 15785 36422 15837 36474
rect 15849 36422 15901 36474
rect 15913 36422 15965 36474
rect 15977 36422 16029 36474
rect 16041 36422 16093 36474
rect 21719 36422 21771 36474
rect 21783 36422 21835 36474
rect 21847 36422 21899 36474
rect 21911 36422 21963 36474
rect 21975 36422 22027 36474
rect 3332 36363 3384 36372
rect 3332 36329 3341 36363
rect 3341 36329 3375 36363
rect 3375 36329 3384 36363
rect 3332 36320 3384 36329
rect 4344 36320 4396 36372
rect 7196 36320 7248 36372
rect 7656 36320 7708 36372
rect 8116 36320 8168 36372
rect 4436 36252 4488 36304
rect 4620 36252 4672 36304
rect 5632 36295 5684 36304
rect 5632 36261 5641 36295
rect 5641 36261 5675 36295
rect 5675 36261 5684 36295
rect 5632 36252 5684 36261
rect 5724 36184 5776 36236
rect 6184 36227 6236 36236
rect 6184 36193 6193 36227
rect 6193 36193 6227 36227
rect 6227 36193 6236 36227
rect 6184 36184 6236 36193
rect 1400 36159 1452 36168
rect 1400 36125 1409 36159
rect 1409 36125 1443 36159
rect 1443 36125 1452 36159
rect 1400 36116 1452 36125
rect 1124 35980 1176 36032
rect 2688 36116 2740 36168
rect 3056 36116 3108 36168
rect 3792 36159 3844 36168
rect 3792 36125 3801 36159
rect 3801 36125 3835 36159
rect 3835 36125 3844 36159
rect 3792 36116 3844 36125
rect 4344 36159 4396 36168
rect 4344 36125 4353 36159
rect 4353 36125 4387 36159
rect 4387 36125 4396 36159
rect 4344 36116 4396 36125
rect 4436 36116 4488 36168
rect 5080 36116 5132 36168
rect 5908 36159 5960 36168
rect 5908 36125 5917 36159
rect 5917 36125 5951 36159
rect 5951 36125 5960 36159
rect 5908 36116 5960 36125
rect 7288 36116 7340 36168
rect 4068 36091 4120 36100
rect 4068 36057 4077 36091
rect 4077 36057 4111 36091
rect 4111 36057 4120 36091
rect 4068 36048 4120 36057
rect 5172 36048 5224 36100
rect 10048 36116 10100 36168
rect 10784 36320 10836 36372
rect 14556 36320 14608 36372
rect 16580 36320 16632 36372
rect 22284 36320 22336 36372
rect 15108 36252 15160 36304
rect 18328 36252 18380 36304
rect 19984 36252 20036 36304
rect 22836 36363 22888 36372
rect 22836 36329 22845 36363
rect 22845 36329 22879 36363
rect 22879 36329 22888 36363
rect 22836 36320 22888 36329
rect 10324 36048 10376 36100
rect 11888 36048 11940 36100
rect 12256 36159 12308 36168
rect 12256 36125 12265 36159
rect 12265 36125 12299 36159
rect 12299 36125 12308 36159
rect 12256 36116 12308 36125
rect 12440 36116 12492 36168
rect 13728 36116 13780 36168
rect 20352 36184 20404 36236
rect 21272 36184 21324 36236
rect 23480 36252 23532 36304
rect 24308 36252 24360 36304
rect 19248 36116 19300 36168
rect 19432 36159 19484 36168
rect 19432 36125 19441 36159
rect 19441 36125 19475 36159
rect 19475 36125 19484 36159
rect 19432 36116 19484 36125
rect 2688 35980 2740 36032
rect 4160 35980 4212 36032
rect 8392 35980 8444 36032
rect 9956 35980 10008 36032
rect 11336 35980 11388 36032
rect 12164 35980 12216 36032
rect 17960 35980 18012 36032
rect 20628 36116 20680 36168
rect 22744 36159 22796 36168
rect 22744 36125 22753 36159
rect 22753 36125 22787 36159
rect 22787 36125 22796 36159
rect 22744 36116 22796 36125
rect 23296 36184 23348 36236
rect 19340 35980 19392 36032
rect 19892 35980 19944 36032
rect 21548 35980 21600 36032
rect 25412 36048 25464 36100
rect 24124 36023 24176 36032
rect 24124 35989 24133 36023
rect 24133 35989 24167 36023
rect 24167 35989 24176 36023
rect 24124 35980 24176 35989
rect 6884 35878 6936 35930
rect 6948 35878 7000 35930
rect 7012 35878 7064 35930
rect 7076 35878 7128 35930
rect 7140 35878 7192 35930
rect 12818 35878 12870 35930
rect 12882 35878 12934 35930
rect 12946 35878 12998 35930
rect 13010 35878 13062 35930
rect 13074 35878 13126 35930
rect 18752 35878 18804 35930
rect 18816 35878 18868 35930
rect 18880 35878 18932 35930
rect 18944 35878 18996 35930
rect 19008 35878 19060 35930
rect 24686 35878 24738 35930
rect 24750 35878 24802 35930
rect 24814 35878 24866 35930
rect 24878 35878 24930 35930
rect 24942 35878 24994 35930
rect 3516 35776 3568 35828
rect 4712 35776 4764 35828
rect 7288 35776 7340 35828
rect 9404 35776 9456 35828
rect 1308 35708 1360 35760
rect 1492 35640 1544 35692
rect 2688 35683 2740 35692
rect 2688 35649 2695 35683
rect 2695 35649 2729 35683
rect 2729 35649 2740 35683
rect 2688 35640 2740 35649
rect 3056 35640 3108 35692
rect 6460 35708 6512 35760
rect 7380 35708 7432 35760
rect 8208 35708 8260 35760
rect 9588 35708 9640 35760
rect 6184 35640 6236 35692
rect 8392 35683 8444 35692
rect 8392 35649 8401 35683
rect 8401 35649 8435 35683
rect 8435 35649 8444 35683
rect 8392 35640 8444 35649
rect 8484 35640 8536 35692
rect 8668 35640 8720 35692
rect 8760 35683 8812 35692
rect 8760 35649 8769 35683
rect 8769 35649 8803 35683
rect 8803 35649 8812 35683
rect 8760 35640 8812 35649
rect 9220 35640 9272 35692
rect 10232 35776 10284 35828
rect 11796 35819 11848 35828
rect 11796 35785 11805 35819
rect 11805 35785 11839 35819
rect 11839 35785 11848 35819
rect 11796 35776 11848 35785
rect 13452 35776 13504 35828
rect 12900 35751 12952 35760
rect 12900 35717 12909 35751
rect 12909 35717 12943 35751
rect 12943 35717 12952 35751
rect 12900 35708 12952 35717
rect 18144 35776 18196 35828
rect 19432 35776 19484 35828
rect 19708 35776 19760 35828
rect 19892 35751 19944 35760
rect 10416 35683 10468 35692
rect 10416 35649 10425 35683
rect 10425 35649 10459 35683
rect 10459 35649 10468 35683
rect 10416 35640 10468 35649
rect 1676 35615 1728 35624
rect 1676 35581 1685 35615
rect 1685 35581 1719 35615
rect 1719 35581 1728 35615
rect 1676 35572 1728 35581
rect 3332 35572 3384 35624
rect 4160 35572 4212 35624
rect 4528 35615 4580 35624
rect 4528 35581 4537 35615
rect 4537 35581 4571 35615
rect 4571 35581 4580 35615
rect 4528 35572 4580 35581
rect 5264 35615 5316 35624
rect 5264 35581 5273 35615
rect 5273 35581 5307 35615
rect 5307 35581 5316 35615
rect 5264 35572 5316 35581
rect 5356 35615 5408 35624
rect 5356 35581 5390 35615
rect 5390 35581 5408 35615
rect 5356 35572 5408 35581
rect 8208 35572 8260 35624
rect 4620 35504 4672 35556
rect 3424 35479 3476 35488
rect 3424 35445 3433 35479
rect 3433 35445 3467 35479
rect 3467 35445 3476 35479
rect 3424 35436 3476 35445
rect 10232 35572 10284 35624
rect 11980 35640 12032 35692
rect 12072 35683 12124 35692
rect 12072 35649 12081 35683
rect 12081 35649 12115 35683
rect 12115 35649 12124 35683
rect 12072 35640 12124 35649
rect 12164 35683 12216 35692
rect 12164 35649 12173 35683
rect 12173 35649 12207 35683
rect 12207 35649 12216 35683
rect 12164 35640 12216 35649
rect 12256 35640 12308 35692
rect 11244 35572 11296 35624
rect 13084 35572 13136 35624
rect 17960 35683 18012 35692
rect 17960 35649 17994 35683
rect 17994 35649 18012 35683
rect 17960 35640 18012 35649
rect 19156 35683 19208 35692
rect 19156 35649 19165 35683
rect 19165 35649 19199 35683
rect 19199 35649 19208 35683
rect 19156 35640 19208 35649
rect 19248 35683 19300 35692
rect 19248 35649 19257 35683
rect 19257 35649 19291 35683
rect 19291 35649 19300 35683
rect 19248 35640 19300 35649
rect 9956 35504 10008 35556
rect 17684 35615 17736 35624
rect 17684 35581 17693 35615
rect 17693 35581 17727 35615
rect 17727 35581 17736 35615
rect 17684 35572 17736 35581
rect 19432 35615 19484 35624
rect 19432 35581 19441 35615
rect 19441 35581 19475 35615
rect 19475 35581 19484 35615
rect 19432 35572 19484 35581
rect 19892 35717 19904 35751
rect 19904 35717 19944 35751
rect 19892 35708 19944 35717
rect 21732 35708 21784 35760
rect 21272 35640 21324 35692
rect 21548 35640 21600 35692
rect 22744 35776 22796 35828
rect 22192 35708 22244 35760
rect 23296 35819 23348 35828
rect 23296 35785 23305 35819
rect 23305 35785 23339 35819
rect 23339 35785 23348 35819
rect 23296 35776 23348 35785
rect 23848 35776 23900 35828
rect 22100 35683 22152 35692
rect 22100 35649 22109 35683
rect 22109 35649 22143 35683
rect 22143 35649 22152 35683
rect 22100 35640 22152 35649
rect 15292 35504 15344 35556
rect 5632 35436 5684 35488
rect 9312 35479 9364 35488
rect 9312 35445 9321 35479
rect 9321 35445 9355 35479
rect 9355 35445 9364 35479
rect 9312 35436 9364 35445
rect 9496 35436 9548 35488
rect 13912 35436 13964 35488
rect 14188 35436 14240 35488
rect 14464 35436 14516 35488
rect 20720 35436 20772 35488
rect 22560 35683 22612 35692
rect 22560 35649 22569 35683
rect 22569 35649 22603 35683
rect 22603 35649 22612 35683
rect 22560 35640 22612 35649
rect 22928 35504 22980 35556
rect 24124 35683 24176 35692
rect 24124 35649 24133 35683
rect 24133 35649 24167 35683
rect 24167 35649 24176 35683
rect 24124 35640 24176 35649
rect 21732 35436 21784 35488
rect 25688 35504 25740 35556
rect 24400 35479 24452 35488
rect 24400 35445 24409 35479
rect 24409 35445 24443 35479
rect 24443 35445 24452 35479
rect 24400 35436 24452 35445
rect 3917 35334 3969 35386
rect 3981 35334 4033 35386
rect 4045 35334 4097 35386
rect 4109 35334 4161 35386
rect 4173 35334 4225 35386
rect 9851 35334 9903 35386
rect 9915 35334 9967 35386
rect 9979 35334 10031 35386
rect 10043 35334 10095 35386
rect 10107 35334 10159 35386
rect 15785 35334 15837 35386
rect 15849 35334 15901 35386
rect 15913 35334 15965 35386
rect 15977 35334 16029 35386
rect 16041 35334 16093 35386
rect 21719 35334 21771 35386
rect 21783 35334 21835 35386
rect 21847 35334 21899 35386
rect 21911 35334 21963 35386
rect 21975 35334 22027 35386
rect 1676 35096 1728 35148
rect 2228 35139 2280 35148
rect 2228 35105 2237 35139
rect 2237 35105 2271 35139
rect 2271 35105 2280 35139
rect 2228 35096 2280 35105
rect 3148 35232 3200 35284
rect 3700 35232 3752 35284
rect 5816 35232 5868 35284
rect 6184 35232 6236 35284
rect 2780 35071 2832 35080
rect 2780 35037 2789 35071
rect 2789 35037 2823 35071
rect 2823 35037 2832 35071
rect 2780 35028 2832 35037
rect 3424 35096 3476 35148
rect 7748 35232 7800 35284
rect 8208 35232 8260 35284
rect 8668 35232 8720 35284
rect 10324 35232 10376 35284
rect 13084 35275 13136 35284
rect 13084 35241 13093 35275
rect 13093 35241 13127 35275
rect 13127 35241 13136 35275
rect 13084 35232 13136 35241
rect 13728 35232 13780 35284
rect 9404 35164 9456 35216
rect 10876 35164 10928 35216
rect 19156 35164 19208 35216
rect 19432 35232 19484 35284
rect 21272 35275 21324 35284
rect 21272 35241 21281 35275
rect 21281 35241 21315 35275
rect 21315 35241 21324 35275
rect 21272 35232 21324 35241
rect 21916 35232 21968 35284
rect 21180 35164 21232 35216
rect 4068 35028 4120 35080
rect 4252 35071 4304 35080
rect 4252 35037 4261 35071
rect 4261 35037 4295 35071
rect 4295 35037 4304 35071
rect 4252 35028 4304 35037
rect 5172 35028 5224 35080
rect 7564 35071 7616 35080
rect 3424 34892 3476 34944
rect 4160 34960 4212 35012
rect 4804 34960 4856 35012
rect 7564 35037 7571 35071
rect 7571 35037 7605 35071
rect 7605 35037 7616 35071
rect 7564 35028 7616 35037
rect 7932 35028 7984 35080
rect 8024 35028 8076 35080
rect 8300 35028 8352 35080
rect 8484 35028 8536 35080
rect 12072 35139 12124 35148
rect 12072 35105 12081 35139
rect 12081 35105 12115 35139
rect 12115 35105 12124 35139
rect 12072 35096 12124 35105
rect 19340 35096 19392 35148
rect 22560 35232 22612 35284
rect 23204 35275 23256 35284
rect 23204 35241 23213 35275
rect 23213 35241 23247 35275
rect 23247 35241 23256 35275
rect 23204 35232 23256 35241
rect 24124 35232 24176 35284
rect 10048 35028 10100 35080
rect 9864 34960 9916 35012
rect 11060 35071 11112 35080
rect 11060 35037 11069 35071
rect 11069 35037 11103 35071
rect 11103 35037 11112 35071
rect 11060 35028 11112 35037
rect 11152 35071 11204 35080
rect 11152 35037 11186 35071
rect 11186 35037 11204 35071
rect 11152 35028 11204 35037
rect 11336 35071 11388 35080
rect 11336 35037 11345 35071
rect 11345 35037 11379 35071
rect 11379 35037 11388 35071
rect 11336 35028 11388 35037
rect 4528 34892 4580 34944
rect 4988 34892 5040 34944
rect 5080 34935 5132 34944
rect 5080 34901 5089 34935
rect 5089 34901 5123 34935
rect 5123 34901 5132 34935
rect 5080 34892 5132 34901
rect 5172 34892 5224 34944
rect 5724 34892 5776 34944
rect 7564 34892 7616 34944
rect 9496 34892 9548 34944
rect 10048 34892 10100 34944
rect 12256 35028 12308 35080
rect 18052 35071 18104 35080
rect 12624 34960 12676 35012
rect 12900 34960 12952 35012
rect 13452 34960 13504 35012
rect 14188 34960 14240 35012
rect 15476 34960 15528 35012
rect 18052 35037 18059 35071
rect 18059 35037 18093 35071
rect 18093 35037 18104 35071
rect 18052 35028 18104 35037
rect 19156 35028 19208 35080
rect 20444 35028 20496 35080
rect 20628 35028 20680 35080
rect 22744 35096 22796 35148
rect 17868 34892 17920 34944
rect 18236 34960 18288 35012
rect 21456 35028 21508 35080
rect 21180 34960 21232 35012
rect 19708 34892 19760 34944
rect 20444 34892 20496 34944
rect 22100 34892 22152 34944
rect 23204 34892 23256 34944
rect 23572 34960 23624 35012
rect 24216 35003 24268 35012
rect 24216 34969 24225 35003
rect 24225 34969 24259 35003
rect 24259 34969 24268 35003
rect 24216 34960 24268 34969
rect 6884 34790 6936 34842
rect 6948 34790 7000 34842
rect 7012 34790 7064 34842
rect 7076 34790 7128 34842
rect 7140 34790 7192 34842
rect 12818 34790 12870 34842
rect 12882 34790 12934 34842
rect 12946 34790 12998 34842
rect 13010 34790 13062 34842
rect 13074 34790 13126 34842
rect 18752 34790 18804 34842
rect 18816 34790 18868 34842
rect 18880 34790 18932 34842
rect 18944 34790 18996 34842
rect 19008 34790 19060 34842
rect 24686 34790 24738 34842
rect 24750 34790 24802 34842
rect 24814 34790 24866 34842
rect 24878 34790 24930 34842
rect 24942 34790 24994 34842
rect 1768 34688 1820 34740
rect 2780 34688 2832 34740
rect 3148 34688 3200 34740
rect 3424 34688 3476 34740
rect 4160 34688 4212 34740
rect 4620 34688 4672 34740
rect 4068 34620 4120 34672
rect 4804 34663 4856 34672
rect 4804 34629 4813 34663
rect 4813 34629 4847 34663
rect 4847 34629 4856 34663
rect 4804 34620 4856 34629
rect 5724 34688 5776 34740
rect 4344 34552 4396 34604
rect 4528 34552 4580 34604
rect 5356 34552 5408 34604
rect 1492 34527 1544 34536
rect 1492 34493 1501 34527
rect 1501 34493 1535 34527
rect 1535 34493 1544 34527
rect 1492 34484 1544 34493
rect 2872 34484 2924 34536
rect 3056 34484 3108 34536
rect 8300 34688 8352 34740
rect 8392 34688 8444 34740
rect 9864 34688 9916 34740
rect 6644 34625 6696 34672
rect 6184 34552 6236 34604
rect 6644 34620 6669 34625
rect 6669 34620 6696 34625
rect 8024 34620 8076 34672
rect 11152 34620 11204 34672
rect 15476 34688 15528 34740
rect 16672 34688 16724 34740
rect 1768 34348 1820 34400
rect 2412 34348 2464 34400
rect 6092 34391 6144 34400
rect 6092 34357 6101 34391
rect 6101 34357 6135 34391
rect 6135 34357 6144 34391
rect 6092 34348 6144 34357
rect 6184 34348 6236 34400
rect 7748 34552 7800 34604
rect 10600 34552 10652 34604
rect 11060 34552 11112 34604
rect 16120 34620 16172 34672
rect 17408 34688 17460 34740
rect 17224 34620 17276 34672
rect 19340 34620 19392 34672
rect 21456 34731 21508 34740
rect 21456 34697 21465 34731
rect 21465 34697 21499 34731
rect 21499 34697 21508 34731
rect 21456 34688 21508 34697
rect 16672 34595 16724 34604
rect 16672 34561 16681 34595
rect 16681 34561 16715 34595
rect 16715 34561 16724 34595
rect 16672 34552 16724 34561
rect 17868 34552 17920 34604
rect 20168 34552 20220 34604
rect 23572 34688 23624 34740
rect 8944 34484 8996 34536
rect 10416 34484 10468 34536
rect 14096 34527 14148 34536
rect 14096 34493 14105 34527
rect 14105 34493 14139 34527
rect 14139 34493 14148 34527
rect 14096 34484 14148 34493
rect 16396 34484 16448 34536
rect 9128 34416 9180 34468
rect 9588 34416 9640 34468
rect 6828 34348 6880 34400
rect 15108 34391 15160 34400
rect 15108 34357 15117 34391
rect 15117 34357 15151 34391
rect 15151 34357 15160 34391
rect 15108 34348 15160 34357
rect 16304 34391 16356 34400
rect 16304 34357 16313 34391
rect 16313 34357 16347 34391
rect 16347 34357 16356 34391
rect 16304 34348 16356 34357
rect 19432 34484 19484 34536
rect 23020 34552 23072 34604
rect 23204 34595 23256 34604
rect 23204 34561 23213 34595
rect 23213 34561 23247 34595
rect 23247 34561 23256 34595
rect 23204 34552 23256 34561
rect 24400 34527 24452 34536
rect 24400 34493 24409 34527
rect 24409 34493 24443 34527
rect 24443 34493 24452 34527
rect 24400 34484 24452 34493
rect 23020 34459 23072 34468
rect 23020 34425 23029 34459
rect 23029 34425 23063 34459
rect 23063 34425 23072 34459
rect 23020 34416 23072 34425
rect 23388 34416 23440 34468
rect 25596 34416 25648 34468
rect 17500 34348 17552 34400
rect 20260 34348 20312 34400
rect 25504 34348 25556 34400
rect 3917 34246 3969 34298
rect 3981 34246 4033 34298
rect 4045 34246 4097 34298
rect 4109 34246 4161 34298
rect 4173 34246 4225 34298
rect 9851 34246 9903 34298
rect 9915 34246 9967 34298
rect 9979 34246 10031 34298
rect 10043 34246 10095 34298
rect 10107 34246 10159 34298
rect 15785 34246 15837 34298
rect 15849 34246 15901 34298
rect 15913 34246 15965 34298
rect 15977 34246 16029 34298
rect 16041 34246 16093 34298
rect 21719 34246 21771 34298
rect 21783 34246 21835 34298
rect 21847 34246 21899 34298
rect 21911 34246 21963 34298
rect 21975 34246 22027 34298
rect 2228 34144 2280 34196
rect 2688 34144 2740 34196
rect 4620 34144 4672 34196
rect 3608 34076 3660 34128
rect 9220 34144 9272 34196
rect 9588 34144 9640 34196
rect 10508 34144 10560 34196
rect 14096 34144 14148 34196
rect 2780 33983 2832 33992
rect 2780 33949 2789 33983
rect 2789 33949 2823 33983
rect 2823 33949 2832 33983
rect 2780 33940 2832 33949
rect 3792 33983 3844 33992
rect 3792 33949 3801 33983
rect 3801 33949 3835 33983
rect 3835 33949 3844 33983
rect 3792 33940 3844 33949
rect 3884 33940 3936 33992
rect 2320 33872 2372 33924
rect 2504 33872 2556 33924
rect 4252 33872 4304 33924
rect 9128 34076 9180 34128
rect 6828 34008 6880 34060
rect 11888 34008 11940 34060
rect 16304 34144 16356 34196
rect 17500 34187 17552 34196
rect 17500 34153 17509 34187
rect 17509 34153 17543 34187
rect 17543 34153 17552 34187
rect 17500 34144 17552 34153
rect 22100 34144 22152 34196
rect 24492 34144 24544 34196
rect 15476 34051 15528 34060
rect 15476 34017 15485 34051
rect 15485 34017 15519 34051
rect 15519 34017 15528 34051
rect 15476 34008 15528 34017
rect 5264 33940 5316 33992
rect 5724 33940 5776 33992
rect 5908 33940 5960 33992
rect 9128 33940 9180 33992
rect 6092 33872 6144 33924
rect 1492 33804 1544 33856
rect 1952 33804 2004 33856
rect 2228 33804 2280 33856
rect 2688 33804 2740 33856
rect 6552 33847 6604 33856
rect 6552 33813 6561 33847
rect 6561 33813 6595 33847
rect 6595 33813 6604 33847
rect 6552 33804 6604 33813
rect 7380 33804 7432 33856
rect 8116 33804 8168 33856
rect 9404 33804 9456 33856
rect 9680 33804 9732 33856
rect 10140 33983 10192 33992
rect 10140 33949 10149 33983
rect 10149 33949 10183 33983
rect 10183 33949 10192 33983
rect 10140 33940 10192 33949
rect 10048 33872 10100 33924
rect 13728 33940 13780 33992
rect 11336 33872 11388 33924
rect 15384 33940 15436 33992
rect 14924 33872 14976 33924
rect 17132 33983 17184 33992
rect 17132 33949 17141 33983
rect 17141 33949 17175 33983
rect 17175 33949 17184 33983
rect 17132 33940 17184 33949
rect 17408 33983 17460 33992
rect 17408 33949 17441 33983
rect 17441 33949 17460 33983
rect 17408 33940 17460 33949
rect 17592 33983 17644 33992
rect 17592 33949 17601 33983
rect 17601 33949 17635 33983
rect 17635 33949 17644 33983
rect 17592 33940 17644 33949
rect 19340 33940 19392 33992
rect 20260 33940 20312 33992
rect 21180 33872 21232 33924
rect 21364 33940 21416 33992
rect 23296 33940 23348 33992
rect 23664 33983 23716 33992
rect 23664 33949 23673 33983
rect 23673 33949 23707 33983
rect 23707 33949 23716 33983
rect 23664 33940 23716 33949
rect 10508 33804 10560 33856
rect 13176 33847 13228 33856
rect 13176 33813 13185 33847
rect 13185 33813 13219 33847
rect 13219 33813 13228 33847
rect 13176 33804 13228 33813
rect 14648 33804 14700 33856
rect 16488 33847 16540 33856
rect 16488 33813 16497 33847
rect 16497 33813 16531 33847
rect 16531 33813 16540 33847
rect 16488 33804 16540 33813
rect 22192 33847 22244 33856
rect 22192 33813 22201 33847
rect 22201 33813 22235 33847
rect 22235 33813 22244 33847
rect 22192 33804 22244 33813
rect 23388 33847 23440 33856
rect 23388 33813 23397 33847
rect 23397 33813 23431 33847
rect 23431 33813 23440 33847
rect 23388 33804 23440 33813
rect 24124 33847 24176 33856
rect 24124 33813 24133 33847
rect 24133 33813 24167 33847
rect 24167 33813 24176 33847
rect 24124 33804 24176 33813
rect 20 33668 72 33720
rect 6884 33702 6936 33754
rect 6948 33702 7000 33754
rect 7012 33702 7064 33754
rect 7076 33702 7128 33754
rect 7140 33702 7192 33754
rect 12818 33702 12870 33754
rect 12882 33702 12934 33754
rect 12946 33702 12998 33754
rect 13010 33702 13062 33754
rect 13074 33702 13126 33754
rect 18752 33702 18804 33754
rect 18816 33702 18868 33754
rect 18880 33702 18932 33754
rect 18944 33702 18996 33754
rect 19008 33702 19060 33754
rect 24686 33702 24738 33754
rect 24750 33702 24802 33754
rect 24814 33702 24866 33754
rect 24878 33702 24930 33754
rect 24942 33702 24994 33754
rect 5724 33600 5776 33652
rect 7656 33600 7708 33652
rect 112 33532 164 33584
rect 2688 33532 2740 33584
rect 848 33464 900 33516
rect 1124 33464 1176 33516
rect 1400 33507 1452 33516
rect 1400 33473 1409 33507
rect 1409 33473 1443 33507
rect 1443 33473 1452 33507
rect 1400 33464 1452 33473
rect 1676 33507 1728 33516
rect 1676 33473 1685 33507
rect 1685 33473 1719 33507
rect 1719 33473 1728 33507
rect 1676 33464 1728 33473
rect 1952 33507 2004 33516
rect 1952 33473 1961 33507
rect 1961 33473 1995 33507
rect 1995 33473 2004 33507
rect 1952 33464 2004 33473
rect 2504 33507 2556 33516
rect 2504 33473 2513 33507
rect 2513 33473 2547 33507
rect 2547 33473 2556 33507
rect 2504 33464 2556 33473
rect 2596 33396 2648 33448
rect 4344 33464 4396 33516
rect 5356 33464 5408 33516
rect 6736 33532 6788 33584
rect 6828 33464 6880 33516
rect 8668 33464 8720 33516
rect 8760 33507 8812 33516
rect 8760 33473 8769 33507
rect 8769 33473 8803 33507
rect 8803 33473 8812 33507
rect 8760 33464 8812 33473
rect 3056 33328 3108 33380
rect 2872 33260 2924 33312
rect 4988 33396 5040 33448
rect 6184 33396 6236 33448
rect 6276 33396 6328 33448
rect 4804 33328 4856 33380
rect 5632 33328 5684 33380
rect 7932 33396 7984 33448
rect 8116 33396 8168 33448
rect 3884 33260 3936 33312
rect 4252 33260 4304 33312
rect 5816 33260 5868 33312
rect 6092 33260 6144 33312
rect 8208 33260 8260 33312
rect 9588 33600 9640 33652
rect 9404 33464 9456 33516
rect 10140 33600 10192 33652
rect 10508 33643 10560 33652
rect 10508 33609 10517 33643
rect 10517 33609 10551 33643
rect 10551 33609 10560 33643
rect 10508 33600 10560 33609
rect 10324 33532 10376 33584
rect 10968 33532 11020 33584
rect 12348 33600 12400 33652
rect 12716 33600 12768 33652
rect 13728 33600 13780 33652
rect 14832 33600 14884 33652
rect 17592 33600 17644 33652
rect 16856 33532 16908 33584
rect 17408 33532 17460 33584
rect 9496 33439 9548 33448
rect 9496 33405 9505 33439
rect 9505 33405 9539 33439
rect 9539 33405 9548 33439
rect 9496 33396 9548 33405
rect 9864 33260 9916 33312
rect 9956 33260 10008 33312
rect 15108 33507 15160 33516
rect 15108 33473 15117 33507
rect 15117 33473 15151 33507
rect 15151 33473 15160 33507
rect 15108 33464 15160 33473
rect 17316 33507 17368 33516
rect 17316 33473 17325 33507
rect 17325 33473 17359 33507
rect 17359 33473 17368 33507
rect 17316 33464 17368 33473
rect 10324 33396 10376 33448
rect 11244 33328 11296 33380
rect 12624 33439 12676 33448
rect 12624 33405 12658 33439
rect 12658 33405 12676 33439
rect 12624 33396 12676 33405
rect 13176 33396 13228 33448
rect 11796 33328 11848 33380
rect 12256 33371 12308 33380
rect 12256 33337 12265 33371
rect 12265 33337 12299 33371
rect 12299 33337 12308 33371
rect 12256 33328 12308 33337
rect 14648 33396 14700 33448
rect 14832 33439 14884 33448
rect 14832 33405 14841 33439
rect 14841 33405 14875 33439
rect 14875 33405 14884 33439
rect 14832 33396 14884 33405
rect 14924 33439 14976 33448
rect 14924 33405 14958 33439
rect 14958 33405 14976 33439
rect 14924 33396 14976 33405
rect 14188 33328 14240 33380
rect 14372 33328 14424 33380
rect 10416 33260 10468 33312
rect 12624 33260 12676 33312
rect 19524 33532 19576 33584
rect 17960 33464 18012 33516
rect 19616 33507 19668 33516
rect 19616 33473 19625 33507
rect 19625 33473 19659 33507
rect 19659 33473 19668 33507
rect 19616 33464 19668 33473
rect 22192 33600 22244 33652
rect 22744 33643 22796 33652
rect 22744 33609 22753 33643
rect 22753 33609 22787 33643
rect 22787 33609 22796 33643
rect 22744 33600 22796 33609
rect 23296 33600 23348 33652
rect 23388 33600 23440 33652
rect 23664 33600 23716 33652
rect 19156 33396 19208 33448
rect 18604 33328 18656 33380
rect 22652 33464 22704 33516
rect 23296 33464 23348 33516
rect 23940 33507 23992 33516
rect 23940 33473 23949 33507
rect 23949 33473 23983 33507
rect 23983 33473 23992 33507
rect 23940 33464 23992 33473
rect 19340 33260 19392 33312
rect 20812 33260 20864 33312
rect 22100 33303 22152 33312
rect 22100 33269 22109 33303
rect 22109 33269 22143 33303
rect 22143 33269 22152 33303
rect 22100 33260 22152 33269
rect 23848 33260 23900 33312
rect 24400 33303 24452 33312
rect 24400 33269 24409 33303
rect 24409 33269 24443 33303
rect 24443 33269 24452 33303
rect 24400 33260 24452 33269
rect 3917 33158 3969 33210
rect 3981 33158 4033 33210
rect 4045 33158 4097 33210
rect 4109 33158 4161 33210
rect 4173 33158 4225 33210
rect 9851 33158 9903 33210
rect 9915 33158 9967 33210
rect 9979 33158 10031 33210
rect 10043 33158 10095 33210
rect 10107 33158 10159 33210
rect 15785 33158 15837 33210
rect 15849 33158 15901 33210
rect 15913 33158 15965 33210
rect 15977 33158 16029 33210
rect 16041 33158 16093 33210
rect 21719 33158 21771 33210
rect 21783 33158 21835 33210
rect 21847 33158 21899 33210
rect 21911 33158 21963 33210
rect 21975 33158 22027 33210
rect 1860 33056 1912 33108
rect 5264 33056 5316 33108
rect 7472 33056 7524 33108
rect 8024 33056 8076 33108
rect 8668 33056 8720 33108
rect 9404 33056 9456 33108
rect 3056 32920 3108 32972
rect 3516 32920 3568 32972
rect 1584 32852 1636 32904
rect 1676 32895 1728 32904
rect 1676 32861 1683 32895
rect 1683 32861 1717 32895
rect 1717 32861 1728 32895
rect 1676 32852 1728 32861
rect 1308 32784 1360 32836
rect 3608 32895 3660 32904
rect 3608 32861 3617 32895
rect 3617 32861 3651 32895
rect 3651 32861 3660 32895
rect 3608 32852 3660 32861
rect 3792 32920 3844 32972
rect 5080 32920 5132 32972
rect 6552 32920 6604 32972
rect 7288 32920 7340 32972
rect 7656 32988 7708 33040
rect 3884 32852 3936 32904
rect 3056 32827 3108 32836
rect 3056 32793 3065 32827
rect 3065 32793 3099 32827
rect 3099 32793 3108 32827
rect 3056 32784 3108 32793
rect 4252 32895 4304 32904
rect 4252 32861 4261 32895
rect 4261 32861 4295 32895
rect 4295 32861 4304 32895
rect 4252 32852 4304 32861
rect 4344 32895 4396 32904
rect 4344 32861 4353 32895
rect 4353 32861 4387 32895
rect 4387 32861 4396 32895
rect 4344 32852 4396 32861
rect 1492 32716 1544 32768
rect 2596 32716 2648 32768
rect 3608 32716 3660 32768
rect 3700 32716 3752 32768
rect 9496 32895 9548 32904
rect 9496 32861 9505 32895
rect 9505 32861 9539 32895
rect 9539 32861 9548 32895
rect 9496 32852 9548 32861
rect 9680 32920 9732 32972
rect 5724 32827 5776 32836
rect 5724 32793 5733 32827
rect 5733 32793 5767 32827
rect 5767 32793 5776 32827
rect 5724 32784 5776 32793
rect 6460 32827 6512 32836
rect 6460 32793 6469 32827
rect 6469 32793 6503 32827
rect 6503 32793 6512 32827
rect 6460 32784 6512 32793
rect 6552 32827 6604 32836
rect 6552 32793 6561 32827
rect 6561 32793 6595 32827
rect 6595 32793 6604 32827
rect 6552 32784 6604 32793
rect 6920 32827 6972 32836
rect 6920 32793 6929 32827
rect 6929 32793 6963 32827
rect 6963 32793 6972 32827
rect 6920 32784 6972 32793
rect 7104 32784 7156 32836
rect 4988 32716 5040 32768
rect 5264 32759 5316 32768
rect 5264 32725 5273 32759
rect 5273 32725 5307 32759
rect 5307 32725 5316 32759
rect 5264 32716 5316 32725
rect 9864 32784 9916 32836
rect 10048 32895 10100 32904
rect 10048 32861 10055 32895
rect 10055 32861 10089 32895
rect 10089 32861 10100 32895
rect 10048 32852 10100 32861
rect 11980 33056 12032 33108
rect 12256 33099 12308 33108
rect 12256 33065 12265 33099
rect 12265 33065 12299 33099
rect 12299 33065 12308 33099
rect 12256 33056 12308 33065
rect 12532 32920 12584 32972
rect 14096 33056 14148 33108
rect 7472 32759 7524 32768
rect 7472 32725 7481 32759
rect 7481 32725 7515 32759
rect 7515 32725 7524 32759
rect 7472 32716 7524 32725
rect 8208 32716 8260 32768
rect 10784 32759 10836 32768
rect 10784 32725 10793 32759
rect 10793 32725 10827 32759
rect 10827 32725 10836 32759
rect 10784 32716 10836 32725
rect 11980 32784 12032 32836
rect 13084 32784 13136 32836
rect 14004 32852 14056 32904
rect 14832 33056 14884 33108
rect 14372 32988 14424 33040
rect 15568 32988 15620 33040
rect 16488 33056 16540 33108
rect 17132 33056 17184 33108
rect 18052 33056 18104 33108
rect 19248 33056 19300 33108
rect 20812 33099 20864 33108
rect 20812 33065 20821 33099
rect 20821 33065 20855 33099
rect 20855 33065 20864 33099
rect 20812 33056 20864 33065
rect 16764 32920 16816 32972
rect 14832 32852 14884 32904
rect 15384 32895 15436 32904
rect 15384 32861 15393 32895
rect 15393 32861 15427 32895
rect 15427 32861 15436 32895
rect 15384 32852 15436 32861
rect 15568 32895 15620 32904
rect 15568 32861 15577 32895
rect 15577 32861 15611 32895
rect 15611 32861 15620 32895
rect 15568 32852 15620 32861
rect 16304 32895 16356 32904
rect 16304 32861 16313 32895
rect 16313 32861 16347 32895
rect 16347 32861 16356 32895
rect 16304 32852 16356 32861
rect 17592 32852 17644 32904
rect 20628 32852 20680 32904
rect 22100 33056 22152 33108
rect 23296 33056 23348 33108
rect 14372 32784 14424 32836
rect 17960 32827 18012 32836
rect 13636 32759 13688 32768
rect 13636 32725 13645 32759
rect 13645 32725 13679 32759
rect 13679 32725 13688 32759
rect 13636 32716 13688 32725
rect 14004 32716 14056 32768
rect 17960 32793 17972 32827
rect 17972 32793 18012 32827
rect 17960 32784 18012 32793
rect 19524 32827 19576 32836
rect 19524 32793 19558 32827
rect 19558 32793 19576 32827
rect 19524 32784 19576 32793
rect 21180 32784 21232 32836
rect 21640 32784 21692 32836
rect 23480 32895 23532 32904
rect 23480 32861 23489 32895
rect 23489 32861 23523 32895
rect 23523 32861 23532 32895
rect 23480 32852 23532 32861
rect 23848 32852 23900 32904
rect 19340 32716 19392 32768
rect 20720 32716 20772 32768
rect 20996 32759 21048 32768
rect 20996 32725 21005 32759
rect 21005 32725 21039 32759
rect 21039 32725 21048 32759
rect 20996 32716 21048 32725
rect 23296 32759 23348 32768
rect 23296 32725 23305 32759
rect 23305 32725 23339 32759
rect 23339 32725 23348 32759
rect 23296 32716 23348 32725
rect 23572 32759 23624 32768
rect 23572 32725 23581 32759
rect 23581 32725 23615 32759
rect 23615 32725 23624 32759
rect 23572 32716 23624 32725
rect 24124 32759 24176 32768
rect 24124 32725 24133 32759
rect 24133 32725 24167 32759
rect 24167 32725 24176 32759
rect 24124 32716 24176 32725
rect 6884 32614 6936 32666
rect 6948 32614 7000 32666
rect 7012 32614 7064 32666
rect 7076 32614 7128 32666
rect 7140 32614 7192 32666
rect 12818 32614 12870 32666
rect 12882 32614 12934 32666
rect 12946 32614 12998 32666
rect 13010 32614 13062 32666
rect 13074 32614 13126 32666
rect 18752 32614 18804 32666
rect 18816 32614 18868 32666
rect 18880 32614 18932 32666
rect 18944 32614 18996 32666
rect 19008 32614 19060 32666
rect 24686 32614 24738 32666
rect 24750 32614 24802 32666
rect 24814 32614 24866 32666
rect 24878 32614 24930 32666
rect 24942 32614 24994 32666
rect 1216 32512 1268 32564
rect 2596 32512 2648 32564
rect 2872 32512 2924 32564
rect 1492 32308 1544 32360
rect 1676 32308 1728 32360
rect 3240 32555 3292 32564
rect 3240 32521 3249 32555
rect 3249 32521 3283 32555
rect 3283 32521 3292 32555
rect 3240 32512 3292 32521
rect 3608 32512 3660 32564
rect 2136 32308 2188 32360
rect 3976 32376 4028 32428
rect 4344 32512 4396 32564
rect 5264 32512 5316 32564
rect 4252 32444 4304 32496
rect 5448 32444 5500 32496
rect 5540 32444 5592 32496
rect 6736 32444 6788 32496
rect 7472 32444 7524 32496
rect 2412 32351 2464 32360
rect 2412 32317 2446 32351
rect 2446 32317 2464 32351
rect 2412 32308 2464 32317
rect 2596 32351 2648 32360
rect 2596 32317 2605 32351
rect 2605 32317 2639 32351
rect 2639 32317 2648 32351
rect 2596 32308 2648 32317
rect 1860 32240 1912 32292
rect 7748 32444 7800 32496
rect 9496 32512 9548 32564
rect 9864 32444 9916 32496
rect 13268 32444 13320 32496
rect 14096 32487 14148 32496
rect 14096 32453 14105 32487
rect 14105 32453 14139 32487
rect 14139 32453 14148 32487
rect 14096 32444 14148 32453
rect 14464 32487 14516 32496
rect 14464 32453 14473 32487
rect 14473 32453 14507 32487
rect 14507 32453 14516 32487
rect 14464 32444 14516 32453
rect 14832 32487 14884 32496
rect 14832 32453 14841 32487
rect 14841 32453 14875 32487
rect 14875 32453 14884 32487
rect 14832 32444 14884 32453
rect 15568 32444 15620 32496
rect 16764 32444 16816 32496
rect 18052 32444 18104 32496
rect 19156 32512 19208 32564
rect 19616 32512 19668 32564
rect 20720 32555 20772 32564
rect 20720 32521 20729 32555
rect 20729 32521 20763 32555
rect 20763 32521 20772 32555
rect 20720 32512 20772 32521
rect 20812 32512 20864 32564
rect 8760 32419 8812 32428
rect 8760 32385 8769 32419
rect 8769 32385 8803 32419
rect 8803 32385 8812 32419
rect 8760 32376 8812 32385
rect 9680 32376 9732 32428
rect 10232 32376 10284 32428
rect 10692 32376 10744 32428
rect 14372 32419 14424 32428
rect 14372 32385 14381 32419
rect 14381 32385 14415 32419
rect 14415 32385 14424 32419
rect 14372 32376 14424 32385
rect 16120 32376 16172 32428
rect 16672 32419 16724 32428
rect 16672 32385 16681 32419
rect 16681 32385 16715 32419
rect 16715 32385 16724 32419
rect 16672 32376 16724 32385
rect 17040 32376 17092 32428
rect 9496 32308 9548 32360
rect 11520 32308 11572 32360
rect 13636 32308 13688 32360
rect 17868 32308 17920 32360
rect 19340 32376 19392 32428
rect 19708 32419 19760 32428
rect 19708 32385 19717 32419
rect 19717 32385 19751 32419
rect 19751 32385 19760 32419
rect 19708 32376 19760 32385
rect 20076 32376 20128 32428
rect 20536 32376 20588 32428
rect 20628 32376 20680 32428
rect 23480 32512 23532 32564
rect 23572 32512 23624 32564
rect 23756 32444 23808 32496
rect 23388 32376 23440 32428
rect 1216 32172 1268 32224
rect 1676 32172 1728 32224
rect 8116 32240 8168 32292
rect 11888 32283 11940 32292
rect 11888 32249 11897 32283
rect 11897 32249 11931 32283
rect 11931 32249 11940 32283
rect 11888 32240 11940 32249
rect 9312 32172 9364 32224
rect 10508 32172 10560 32224
rect 11060 32215 11112 32224
rect 11060 32181 11069 32215
rect 11069 32181 11103 32215
rect 11103 32181 11112 32215
rect 11060 32172 11112 32181
rect 15568 32172 15620 32224
rect 16948 32172 17000 32224
rect 19432 32308 19484 32360
rect 23572 32308 23624 32360
rect 23112 32240 23164 32292
rect 21456 32215 21508 32224
rect 21456 32181 21465 32215
rect 21465 32181 21499 32215
rect 21499 32181 21508 32215
rect 21456 32172 21508 32181
rect 23480 32215 23532 32224
rect 23480 32181 23489 32215
rect 23489 32181 23523 32215
rect 23523 32181 23532 32215
rect 23480 32172 23532 32181
rect 24400 32215 24452 32224
rect 24400 32181 24409 32215
rect 24409 32181 24443 32215
rect 24443 32181 24452 32215
rect 24400 32172 24452 32181
rect 3917 32070 3969 32122
rect 3981 32070 4033 32122
rect 4045 32070 4097 32122
rect 4109 32070 4161 32122
rect 4173 32070 4225 32122
rect 9851 32070 9903 32122
rect 9915 32070 9967 32122
rect 9979 32070 10031 32122
rect 10043 32070 10095 32122
rect 10107 32070 10159 32122
rect 15785 32070 15837 32122
rect 15849 32070 15901 32122
rect 15913 32070 15965 32122
rect 15977 32070 16029 32122
rect 16041 32070 16093 32122
rect 21719 32070 21771 32122
rect 21783 32070 21835 32122
rect 21847 32070 21899 32122
rect 21911 32070 21963 32122
rect 21975 32070 22027 32122
rect 2596 31968 2648 32020
rect 6460 31968 6512 32020
rect 6552 31968 6604 32020
rect 8760 31968 8812 32020
rect 10232 31968 10284 32020
rect 10784 31968 10836 32020
rect 14004 31968 14056 32020
rect 14096 31968 14148 32020
rect 14924 31968 14976 32020
rect 16672 31968 16724 32020
rect 17316 31968 17368 32020
rect 18420 31968 18472 32020
rect 19156 31968 19208 32020
rect 21456 31968 21508 32020
rect 5080 31832 5132 31884
rect 5356 31832 5408 31884
rect 480 31628 532 31680
rect 664 31628 716 31680
rect 1768 31764 1820 31816
rect 2780 31807 2832 31816
rect 2780 31773 2789 31807
rect 2789 31773 2823 31807
rect 2823 31773 2832 31807
rect 2780 31764 2832 31773
rect 1584 31628 1636 31680
rect 1768 31628 1820 31680
rect 2228 31628 2280 31680
rect 3240 31628 3292 31680
rect 4344 31696 4396 31748
rect 4620 31696 4672 31748
rect 4804 31696 4856 31748
rect 6920 31832 6972 31884
rect 7472 31875 7524 31884
rect 7472 31841 7481 31875
rect 7481 31841 7515 31875
rect 7515 31841 7524 31875
rect 7472 31832 7524 31841
rect 16396 31900 16448 31952
rect 18144 31900 18196 31952
rect 21364 31900 21416 31952
rect 6184 31696 6236 31748
rect 6460 31764 6512 31816
rect 6828 31764 6880 31816
rect 7656 31764 7708 31816
rect 10416 31832 10468 31884
rect 10692 31875 10744 31884
rect 10692 31841 10726 31875
rect 10726 31841 10744 31875
rect 10692 31832 10744 31841
rect 11060 31832 11112 31884
rect 11244 31832 11296 31884
rect 7564 31696 7616 31748
rect 10600 31807 10652 31816
rect 10600 31773 10609 31807
rect 10609 31773 10643 31807
rect 10643 31773 10652 31807
rect 10600 31764 10652 31773
rect 13176 31832 13228 31884
rect 16856 31875 16908 31884
rect 16856 31841 16865 31875
rect 16865 31841 16899 31875
rect 16899 31841 16908 31875
rect 16856 31832 16908 31841
rect 12072 31764 12124 31816
rect 12532 31764 12584 31816
rect 15568 31764 15620 31816
rect 5080 31628 5132 31680
rect 5908 31628 5960 31680
rect 8852 31628 8904 31680
rect 9404 31628 9456 31680
rect 9588 31628 9640 31680
rect 11796 31628 11848 31680
rect 12072 31628 12124 31680
rect 12716 31696 12768 31748
rect 14832 31696 14884 31748
rect 13268 31628 13320 31680
rect 14188 31628 14240 31680
rect 15108 31628 15160 31680
rect 16672 31807 16724 31816
rect 16672 31773 16706 31807
rect 16706 31773 16724 31807
rect 16672 31764 16724 31773
rect 17500 31764 17552 31816
rect 17776 31764 17828 31816
rect 24492 31900 24544 31952
rect 23480 31832 23532 31884
rect 16764 31628 16816 31680
rect 22836 31628 22888 31680
rect 23296 31696 23348 31748
rect 23572 31764 23624 31816
rect 23664 31807 23716 31816
rect 23664 31773 23673 31807
rect 23673 31773 23707 31807
rect 23707 31773 23716 31807
rect 23664 31764 23716 31773
rect 24216 31807 24268 31816
rect 24216 31773 24225 31807
rect 24225 31773 24259 31807
rect 24259 31773 24268 31807
rect 24216 31764 24268 31773
rect 6884 31526 6936 31578
rect 6948 31526 7000 31578
rect 7012 31526 7064 31578
rect 7076 31526 7128 31578
rect 7140 31526 7192 31578
rect 12818 31526 12870 31578
rect 12882 31526 12934 31578
rect 12946 31526 12998 31578
rect 13010 31526 13062 31578
rect 13074 31526 13126 31578
rect 18752 31526 18804 31578
rect 18816 31526 18868 31578
rect 18880 31526 18932 31578
rect 18944 31526 18996 31578
rect 19008 31526 19060 31578
rect 24686 31526 24738 31578
rect 24750 31526 24802 31578
rect 24814 31526 24866 31578
rect 24878 31526 24930 31578
rect 24942 31526 24994 31578
rect 1124 31356 1176 31408
rect 1584 31288 1636 31340
rect 2044 31288 2096 31340
rect 2596 31288 2648 31340
rect 3884 31424 3936 31476
rect 4620 31424 4672 31476
rect 1768 31220 1820 31272
rect 2780 31220 2832 31272
rect 5540 31424 5592 31476
rect 12716 31424 12768 31476
rect 12900 31424 12952 31476
rect 7564 31356 7616 31408
rect 11888 31356 11940 31408
rect 14372 31424 14424 31476
rect 18052 31424 18104 31476
rect 18604 31424 18656 31476
rect 4804 31288 4856 31340
rect 5264 31288 5316 31340
rect 5540 31288 5592 31340
rect 5724 31288 5776 31340
rect 7472 31288 7524 31340
rect 8944 31288 8996 31340
rect 12900 31288 12952 31340
rect 13084 31331 13136 31340
rect 13084 31297 13093 31331
rect 13093 31297 13127 31331
rect 13127 31297 13136 31331
rect 13084 31288 13136 31297
rect 13452 31288 13504 31340
rect 13912 31399 13964 31408
rect 13912 31365 13921 31399
rect 13921 31365 13955 31399
rect 13955 31365 13964 31399
rect 13912 31356 13964 31365
rect 22836 31467 22888 31476
rect 22836 31433 22845 31467
rect 22845 31433 22879 31467
rect 22879 31433 22888 31467
rect 22836 31424 22888 31433
rect 23480 31424 23532 31476
rect 23940 31424 23992 31476
rect 23020 31356 23072 31408
rect 16028 31288 16080 31340
rect 18144 31331 18196 31340
rect 18144 31297 18153 31331
rect 18153 31297 18187 31331
rect 18187 31297 18196 31331
rect 18144 31288 18196 31297
rect 22192 31288 22244 31340
rect 9036 31220 9088 31272
rect 12440 31220 12492 31272
rect 13268 31220 13320 31272
rect 14188 31220 14240 31272
rect 19708 31220 19760 31272
rect 21824 31263 21876 31272
rect 21824 31229 21833 31263
rect 21833 31229 21867 31263
rect 21867 31229 21876 31263
rect 21824 31220 21876 31229
rect 4620 31152 4672 31204
rect 3056 31084 3108 31136
rect 4528 31084 4580 31136
rect 4804 31084 4856 31136
rect 6368 31152 6420 31204
rect 12256 31152 12308 31204
rect 5908 31127 5960 31136
rect 5908 31093 5917 31127
rect 5917 31093 5951 31127
rect 5951 31093 5960 31127
rect 5908 31084 5960 31093
rect 8576 31084 8628 31136
rect 9220 31084 9272 31136
rect 9680 31084 9732 31136
rect 10692 31084 10744 31136
rect 10968 31084 11020 31136
rect 12624 31084 12676 31136
rect 18696 31152 18748 31204
rect 25044 31288 25096 31340
rect 16488 31084 16540 31136
rect 18604 31084 18656 31136
rect 20536 31084 20588 31136
rect 23204 31127 23256 31136
rect 23204 31093 23213 31127
rect 23213 31093 23247 31127
rect 23247 31093 23256 31127
rect 23204 31084 23256 31093
rect 24400 31127 24452 31136
rect 24400 31093 24409 31127
rect 24409 31093 24443 31127
rect 24443 31093 24452 31127
rect 24400 31084 24452 31093
rect 3917 30982 3969 31034
rect 3981 30982 4033 31034
rect 4045 30982 4097 31034
rect 4109 30982 4161 31034
rect 4173 30982 4225 31034
rect 9851 30982 9903 31034
rect 9915 30982 9967 31034
rect 9979 30982 10031 31034
rect 10043 30982 10095 31034
rect 10107 30982 10159 31034
rect 15785 30982 15837 31034
rect 15849 30982 15901 31034
rect 15913 30982 15965 31034
rect 15977 30982 16029 31034
rect 16041 30982 16093 31034
rect 21719 30982 21771 31034
rect 21783 30982 21835 31034
rect 21847 30982 21899 31034
rect 21911 30982 21963 31034
rect 21975 30982 22027 31034
rect 3608 30880 3660 30932
rect 4804 30880 4856 30932
rect 6092 30923 6144 30932
rect 6092 30889 6101 30923
rect 6101 30889 6135 30923
rect 6135 30889 6144 30923
rect 6092 30880 6144 30889
rect 6460 30880 6512 30932
rect 7380 30880 7432 30932
rect 9680 30880 9732 30932
rect 480 30812 532 30864
rect 10508 30880 10560 30932
rect 12256 30923 12308 30932
rect 12256 30889 12265 30923
rect 12265 30889 12299 30923
rect 12299 30889 12308 30923
rect 12256 30880 12308 30889
rect 12440 30880 12492 30932
rect 1400 30719 1452 30728
rect 1400 30685 1409 30719
rect 1409 30685 1443 30719
rect 1443 30685 1452 30719
rect 1400 30676 1452 30685
rect 1768 30676 1820 30728
rect 1952 30676 2004 30728
rect 2504 30676 2556 30728
rect 2688 30676 2740 30728
rect 5080 30744 5132 30796
rect 5908 30744 5960 30796
rect 7472 30787 7524 30796
rect 7472 30753 7481 30787
rect 7481 30753 7515 30787
rect 7515 30753 7524 30787
rect 7472 30744 7524 30753
rect 3976 30676 4028 30728
rect 4896 30676 4948 30728
rect 7288 30676 7340 30728
rect 9956 30744 10008 30796
rect 3332 30583 3384 30592
rect 3332 30549 3341 30583
rect 3341 30549 3375 30583
rect 3375 30549 3384 30583
rect 3332 30540 3384 30549
rect 3516 30540 3568 30592
rect 4068 30540 4120 30592
rect 4804 30583 4856 30592
rect 4804 30549 4813 30583
rect 4813 30549 4847 30583
rect 4847 30549 4856 30583
rect 4804 30540 4856 30549
rect 5080 30651 5132 30660
rect 5080 30617 5089 30651
rect 5089 30617 5123 30651
rect 5123 30617 5132 30651
rect 5080 30608 5132 30617
rect 5724 30608 5776 30660
rect 8668 30676 8720 30728
rect 11704 30676 11756 30728
rect 13452 30880 13504 30932
rect 14832 30880 14884 30932
rect 16304 30880 16356 30932
rect 18604 30880 18656 30932
rect 23020 30923 23072 30932
rect 23020 30889 23029 30923
rect 23029 30889 23063 30923
rect 23063 30889 23072 30923
rect 23020 30880 23072 30889
rect 23204 30880 23256 30932
rect 23388 30880 23440 30932
rect 12532 30744 12584 30796
rect 13452 30744 13504 30796
rect 13820 30744 13872 30796
rect 14464 30744 14516 30796
rect 15016 30744 15068 30796
rect 15568 30744 15620 30796
rect 15936 30787 15988 30796
rect 15936 30753 15945 30787
rect 15945 30753 15979 30787
rect 15979 30753 15988 30787
rect 15936 30744 15988 30753
rect 16304 30787 16356 30796
rect 16304 30753 16338 30787
rect 16338 30753 16356 30787
rect 16304 30744 16356 30753
rect 16488 30787 16540 30796
rect 16488 30753 16497 30787
rect 16497 30753 16531 30787
rect 16531 30753 16540 30787
rect 16488 30744 16540 30753
rect 17500 30787 17552 30796
rect 17500 30753 17509 30787
rect 17509 30753 17543 30787
rect 17543 30753 17552 30787
rect 17500 30744 17552 30753
rect 14740 30676 14792 30728
rect 15292 30719 15344 30728
rect 15292 30685 15301 30719
rect 15301 30685 15335 30719
rect 15335 30685 15344 30719
rect 15292 30676 15344 30685
rect 15476 30719 15528 30728
rect 15476 30685 15485 30719
rect 15485 30685 15519 30719
rect 15519 30685 15528 30719
rect 15476 30676 15528 30685
rect 15660 30676 15712 30728
rect 18144 30676 18196 30728
rect 18972 30812 19024 30864
rect 20076 30812 20128 30864
rect 5908 30583 5960 30592
rect 5908 30549 5917 30583
rect 5917 30549 5951 30583
rect 5951 30549 5960 30583
rect 5908 30540 5960 30549
rect 8944 30608 8996 30660
rect 9036 30608 9088 30660
rect 18972 30608 19024 30660
rect 7564 30540 7616 30592
rect 7748 30540 7800 30592
rect 7932 30540 7984 30592
rect 8116 30540 8168 30592
rect 9496 30540 9548 30592
rect 10508 30540 10560 30592
rect 11060 30583 11112 30592
rect 11060 30549 11069 30583
rect 11069 30549 11103 30583
rect 11103 30549 11112 30583
rect 11060 30540 11112 30549
rect 11612 30583 11664 30592
rect 11612 30549 11621 30583
rect 11621 30549 11655 30583
rect 11655 30549 11664 30583
rect 11612 30540 11664 30549
rect 14832 30540 14884 30592
rect 19248 30540 19300 30592
rect 19340 30583 19392 30592
rect 19340 30549 19349 30583
rect 19349 30549 19383 30583
rect 19383 30549 19392 30583
rect 19340 30540 19392 30549
rect 19616 30583 19668 30592
rect 19616 30549 19625 30583
rect 19625 30549 19659 30583
rect 19659 30549 19668 30583
rect 19616 30540 19668 30549
rect 21456 30676 21508 30728
rect 23204 30719 23256 30728
rect 23204 30685 23213 30719
rect 23213 30685 23247 30719
rect 23247 30685 23256 30719
rect 23204 30676 23256 30685
rect 23848 30651 23900 30660
rect 23848 30617 23857 30651
rect 23857 30617 23891 30651
rect 23891 30617 23900 30651
rect 23848 30608 23900 30617
rect 24216 30651 24268 30660
rect 24216 30617 24225 30651
rect 24225 30617 24259 30651
rect 24259 30617 24268 30651
rect 24216 30608 24268 30617
rect 20352 30540 20404 30592
rect 20812 30540 20864 30592
rect 20904 30540 20956 30592
rect 21088 30583 21140 30592
rect 21088 30549 21097 30583
rect 21097 30549 21131 30583
rect 21131 30549 21140 30583
rect 21088 30540 21140 30549
rect 22836 30540 22888 30592
rect 23572 30540 23624 30592
rect 6884 30438 6936 30490
rect 6948 30438 7000 30490
rect 7012 30438 7064 30490
rect 7076 30438 7128 30490
rect 7140 30438 7192 30490
rect 12818 30438 12870 30490
rect 12882 30438 12934 30490
rect 12946 30438 12998 30490
rect 13010 30438 13062 30490
rect 13074 30438 13126 30490
rect 18752 30438 18804 30490
rect 18816 30438 18868 30490
rect 18880 30438 18932 30490
rect 18944 30438 18996 30490
rect 19008 30438 19060 30490
rect 24686 30438 24738 30490
rect 24750 30438 24802 30490
rect 24814 30438 24866 30490
rect 24878 30438 24930 30490
rect 24942 30438 24994 30490
rect 1308 30336 1360 30388
rect 2780 30336 2832 30388
rect 2688 30311 2740 30320
rect 2688 30277 2697 30311
rect 2697 30277 2731 30311
rect 2731 30277 2740 30311
rect 2688 30268 2740 30277
rect 3332 30336 3384 30388
rect 3976 30379 4028 30388
rect 3976 30345 3985 30379
rect 3985 30345 4019 30379
rect 4019 30345 4028 30379
rect 3976 30336 4028 30345
rect 1492 30200 1544 30252
rect 1676 30200 1728 30252
rect 2780 30200 2832 30252
rect 3240 30200 3292 30252
rect 3424 30243 3476 30252
rect 3424 30209 3433 30243
rect 3433 30209 3467 30243
rect 3467 30209 3476 30243
rect 4252 30268 4304 30320
rect 6184 30336 6236 30388
rect 8024 30336 8076 30388
rect 9680 30336 9732 30388
rect 3424 30200 3476 30209
rect 5172 30243 5224 30252
rect 5172 30209 5181 30243
rect 5181 30209 5224 30243
rect 1584 30175 1636 30184
rect 1584 30141 1593 30175
rect 1593 30141 1627 30175
rect 1627 30141 1636 30175
rect 1584 30132 1636 30141
rect 2136 30132 2188 30184
rect 3056 30132 3108 30184
rect 5172 30200 5224 30209
rect 5540 30200 5592 30252
rect 6276 30200 6328 30252
rect 1492 30064 1544 30116
rect 4804 30107 4856 30116
rect 4804 30073 4813 30107
rect 4813 30073 4847 30107
rect 4847 30073 4856 30107
rect 4804 30064 4856 30073
rect 2136 30039 2188 30048
rect 2136 30005 2145 30039
rect 2145 30005 2179 30039
rect 2179 30005 2188 30039
rect 2136 29996 2188 30005
rect 4712 29996 4764 30048
rect 5356 29996 5408 30048
rect 6184 30132 6236 30184
rect 8208 30311 8260 30320
rect 8208 30277 8217 30311
rect 8217 30277 8251 30311
rect 8251 30277 8260 30311
rect 8208 30268 8260 30277
rect 8576 30268 8628 30320
rect 9036 30311 9088 30320
rect 9036 30277 9045 30311
rect 9045 30277 9079 30311
rect 9079 30277 9088 30311
rect 9036 30268 9088 30277
rect 11520 30268 11572 30320
rect 15936 30336 15988 30388
rect 7656 30200 7708 30252
rect 8668 30243 8720 30252
rect 8668 30209 8677 30243
rect 8677 30209 8711 30243
rect 8711 30209 8720 30243
rect 8668 30200 8720 30209
rect 8852 30200 8904 30252
rect 8116 30132 8168 30184
rect 9036 30132 9088 30184
rect 9864 30200 9916 30252
rect 9680 30175 9732 30184
rect 9680 30141 9689 30175
rect 9689 30141 9723 30175
rect 9723 30141 9732 30175
rect 9680 30132 9732 30141
rect 10048 30132 10100 30184
rect 12072 30243 12124 30252
rect 12072 30209 12081 30243
rect 12081 30209 12115 30243
rect 12115 30209 12124 30243
rect 12072 30200 12124 30209
rect 10508 30175 10560 30184
rect 10508 30141 10542 30175
rect 10542 30141 10560 30175
rect 10508 30132 10560 30141
rect 11060 30132 11112 30184
rect 10232 30064 10284 30116
rect 17316 30268 17368 30320
rect 19248 30336 19300 30388
rect 20444 30268 20496 30320
rect 21456 30379 21508 30388
rect 21456 30345 21465 30379
rect 21465 30345 21499 30379
rect 21499 30345 21508 30379
rect 21456 30336 21508 30345
rect 23572 30379 23624 30388
rect 23572 30345 23581 30379
rect 23581 30345 23615 30379
rect 23615 30345 23624 30379
rect 23572 30336 23624 30345
rect 17960 30243 18012 30252
rect 17960 30209 17969 30243
rect 17969 30209 18003 30243
rect 18003 30209 18012 30243
rect 17960 30200 18012 30209
rect 18236 30243 18288 30252
rect 18236 30209 18243 30243
rect 18243 30209 18277 30243
rect 18277 30209 18288 30243
rect 18236 30200 18288 30209
rect 19064 30200 19116 30252
rect 20904 30200 20956 30252
rect 21088 30205 21140 30250
rect 21088 30198 21097 30205
rect 21097 30198 21131 30205
rect 21131 30198 21140 30205
rect 21180 30243 21232 30252
rect 21180 30209 21189 30243
rect 21189 30209 21223 30243
rect 21223 30209 21232 30243
rect 21180 30200 21232 30209
rect 22836 30268 22888 30320
rect 14188 30132 14240 30184
rect 5908 30039 5960 30048
rect 5908 30005 5917 30039
rect 5917 30005 5951 30039
rect 5951 30005 5960 30039
rect 5908 29996 5960 30005
rect 7380 30039 7432 30048
rect 7380 30005 7389 30039
rect 7389 30005 7423 30039
rect 7423 30005 7432 30039
rect 7380 29996 7432 30005
rect 7932 29996 7984 30048
rect 9220 30039 9272 30048
rect 9220 30005 9229 30039
rect 9229 30005 9263 30039
rect 9263 30005 9272 30039
rect 9220 29996 9272 30005
rect 11336 30039 11388 30048
rect 11336 30005 11345 30039
rect 11345 30005 11379 30039
rect 11379 30005 11388 30039
rect 11336 29996 11388 30005
rect 12716 29996 12768 30048
rect 14464 30064 14516 30116
rect 15476 29996 15528 30048
rect 17960 29996 18012 30048
rect 18236 29996 18288 30048
rect 23020 30200 23072 30252
rect 23388 30200 23440 30252
rect 23572 30200 23624 30252
rect 20628 29996 20680 30048
rect 20996 30039 21048 30048
rect 20996 30005 21005 30039
rect 21005 30005 21039 30039
rect 21039 30005 21048 30039
rect 20996 29996 21048 30005
rect 22560 29996 22612 30048
rect 23848 29996 23900 30048
rect 24400 30039 24452 30048
rect 24400 30005 24409 30039
rect 24409 30005 24443 30039
rect 24443 30005 24452 30039
rect 24400 29996 24452 30005
rect 3917 29894 3969 29946
rect 3981 29894 4033 29946
rect 4045 29894 4097 29946
rect 4109 29894 4161 29946
rect 4173 29894 4225 29946
rect 9851 29894 9903 29946
rect 9915 29894 9967 29946
rect 9979 29894 10031 29946
rect 10043 29894 10095 29946
rect 10107 29894 10159 29946
rect 15785 29894 15837 29946
rect 15849 29894 15901 29946
rect 15913 29894 15965 29946
rect 15977 29894 16029 29946
rect 16041 29894 16093 29946
rect 21719 29894 21771 29946
rect 21783 29894 21835 29946
rect 21847 29894 21899 29946
rect 21911 29894 21963 29946
rect 21975 29894 22027 29946
rect 1400 29588 1452 29640
rect 1952 29792 2004 29844
rect 2320 29792 2372 29844
rect 2412 29792 2464 29844
rect 3608 29792 3660 29844
rect 3792 29792 3844 29844
rect 2228 29588 2280 29640
rect 2688 29724 2740 29776
rect 3516 29656 3568 29708
rect 5080 29767 5132 29776
rect 5080 29733 5089 29767
rect 5089 29733 5123 29767
rect 5123 29733 5132 29767
rect 5080 29724 5132 29733
rect 4068 29699 4120 29708
rect 4068 29665 4077 29699
rect 4077 29665 4111 29699
rect 4111 29665 4120 29699
rect 4068 29656 4120 29665
rect 3056 29588 3108 29640
rect 1308 29520 1360 29572
rect 4252 29588 4304 29640
rect 4896 29588 4948 29640
rect 5908 29656 5960 29708
rect 5356 29520 5408 29572
rect 6644 29588 6696 29640
rect 7380 29588 7432 29640
rect 7196 29520 7248 29572
rect 11520 29792 11572 29844
rect 12072 29792 12124 29844
rect 8208 29724 8260 29776
rect 9496 29724 9548 29776
rect 8576 29588 8628 29640
rect 9496 29588 9548 29640
rect 9772 29724 9824 29776
rect 10140 29656 10192 29708
rect 12532 29724 12584 29776
rect 15200 29792 15252 29844
rect 15752 29792 15804 29844
rect 19340 29835 19392 29844
rect 19340 29801 19349 29835
rect 19349 29801 19383 29835
rect 19383 29801 19392 29835
rect 19340 29792 19392 29801
rect 19616 29792 19668 29844
rect 10876 29656 10928 29708
rect 15476 29724 15528 29776
rect 16488 29767 16540 29776
rect 16488 29733 16497 29767
rect 16497 29733 16531 29767
rect 16531 29733 16540 29767
rect 16488 29724 16540 29733
rect 19800 29724 19852 29776
rect 2596 29452 2648 29504
rect 2688 29452 2740 29504
rect 3700 29452 3752 29504
rect 5908 29452 5960 29504
rect 9404 29520 9456 29572
rect 9864 29588 9916 29640
rect 10968 29631 11020 29640
rect 10968 29597 10977 29631
rect 10977 29597 11011 29631
rect 11011 29597 11020 29631
rect 10968 29588 11020 29597
rect 11612 29588 11664 29640
rect 11980 29631 12032 29640
rect 11980 29597 11987 29631
rect 11987 29597 12021 29631
rect 12021 29597 12032 29631
rect 11980 29588 12032 29597
rect 12716 29588 12768 29640
rect 14004 29588 14056 29640
rect 13636 29563 13688 29572
rect 13636 29529 13645 29563
rect 13645 29529 13679 29563
rect 13679 29529 13688 29563
rect 13636 29520 13688 29529
rect 14832 29588 14884 29640
rect 14556 29520 14608 29572
rect 15752 29631 15804 29640
rect 15752 29597 15759 29631
rect 15759 29597 15793 29631
rect 15793 29597 15804 29631
rect 15752 29588 15804 29597
rect 16304 29588 16356 29640
rect 19248 29631 19300 29640
rect 19248 29597 19257 29631
rect 19257 29597 19291 29631
rect 19291 29597 19300 29631
rect 19248 29588 19300 29597
rect 19432 29588 19484 29640
rect 20904 29835 20956 29844
rect 20904 29801 20913 29835
rect 20913 29801 20947 29835
rect 20947 29801 20956 29835
rect 20904 29792 20956 29801
rect 22560 29792 22612 29844
rect 23572 29792 23624 29844
rect 23388 29724 23440 29776
rect 21088 29656 21140 29708
rect 22284 29656 22336 29708
rect 20168 29631 20220 29640
rect 17040 29520 17092 29572
rect 19064 29520 19116 29572
rect 20168 29597 20175 29631
rect 20175 29597 20209 29631
rect 20209 29597 20220 29631
rect 20168 29588 20220 29597
rect 21180 29588 21232 29640
rect 21640 29631 21692 29640
rect 21640 29597 21647 29631
rect 21647 29597 21681 29631
rect 21681 29597 21692 29631
rect 21640 29588 21692 29597
rect 7748 29452 7800 29504
rect 8852 29452 8904 29504
rect 10876 29452 10928 29504
rect 14372 29452 14424 29504
rect 14648 29452 14700 29504
rect 19248 29452 19300 29504
rect 19524 29495 19576 29504
rect 19524 29461 19533 29495
rect 19533 29461 19567 29495
rect 19567 29461 19576 29495
rect 19524 29452 19576 29461
rect 21824 29520 21876 29572
rect 22928 29520 22980 29572
rect 25320 29588 25372 29640
rect 22376 29495 22428 29504
rect 22376 29461 22385 29495
rect 22385 29461 22419 29495
rect 22419 29461 22428 29495
rect 22376 29452 22428 29461
rect 24216 29563 24268 29572
rect 24216 29529 24225 29563
rect 24225 29529 24259 29563
rect 24259 29529 24268 29563
rect 24216 29520 24268 29529
rect 6884 29350 6936 29402
rect 6948 29350 7000 29402
rect 7012 29350 7064 29402
rect 7076 29350 7128 29402
rect 7140 29350 7192 29402
rect 12818 29350 12870 29402
rect 12882 29350 12934 29402
rect 12946 29350 12998 29402
rect 13010 29350 13062 29402
rect 13074 29350 13126 29402
rect 18752 29350 18804 29402
rect 18816 29350 18868 29402
rect 18880 29350 18932 29402
rect 18944 29350 18996 29402
rect 19008 29350 19060 29402
rect 24686 29350 24738 29402
rect 24750 29350 24802 29402
rect 24814 29350 24866 29402
rect 24878 29350 24930 29402
rect 24942 29350 24994 29402
rect 1124 29248 1176 29300
rect 2320 29155 2372 29164
rect 2320 29121 2329 29155
rect 2329 29121 2363 29155
rect 2363 29121 2372 29155
rect 2320 29112 2372 29121
rect 2596 29155 2648 29164
rect 2596 29121 2605 29155
rect 2605 29121 2639 29155
rect 2639 29121 2648 29155
rect 2596 29112 2648 29121
rect 4712 29248 4764 29300
rect 7748 29248 7800 29300
rect 1400 29087 1452 29096
rect 1400 29053 1409 29087
rect 1409 29053 1443 29087
rect 1443 29053 1452 29087
rect 1400 29044 1452 29053
rect 3884 29112 3936 29164
rect 4896 29112 4948 29164
rect 6092 29112 6144 29164
rect 9588 29248 9640 29300
rect 10140 29291 10192 29300
rect 10140 29257 10149 29291
rect 10149 29257 10183 29291
rect 10183 29257 10192 29291
rect 10140 29248 10192 29257
rect 10784 29248 10836 29300
rect 11336 29248 11388 29300
rect 8852 29112 8904 29164
rect 9680 29180 9732 29232
rect 9588 29122 9640 29174
rect 13636 29248 13688 29300
rect 14372 29248 14424 29300
rect 1860 28976 1912 29028
rect 2044 29019 2096 29028
rect 2044 28985 2053 29019
rect 2053 28985 2087 29019
rect 2087 28985 2096 29019
rect 2044 28976 2096 28985
rect 4160 29044 4212 29096
rect 4528 29044 4580 29096
rect 6644 29044 6696 29096
rect 7380 29044 7432 29096
rect 9036 29044 9088 29096
rect 12532 29112 12584 29164
rect 13176 29180 13228 29232
rect 22284 29180 22336 29232
rect 12992 29155 13044 29164
rect 12992 29121 12999 29155
rect 12999 29121 13033 29155
rect 13033 29121 13044 29155
rect 12992 29112 13044 29121
rect 13728 29112 13780 29164
rect 1584 28908 1636 28960
rect 3516 28908 3568 28960
rect 3608 28908 3660 28960
rect 5540 28908 5592 28960
rect 7288 28976 7340 29028
rect 7748 28976 7800 29028
rect 8392 28976 8444 29028
rect 10232 28976 10284 29028
rect 12256 28976 12308 29028
rect 13912 29044 13964 29096
rect 8300 28908 8352 28960
rect 8852 28908 8904 28960
rect 9864 28908 9916 28960
rect 14004 28976 14056 29028
rect 15108 29019 15160 29028
rect 15108 28985 15117 29019
rect 15117 28985 15151 29019
rect 15151 28985 15160 29019
rect 15108 28976 15160 28985
rect 16948 29112 17000 29164
rect 17408 29112 17460 29164
rect 17868 29112 17920 29164
rect 20720 29112 20772 29164
rect 21364 29155 21416 29164
rect 21364 29121 21373 29155
rect 21373 29121 21407 29155
rect 21407 29121 21416 29155
rect 21364 29112 21416 29121
rect 17040 29087 17092 29096
rect 17040 29053 17049 29087
rect 17049 29053 17083 29087
rect 17083 29053 17092 29087
rect 17040 29044 17092 29053
rect 21824 29112 21876 29164
rect 22376 29155 22428 29164
rect 22376 29121 22385 29155
rect 22385 29121 22419 29155
rect 22419 29121 22428 29155
rect 22376 29112 22428 29121
rect 22560 29155 22612 29164
rect 22560 29121 22569 29155
rect 22569 29121 22603 29155
rect 22603 29121 22612 29155
rect 22560 29112 22612 29121
rect 14832 28908 14884 28960
rect 22100 28976 22152 29028
rect 22928 29019 22980 29028
rect 22928 28985 22937 29019
rect 22937 28985 22971 29019
rect 22971 28985 22980 29019
rect 22928 28976 22980 28985
rect 23388 28976 23440 29028
rect 24124 29155 24176 29164
rect 24124 29121 24133 29155
rect 24133 29121 24167 29155
rect 24167 29121 24176 29155
rect 24124 29112 24176 29121
rect 24400 29019 24452 29028
rect 24400 28985 24409 29019
rect 24409 28985 24443 29019
rect 24443 28985 24452 29019
rect 24400 28976 24452 28985
rect 18420 28908 18472 28960
rect 18604 28908 18656 28960
rect 21732 28908 21784 28960
rect 22468 28951 22520 28960
rect 22468 28917 22477 28951
rect 22477 28917 22511 28951
rect 22511 28917 22520 28951
rect 22468 28908 22520 28917
rect 23940 28908 23992 28960
rect 3917 28806 3969 28858
rect 3981 28806 4033 28858
rect 4045 28806 4097 28858
rect 4109 28806 4161 28858
rect 4173 28806 4225 28858
rect 9851 28806 9903 28858
rect 9915 28806 9967 28858
rect 9979 28806 10031 28858
rect 10043 28806 10095 28858
rect 10107 28806 10159 28858
rect 15785 28806 15837 28858
rect 15849 28806 15901 28858
rect 15913 28806 15965 28858
rect 15977 28806 16029 28858
rect 16041 28806 16093 28858
rect 21719 28806 21771 28858
rect 21783 28806 21835 28858
rect 21847 28806 21899 28858
rect 21911 28806 21963 28858
rect 21975 28806 22027 28858
rect 1952 28704 2004 28756
rect 3608 28704 3660 28756
rect 5908 28704 5960 28756
rect 8024 28704 8076 28756
rect 10600 28704 10652 28756
rect 18604 28704 18656 28756
rect 19248 28704 19300 28756
rect 19340 28704 19392 28756
rect 1216 28500 1268 28552
rect 2320 28543 2372 28552
rect 2320 28509 2329 28543
rect 2329 28509 2363 28543
rect 2363 28509 2372 28543
rect 2320 28500 2372 28509
rect 2504 28500 2556 28552
rect 2688 28500 2740 28552
rect 756 28432 808 28484
rect 3884 28432 3936 28484
rect 1952 28407 2004 28416
rect 1952 28373 1961 28407
rect 1961 28373 1995 28407
rect 1995 28373 2004 28407
rect 1952 28364 2004 28373
rect 2596 28364 2648 28416
rect 3792 28364 3844 28416
rect 5540 28500 5592 28552
rect 5908 28500 5960 28552
rect 4344 28475 4396 28484
rect 4344 28441 4353 28475
rect 4353 28441 4387 28475
rect 4387 28441 4396 28475
rect 4344 28432 4396 28441
rect 5172 28432 5224 28484
rect 5264 28432 5316 28484
rect 8668 28636 8720 28688
rect 15476 28636 15528 28688
rect 7472 28568 7524 28620
rect 6276 28543 6328 28552
rect 6276 28509 6285 28543
rect 6285 28509 6319 28543
rect 6319 28509 6328 28543
rect 6276 28500 6328 28509
rect 6552 28543 6604 28552
rect 6552 28509 6561 28543
rect 6561 28509 6604 28543
rect 6552 28500 6604 28509
rect 6644 28500 6696 28552
rect 11612 28568 11664 28620
rect 11888 28568 11940 28620
rect 12164 28568 12216 28620
rect 15936 28611 15988 28620
rect 15936 28577 15945 28611
rect 15945 28577 15979 28611
rect 15979 28577 15988 28611
rect 15936 28568 15988 28577
rect 17868 28679 17920 28688
rect 17868 28645 17877 28679
rect 17877 28645 17911 28679
rect 17911 28645 17920 28679
rect 17868 28636 17920 28645
rect 21364 28704 21416 28756
rect 22560 28704 22612 28756
rect 23388 28747 23440 28756
rect 23388 28713 23397 28747
rect 23397 28713 23431 28747
rect 23431 28713 23440 28747
rect 23388 28704 23440 28713
rect 16488 28611 16540 28620
rect 16488 28577 16497 28611
rect 16497 28577 16531 28611
rect 16531 28577 16540 28611
rect 16488 28568 16540 28577
rect 8208 28500 8260 28552
rect 4896 28364 4948 28416
rect 12440 28432 12492 28484
rect 15292 28543 15344 28552
rect 15292 28509 15301 28543
rect 15301 28509 15335 28543
rect 15335 28509 15344 28543
rect 15292 28500 15344 28509
rect 15660 28500 15712 28552
rect 16212 28543 16264 28552
rect 16212 28509 16221 28543
rect 16221 28509 16255 28543
rect 16255 28509 16264 28543
rect 16212 28500 16264 28509
rect 17500 28568 17552 28620
rect 18144 28611 18196 28620
rect 18144 28577 18153 28611
rect 18153 28577 18187 28611
rect 18187 28577 18196 28611
rect 18144 28568 18196 28577
rect 18604 28568 18656 28620
rect 20444 28636 20496 28688
rect 7288 28407 7340 28416
rect 7288 28373 7297 28407
rect 7297 28373 7331 28407
rect 7331 28373 7340 28407
rect 7288 28364 7340 28373
rect 8024 28364 8076 28416
rect 12624 28364 12676 28416
rect 12716 28364 12768 28416
rect 18236 28543 18288 28552
rect 18236 28509 18270 28543
rect 18270 28509 18288 28543
rect 18236 28500 18288 28509
rect 18420 28543 18472 28552
rect 18420 28509 18429 28543
rect 18429 28509 18463 28543
rect 18463 28509 18472 28543
rect 18420 28500 18472 28509
rect 19800 28500 19852 28552
rect 19892 28543 19944 28552
rect 19892 28509 19901 28543
rect 19901 28509 19935 28543
rect 19935 28509 19944 28543
rect 19892 28500 19944 28509
rect 20444 28500 20496 28552
rect 20628 28543 20680 28552
rect 20628 28509 20637 28543
rect 20637 28509 20671 28543
rect 20671 28509 20680 28543
rect 20628 28500 20680 28509
rect 22192 28636 22244 28688
rect 23848 28636 23900 28688
rect 22468 28611 22520 28620
rect 22468 28577 22477 28611
rect 22477 28577 22511 28611
rect 22511 28577 22520 28611
rect 22468 28568 22520 28577
rect 13268 28364 13320 28416
rect 13912 28364 13964 28416
rect 16212 28364 16264 28416
rect 16488 28364 16540 28416
rect 16580 28364 16632 28416
rect 18420 28364 18472 28416
rect 18880 28364 18932 28416
rect 19248 28364 19300 28416
rect 22376 28500 22428 28552
rect 22560 28543 22612 28552
rect 22560 28509 22569 28543
rect 22569 28509 22603 28543
rect 22603 28509 22612 28543
rect 22560 28500 22612 28509
rect 20076 28407 20128 28416
rect 20076 28373 20085 28407
rect 20085 28373 20119 28407
rect 20119 28373 20128 28407
rect 20076 28364 20128 28373
rect 20536 28364 20588 28416
rect 23296 28543 23348 28552
rect 23296 28509 23305 28543
rect 23305 28509 23339 28543
rect 23339 28509 23348 28543
rect 23296 28500 23348 28509
rect 23664 28500 23716 28552
rect 23940 28543 23992 28552
rect 23940 28509 23949 28543
rect 23949 28509 23983 28543
rect 23983 28509 23992 28543
rect 23940 28500 23992 28509
rect 23664 28407 23716 28416
rect 23664 28373 23673 28407
rect 23673 28373 23707 28407
rect 23707 28373 23716 28407
rect 23664 28364 23716 28373
rect 24124 28407 24176 28416
rect 24124 28373 24133 28407
rect 24133 28373 24167 28407
rect 24167 28373 24176 28407
rect 24124 28364 24176 28373
rect 6884 28262 6936 28314
rect 6948 28262 7000 28314
rect 7012 28262 7064 28314
rect 7076 28262 7128 28314
rect 7140 28262 7192 28314
rect 12818 28262 12870 28314
rect 12882 28262 12934 28314
rect 12946 28262 12998 28314
rect 13010 28262 13062 28314
rect 13074 28262 13126 28314
rect 18752 28262 18804 28314
rect 18816 28262 18868 28314
rect 18880 28262 18932 28314
rect 18944 28262 18996 28314
rect 19008 28262 19060 28314
rect 24686 28262 24738 28314
rect 24750 28262 24802 28314
rect 24814 28262 24866 28314
rect 24878 28262 24930 28314
rect 24942 28262 24994 28314
rect 2044 28160 2096 28212
rect 3516 28160 3568 28212
rect 4344 28160 4396 28212
rect 4620 28203 4672 28212
rect 4620 28169 4629 28203
rect 4629 28169 4663 28203
rect 4663 28169 4672 28203
rect 4620 28160 4672 28169
rect 2228 28092 2280 28144
rect 3056 28092 3108 28144
rect 5172 28092 5224 28144
rect 6552 28160 6604 28212
rect 7380 28092 7432 28144
rect 1768 28024 1820 28076
rect 2504 28024 2556 28076
rect 2780 28067 2832 28076
rect 2780 28033 2789 28067
rect 2789 28033 2823 28067
rect 2823 28033 2832 28067
rect 2780 28024 2832 28033
rect 1400 27999 1452 28008
rect 1400 27965 1409 27999
rect 1409 27965 1443 27999
rect 1443 27965 1452 27999
rect 1400 27956 1452 27965
rect 2136 27956 2188 28008
rect 2412 27956 2464 28008
rect 2596 27888 2648 27940
rect 2136 27820 2188 27872
rect 2320 27820 2372 27872
rect 5908 28024 5960 28076
rect 10968 28160 11020 28212
rect 8668 28092 8720 28144
rect 5080 27956 5132 28008
rect 6644 27956 6696 28008
rect 8208 28024 8260 28076
rect 10600 28092 10652 28144
rect 11244 28160 11296 28212
rect 12440 28160 12492 28212
rect 15752 28160 15804 28212
rect 17868 28160 17920 28212
rect 18420 28160 18472 28212
rect 19892 28160 19944 28212
rect 20536 28160 20588 28212
rect 21640 28160 21692 28212
rect 22192 28160 22244 28212
rect 23572 28160 23624 28212
rect 23664 28160 23716 28212
rect 11520 28067 11572 28076
rect 11520 28033 11529 28067
rect 11529 28033 11563 28067
rect 11563 28033 11572 28067
rect 11520 28024 11572 28033
rect 11612 28024 11664 28076
rect 5908 27931 5960 27940
rect 5908 27897 5917 27931
rect 5917 27897 5951 27931
rect 5951 27897 5960 27931
rect 5908 27888 5960 27897
rect 4252 27820 4304 27872
rect 4436 27820 4488 27872
rect 8300 27863 8352 27872
rect 8300 27829 8309 27863
rect 8309 27829 8343 27863
rect 8343 27829 8352 27863
rect 8300 27820 8352 27829
rect 9128 27820 9180 27872
rect 9680 27863 9732 27872
rect 9680 27829 9689 27863
rect 9689 27829 9723 27863
rect 9723 27829 9732 27863
rect 9680 27820 9732 27829
rect 11796 27999 11848 28008
rect 11796 27965 11805 27999
rect 11805 27965 11839 27999
rect 11839 27965 11848 27999
rect 11796 27956 11848 27965
rect 10324 27820 10376 27872
rect 11244 27820 11296 27872
rect 14740 28024 14792 28076
rect 15936 28024 15988 28076
rect 17040 28092 17092 28144
rect 18696 28092 18748 28144
rect 18788 28092 18840 28144
rect 19616 28092 19668 28144
rect 16856 28024 16908 28076
rect 20260 28024 20312 28076
rect 22100 28067 22152 28076
rect 22100 28033 22109 28067
rect 22109 28033 22143 28067
rect 22143 28033 22152 28067
rect 22100 28024 22152 28033
rect 14832 27999 14884 28008
rect 14832 27965 14841 27999
rect 14841 27965 14875 27999
rect 14875 27965 14884 27999
rect 14832 27956 14884 27965
rect 17868 27888 17920 27940
rect 19432 27956 19484 28008
rect 22560 28024 22612 28076
rect 23848 28067 23900 28076
rect 23848 28033 23857 28067
rect 23857 28033 23891 28067
rect 23891 28033 23900 28067
rect 23848 28024 23900 28033
rect 19340 27820 19392 27872
rect 19800 27820 19852 27872
rect 23664 27863 23716 27872
rect 23664 27829 23673 27863
rect 23673 27829 23707 27863
rect 23707 27829 23716 27863
rect 23664 27820 23716 27829
rect 24400 27863 24452 27872
rect 24400 27829 24409 27863
rect 24409 27829 24443 27863
rect 24443 27829 24452 27863
rect 24400 27820 24452 27829
rect 3917 27718 3969 27770
rect 3981 27718 4033 27770
rect 4045 27718 4097 27770
rect 4109 27718 4161 27770
rect 4173 27718 4225 27770
rect 9851 27718 9903 27770
rect 9915 27718 9967 27770
rect 9979 27718 10031 27770
rect 10043 27718 10095 27770
rect 10107 27718 10159 27770
rect 15785 27718 15837 27770
rect 15849 27718 15901 27770
rect 15913 27718 15965 27770
rect 15977 27718 16029 27770
rect 16041 27718 16093 27770
rect 21719 27718 21771 27770
rect 21783 27718 21835 27770
rect 21847 27718 21899 27770
rect 21911 27718 21963 27770
rect 21975 27718 22027 27770
rect 1860 27616 1912 27668
rect 3608 27616 3660 27668
rect 3700 27616 3752 27668
rect 2872 27548 2924 27600
rect 4620 27548 4672 27600
rect 4160 27480 4212 27532
rect 4344 27480 4396 27532
rect 5540 27616 5592 27668
rect 6092 27616 6144 27668
rect 11244 27659 11296 27668
rect 11244 27625 11253 27659
rect 11253 27625 11287 27659
rect 11287 27625 11296 27659
rect 11244 27616 11296 27625
rect 11796 27616 11848 27668
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 2228 27412 2280 27464
rect 2964 27412 3016 27464
rect 1584 27344 1636 27396
rect 3792 27455 3844 27464
rect 3792 27421 3801 27455
rect 3801 27421 3835 27455
rect 3835 27421 3844 27455
rect 3792 27412 3844 27421
rect 4804 27412 4856 27464
rect 5908 27480 5960 27532
rect 13544 27548 13596 27600
rect 17684 27616 17736 27668
rect 22100 27616 22152 27668
rect 7840 27480 7892 27532
rect 8208 27480 8260 27532
rect 9680 27480 9732 27532
rect 10968 27480 11020 27532
rect 5448 27412 5500 27464
rect 6460 27455 6512 27464
rect 6460 27421 6469 27455
rect 6469 27421 6503 27455
rect 6503 27421 6512 27455
rect 6460 27412 6512 27421
rect 7288 27412 7340 27464
rect 7564 27412 7616 27464
rect 8024 27412 8076 27464
rect 2412 27319 2464 27328
rect 2412 27285 2421 27319
rect 2421 27285 2455 27319
rect 2455 27285 2464 27319
rect 2412 27276 2464 27285
rect 2596 27276 2648 27328
rect 5448 27276 5500 27328
rect 6920 27387 6972 27396
rect 6920 27353 6929 27387
rect 6929 27353 6963 27387
rect 6963 27353 6972 27387
rect 6920 27344 6972 27353
rect 9588 27387 9640 27396
rect 9588 27353 9597 27387
rect 9597 27353 9631 27387
rect 9631 27353 9640 27387
rect 9588 27344 9640 27353
rect 9680 27387 9732 27396
rect 9680 27353 9689 27387
rect 9689 27353 9723 27387
rect 9723 27353 9732 27387
rect 9680 27344 9732 27353
rect 10048 27387 10100 27396
rect 10048 27353 10057 27387
rect 10057 27353 10091 27387
rect 10091 27353 10100 27387
rect 10048 27344 10100 27353
rect 11152 27455 11204 27464
rect 11152 27421 11161 27455
rect 11161 27421 11195 27455
rect 11195 27421 11204 27455
rect 11152 27412 11204 27421
rect 11520 27412 11572 27464
rect 11612 27455 11664 27464
rect 11612 27421 11621 27455
rect 11621 27421 11655 27455
rect 11655 27421 11664 27455
rect 11612 27412 11664 27421
rect 11888 27523 11940 27532
rect 11888 27489 11897 27523
rect 11897 27489 11931 27523
rect 11931 27489 11940 27523
rect 11888 27480 11940 27489
rect 13176 27480 13228 27532
rect 17316 27548 17368 27600
rect 18236 27548 18288 27600
rect 17040 27480 17092 27532
rect 17408 27480 17460 27532
rect 17592 27480 17644 27532
rect 18696 27480 18748 27532
rect 12532 27412 12584 27464
rect 14188 27455 14240 27464
rect 14188 27421 14197 27455
rect 14197 27421 14231 27455
rect 14231 27421 14240 27455
rect 14188 27412 14240 27421
rect 14372 27412 14424 27464
rect 14832 27412 14884 27464
rect 14556 27344 14608 27396
rect 19800 27455 19852 27464
rect 19800 27421 19809 27455
rect 19809 27421 19843 27455
rect 19843 27421 19852 27455
rect 19800 27412 19852 27421
rect 20076 27523 20128 27532
rect 20076 27489 20085 27523
rect 20085 27489 20119 27523
rect 20119 27489 20128 27523
rect 20076 27480 20128 27489
rect 23848 27616 23900 27668
rect 7380 27276 7432 27328
rect 7472 27319 7524 27328
rect 7472 27285 7481 27319
rect 7481 27285 7515 27319
rect 7515 27285 7524 27319
rect 7472 27276 7524 27285
rect 7840 27276 7892 27328
rect 8392 27276 8444 27328
rect 10324 27276 10376 27328
rect 10416 27319 10468 27328
rect 10416 27285 10425 27319
rect 10425 27285 10459 27319
rect 10459 27285 10468 27319
rect 10416 27276 10468 27285
rect 11888 27276 11940 27328
rect 12348 27276 12400 27328
rect 12716 27276 12768 27328
rect 14740 27276 14792 27328
rect 20904 27344 20956 27396
rect 22744 27412 22796 27464
rect 23664 27412 23716 27464
rect 23756 27412 23808 27464
rect 21916 27276 21968 27328
rect 25136 27344 25188 27396
rect 22836 27319 22888 27328
rect 22836 27285 22845 27319
rect 22845 27285 22879 27319
rect 22879 27285 22888 27319
rect 22836 27276 22888 27285
rect 23572 27319 23624 27328
rect 23572 27285 23581 27319
rect 23581 27285 23615 27319
rect 23615 27285 23624 27319
rect 23572 27276 23624 27285
rect 6884 27174 6936 27226
rect 6948 27174 7000 27226
rect 7012 27174 7064 27226
rect 7076 27174 7128 27226
rect 7140 27174 7192 27226
rect 12818 27174 12870 27226
rect 12882 27174 12934 27226
rect 12946 27174 12998 27226
rect 13010 27174 13062 27226
rect 13074 27174 13126 27226
rect 18752 27174 18804 27226
rect 18816 27174 18868 27226
rect 18880 27174 18932 27226
rect 18944 27174 18996 27226
rect 19008 27174 19060 27226
rect 24686 27174 24738 27226
rect 24750 27174 24802 27226
rect 24814 27174 24866 27226
rect 24878 27174 24930 27226
rect 24942 27174 24994 27226
rect 2136 27072 2188 27124
rect 3056 27115 3108 27124
rect 3056 27081 3065 27115
rect 3065 27081 3099 27115
rect 3099 27081 3108 27115
rect 3056 27072 3108 27081
rect 1308 27004 1360 27056
rect 480 26936 532 26988
rect 2044 26979 2096 26988
rect 2044 26945 2053 26979
rect 2053 26945 2087 26979
rect 2087 26945 2096 26979
rect 2044 26936 2096 26945
rect 2136 26979 2188 26988
rect 2136 26945 2145 26979
rect 2145 26945 2179 26979
rect 2179 26945 2188 26979
rect 2136 26936 2188 26945
rect 2504 26979 2556 26988
rect 2504 26945 2513 26979
rect 2513 26945 2547 26979
rect 2547 26945 2556 26979
rect 2504 26936 2556 26945
rect 296 26868 348 26920
rect 2412 26868 2464 26920
rect 20 26596 72 26648
rect 848 26596 900 26648
rect 1584 26732 1636 26784
rect 4344 27004 4396 27056
rect 4528 27004 4580 27056
rect 4804 27004 4856 27056
rect 6276 27004 6328 27056
rect 7564 27004 7616 27056
rect 7840 27004 7892 27056
rect 8300 27004 8352 27056
rect 9680 27072 9732 27124
rect 11152 27072 11204 27124
rect 11612 27115 11664 27124
rect 11612 27081 11621 27115
rect 11621 27081 11655 27115
rect 11655 27081 11664 27115
rect 11612 27072 11664 27081
rect 4160 26936 4212 26988
rect 4620 26936 4672 26988
rect 8852 26979 8904 26988
rect 8852 26945 8875 26979
rect 8875 26945 8904 26979
rect 11060 27004 11112 27056
rect 12440 27072 12492 27124
rect 18236 27072 18288 27124
rect 8852 26936 8904 26945
rect 9036 26936 9088 26988
rect 9220 26936 9272 26988
rect 10140 26936 10192 26988
rect 11612 26936 11664 26988
rect 8300 26868 8352 26920
rect 9128 26868 9180 26920
rect 10416 26868 10468 26920
rect 20904 27004 20956 27056
rect 21916 27072 21968 27124
rect 12072 26979 12124 26988
rect 12072 26945 12081 26979
rect 12081 26945 12115 26979
rect 12115 26945 12124 26979
rect 12072 26936 12124 26945
rect 12348 26936 12400 26988
rect 13636 26936 13688 26988
rect 13728 26979 13780 26988
rect 13728 26945 13737 26979
rect 13737 26945 13771 26979
rect 13771 26945 13780 26979
rect 13728 26936 13780 26945
rect 14556 26979 14608 26988
rect 14556 26945 14590 26979
rect 14590 26945 14608 26979
rect 14556 26936 14608 26945
rect 14740 26979 14792 26988
rect 14740 26945 14749 26979
rect 14749 26945 14783 26979
rect 14783 26945 14792 26979
rect 14740 26936 14792 26945
rect 17408 26936 17460 26988
rect 19984 26936 20036 26988
rect 21364 26936 21416 26988
rect 22192 26936 22244 26988
rect 22744 27004 22796 27056
rect 12164 26911 12216 26920
rect 12164 26877 12173 26911
rect 12173 26877 12207 26911
rect 12207 26877 12216 26911
rect 12164 26868 12216 26877
rect 13544 26911 13596 26920
rect 4804 26775 4856 26784
rect 4804 26741 4813 26775
rect 4813 26741 4847 26775
rect 4847 26741 4856 26775
rect 4804 26732 4856 26741
rect 11060 26732 11112 26784
rect 12256 26732 12308 26784
rect 12440 26732 12492 26784
rect 13544 26877 13553 26911
rect 13553 26877 13587 26911
rect 13587 26877 13596 26911
rect 13544 26868 13596 26877
rect 13912 26868 13964 26920
rect 13176 26775 13228 26784
rect 13176 26741 13185 26775
rect 13185 26741 13219 26775
rect 13219 26741 13228 26775
rect 13176 26732 13228 26741
rect 14188 26732 14240 26784
rect 20076 26868 20128 26920
rect 20628 26868 20680 26920
rect 14464 26732 14516 26784
rect 14740 26732 14792 26784
rect 19248 26800 19300 26852
rect 16672 26732 16724 26784
rect 17408 26732 17460 26784
rect 17684 26775 17736 26784
rect 17684 26741 17693 26775
rect 17693 26741 17727 26775
rect 17727 26741 17736 26775
rect 17684 26732 17736 26741
rect 22192 26775 22244 26784
rect 22192 26741 22201 26775
rect 22201 26741 22235 26775
rect 22235 26741 22244 26775
rect 22192 26732 22244 26741
rect 23020 26732 23072 26784
rect 23756 26775 23808 26784
rect 23756 26741 23765 26775
rect 23765 26741 23799 26775
rect 23799 26741 23808 26775
rect 23756 26732 23808 26741
rect 24216 26775 24268 26784
rect 24216 26741 24225 26775
rect 24225 26741 24259 26775
rect 24259 26741 24268 26775
rect 24216 26732 24268 26741
rect 3917 26630 3969 26682
rect 3981 26630 4033 26682
rect 4045 26630 4097 26682
rect 4109 26630 4161 26682
rect 4173 26630 4225 26682
rect 9851 26630 9903 26682
rect 9915 26630 9967 26682
rect 9979 26630 10031 26682
rect 10043 26630 10095 26682
rect 10107 26630 10159 26682
rect 15785 26630 15837 26682
rect 15849 26630 15901 26682
rect 15913 26630 15965 26682
rect 15977 26630 16029 26682
rect 16041 26630 16093 26682
rect 21719 26630 21771 26682
rect 21783 26630 21835 26682
rect 21847 26630 21899 26682
rect 21911 26630 21963 26682
rect 21975 26630 22027 26682
rect 1400 26528 1452 26580
rect 112 26460 164 26512
rect 2136 26528 2188 26580
rect 2872 26528 2924 26580
rect 1584 26503 1636 26512
rect 1584 26469 1593 26503
rect 1593 26469 1627 26503
rect 1627 26469 1636 26503
rect 1584 26460 1636 26469
rect 5448 26528 5500 26580
rect 6460 26460 6512 26512
rect 7196 26460 7248 26512
rect 8300 26571 8352 26580
rect 8300 26537 8309 26571
rect 8309 26537 8343 26571
rect 8343 26537 8352 26571
rect 8300 26528 8352 26537
rect 13084 26528 13136 26580
rect 13176 26528 13228 26580
rect 14004 26528 14056 26580
rect 15292 26528 15344 26580
rect 15476 26528 15528 26580
rect 15844 26528 15896 26580
rect 17684 26528 17736 26580
rect 8668 26460 8720 26512
rect 9220 26460 9272 26512
rect 11520 26460 11572 26512
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 2780 26392 2832 26444
rect 3332 26392 3384 26444
rect 4988 26392 5040 26444
rect 5448 26392 5500 26444
rect 6644 26392 6696 26444
rect 12256 26392 12308 26444
rect 13544 26392 13596 26444
rect 14372 26392 14424 26444
rect 1676 26324 1728 26376
rect 4344 26256 4396 26308
rect 8024 26324 8076 26376
rect 8576 26324 8628 26376
rect 7196 26256 7248 26308
rect 7748 26256 7800 26308
rect 7840 26256 7892 26308
rect 9128 26256 9180 26308
rect 11888 26324 11940 26376
rect 12164 26324 12216 26376
rect 14464 26324 14516 26376
rect 15292 26435 15344 26444
rect 15292 26401 15301 26435
rect 15301 26401 15335 26435
rect 15335 26401 15344 26435
rect 15292 26392 15344 26401
rect 15476 26392 15528 26444
rect 16580 26460 16632 26512
rect 16120 26392 16172 26444
rect 16304 26392 16356 26444
rect 16672 26435 16724 26444
rect 16672 26401 16681 26435
rect 16681 26401 16715 26435
rect 16715 26401 16724 26435
rect 16672 26392 16724 26401
rect 16764 26392 16816 26444
rect 21364 26571 21416 26580
rect 21364 26537 21373 26571
rect 21373 26537 21407 26571
rect 21407 26537 21416 26571
rect 21364 26528 21416 26537
rect 15108 26367 15160 26376
rect 15108 26333 15142 26367
rect 15142 26333 15160 26367
rect 15108 26324 15160 26333
rect 17040 26367 17092 26376
rect 17040 26333 17074 26367
rect 17074 26333 17092 26367
rect 17040 26324 17092 26333
rect 17868 26367 17920 26376
rect 17868 26333 17877 26367
rect 17877 26333 17911 26367
rect 17911 26333 17920 26367
rect 21088 26392 21140 26444
rect 22284 26528 22336 26580
rect 22468 26392 22520 26444
rect 17868 26324 17920 26333
rect 20076 26324 20128 26376
rect 1676 26188 1728 26240
rect 4528 26188 4580 26240
rect 5356 26188 5408 26240
rect 6276 26188 6328 26240
rect 12440 26188 12492 26240
rect 12532 26231 12584 26240
rect 12532 26197 12541 26231
rect 12541 26197 12575 26231
rect 12575 26197 12584 26231
rect 12532 26188 12584 26197
rect 20260 26299 20312 26308
rect 15108 26188 15160 26240
rect 20260 26265 20272 26299
rect 20272 26265 20312 26299
rect 20260 26256 20312 26265
rect 21364 26256 21416 26308
rect 23112 26367 23164 26376
rect 23112 26333 23119 26367
rect 23119 26333 23153 26367
rect 23153 26333 23164 26367
rect 23112 26324 23164 26333
rect 18512 26231 18564 26240
rect 18512 26197 18521 26231
rect 18521 26197 18555 26231
rect 18555 26197 18564 26231
rect 18512 26188 18564 26197
rect 23848 26231 23900 26240
rect 23848 26197 23857 26231
rect 23857 26197 23891 26231
rect 23891 26197 23900 26231
rect 23848 26188 23900 26197
rect 6884 26086 6936 26138
rect 6948 26086 7000 26138
rect 7012 26086 7064 26138
rect 7076 26086 7128 26138
rect 7140 26086 7192 26138
rect 12818 26086 12870 26138
rect 12882 26086 12934 26138
rect 12946 26086 12998 26138
rect 13010 26086 13062 26138
rect 13074 26086 13126 26138
rect 18752 26086 18804 26138
rect 18816 26086 18868 26138
rect 18880 26086 18932 26138
rect 18944 26086 18996 26138
rect 19008 26086 19060 26138
rect 24686 26086 24738 26138
rect 24750 26086 24802 26138
rect 24814 26086 24866 26138
rect 24878 26086 24930 26138
rect 24942 26086 24994 26138
rect 940 25984 992 26036
rect 848 25916 900 25968
rect 1492 25848 1544 25900
rect 2136 26027 2188 26036
rect 2136 25993 2145 26027
rect 2145 25993 2179 26027
rect 2179 25993 2188 26027
rect 2136 25984 2188 25993
rect 2688 26027 2740 26036
rect 2688 25993 2697 26027
rect 2697 25993 2731 26027
rect 2731 25993 2740 26027
rect 2688 25984 2740 25993
rect 4068 25916 4120 25968
rect 4252 25916 4304 25968
rect 4528 25959 4580 25968
rect 4528 25925 4537 25959
rect 4537 25925 4571 25959
rect 4571 25925 4580 25959
rect 4528 25916 4580 25925
rect 6552 25984 6604 26036
rect 7656 25984 7708 26036
rect 8116 25984 8168 26036
rect 9496 25984 9548 26036
rect 9772 25984 9824 26036
rect 10692 25984 10744 26036
rect 11520 25984 11572 26036
rect 14832 25984 14884 26036
rect 16672 25984 16724 26036
rect 2228 25891 2280 25900
rect 2228 25857 2237 25891
rect 2237 25857 2271 25891
rect 2271 25857 2280 25891
rect 2228 25848 2280 25857
rect 2504 25891 2556 25900
rect 2504 25857 2513 25891
rect 2513 25857 2547 25891
rect 2547 25857 2556 25891
rect 2504 25848 2556 25857
rect 3792 25848 3844 25900
rect 5080 25848 5132 25900
rect 15200 25916 15252 25968
rect 15384 25916 15436 25968
rect 17868 25959 17920 25968
rect 17868 25925 17902 25959
rect 17902 25925 17920 25959
rect 17868 25916 17920 25925
rect 18512 25916 18564 25968
rect 4804 25780 4856 25832
rect 5448 25848 5500 25900
rect 5632 25780 5684 25832
rect 2412 25755 2464 25764
rect 2412 25721 2421 25755
rect 2421 25721 2455 25755
rect 2455 25721 2464 25755
rect 2412 25712 2464 25721
rect 1584 25687 1636 25696
rect 1584 25653 1593 25687
rect 1593 25653 1627 25687
rect 1627 25653 1636 25687
rect 1584 25644 1636 25653
rect 2228 25644 2280 25696
rect 2320 25644 2372 25696
rect 2872 25644 2924 25696
rect 6092 25644 6144 25696
rect 7840 25644 7892 25696
rect 8024 25644 8076 25696
rect 9220 25780 9272 25832
rect 10140 25848 10192 25900
rect 11980 25848 12032 25900
rect 20260 25984 20312 26036
rect 22836 25984 22888 26036
rect 23848 25984 23900 26036
rect 14740 25780 14792 25832
rect 10876 25644 10928 25696
rect 11888 25644 11940 25696
rect 13268 25644 13320 25696
rect 15660 25644 15712 25696
rect 22284 25848 22336 25900
rect 23388 25891 23440 25900
rect 23388 25857 23397 25891
rect 23397 25857 23431 25891
rect 23431 25857 23440 25891
rect 23388 25848 23440 25857
rect 23940 25916 23992 25968
rect 22192 25780 22244 25832
rect 25136 25780 25188 25832
rect 25320 25780 25372 25832
rect 17960 25644 18012 25696
rect 18512 25644 18564 25696
rect 18604 25644 18656 25696
rect 19248 25687 19300 25696
rect 19248 25653 19257 25687
rect 19257 25653 19291 25687
rect 19291 25653 19300 25687
rect 19248 25644 19300 25653
rect 22560 25644 22612 25696
rect 23848 25687 23900 25696
rect 23848 25653 23857 25687
rect 23857 25653 23891 25687
rect 23891 25653 23900 25687
rect 23848 25644 23900 25653
rect 24400 25687 24452 25696
rect 24400 25653 24409 25687
rect 24409 25653 24443 25687
rect 24443 25653 24452 25687
rect 24400 25644 24452 25653
rect 3917 25542 3969 25594
rect 3981 25542 4033 25594
rect 4045 25542 4097 25594
rect 4109 25542 4161 25594
rect 4173 25542 4225 25594
rect 9851 25542 9903 25594
rect 9915 25542 9967 25594
rect 9979 25542 10031 25594
rect 10043 25542 10095 25594
rect 10107 25542 10159 25594
rect 15785 25542 15837 25594
rect 15849 25542 15901 25594
rect 15913 25542 15965 25594
rect 15977 25542 16029 25594
rect 16041 25542 16093 25594
rect 21719 25542 21771 25594
rect 21783 25542 21835 25594
rect 21847 25542 21899 25594
rect 21911 25542 21963 25594
rect 21975 25542 22027 25594
rect 1584 25440 1636 25492
rect 6276 25440 6328 25492
rect 7472 25440 7524 25492
rect 2136 25415 2188 25424
rect 2136 25381 2145 25415
rect 2145 25381 2179 25415
rect 2179 25381 2188 25415
rect 2136 25372 2188 25381
rect 2320 25372 2372 25424
rect 940 25100 992 25152
rect 1676 25279 1728 25288
rect 1676 25245 1685 25279
rect 1685 25245 1719 25279
rect 1719 25245 1728 25279
rect 1676 25236 1728 25245
rect 1952 25279 2004 25288
rect 1952 25245 1961 25279
rect 1961 25245 1995 25279
rect 1995 25245 2004 25279
rect 1952 25236 2004 25245
rect 3240 25304 3292 25356
rect 3608 25304 3660 25356
rect 4344 25304 4396 25356
rect 10048 25304 10100 25356
rect 10416 25304 10468 25356
rect 10692 25347 10744 25356
rect 10692 25313 10726 25347
rect 10726 25313 10744 25347
rect 10692 25304 10744 25313
rect 10876 25347 10928 25356
rect 10876 25313 10885 25347
rect 10885 25313 10919 25347
rect 10919 25313 10928 25347
rect 10876 25304 10928 25313
rect 12072 25440 12124 25492
rect 15200 25440 15252 25492
rect 12532 25415 12584 25424
rect 12532 25381 12541 25415
rect 12541 25381 12575 25415
rect 12575 25381 12584 25415
rect 12532 25372 12584 25381
rect 18604 25483 18656 25492
rect 18604 25449 18613 25483
rect 18613 25449 18647 25483
rect 18647 25449 18656 25483
rect 18604 25440 18656 25449
rect 19248 25440 19300 25492
rect 11612 25304 11664 25356
rect 13728 25304 13780 25356
rect 14464 25304 14516 25356
rect 14648 25304 14700 25356
rect 19892 25372 19944 25424
rect 20168 25372 20220 25424
rect 21088 25372 21140 25424
rect 23388 25440 23440 25492
rect 25872 25440 25924 25492
rect 15108 25347 15160 25356
rect 15108 25313 15142 25347
rect 15142 25313 15160 25347
rect 15108 25304 15160 25313
rect 15292 25347 15344 25356
rect 15292 25313 15301 25347
rect 15301 25313 15335 25347
rect 15335 25313 15344 25347
rect 15292 25304 15344 25313
rect 16304 25304 16356 25356
rect 16580 25304 16632 25356
rect 23480 25304 23532 25356
rect 23940 25304 23992 25356
rect 2688 25236 2740 25288
rect 3056 25236 3108 25288
rect 5632 25236 5684 25288
rect 1584 25143 1636 25152
rect 1584 25109 1593 25143
rect 1593 25109 1627 25143
rect 1627 25109 1636 25143
rect 1584 25100 1636 25109
rect 5172 25168 5224 25220
rect 6092 25168 6144 25220
rect 3332 25143 3384 25152
rect 3332 25109 3341 25143
rect 3341 25109 3375 25143
rect 3375 25109 3384 25143
rect 3332 25100 3384 25109
rect 4896 25100 4948 25152
rect 6276 25143 6328 25152
rect 6276 25109 6285 25143
rect 6285 25109 6319 25143
rect 6319 25109 6328 25143
rect 6276 25100 6328 25109
rect 6460 25100 6512 25152
rect 7196 25168 7248 25220
rect 7380 25211 7432 25220
rect 7380 25177 7389 25211
rect 7389 25177 7423 25211
rect 7423 25177 7432 25211
rect 7380 25168 7432 25177
rect 7288 25100 7340 25152
rect 7564 25143 7616 25152
rect 7564 25109 7573 25143
rect 7573 25109 7607 25143
rect 7607 25109 7616 25143
rect 7564 25100 7616 25109
rect 10600 25279 10652 25288
rect 10600 25245 10609 25279
rect 10609 25245 10643 25279
rect 10643 25245 10652 25279
rect 10600 25236 10652 25245
rect 11980 25100 12032 25152
rect 12256 25236 12308 25288
rect 12900 25279 12952 25288
rect 12900 25245 12934 25279
rect 12934 25245 12952 25279
rect 12900 25236 12952 25245
rect 13084 25279 13136 25288
rect 13084 25245 13093 25279
rect 13093 25245 13127 25279
rect 13127 25245 13136 25279
rect 13084 25236 13136 25245
rect 17500 25236 17552 25288
rect 12440 25100 12492 25152
rect 12624 25100 12676 25152
rect 12900 25100 12952 25152
rect 17960 25168 18012 25220
rect 15936 25143 15988 25152
rect 15936 25109 15945 25143
rect 15945 25109 15979 25143
rect 15979 25109 15988 25143
rect 15936 25100 15988 25109
rect 16580 25100 16632 25152
rect 19984 25236 20036 25288
rect 20444 25236 20496 25288
rect 23756 25236 23808 25288
rect 21180 25168 21232 25220
rect 20352 25100 20404 25152
rect 24124 25143 24176 25152
rect 24124 25109 24133 25143
rect 24133 25109 24167 25143
rect 24167 25109 24176 25143
rect 24124 25100 24176 25109
rect 296 24964 348 25016
rect 664 24964 716 25016
rect 6884 24998 6936 25050
rect 6948 24998 7000 25050
rect 7012 24998 7064 25050
rect 7076 24998 7128 25050
rect 7140 24998 7192 25050
rect 12818 24998 12870 25050
rect 12882 24998 12934 25050
rect 12946 24998 12998 25050
rect 13010 24998 13062 25050
rect 13074 24998 13126 25050
rect 18752 24998 18804 25050
rect 18816 24998 18868 25050
rect 18880 24998 18932 25050
rect 18944 24998 18996 25050
rect 19008 24998 19060 25050
rect 24686 24998 24738 25050
rect 24750 24998 24802 25050
rect 24814 24998 24866 25050
rect 24878 24998 24930 25050
rect 24942 24998 24994 25050
rect 1584 24896 1636 24948
rect 1860 24896 1912 24948
rect 2228 24896 2280 24948
rect 3792 24896 3844 24948
rect 7288 24896 7340 24948
rect 112 24828 164 24880
rect 3056 24828 3108 24880
rect 3424 24871 3476 24880
rect 3424 24837 3433 24871
rect 3433 24837 3467 24871
rect 3467 24837 3476 24871
rect 3424 24828 3476 24837
rect 1400 24803 1452 24812
rect 1400 24769 1409 24803
rect 1409 24769 1443 24803
rect 1443 24769 1452 24803
rect 1400 24760 1452 24769
rect 2228 24760 2280 24812
rect 3700 24803 3752 24812
rect 3700 24769 3709 24803
rect 3709 24769 3743 24803
rect 3743 24769 3752 24803
rect 3700 24760 3752 24769
rect 3792 24803 3844 24812
rect 3792 24769 3801 24803
rect 3801 24769 3835 24803
rect 3835 24769 3844 24803
rect 3792 24760 3844 24769
rect 4252 24828 4304 24880
rect 4344 24828 4396 24880
rect 5448 24760 5500 24812
rect 3332 24692 3384 24744
rect 5908 24760 5960 24812
rect 10508 24896 10560 24948
rect 10600 24896 10652 24948
rect 12256 24896 12308 24948
rect 13176 24939 13228 24948
rect 13176 24905 13185 24939
rect 13185 24905 13219 24939
rect 13219 24905 13228 24939
rect 13176 24896 13228 24905
rect 15936 24896 15988 24948
rect 19984 24896 20036 24948
rect 8208 24760 8260 24812
rect 8392 24803 8444 24812
rect 8392 24769 8401 24803
rect 8401 24769 8435 24803
rect 8435 24769 8444 24803
rect 8392 24760 8444 24769
rect 8944 24760 8996 24812
rect 1308 24556 1360 24608
rect 4712 24667 4764 24676
rect 4712 24633 4721 24667
rect 4721 24633 4755 24667
rect 4755 24633 4764 24667
rect 4712 24624 4764 24633
rect 5356 24624 5408 24676
rect 6092 24624 6144 24676
rect 2412 24599 2464 24608
rect 2412 24565 2421 24599
rect 2421 24565 2455 24599
rect 2455 24565 2464 24599
rect 2412 24556 2464 24565
rect 8024 24692 8076 24744
rect 9128 24692 9180 24744
rect 9496 24735 9548 24744
rect 9496 24701 9505 24735
rect 9505 24701 9539 24735
rect 9539 24701 9548 24735
rect 9496 24692 9548 24701
rect 9680 24735 9732 24744
rect 9680 24701 9689 24735
rect 9689 24701 9723 24735
rect 9723 24701 9732 24735
rect 9680 24692 9732 24701
rect 10508 24803 10560 24812
rect 10508 24769 10542 24803
rect 10542 24769 10560 24803
rect 10508 24760 10560 24769
rect 10048 24692 10100 24744
rect 10416 24735 10468 24744
rect 10416 24701 10425 24735
rect 10425 24701 10459 24735
rect 10459 24701 10468 24735
rect 10416 24692 10468 24701
rect 11520 24760 11572 24812
rect 13268 24760 13320 24812
rect 14832 24760 14884 24812
rect 15476 24760 15528 24812
rect 17960 24828 18012 24880
rect 19248 24828 19300 24880
rect 20260 24896 20312 24948
rect 18788 24803 18840 24812
rect 18788 24769 18811 24803
rect 18811 24769 18840 24803
rect 10876 24692 10928 24744
rect 12164 24735 12216 24744
rect 12164 24701 12173 24735
rect 12173 24701 12207 24735
rect 12207 24701 12216 24735
rect 12164 24692 12216 24701
rect 16120 24692 16172 24744
rect 18788 24760 18840 24769
rect 18512 24735 18564 24744
rect 18512 24701 18521 24735
rect 18521 24701 18555 24735
rect 18555 24701 18564 24735
rect 18512 24692 18564 24701
rect 14556 24624 14608 24676
rect 14924 24624 14976 24676
rect 16856 24624 16908 24676
rect 17500 24624 17552 24676
rect 20168 24760 20220 24812
rect 20260 24803 20312 24812
rect 20260 24769 20267 24803
rect 20267 24769 20301 24803
rect 20301 24769 20312 24803
rect 20260 24760 20312 24769
rect 20996 24760 21048 24812
rect 21640 24760 21692 24812
rect 23204 24803 23256 24812
rect 23204 24769 23213 24803
rect 23213 24769 23247 24803
rect 23247 24769 23256 24803
rect 23204 24760 23256 24769
rect 23388 24760 23440 24812
rect 23480 24760 23532 24812
rect 6736 24556 6788 24608
rect 10692 24556 10744 24608
rect 10876 24556 10928 24608
rect 12992 24556 13044 24608
rect 14188 24556 14240 24608
rect 15108 24556 15160 24608
rect 16212 24599 16264 24608
rect 16212 24565 16221 24599
rect 16221 24565 16255 24599
rect 16255 24565 16264 24599
rect 16212 24556 16264 24565
rect 17776 24556 17828 24608
rect 22284 24624 22336 24676
rect 19984 24556 20036 24608
rect 20444 24556 20496 24608
rect 22376 24556 22428 24608
rect 22928 24556 22980 24608
rect 23572 24556 23624 24608
rect 23664 24599 23716 24608
rect 23664 24565 23673 24599
rect 23673 24565 23707 24599
rect 23707 24565 23716 24599
rect 23664 24556 23716 24565
rect 24400 24599 24452 24608
rect 24400 24565 24409 24599
rect 24409 24565 24443 24599
rect 24443 24565 24452 24599
rect 24400 24556 24452 24565
rect 388 24488 440 24540
rect 3917 24454 3969 24506
rect 3981 24454 4033 24506
rect 4045 24454 4097 24506
rect 4109 24454 4161 24506
rect 4173 24454 4225 24506
rect 9851 24454 9903 24506
rect 9915 24454 9967 24506
rect 9979 24454 10031 24506
rect 10043 24454 10095 24506
rect 10107 24454 10159 24506
rect 15785 24454 15837 24506
rect 15849 24454 15901 24506
rect 15913 24454 15965 24506
rect 15977 24454 16029 24506
rect 16041 24454 16093 24506
rect 21719 24454 21771 24506
rect 21783 24454 21835 24506
rect 21847 24454 21899 24506
rect 21911 24454 21963 24506
rect 21975 24454 22027 24506
rect 3056 24395 3108 24404
rect 3056 24361 3065 24395
rect 3065 24361 3099 24395
rect 3099 24361 3108 24395
rect 3056 24352 3108 24361
rect 3148 24352 3200 24404
rect 3700 24352 3752 24404
rect 3792 24352 3844 24404
rect 388 24284 440 24336
rect 2412 24216 2464 24268
rect 2872 24216 2924 24268
rect 2228 24148 2280 24200
rect 1860 24080 1912 24132
rect 2136 24123 2188 24132
rect 2136 24089 2145 24123
rect 2145 24089 2179 24123
rect 2179 24089 2188 24123
rect 2136 24080 2188 24089
rect 2964 24080 3016 24132
rect 4160 24148 4212 24200
rect 6460 24148 6512 24200
rect 8576 24352 8628 24404
rect 9496 24352 9548 24404
rect 10232 24395 10284 24404
rect 10232 24361 10241 24395
rect 10241 24361 10275 24395
rect 10275 24361 10284 24395
rect 10232 24352 10284 24361
rect 8576 24216 8628 24268
rect 9220 24259 9272 24268
rect 9220 24225 9229 24259
rect 9229 24225 9263 24259
rect 9263 24225 9272 24259
rect 9220 24216 9272 24225
rect 11612 24259 11664 24268
rect 11612 24225 11621 24259
rect 11621 24225 11655 24259
rect 11655 24225 11664 24259
rect 11612 24216 11664 24225
rect 11980 24216 12032 24268
rect 12256 24259 12308 24268
rect 12256 24225 12265 24259
rect 12265 24225 12299 24259
rect 12299 24225 12308 24259
rect 12256 24216 12308 24225
rect 16120 24352 16172 24404
rect 16212 24352 16264 24404
rect 17500 24352 17552 24404
rect 14648 24284 14700 24336
rect 12992 24216 13044 24268
rect 13176 24216 13228 24268
rect 12808 24191 12860 24200
rect 12808 24157 12817 24191
rect 12817 24157 12851 24191
rect 12851 24157 12860 24191
rect 12808 24148 12860 24157
rect 13728 24148 13780 24200
rect 14188 24148 14240 24200
rect 6920 24080 6972 24132
rect 7656 24080 7708 24132
rect 9772 24080 9824 24132
rect 11704 24080 11756 24132
rect 14372 24216 14424 24268
rect 14832 24216 14884 24268
rect 15108 24259 15160 24268
rect 15108 24225 15142 24259
rect 15142 24225 15160 24259
rect 15108 24216 15160 24225
rect 15292 24259 15344 24268
rect 15292 24225 15301 24259
rect 15301 24225 15335 24259
rect 15335 24225 15344 24259
rect 15292 24216 15344 24225
rect 16304 24148 16356 24200
rect 16856 24216 16908 24268
rect 20352 24352 20404 24404
rect 21364 24352 21416 24404
rect 21640 24352 21692 24404
rect 22928 24352 22980 24404
rect 23204 24352 23256 24404
rect 23572 24352 23624 24404
rect 25780 24352 25832 24404
rect 20168 24284 20220 24336
rect 17960 24148 18012 24200
rect 18328 24148 18380 24200
rect 18788 24148 18840 24200
rect 19892 24148 19944 24200
rect 19984 24191 20036 24200
rect 19984 24157 19993 24191
rect 19993 24157 20027 24191
rect 20027 24157 20036 24191
rect 19984 24148 20036 24157
rect 20168 24148 20220 24200
rect 22284 24191 22336 24200
rect 22284 24157 22307 24191
rect 22307 24157 22336 24191
rect 22284 24148 22336 24157
rect 23940 24191 23992 24200
rect 23940 24157 23949 24191
rect 23949 24157 23983 24191
rect 23983 24157 23992 24191
rect 23940 24148 23992 24157
rect 20628 24123 20680 24132
rect 2228 24012 2280 24064
rect 3240 24012 3292 24064
rect 9680 24012 9732 24064
rect 10600 24012 10652 24064
rect 16856 24055 16908 24064
rect 16856 24021 16865 24055
rect 16865 24021 16899 24055
rect 16899 24021 16908 24055
rect 16856 24012 16908 24021
rect 18052 24055 18104 24064
rect 18052 24021 18061 24055
rect 18061 24021 18095 24055
rect 18095 24021 18104 24055
rect 18052 24012 18104 24021
rect 20628 24089 20640 24123
rect 20640 24089 20680 24123
rect 20628 24080 20680 24089
rect 21180 24080 21232 24132
rect 23572 24055 23624 24064
rect 23572 24021 23581 24055
rect 23581 24021 23615 24055
rect 23615 24021 23624 24055
rect 23572 24012 23624 24021
rect 24124 24055 24176 24064
rect 24124 24021 24133 24055
rect 24133 24021 24167 24055
rect 24167 24021 24176 24055
rect 24124 24012 24176 24021
rect 6884 23910 6936 23962
rect 6948 23910 7000 23962
rect 7012 23910 7064 23962
rect 7076 23910 7128 23962
rect 7140 23910 7192 23962
rect 12818 23910 12870 23962
rect 12882 23910 12934 23962
rect 12946 23910 12998 23962
rect 13010 23910 13062 23962
rect 13074 23910 13126 23962
rect 18752 23910 18804 23962
rect 18816 23910 18868 23962
rect 18880 23910 18932 23962
rect 18944 23910 18996 23962
rect 19008 23910 19060 23962
rect 24686 23910 24738 23962
rect 24750 23910 24802 23962
rect 24814 23910 24866 23962
rect 24878 23910 24930 23962
rect 24942 23910 24994 23962
rect 2136 23808 2188 23860
rect 3424 23808 3476 23860
rect 3516 23808 3568 23860
rect 1308 23740 1360 23792
rect 1492 23715 1544 23724
rect 1492 23681 1501 23715
rect 1501 23681 1535 23715
rect 1535 23681 1544 23715
rect 1492 23672 1544 23681
rect 1676 23672 1728 23724
rect 2596 23672 2648 23724
rect 3424 23715 3476 23724
rect 3424 23681 3433 23715
rect 3433 23681 3467 23715
rect 3467 23681 3476 23715
rect 3424 23672 3476 23681
rect 1400 23604 1452 23656
rect 4988 23808 5040 23860
rect 5080 23808 5132 23860
rect 5356 23808 5408 23860
rect 8392 23808 8444 23860
rect 12256 23808 12308 23860
rect 13452 23808 13504 23860
rect 14924 23808 14976 23860
rect 16580 23808 16632 23860
rect 16856 23808 16908 23860
rect 4252 23672 4304 23724
rect 4528 23715 4580 23724
rect 4528 23681 4537 23715
rect 4537 23681 4571 23715
rect 4571 23681 4580 23715
rect 4528 23672 4580 23681
rect 5264 23715 5316 23724
rect 5264 23681 5273 23715
rect 5273 23681 5307 23715
rect 5307 23681 5316 23715
rect 5264 23672 5316 23681
rect 5540 23647 5592 23656
rect 5540 23613 5549 23647
rect 5549 23613 5583 23647
rect 5583 23613 5592 23647
rect 5540 23604 5592 23613
rect 4988 23579 5040 23588
rect 4988 23545 4997 23579
rect 4997 23545 5031 23579
rect 5031 23545 5040 23579
rect 4988 23536 5040 23545
rect 8944 23740 8996 23792
rect 7840 23604 7892 23656
rect 8024 23604 8076 23656
rect 2780 23468 2832 23520
rect 6184 23511 6236 23520
rect 6184 23477 6193 23511
rect 6193 23477 6227 23511
rect 6227 23477 6236 23511
rect 6184 23468 6236 23477
rect 11244 23672 11296 23724
rect 11060 23604 11112 23656
rect 11704 23672 11756 23724
rect 12348 23672 12400 23724
rect 13636 23672 13688 23724
rect 15292 23715 15344 23724
rect 15292 23681 15301 23715
rect 15301 23681 15344 23715
rect 15292 23672 15344 23681
rect 18052 23715 18104 23724
rect 18052 23681 18061 23715
rect 18061 23681 18095 23715
rect 18095 23681 18104 23715
rect 18052 23672 18104 23681
rect 20628 23808 20680 23860
rect 18604 23715 18656 23724
rect 18604 23681 18613 23715
rect 18613 23681 18647 23715
rect 18647 23681 18656 23715
rect 18604 23672 18656 23681
rect 23480 23851 23532 23860
rect 23480 23817 23489 23851
rect 23489 23817 23523 23851
rect 23523 23817 23532 23851
rect 23480 23808 23532 23817
rect 14648 23604 14700 23656
rect 13268 23468 13320 23520
rect 13636 23468 13688 23520
rect 17500 23604 17552 23656
rect 23112 23740 23164 23792
rect 22376 23715 22428 23724
rect 22376 23681 22385 23715
rect 22385 23681 22419 23715
rect 22419 23681 22428 23715
rect 22376 23672 22428 23681
rect 22468 23715 22520 23724
rect 22468 23681 22477 23715
rect 22477 23681 22511 23715
rect 22511 23681 22520 23715
rect 22468 23672 22520 23681
rect 22836 23672 22888 23724
rect 24032 23672 24084 23724
rect 18328 23579 18380 23588
rect 18328 23545 18337 23579
rect 18337 23545 18371 23579
rect 18371 23545 18380 23579
rect 18328 23536 18380 23545
rect 19800 23536 19852 23588
rect 21640 23536 21692 23588
rect 16120 23468 16172 23520
rect 16580 23468 16632 23520
rect 18788 23468 18840 23520
rect 23940 23468 23992 23520
rect 24400 23511 24452 23520
rect 24400 23477 24409 23511
rect 24409 23477 24443 23511
rect 24443 23477 24452 23511
rect 24400 23468 24452 23477
rect 3917 23366 3969 23418
rect 3981 23366 4033 23418
rect 4045 23366 4097 23418
rect 4109 23366 4161 23418
rect 4173 23366 4225 23418
rect 9851 23366 9903 23418
rect 9915 23366 9967 23418
rect 9979 23366 10031 23418
rect 10043 23366 10095 23418
rect 10107 23366 10159 23418
rect 15785 23366 15837 23418
rect 15849 23366 15901 23418
rect 15913 23366 15965 23418
rect 15977 23366 16029 23418
rect 16041 23366 16093 23418
rect 21719 23366 21771 23418
rect 21783 23366 21835 23418
rect 21847 23366 21899 23418
rect 21911 23366 21963 23418
rect 21975 23366 22027 23418
rect 2504 23264 2556 23316
rect 1400 23171 1452 23180
rect 1400 23137 1409 23171
rect 1409 23137 1443 23171
rect 1443 23137 1452 23171
rect 1400 23128 1452 23137
rect 5540 23264 5592 23316
rect 7196 23264 7248 23316
rect 9220 23264 9272 23316
rect 8668 23196 8720 23248
rect 12072 23196 12124 23248
rect 12532 23196 12584 23248
rect 16120 23196 16172 23248
rect 18604 23264 18656 23316
rect 19340 23264 19392 23316
rect 21640 23264 21692 23316
rect 23480 23264 23532 23316
rect 23572 23264 23624 23316
rect 24032 23307 24084 23316
rect 24032 23273 24041 23307
rect 24041 23273 24075 23307
rect 24075 23273 24084 23307
rect 24032 23264 24084 23273
rect 6736 23128 6788 23180
rect 2688 23060 2740 23112
rect 1308 22992 1360 23044
rect 4344 22992 4396 23044
rect 5448 23060 5500 23112
rect 6184 23060 6236 23112
rect 7104 23103 7156 23112
rect 7104 23069 7113 23103
rect 7113 23069 7147 23103
rect 7147 23069 7156 23103
rect 7104 23060 7156 23069
rect 11704 23128 11756 23180
rect 13544 23128 13596 23180
rect 13912 23128 13964 23180
rect 7564 23060 7616 23112
rect 2412 22967 2464 22976
rect 2412 22933 2421 22967
rect 2421 22933 2455 22967
rect 2455 22933 2464 22967
rect 2412 22924 2464 22933
rect 4620 22924 4672 22976
rect 5448 22924 5500 22976
rect 6184 22924 6236 22976
rect 8300 22992 8352 23044
rect 9128 23103 9180 23112
rect 9128 23069 9137 23103
rect 9137 23069 9171 23103
rect 9171 23069 9180 23103
rect 9128 23060 9180 23069
rect 9772 23060 9824 23112
rect 10140 23060 10192 23112
rect 14832 23060 14884 23112
rect 15016 23060 15068 23112
rect 22744 23196 22796 23248
rect 7472 22924 7524 22976
rect 7564 22924 7616 22976
rect 8392 22967 8444 22976
rect 8392 22933 8401 22967
rect 8401 22933 8435 22967
rect 8435 22933 8444 22967
rect 8392 22924 8444 22933
rect 9772 22924 9824 22976
rect 10968 22967 11020 22976
rect 10968 22933 10977 22967
rect 10977 22933 11011 22967
rect 11011 22933 11020 22967
rect 10968 22924 11020 22933
rect 11336 22992 11388 23044
rect 12440 22992 12492 23044
rect 15200 22992 15252 23044
rect 16304 23103 16356 23112
rect 16304 23069 16313 23103
rect 16313 23069 16347 23103
rect 16347 23069 16356 23103
rect 16304 23060 16356 23069
rect 16580 23103 16632 23112
rect 16580 23069 16589 23103
rect 16589 23069 16623 23103
rect 16623 23069 16632 23103
rect 16580 23060 16632 23069
rect 17776 23060 17828 23112
rect 18052 23060 18104 23112
rect 20444 23060 20496 23112
rect 19524 22992 19576 23044
rect 20628 22992 20680 23044
rect 22468 23128 22520 23180
rect 23664 23196 23716 23248
rect 20812 23060 20864 23112
rect 23388 23103 23440 23112
rect 23388 23069 23397 23103
rect 23397 23069 23431 23103
rect 23431 23069 23440 23103
rect 23388 23060 23440 23069
rect 22560 22992 22612 23044
rect 13360 22924 13412 22976
rect 20904 22924 20956 22976
rect 23204 22967 23256 22976
rect 23204 22933 23213 22967
rect 23213 22933 23247 22967
rect 23247 22933 23256 22967
rect 23204 22924 23256 22933
rect 23664 22967 23716 22976
rect 23664 22933 23673 22967
rect 23673 22933 23707 22967
rect 23707 22933 23716 22967
rect 23664 22924 23716 22933
rect 6884 22822 6936 22874
rect 6948 22822 7000 22874
rect 7012 22822 7064 22874
rect 7076 22822 7128 22874
rect 7140 22822 7192 22874
rect 12818 22822 12870 22874
rect 12882 22822 12934 22874
rect 12946 22822 12998 22874
rect 13010 22822 13062 22874
rect 13074 22822 13126 22874
rect 18752 22822 18804 22874
rect 18816 22822 18868 22874
rect 18880 22822 18932 22874
rect 18944 22822 18996 22874
rect 19008 22822 19060 22874
rect 24686 22822 24738 22874
rect 24750 22822 24802 22874
rect 24814 22822 24866 22874
rect 24878 22822 24930 22874
rect 24942 22822 24994 22874
rect 1216 22720 1268 22772
rect 9128 22720 9180 22772
rect 9220 22763 9272 22772
rect 9220 22729 9229 22763
rect 9229 22729 9263 22763
rect 9263 22729 9272 22763
rect 9220 22720 9272 22729
rect 1400 22627 1452 22636
rect 1400 22593 1409 22627
rect 1409 22593 1443 22627
rect 1443 22593 1452 22627
rect 1400 22584 1452 22593
rect 4252 22652 4304 22704
rect 2780 22627 2832 22636
rect 2780 22593 2789 22627
rect 2789 22593 2823 22627
rect 2823 22593 2832 22627
rect 2780 22584 2832 22593
rect 3148 22584 3200 22636
rect 4068 22584 4120 22636
rect 4436 22584 4488 22636
rect 4252 22516 4304 22568
rect 2964 22491 3016 22500
rect 2964 22457 2973 22491
rect 2973 22457 3007 22491
rect 3007 22457 3016 22491
rect 2964 22448 3016 22457
rect 5356 22627 5408 22636
rect 5356 22593 5390 22627
rect 5390 22593 5408 22627
rect 5356 22584 5408 22593
rect 4896 22516 4948 22568
rect 4988 22559 5040 22568
rect 4988 22525 4997 22559
rect 4997 22525 5031 22559
rect 5031 22525 5040 22559
rect 4988 22516 5040 22525
rect 4804 22448 4856 22500
rect 5540 22559 5592 22568
rect 5540 22525 5549 22559
rect 5549 22525 5583 22559
rect 5583 22525 5592 22559
rect 5540 22516 5592 22525
rect 2412 22423 2464 22432
rect 2412 22389 2421 22423
rect 2421 22389 2455 22423
rect 2455 22389 2464 22423
rect 2412 22380 2464 22389
rect 3976 22423 4028 22432
rect 3976 22389 3985 22423
rect 3985 22389 4019 22423
rect 4019 22389 4028 22423
rect 3976 22380 4028 22389
rect 5540 22380 5592 22432
rect 10232 22695 10284 22704
rect 10232 22661 10241 22695
rect 10241 22661 10275 22695
rect 10275 22661 10284 22695
rect 10232 22652 10284 22661
rect 10968 22652 11020 22704
rect 11152 22652 11204 22704
rect 13268 22720 13320 22772
rect 13820 22720 13872 22772
rect 16672 22720 16724 22772
rect 17040 22720 17092 22772
rect 7840 22584 7892 22636
rect 8300 22627 8352 22636
rect 8300 22593 8309 22627
rect 8309 22593 8343 22627
rect 8343 22593 8352 22627
rect 8300 22584 8352 22593
rect 8668 22627 8720 22636
rect 8668 22593 8677 22627
rect 8677 22593 8711 22627
rect 8711 22593 8720 22627
rect 8668 22584 8720 22593
rect 9128 22584 9180 22636
rect 10416 22584 10468 22636
rect 10692 22627 10744 22636
rect 10692 22593 10701 22627
rect 10701 22593 10735 22627
rect 10735 22593 10744 22627
rect 10692 22584 10744 22593
rect 11888 22584 11940 22636
rect 11980 22584 12032 22636
rect 18236 22652 18288 22704
rect 23204 22720 23256 22772
rect 23756 22720 23808 22772
rect 15660 22584 15712 22636
rect 16304 22584 16356 22636
rect 19248 22584 19300 22636
rect 19616 22627 19668 22636
rect 19616 22593 19625 22627
rect 19625 22593 19659 22627
rect 19659 22593 19668 22627
rect 19616 22584 19668 22593
rect 20444 22652 20496 22704
rect 21272 22652 21324 22704
rect 6184 22516 6236 22568
rect 6184 22423 6236 22432
rect 6184 22389 6193 22423
rect 6193 22389 6227 22423
rect 6227 22389 6236 22423
rect 6184 22380 6236 22389
rect 8392 22516 8444 22568
rect 10508 22516 10560 22568
rect 11336 22448 11388 22500
rect 12716 22559 12768 22568
rect 12716 22525 12725 22559
rect 12725 22525 12759 22559
rect 12759 22525 12768 22559
rect 12716 22516 12768 22525
rect 6644 22380 6696 22432
rect 7196 22380 7248 22432
rect 7380 22423 7432 22432
rect 7380 22389 7389 22423
rect 7389 22389 7423 22423
rect 7423 22389 7432 22423
rect 7380 22380 7432 22389
rect 9404 22380 9456 22432
rect 9772 22380 9824 22432
rect 11888 22423 11940 22432
rect 11888 22389 11897 22423
rect 11897 22389 11931 22423
rect 11931 22389 11940 22423
rect 11888 22380 11940 22389
rect 13728 22423 13780 22432
rect 13728 22389 13737 22423
rect 13737 22389 13771 22423
rect 13771 22389 13780 22423
rect 13728 22380 13780 22389
rect 14648 22380 14700 22432
rect 15108 22380 15160 22432
rect 15384 22380 15436 22432
rect 19892 22448 19944 22500
rect 23572 22627 23624 22636
rect 23572 22593 23581 22627
rect 23581 22593 23615 22627
rect 23615 22593 23624 22627
rect 23572 22584 23624 22593
rect 23664 22516 23716 22568
rect 20628 22448 20680 22500
rect 18512 22380 18564 22432
rect 19248 22380 19300 22432
rect 19708 22423 19760 22432
rect 19708 22389 19717 22423
rect 19717 22389 19751 22423
rect 19751 22389 19760 22423
rect 19708 22380 19760 22389
rect 20260 22423 20312 22432
rect 20260 22389 20269 22423
rect 20269 22389 20303 22423
rect 20303 22389 20312 22423
rect 20260 22380 20312 22389
rect 23480 22423 23532 22432
rect 23480 22389 23489 22423
rect 23489 22389 23523 22423
rect 23523 22389 23532 22423
rect 23480 22380 23532 22389
rect 24400 22423 24452 22432
rect 24400 22389 24409 22423
rect 24409 22389 24443 22423
rect 24443 22389 24452 22423
rect 24400 22380 24452 22389
rect 3917 22278 3969 22330
rect 3981 22278 4033 22330
rect 4045 22278 4097 22330
rect 4109 22278 4161 22330
rect 4173 22278 4225 22330
rect 9851 22278 9903 22330
rect 9915 22278 9967 22330
rect 9979 22278 10031 22330
rect 10043 22278 10095 22330
rect 10107 22278 10159 22330
rect 15785 22278 15837 22330
rect 15849 22278 15901 22330
rect 15913 22278 15965 22330
rect 15977 22278 16029 22330
rect 16041 22278 16093 22330
rect 21719 22278 21771 22330
rect 21783 22278 21835 22330
rect 21847 22278 21899 22330
rect 21911 22278 21963 22330
rect 21975 22278 22027 22330
rect 20 22176 72 22228
rect 1308 22176 1360 22228
rect 2780 22176 2832 22228
rect 4344 22176 4396 22228
rect 4988 22176 5040 22228
rect 5172 22176 5224 22228
rect 7380 22151 7432 22160
rect 7380 22117 7389 22151
rect 7389 22117 7423 22151
rect 7423 22117 7432 22151
rect 7380 22108 7432 22117
rect 2320 22040 2372 22092
rect 3884 22083 3936 22092
rect 3884 22049 3893 22083
rect 3893 22049 3927 22083
rect 3927 22049 3936 22083
rect 3884 22040 3936 22049
rect 4896 22040 4948 22092
rect 5540 22040 5592 22092
rect 6000 22040 6052 22092
rect 7196 22083 7248 22092
rect 7196 22049 7205 22083
rect 7205 22049 7239 22083
rect 7239 22049 7248 22083
rect 7196 22040 7248 22049
rect 7564 22219 7616 22228
rect 7564 22185 7573 22219
rect 7573 22185 7607 22219
rect 7607 22185 7616 22219
rect 7564 22176 7616 22185
rect 10508 22219 10560 22228
rect 10508 22185 10517 22219
rect 10517 22185 10551 22219
rect 10551 22185 10560 22219
rect 10508 22176 10560 22185
rect 11980 22176 12032 22228
rect 12716 22176 12768 22228
rect 11060 22108 11112 22160
rect 8576 22040 8628 22092
rect 9220 22040 9272 22092
rect 9404 22040 9456 22092
rect 2412 21972 2464 22024
rect 1860 21947 1912 21956
rect 1860 21913 1869 21947
rect 1869 21913 1903 21947
rect 1903 21913 1912 21947
rect 1860 21904 1912 21913
rect 2044 21904 2096 21956
rect 3608 21904 3660 21956
rect 5632 21972 5684 22024
rect 7288 21972 7340 22024
rect 7472 22015 7524 22024
rect 7472 21981 7481 22015
rect 7481 21981 7515 22015
rect 7515 21981 7524 22015
rect 7472 21972 7524 21981
rect 4436 21904 4488 21956
rect 6000 21904 6052 21956
rect 6184 21904 6236 21956
rect 8668 21972 8720 22024
rect 9312 21972 9364 22024
rect 10232 21972 10284 22024
rect 10416 21972 10468 22024
rect 8208 21904 8260 21956
rect 12440 21972 12492 22024
rect 15108 22151 15160 22160
rect 15108 22117 15117 22151
rect 15117 22117 15151 22151
rect 15151 22117 15160 22151
rect 15108 22108 15160 22117
rect 17868 22108 17920 22160
rect 18420 22108 18472 22160
rect 15384 22083 15436 22092
rect 15384 22049 15393 22083
rect 15393 22049 15427 22083
rect 15427 22049 15436 22083
rect 15384 22040 15436 22049
rect 16028 22040 16080 22092
rect 19708 22176 19760 22228
rect 20260 22176 20312 22228
rect 11520 21951 11545 21956
rect 11545 21951 11572 21956
rect 11520 21904 11572 21951
rect 2412 21836 2464 21888
rect 2964 21836 3016 21888
rect 12164 21836 12216 21888
rect 12256 21879 12308 21888
rect 12256 21845 12265 21879
rect 12265 21845 12299 21879
rect 12299 21845 12308 21879
rect 12256 21836 12308 21845
rect 13544 21836 13596 21888
rect 13820 21836 13872 21888
rect 15660 22015 15712 22024
rect 15660 21981 15669 22015
rect 15669 21981 15703 22015
rect 15703 21981 15712 22015
rect 15660 21972 15712 21981
rect 17316 21972 17368 22024
rect 17684 21972 17736 22024
rect 18236 21972 18288 22024
rect 19524 21972 19576 22024
rect 19892 22040 19944 22092
rect 20168 22040 20220 22092
rect 21824 22151 21876 22160
rect 21824 22117 21833 22151
rect 21833 22117 21867 22151
rect 21867 22117 21876 22151
rect 21824 22108 21876 22117
rect 22284 21972 22336 22024
rect 25688 21972 25740 22024
rect 20536 21947 20588 21956
rect 19616 21836 19668 21888
rect 19984 21879 20036 21888
rect 19984 21845 19993 21879
rect 19993 21845 20027 21879
rect 20027 21845 20036 21879
rect 19984 21836 20036 21845
rect 20536 21913 20570 21947
rect 20570 21913 20588 21947
rect 20536 21904 20588 21913
rect 22652 21947 22704 21956
rect 22652 21913 22664 21947
rect 22664 21913 22704 21947
rect 22652 21904 22704 21913
rect 23756 21879 23808 21888
rect 23756 21845 23765 21879
rect 23765 21845 23799 21879
rect 23799 21845 23808 21879
rect 23756 21836 23808 21845
rect 24124 21879 24176 21888
rect 24124 21845 24133 21879
rect 24133 21845 24167 21879
rect 24167 21845 24176 21879
rect 24124 21836 24176 21845
rect 6884 21734 6936 21786
rect 6948 21734 7000 21786
rect 7012 21734 7064 21786
rect 7076 21734 7128 21786
rect 7140 21734 7192 21786
rect 12818 21734 12870 21786
rect 12882 21734 12934 21786
rect 12946 21734 12998 21786
rect 13010 21734 13062 21786
rect 13074 21734 13126 21786
rect 18752 21734 18804 21786
rect 18816 21734 18868 21786
rect 18880 21734 18932 21786
rect 18944 21734 18996 21786
rect 19008 21734 19060 21786
rect 24686 21734 24738 21786
rect 24750 21734 24802 21786
rect 24814 21734 24866 21786
rect 24878 21734 24930 21786
rect 24942 21734 24994 21786
rect 1032 21564 1084 21616
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 2136 21564 2188 21616
rect 848 21428 900 21480
rect 2044 21496 2096 21548
rect 3884 21632 3936 21684
rect 6736 21632 6788 21684
rect 8208 21632 8260 21684
rect 8392 21632 8444 21684
rect 12164 21632 12216 21684
rect 2596 21564 2648 21616
rect 2504 21539 2556 21548
rect 2504 21505 2511 21539
rect 2511 21505 2545 21539
rect 2545 21505 2556 21539
rect 2504 21496 2556 21505
rect 3056 21496 3108 21548
rect 2136 21335 2188 21344
rect 2136 21301 2145 21335
rect 2145 21301 2179 21335
rect 2179 21301 2188 21335
rect 2136 21292 2188 21301
rect 2320 21292 2372 21344
rect 3240 21335 3292 21344
rect 3240 21301 3249 21335
rect 3249 21301 3283 21335
rect 3283 21301 3292 21335
rect 3240 21292 3292 21301
rect 3792 21496 3844 21548
rect 4252 21564 4304 21616
rect 7656 21564 7708 21616
rect 7564 21496 7616 21548
rect 7748 21496 7800 21548
rect 8576 21564 8628 21616
rect 13544 21607 13596 21616
rect 13544 21573 13553 21607
rect 13553 21573 13587 21607
rect 13587 21573 13596 21607
rect 13544 21564 13596 21573
rect 8392 21496 8444 21548
rect 9312 21496 9364 21548
rect 12348 21496 12400 21548
rect 13268 21496 13320 21548
rect 14188 21632 14240 21684
rect 15660 21632 15712 21684
rect 19892 21675 19944 21684
rect 19892 21641 19901 21675
rect 19901 21641 19935 21675
rect 19935 21641 19944 21675
rect 19892 21632 19944 21641
rect 19984 21632 20036 21684
rect 20996 21632 21048 21684
rect 13820 21496 13872 21548
rect 14004 21496 14056 21548
rect 14924 21496 14976 21548
rect 16672 21539 16724 21548
rect 16672 21505 16681 21539
rect 16681 21505 16715 21539
rect 16715 21505 16724 21539
rect 16672 21496 16724 21505
rect 17684 21539 17736 21548
rect 17684 21505 17718 21539
rect 17718 21505 17736 21539
rect 17684 21496 17736 21505
rect 3516 21428 3568 21480
rect 6184 21428 6236 21480
rect 6644 21471 6696 21480
rect 6644 21437 6653 21471
rect 6653 21437 6687 21471
rect 6687 21437 6696 21471
rect 6644 21428 6696 21437
rect 11060 21428 11112 21480
rect 13728 21428 13780 21480
rect 14740 21471 14792 21480
rect 14740 21437 14749 21471
rect 14749 21437 14783 21471
rect 14783 21437 14792 21471
rect 14740 21428 14792 21437
rect 16396 21428 16448 21480
rect 16856 21471 16908 21480
rect 16856 21437 16865 21471
rect 16865 21437 16899 21471
rect 16899 21437 16908 21471
rect 16856 21428 16908 21437
rect 4436 21360 4488 21412
rect 17868 21471 17920 21480
rect 17868 21437 17877 21471
rect 17877 21437 17911 21471
rect 17911 21437 17920 21471
rect 17868 21428 17920 21437
rect 18052 21428 18104 21480
rect 18604 21428 18656 21480
rect 4528 21292 4580 21344
rect 7656 21335 7708 21344
rect 7656 21301 7665 21335
rect 7665 21301 7699 21335
rect 7699 21301 7708 21335
rect 7656 21292 7708 21301
rect 20536 21496 20588 21548
rect 9036 21292 9088 21344
rect 12532 21335 12584 21344
rect 12532 21301 12541 21335
rect 12541 21301 12575 21335
rect 12575 21301 12584 21335
rect 12532 21292 12584 21301
rect 15108 21292 15160 21344
rect 15660 21292 15712 21344
rect 16488 21292 16540 21344
rect 17040 21292 17092 21344
rect 17684 21292 17736 21344
rect 18512 21335 18564 21344
rect 18512 21301 18521 21335
rect 18521 21301 18555 21335
rect 18555 21301 18564 21335
rect 18512 21292 18564 21301
rect 19892 21292 19944 21344
rect 21180 21360 21232 21412
rect 21916 21564 21968 21616
rect 22008 21496 22060 21548
rect 22652 21632 22704 21684
rect 23664 21632 23716 21684
rect 22468 21496 22520 21548
rect 23020 21535 23045 21548
rect 23045 21535 23072 21548
rect 23020 21496 23072 21535
rect 24492 21496 24544 21548
rect 25320 21496 25372 21548
rect 23480 21428 23532 21480
rect 22652 21360 22704 21412
rect 24124 21360 24176 21412
rect 22468 21335 22520 21344
rect 22468 21301 22477 21335
rect 22477 21301 22511 21335
rect 22511 21301 22520 21335
rect 22468 21292 22520 21301
rect 24216 21335 24268 21344
rect 24216 21301 24225 21335
rect 24225 21301 24259 21335
rect 24259 21301 24268 21335
rect 24216 21292 24268 21301
rect 3917 21190 3969 21242
rect 3981 21190 4033 21242
rect 4045 21190 4097 21242
rect 4109 21190 4161 21242
rect 4173 21190 4225 21242
rect 9851 21190 9903 21242
rect 9915 21190 9967 21242
rect 9979 21190 10031 21242
rect 10043 21190 10095 21242
rect 10107 21190 10159 21242
rect 15785 21190 15837 21242
rect 15849 21190 15901 21242
rect 15913 21190 15965 21242
rect 15977 21190 16029 21242
rect 16041 21190 16093 21242
rect 21719 21190 21771 21242
rect 21783 21190 21835 21242
rect 21847 21190 21899 21242
rect 21911 21190 21963 21242
rect 21975 21190 22027 21242
rect 1676 21088 1728 21140
rect 4436 21088 4488 21140
rect 2044 21020 2096 21072
rect 2872 20952 2924 21004
rect 3516 20952 3568 21004
rect 3700 20952 3752 21004
rect 4988 21088 5040 21140
rect 7380 21088 7432 21140
rect 9036 21088 9088 21140
rect 11336 21088 11388 21140
rect 940 20884 992 20936
rect 2044 20884 2096 20936
rect 3792 20884 3844 20936
rect 6276 20884 6328 20936
rect 7288 21020 7340 21072
rect 7656 20952 7708 21004
rect 9220 20952 9272 21004
rect 11152 20952 11204 21004
rect 12532 21088 12584 21140
rect 14740 21088 14792 21140
rect 16672 21088 16724 21140
rect 18604 21088 18656 21140
rect 19064 21088 19116 21140
rect 17040 21063 17092 21072
rect 17040 21029 17049 21063
rect 17049 21029 17083 21063
rect 17083 21029 17092 21063
rect 17040 21020 17092 21029
rect 12256 20952 12308 21004
rect 7288 20884 7340 20936
rect 1492 20859 1544 20868
rect 1492 20825 1501 20859
rect 1501 20825 1535 20859
rect 1535 20825 1544 20859
rect 1492 20816 1544 20825
rect 2596 20816 2648 20868
rect 2688 20816 2740 20868
rect 7472 20884 7524 20936
rect 7564 20884 7616 20936
rect 2136 20748 2188 20800
rect 2504 20748 2556 20800
rect 3056 20748 3108 20800
rect 3516 20748 3568 20800
rect 5448 20748 5500 20800
rect 7748 20859 7800 20868
rect 7748 20825 7757 20859
rect 7757 20825 7791 20859
rect 7791 20825 7800 20859
rect 7748 20816 7800 20825
rect 8300 20816 8352 20868
rect 8944 20816 8996 20868
rect 9036 20748 9088 20800
rect 10416 20791 10468 20800
rect 10416 20757 10425 20791
rect 10425 20757 10459 20791
rect 10459 20757 10468 20791
rect 10416 20748 10468 20757
rect 12440 20927 12492 20936
rect 12440 20893 12449 20927
rect 12449 20893 12483 20927
rect 12483 20893 12492 20927
rect 12440 20884 12492 20893
rect 12532 20927 12584 20936
rect 14556 20952 14608 21004
rect 15016 20995 15068 21004
rect 15016 20961 15025 20995
rect 15025 20961 15059 20995
rect 15059 20961 15068 20995
rect 15016 20952 15068 20961
rect 12532 20893 12566 20927
rect 12566 20893 12584 20927
rect 12532 20884 12584 20893
rect 18236 20952 18288 21004
rect 15568 20816 15620 20868
rect 16764 20884 16816 20936
rect 17316 20927 17368 20936
rect 17316 20893 17325 20927
rect 17325 20893 17359 20927
rect 17359 20893 17368 20927
rect 17316 20884 17368 20893
rect 17408 20927 17460 20936
rect 17408 20893 17442 20927
rect 17442 20893 17460 20927
rect 17408 20884 17460 20893
rect 17592 20927 17644 20936
rect 17592 20893 17601 20927
rect 17601 20893 17635 20927
rect 17635 20893 17644 20927
rect 17592 20884 17644 20893
rect 18512 20923 18564 20936
rect 19524 21020 19576 21072
rect 19984 21020 20036 21072
rect 22100 21088 22152 21140
rect 22468 21088 22520 21140
rect 22652 21088 22704 21140
rect 24216 21088 24268 21140
rect 18972 20952 19024 21004
rect 18512 20889 18529 20923
rect 18529 20889 18563 20923
rect 18563 20889 18564 20923
rect 18512 20884 18564 20889
rect 18512 20748 18564 20800
rect 19432 20748 19484 20800
rect 19524 20748 19576 20800
rect 21180 20995 21232 21004
rect 21180 20961 21189 20995
rect 21189 20961 21223 20995
rect 21223 20961 21232 20995
rect 21180 20952 21232 20961
rect 22836 20816 22888 20868
rect 19708 20791 19760 20800
rect 19708 20757 19717 20791
rect 19717 20757 19751 20791
rect 19751 20757 19760 20791
rect 19708 20748 19760 20757
rect 23940 20791 23992 20800
rect 23940 20757 23949 20791
rect 23949 20757 23983 20791
rect 23983 20757 23992 20791
rect 23940 20748 23992 20757
rect 6884 20646 6936 20698
rect 6948 20646 7000 20698
rect 7012 20646 7064 20698
rect 7076 20646 7128 20698
rect 7140 20646 7192 20698
rect 12818 20646 12870 20698
rect 12882 20646 12934 20698
rect 12946 20646 12998 20698
rect 13010 20646 13062 20698
rect 13074 20646 13126 20698
rect 18752 20646 18804 20698
rect 18816 20646 18868 20698
rect 18880 20646 18932 20698
rect 18944 20646 18996 20698
rect 19008 20646 19060 20698
rect 24686 20646 24738 20698
rect 24750 20646 24802 20698
rect 24814 20646 24866 20698
rect 24878 20646 24930 20698
rect 24942 20646 24994 20698
rect 1216 20544 1268 20596
rect 2596 20544 2648 20596
rect 7380 20544 7432 20596
rect 7748 20544 7800 20596
rect 10324 20544 10376 20596
rect 10784 20544 10836 20596
rect 11520 20544 11572 20596
rect 12072 20544 12124 20596
rect 12440 20544 12492 20596
rect 16488 20544 16540 20596
rect 17500 20544 17552 20596
rect 17592 20544 17644 20596
rect 17868 20544 17920 20596
rect 18512 20544 18564 20596
rect 2780 20476 2832 20528
rect 1400 20451 1452 20460
rect 1400 20417 1409 20451
rect 1409 20417 1443 20451
rect 1443 20417 1452 20451
rect 1400 20408 1452 20417
rect 1216 20340 1268 20392
rect 3332 20476 3384 20528
rect 4252 20476 4304 20528
rect 4620 20476 4672 20528
rect 6184 20476 6236 20528
rect 2964 20408 3016 20460
rect 3148 20451 3200 20460
rect 3148 20417 3157 20451
rect 3157 20417 3191 20451
rect 3191 20417 3200 20451
rect 3148 20408 3200 20417
rect 3240 20451 3292 20460
rect 3240 20417 3249 20451
rect 3249 20417 3283 20451
rect 3283 20417 3292 20451
rect 3240 20408 3292 20417
rect 4712 20408 4764 20460
rect 4896 20408 4948 20460
rect 5172 20451 5224 20460
rect 5172 20417 5181 20451
rect 5181 20417 5215 20451
rect 5215 20417 5224 20451
rect 5172 20408 5224 20417
rect 5356 20408 5408 20460
rect 6644 20408 6696 20460
rect 7472 20408 7524 20460
rect 10416 20476 10468 20528
rect 10508 20519 10560 20528
rect 10508 20485 10517 20519
rect 10517 20485 10551 20519
rect 10551 20485 10560 20519
rect 10508 20476 10560 20485
rect 9036 20408 9088 20460
rect 9588 20408 9640 20460
rect 9680 20451 9732 20460
rect 9680 20417 9689 20451
rect 9689 20417 9723 20451
rect 9723 20417 9732 20451
rect 9680 20408 9732 20417
rect 10968 20408 11020 20460
rect 15292 20476 15344 20528
rect 19524 20544 19576 20596
rect 22744 20544 22796 20596
rect 23572 20544 23624 20596
rect 24400 20544 24452 20596
rect 3056 20340 3108 20392
rect 5448 20340 5500 20392
rect 5908 20340 5960 20392
rect 6736 20340 6788 20392
rect 12164 20340 12216 20392
rect 14004 20408 14056 20460
rect 14372 20408 14424 20460
rect 15016 20408 15068 20460
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 13544 20340 13596 20392
rect 10968 20272 11020 20324
rect 11980 20272 12032 20324
rect 12532 20272 12584 20324
rect 15292 20340 15344 20392
rect 14556 20272 14608 20324
rect 16948 20272 17000 20324
rect 4160 20247 4212 20256
rect 4160 20213 4169 20247
rect 4169 20213 4203 20247
rect 4203 20213 4212 20247
rect 4160 20204 4212 20213
rect 6092 20247 6144 20256
rect 6092 20213 6101 20247
rect 6101 20213 6135 20247
rect 6135 20213 6144 20247
rect 6092 20204 6144 20213
rect 6184 20204 6236 20256
rect 7840 20204 7892 20256
rect 10692 20247 10744 20256
rect 10692 20213 10701 20247
rect 10701 20213 10735 20247
rect 10735 20213 10744 20247
rect 10692 20204 10744 20213
rect 11520 20204 11572 20256
rect 12716 20204 12768 20256
rect 18512 20451 18564 20460
rect 18512 20417 18521 20451
rect 18521 20417 18555 20451
rect 18555 20417 18564 20451
rect 18512 20408 18564 20417
rect 18604 20451 18656 20460
rect 18604 20417 18613 20451
rect 18613 20417 18647 20451
rect 18647 20417 18656 20451
rect 18604 20408 18656 20417
rect 19248 20408 19300 20460
rect 19708 20408 19760 20460
rect 22560 20408 22612 20460
rect 23756 20476 23808 20528
rect 23848 20476 23900 20528
rect 25872 20408 25924 20460
rect 19064 20272 19116 20324
rect 20260 20204 20312 20256
rect 20720 20247 20772 20256
rect 20720 20213 20729 20247
rect 20729 20213 20763 20247
rect 20763 20213 20772 20247
rect 20720 20204 20772 20213
rect 21364 20204 21416 20256
rect 22744 20204 22796 20256
rect 22836 20204 22888 20256
rect 23756 20247 23808 20256
rect 23756 20213 23765 20247
rect 23765 20213 23799 20247
rect 23799 20213 23808 20247
rect 23756 20204 23808 20213
rect 3917 20102 3969 20154
rect 3981 20102 4033 20154
rect 4045 20102 4097 20154
rect 4109 20102 4161 20154
rect 4173 20102 4225 20154
rect 9851 20102 9903 20154
rect 9915 20102 9967 20154
rect 9979 20102 10031 20154
rect 10043 20102 10095 20154
rect 10107 20102 10159 20154
rect 15785 20102 15837 20154
rect 15849 20102 15901 20154
rect 15913 20102 15965 20154
rect 15977 20102 16029 20154
rect 16041 20102 16093 20154
rect 21719 20102 21771 20154
rect 21783 20102 21835 20154
rect 21847 20102 21899 20154
rect 21911 20102 21963 20154
rect 21975 20102 22027 20154
rect 1768 20000 1820 20052
rect 1952 20000 2004 20052
rect 2688 19975 2740 19984
rect 2688 19941 2697 19975
rect 2697 19941 2731 19975
rect 2731 19941 2740 19975
rect 2688 19932 2740 19941
rect 3516 20043 3568 20052
rect 3516 20009 3525 20043
rect 3525 20009 3559 20043
rect 3559 20009 3568 20043
rect 3516 20000 3568 20009
rect 5172 20000 5224 20052
rect 7564 20000 7616 20052
rect 8024 20000 8076 20052
rect 4712 19932 4764 19984
rect 1584 19796 1636 19848
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 4988 19864 5040 19916
rect 9036 19864 9088 19916
rect 9220 19864 9272 19916
rect 9404 19864 9456 19916
rect 1308 19728 1360 19780
rect 3332 19839 3384 19848
rect 3332 19805 3341 19839
rect 3341 19805 3375 19839
rect 3375 19805 3384 19839
rect 3332 19796 3384 19805
rect 3516 19796 3568 19848
rect 3792 19839 3844 19848
rect 3792 19805 3801 19839
rect 3801 19805 3835 19839
rect 3835 19805 3844 19839
rect 3792 19796 3844 19805
rect 10968 20000 11020 20052
rect 11612 20000 11664 20052
rect 11152 19864 11204 19916
rect 11336 19864 11388 19916
rect 11980 20000 12032 20052
rect 12072 20000 12124 20052
rect 14556 20000 14608 20052
rect 14740 20000 14792 20052
rect 18512 20000 18564 20052
rect 14372 19864 14424 19916
rect 17040 19864 17092 19916
rect 204 19660 256 19712
rect 1584 19660 1636 19712
rect 1676 19660 1728 19712
rect 5356 19728 5408 19780
rect 7656 19728 7708 19780
rect 8024 19728 8076 19780
rect 9496 19728 9548 19780
rect 3608 19660 3660 19712
rect 3884 19660 3936 19712
rect 8576 19660 8628 19712
rect 8944 19660 8996 19712
rect 9220 19660 9272 19712
rect 11980 19839 12032 19848
rect 11980 19805 11989 19839
rect 11989 19805 12023 19839
rect 12023 19805 12032 19839
rect 11980 19796 12032 19805
rect 12256 19839 12308 19848
rect 12256 19805 12263 19839
rect 12263 19805 12297 19839
rect 12297 19805 12308 19839
rect 12256 19796 12308 19805
rect 13820 19796 13872 19848
rect 14740 19839 14792 19848
rect 14740 19805 14747 19839
rect 14747 19805 14781 19839
rect 14781 19805 14792 19839
rect 14740 19796 14792 19805
rect 9956 19775 9981 19780
rect 9981 19775 10008 19780
rect 9956 19728 10008 19775
rect 11060 19728 11112 19780
rect 11152 19728 11204 19780
rect 13636 19728 13688 19780
rect 16488 19796 16540 19848
rect 14924 19728 14976 19780
rect 17500 19728 17552 19780
rect 19064 20000 19116 20052
rect 19892 20000 19944 20052
rect 20720 20000 20772 20052
rect 21364 20000 21416 20052
rect 21548 20000 21600 20052
rect 23848 20000 23900 20052
rect 20720 19864 20772 19916
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 19616 19796 19668 19848
rect 21824 19839 21876 19848
rect 21824 19805 21833 19839
rect 21833 19805 21867 19839
rect 21867 19805 21876 19839
rect 21824 19796 21876 19805
rect 22284 19796 22336 19848
rect 12072 19660 12124 19712
rect 13176 19660 13228 19712
rect 15476 19703 15528 19712
rect 15476 19669 15485 19703
rect 15485 19669 15519 19703
rect 15519 19669 15528 19703
rect 15476 19660 15528 19669
rect 15752 19660 15804 19712
rect 20076 19660 20128 19712
rect 20168 19660 20220 19712
rect 22560 19728 22612 19780
rect 23296 19796 23348 19848
rect 24216 19771 24268 19780
rect 24216 19737 24225 19771
rect 24225 19737 24259 19771
rect 24259 19737 24268 19771
rect 24216 19728 24268 19737
rect 22652 19660 22704 19712
rect 23572 19703 23624 19712
rect 23572 19669 23581 19703
rect 23581 19669 23615 19703
rect 23615 19669 23624 19703
rect 23572 19660 23624 19669
rect 6884 19558 6936 19610
rect 6948 19558 7000 19610
rect 7012 19558 7064 19610
rect 7076 19558 7128 19610
rect 7140 19558 7192 19610
rect 12818 19558 12870 19610
rect 12882 19558 12934 19610
rect 12946 19558 12998 19610
rect 13010 19558 13062 19610
rect 13074 19558 13126 19610
rect 18752 19558 18804 19610
rect 18816 19558 18868 19610
rect 18880 19558 18932 19610
rect 18944 19558 18996 19610
rect 19008 19558 19060 19610
rect 24686 19558 24738 19610
rect 24750 19558 24802 19610
rect 24814 19558 24866 19610
rect 24878 19558 24930 19610
rect 24942 19558 24994 19610
rect 1308 19456 1360 19508
rect 3792 19456 3844 19508
rect 3884 19456 3936 19508
rect 6644 19456 6696 19508
rect 7564 19456 7616 19508
rect 7656 19456 7708 19508
rect 7748 19456 7800 19508
rect 9218 19456 9270 19508
rect 1584 19320 1636 19372
rect 1768 19320 1820 19372
rect 3148 19388 3200 19440
rect 2872 19363 2924 19372
rect 2872 19329 2881 19363
rect 2881 19329 2915 19363
rect 2915 19329 2924 19363
rect 2872 19320 2924 19329
rect 3516 19320 3568 19372
rect 2320 19116 2372 19168
rect 2412 19159 2464 19168
rect 2412 19125 2421 19159
rect 2421 19125 2455 19159
rect 2455 19125 2464 19159
rect 2412 19116 2464 19125
rect 3056 19184 3108 19236
rect 5540 19252 5592 19304
rect 8944 19363 8996 19372
rect 8944 19329 8953 19363
rect 8953 19329 8987 19363
rect 8987 19329 8996 19363
rect 8944 19320 8996 19329
rect 9404 19456 9456 19508
rect 9496 19456 9548 19508
rect 12164 19456 12216 19508
rect 12256 19456 12308 19508
rect 12900 19456 12952 19508
rect 11520 19363 11572 19372
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 11520 19320 11572 19329
rect 12992 19388 13044 19440
rect 13544 19388 13596 19440
rect 13728 19388 13780 19440
rect 12532 19320 12584 19372
rect 12716 19320 12768 19372
rect 3240 19116 3292 19168
rect 8852 19184 8904 19236
rect 16856 19456 16908 19508
rect 20812 19456 20864 19508
rect 16488 19388 16540 19440
rect 15476 19363 15528 19372
rect 15476 19329 15485 19363
rect 15485 19329 15519 19363
rect 15519 19329 15528 19363
rect 15476 19320 15528 19329
rect 19616 19320 19668 19372
rect 20444 19320 20496 19372
rect 21088 19320 21140 19372
rect 21824 19320 21876 19372
rect 22376 19320 22428 19372
rect 24032 19388 24084 19440
rect 25872 19320 25924 19372
rect 14832 19252 14884 19304
rect 15200 19295 15252 19304
rect 15200 19261 15209 19295
rect 15209 19261 15243 19295
rect 15243 19261 15252 19295
rect 15200 19252 15252 19261
rect 15292 19295 15344 19304
rect 15292 19261 15326 19295
rect 15326 19261 15344 19295
rect 15292 19252 15344 19261
rect 16672 19295 16724 19304
rect 16672 19261 16681 19295
rect 16681 19261 16715 19295
rect 16715 19261 16724 19295
rect 16672 19252 16724 19261
rect 8576 19116 8628 19168
rect 14924 19227 14976 19236
rect 14924 19193 14933 19227
rect 14933 19193 14967 19227
rect 14967 19193 14976 19227
rect 14924 19184 14976 19193
rect 14004 19116 14056 19168
rect 14740 19116 14792 19168
rect 16120 19159 16172 19168
rect 16120 19125 16129 19159
rect 16129 19125 16163 19159
rect 16163 19125 16172 19159
rect 16120 19116 16172 19125
rect 16488 19159 16540 19168
rect 16488 19125 16497 19159
rect 16497 19125 16531 19159
rect 16531 19125 16540 19159
rect 16488 19116 16540 19125
rect 17684 19159 17736 19168
rect 17684 19125 17693 19159
rect 17693 19125 17727 19159
rect 17727 19125 17736 19159
rect 17684 19116 17736 19125
rect 18604 19116 18656 19168
rect 23480 19159 23532 19168
rect 23480 19125 23489 19159
rect 23489 19125 23523 19159
rect 23523 19125 23532 19159
rect 23480 19116 23532 19125
rect 24400 19159 24452 19168
rect 24400 19125 24409 19159
rect 24409 19125 24443 19159
rect 24443 19125 24452 19159
rect 24400 19116 24452 19125
rect 3917 19014 3969 19066
rect 3981 19014 4033 19066
rect 4045 19014 4097 19066
rect 4109 19014 4161 19066
rect 4173 19014 4225 19066
rect 9851 19014 9903 19066
rect 9915 19014 9967 19066
rect 9979 19014 10031 19066
rect 10043 19014 10095 19066
rect 10107 19014 10159 19066
rect 15785 19014 15837 19066
rect 15849 19014 15901 19066
rect 15913 19014 15965 19066
rect 15977 19014 16029 19066
rect 16041 19014 16093 19066
rect 21719 19014 21771 19066
rect 21783 19014 21835 19066
rect 21847 19014 21899 19066
rect 21911 19014 21963 19066
rect 21975 19014 22027 19066
rect 1492 18912 1544 18964
rect 6644 18912 6696 18964
rect 8852 18912 8904 18964
rect 10508 18912 10560 18964
rect 1952 18887 2004 18896
rect 1952 18853 1961 18887
rect 1961 18853 1995 18887
rect 1995 18853 2004 18887
rect 1952 18844 2004 18853
rect 940 18776 992 18828
rect 756 18708 808 18760
rect 1584 18615 1636 18624
rect 1584 18581 1593 18615
rect 1593 18581 1627 18615
rect 1627 18581 1636 18615
rect 1584 18572 1636 18581
rect 3700 18776 3752 18828
rect 4620 18708 4672 18760
rect 5540 18708 5592 18760
rect 2596 18687 2621 18692
rect 2621 18687 2648 18692
rect 2596 18640 2648 18687
rect 3608 18640 3660 18692
rect 7288 18708 7340 18760
rect 7564 18708 7616 18760
rect 7656 18751 7708 18760
rect 7656 18717 7665 18751
rect 7665 18717 7699 18751
rect 7699 18717 7708 18751
rect 7656 18708 7708 18717
rect 7748 18751 7800 18760
rect 7748 18717 7757 18751
rect 7757 18717 7791 18751
rect 7791 18717 7800 18751
rect 7748 18708 7800 18717
rect 8208 18708 8260 18760
rect 9036 18776 9088 18828
rect 10232 18776 10284 18828
rect 10968 18776 11020 18828
rect 9588 18708 9640 18760
rect 12440 18819 12492 18828
rect 12440 18785 12449 18819
rect 12449 18785 12483 18819
rect 12483 18785 12492 18819
rect 12440 18776 12492 18785
rect 14924 18912 14976 18964
rect 15476 18912 15528 18964
rect 16396 18912 16448 18964
rect 16488 18912 16540 18964
rect 20996 18912 21048 18964
rect 15292 18776 15344 18828
rect 16396 18819 16448 18828
rect 16396 18785 16405 18819
rect 16405 18785 16439 18819
rect 16439 18785 16448 18819
rect 16396 18776 16448 18785
rect 17684 18776 17736 18828
rect 2780 18572 2832 18624
rect 4344 18572 4396 18624
rect 4988 18572 5040 18624
rect 5172 18572 5224 18624
rect 6184 18572 6236 18624
rect 11060 18640 11112 18692
rect 12072 18640 12124 18692
rect 12532 18640 12584 18692
rect 12900 18640 12952 18692
rect 12992 18640 13044 18692
rect 13728 18640 13780 18692
rect 14740 18708 14792 18760
rect 14832 18708 14884 18760
rect 16856 18708 16908 18760
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 19800 18751 19852 18760
rect 19800 18717 19809 18751
rect 19809 18717 19843 18751
rect 19843 18717 19852 18751
rect 19800 18708 19852 18717
rect 23664 18819 23716 18828
rect 23664 18785 23673 18819
rect 23673 18785 23707 18819
rect 23707 18785 23716 18819
rect 23664 18776 23716 18785
rect 8576 18572 8628 18624
rect 8668 18615 8720 18624
rect 8668 18581 8677 18615
rect 8677 18581 8711 18615
rect 8711 18581 8720 18615
rect 8668 18572 8720 18581
rect 9680 18572 9732 18624
rect 11980 18572 12032 18624
rect 12440 18572 12492 18624
rect 17684 18640 17736 18692
rect 20352 18640 20404 18692
rect 22744 18708 22796 18760
rect 23480 18708 23532 18760
rect 23572 18708 23624 18760
rect 24124 18708 24176 18760
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 14372 18572 14424 18624
rect 15016 18572 15068 18624
rect 16672 18572 16724 18624
rect 17500 18572 17552 18624
rect 18052 18572 18104 18624
rect 19708 18615 19760 18624
rect 19708 18581 19717 18615
rect 19717 18581 19751 18615
rect 19751 18581 19760 18615
rect 19708 18572 19760 18581
rect 21916 18572 21968 18624
rect 23480 18572 23532 18624
rect 23572 18572 23624 18624
rect 24124 18615 24176 18624
rect 24124 18581 24133 18615
rect 24133 18581 24167 18615
rect 24167 18581 24176 18615
rect 24124 18572 24176 18581
rect 24216 18572 24268 18624
rect 6884 18470 6936 18522
rect 6948 18470 7000 18522
rect 7012 18470 7064 18522
rect 7076 18470 7128 18522
rect 7140 18470 7192 18522
rect 12818 18470 12870 18522
rect 12882 18470 12934 18522
rect 12946 18470 12998 18522
rect 13010 18470 13062 18522
rect 13074 18470 13126 18522
rect 18752 18470 18804 18522
rect 18816 18470 18868 18522
rect 18880 18470 18932 18522
rect 18944 18470 18996 18522
rect 19008 18470 19060 18522
rect 24686 18470 24738 18522
rect 24750 18470 24802 18522
rect 24814 18470 24866 18522
rect 24878 18470 24930 18522
rect 24942 18470 24994 18522
rect 3516 18368 3568 18420
rect 5908 18368 5960 18420
rect 6552 18411 6604 18420
rect 6552 18377 6561 18411
rect 6561 18377 6595 18411
rect 6595 18377 6604 18411
rect 6552 18368 6604 18377
rect 6736 18368 6788 18420
rect 756 18300 808 18352
rect 1676 18343 1728 18352
rect 1676 18309 1685 18343
rect 1685 18309 1719 18343
rect 1719 18309 1728 18343
rect 1676 18300 1728 18309
rect 1860 18232 1912 18284
rect 1952 18275 2004 18284
rect 1952 18241 1961 18275
rect 1961 18241 1995 18275
rect 1995 18241 2004 18275
rect 1952 18232 2004 18241
rect 2228 18300 2280 18352
rect 3240 18275 3292 18284
rect 3240 18241 3249 18275
rect 3249 18241 3283 18275
rect 3283 18241 3292 18275
rect 3240 18232 3292 18241
rect 2320 18164 2372 18216
rect 3792 18164 3844 18216
rect 4344 18232 4396 18284
rect 4988 18275 5040 18284
rect 4988 18241 5022 18275
rect 5022 18241 5040 18275
rect 4988 18232 5040 18241
rect 5172 18275 5224 18284
rect 5172 18241 5181 18275
rect 5181 18241 5215 18275
rect 5215 18241 5224 18275
rect 5172 18232 5224 18241
rect 6644 18300 6696 18352
rect 6920 18275 6972 18284
rect 6920 18241 6929 18275
rect 6929 18241 6963 18275
rect 6963 18241 6972 18275
rect 6920 18232 6972 18241
rect 7288 18275 7340 18284
rect 7288 18241 7297 18275
rect 7297 18241 7331 18275
rect 7331 18241 7340 18275
rect 7288 18232 7340 18241
rect 7472 18300 7524 18352
rect 2780 18096 2832 18148
rect 3056 18028 3108 18080
rect 3332 18028 3384 18080
rect 4160 18207 4212 18216
rect 4160 18173 4169 18207
rect 4169 18173 4203 18207
rect 4203 18173 4212 18207
rect 4160 18164 4212 18173
rect 4528 18164 4580 18216
rect 6736 18164 6788 18216
rect 9036 18232 9088 18284
rect 7748 18164 7800 18216
rect 10232 18368 10284 18420
rect 10600 18368 10652 18420
rect 11980 18300 12032 18352
rect 12900 18300 12952 18352
rect 13728 18368 13780 18420
rect 15476 18368 15528 18420
rect 16396 18368 16448 18420
rect 9680 18232 9732 18284
rect 10600 18275 10652 18284
rect 10600 18241 10609 18275
rect 10609 18241 10643 18275
rect 10643 18241 10652 18275
rect 10600 18232 10652 18241
rect 10968 18232 11020 18284
rect 11060 18232 11112 18284
rect 12256 18232 12308 18284
rect 12624 18232 12676 18284
rect 13728 18275 13780 18284
rect 13728 18241 13737 18275
rect 13737 18241 13771 18275
rect 13771 18241 13780 18275
rect 13728 18232 13780 18241
rect 14004 18275 14056 18284
rect 14004 18241 14013 18275
rect 14013 18241 14047 18275
rect 14047 18241 14056 18275
rect 14004 18232 14056 18241
rect 15016 18232 15068 18284
rect 18052 18232 18104 18284
rect 19340 18232 19392 18284
rect 19432 18275 19484 18284
rect 19432 18241 19441 18275
rect 19441 18241 19475 18275
rect 19475 18241 19484 18275
rect 19432 18232 19484 18241
rect 19800 18368 19852 18420
rect 22284 18368 22336 18420
rect 20352 18343 20404 18352
rect 20352 18309 20375 18343
rect 20375 18309 20404 18343
rect 20352 18300 20404 18309
rect 22100 18343 22152 18352
rect 22100 18309 22109 18343
rect 22109 18309 22143 18343
rect 22143 18309 22152 18343
rect 22100 18300 22152 18309
rect 21640 18232 21692 18284
rect 21916 18275 21968 18284
rect 21916 18241 21925 18275
rect 21925 18241 21959 18275
rect 21959 18241 21968 18275
rect 21916 18232 21968 18241
rect 23388 18368 23440 18420
rect 23480 18368 23532 18420
rect 23664 18368 23716 18420
rect 24400 18411 24452 18420
rect 24400 18377 24409 18411
rect 24409 18377 24443 18411
rect 24443 18377 24452 18411
rect 24400 18368 24452 18377
rect 4896 18028 4948 18080
rect 5264 18028 5316 18080
rect 5540 18028 5592 18080
rect 5908 18028 5960 18080
rect 6368 18028 6420 18080
rect 12440 18096 12492 18148
rect 13452 18207 13504 18216
rect 13452 18173 13461 18207
rect 13461 18173 13495 18207
rect 13495 18173 13504 18207
rect 13452 18164 13504 18173
rect 14648 18139 14700 18148
rect 14648 18105 14657 18139
rect 14657 18105 14691 18139
rect 14691 18105 14700 18139
rect 14648 18096 14700 18105
rect 10968 18028 11020 18080
rect 11888 18028 11940 18080
rect 11980 18071 12032 18080
rect 11980 18037 11989 18071
rect 11989 18037 12023 18071
rect 12023 18037 12032 18071
rect 11980 18028 12032 18037
rect 12348 18028 12400 18080
rect 17960 18096 18012 18148
rect 15936 18028 15988 18080
rect 19524 18071 19576 18080
rect 19524 18037 19533 18071
rect 19533 18037 19567 18071
rect 19567 18037 19576 18071
rect 19524 18028 19576 18037
rect 23756 18275 23808 18284
rect 23756 18241 23765 18275
rect 23765 18241 23799 18275
rect 23799 18241 23808 18275
rect 23756 18232 23808 18241
rect 24216 18275 24268 18284
rect 24216 18241 24225 18275
rect 24225 18241 24259 18275
rect 24259 18241 24268 18275
rect 24216 18232 24268 18241
rect 22744 18028 22796 18080
rect 23940 18028 23992 18080
rect 24032 18071 24084 18080
rect 24032 18037 24041 18071
rect 24041 18037 24075 18071
rect 24075 18037 24084 18071
rect 24032 18028 24084 18037
rect 3917 17926 3969 17978
rect 3981 17926 4033 17978
rect 4045 17926 4097 17978
rect 4109 17926 4161 17978
rect 4173 17926 4225 17978
rect 9851 17926 9903 17978
rect 9915 17926 9967 17978
rect 9979 17926 10031 17978
rect 10043 17926 10095 17978
rect 10107 17926 10159 17978
rect 15785 17926 15837 17978
rect 15849 17926 15901 17978
rect 15913 17926 15965 17978
rect 15977 17926 16029 17978
rect 16041 17926 16093 17978
rect 21719 17926 21771 17978
rect 21783 17926 21835 17978
rect 21847 17926 21899 17978
rect 21911 17926 21963 17978
rect 21975 17926 22027 17978
rect 3332 17824 3384 17876
rect 6736 17824 6788 17876
rect 6920 17824 6972 17876
rect 10692 17824 10744 17876
rect 12900 17824 12952 17876
rect 15200 17824 15252 17876
rect 17316 17824 17368 17876
rect 18052 17824 18104 17876
rect 19340 17824 19392 17876
rect 19616 17824 19668 17876
rect 21640 17824 21692 17876
rect 22284 17824 22336 17876
rect 1860 17756 1912 17808
rect 2412 17756 2464 17808
rect 9680 17799 9732 17808
rect 9680 17765 9689 17799
rect 9689 17765 9723 17799
rect 9723 17765 9732 17799
rect 9680 17756 9732 17765
rect 2872 17731 2924 17740
rect 2872 17697 2881 17731
rect 2881 17697 2915 17731
rect 2915 17697 2924 17731
rect 2872 17688 2924 17697
rect 7656 17688 7708 17740
rect 1768 17620 1820 17672
rect 2780 17620 2832 17672
rect 5172 17620 5224 17672
rect 5816 17663 5868 17672
rect 5816 17629 5825 17663
rect 5825 17629 5859 17663
rect 5859 17629 5868 17663
rect 5816 17620 5868 17629
rect 6092 17663 6144 17672
rect 6092 17629 6099 17663
rect 6099 17629 6133 17663
rect 6133 17629 6144 17663
rect 6092 17620 6144 17629
rect 6460 17620 6512 17672
rect 9036 17663 9088 17672
rect 9036 17629 9045 17663
rect 9045 17629 9079 17663
rect 9079 17629 9088 17663
rect 9036 17620 9088 17629
rect 1584 17484 1636 17536
rect 2228 17484 2280 17536
rect 2412 17484 2464 17536
rect 2964 17484 3016 17536
rect 3516 17527 3568 17536
rect 3516 17493 3525 17527
rect 3525 17493 3559 17527
rect 3559 17493 3568 17527
rect 3516 17484 3568 17493
rect 9128 17484 9180 17536
rect 10140 17620 10192 17672
rect 10232 17663 10284 17672
rect 10232 17629 10241 17663
rect 10241 17629 10275 17663
rect 10275 17629 10284 17663
rect 10232 17620 10284 17629
rect 11704 17688 11756 17740
rect 19064 17756 19116 17808
rect 11980 17620 12032 17672
rect 12256 17663 12308 17672
rect 12256 17629 12265 17663
rect 12265 17629 12299 17663
rect 12299 17629 12308 17663
rect 12256 17620 12308 17629
rect 11520 17595 11572 17604
rect 11520 17561 11529 17595
rect 11529 17561 11563 17595
rect 11563 17561 11572 17595
rect 11520 17552 11572 17561
rect 11888 17595 11940 17604
rect 11888 17561 11897 17595
rect 11897 17561 11931 17595
rect 11931 17561 11940 17595
rect 11888 17552 11940 17561
rect 15200 17620 15252 17672
rect 17316 17620 17368 17672
rect 17960 17620 18012 17672
rect 13452 17552 13504 17604
rect 19892 17620 19944 17672
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21048 17663
rect 20996 17620 21048 17629
rect 22652 17663 22704 17672
rect 22652 17629 22661 17663
rect 22661 17629 22695 17663
rect 22695 17629 22704 17663
rect 22652 17620 22704 17629
rect 22744 17620 22796 17672
rect 12440 17484 12492 17536
rect 14648 17484 14700 17536
rect 16580 17484 16632 17536
rect 16764 17484 16816 17536
rect 17040 17484 17092 17536
rect 17132 17527 17184 17536
rect 17132 17493 17141 17527
rect 17141 17493 17175 17527
rect 17175 17493 17184 17527
rect 17132 17484 17184 17493
rect 19064 17484 19116 17536
rect 20720 17484 20772 17536
rect 22376 17527 22428 17536
rect 22376 17493 22385 17527
rect 22385 17493 22419 17527
rect 22419 17493 22428 17527
rect 22376 17484 22428 17493
rect 22560 17484 22612 17536
rect 6884 17382 6936 17434
rect 6948 17382 7000 17434
rect 7012 17382 7064 17434
rect 7076 17382 7128 17434
rect 7140 17382 7192 17434
rect 12818 17382 12870 17434
rect 12882 17382 12934 17434
rect 12946 17382 12998 17434
rect 13010 17382 13062 17434
rect 13074 17382 13126 17434
rect 18752 17382 18804 17434
rect 18816 17382 18868 17434
rect 18880 17382 18932 17434
rect 18944 17382 18996 17434
rect 19008 17382 19060 17434
rect 24686 17382 24738 17434
rect 24750 17382 24802 17434
rect 24814 17382 24866 17434
rect 24878 17382 24930 17434
rect 24942 17382 24994 17434
rect 25504 17416 25556 17468
rect 940 17280 992 17332
rect 1860 17280 1912 17332
rect 1308 17212 1360 17264
rect 6276 17280 6328 17332
rect 6552 17280 6604 17332
rect 7748 17280 7800 17332
rect 9220 17280 9272 17332
rect 3056 17212 3108 17264
rect 5908 17212 5960 17264
rect 296 17076 348 17128
rect 664 17076 716 17128
rect 2228 17187 2280 17196
rect 2228 17153 2237 17187
rect 2237 17153 2271 17187
rect 2271 17153 2280 17187
rect 2228 17144 2280 17153
rect 6736 17144 6788 17196
rect 7564 17144 7616 17196
rect 7840 17144 7892 17196
rect 1308 17008 1360 17060
rect 1768 16940 1820 16992
rect 5448 17076 5500 17128
rect 7196 17076 7248 17128
rect 7748 17076 7800 17128
rect 8852 16940 8904 16992
rect 9680 17280 9732 17332
rect 10232 17280 10284 17332
rect 11888 17280 11940 17332
rect 13544 17280 13596 17332
rect 20996 17280 21048 17332
rect 22100 17280 22152 17332
rect 23020 17280 23072 17332
rect 23756 17280 23808 17332
rect 9588 17212 9640 17264
rect 10324 17212 10376 17264
rect 9680 17144 9732 17196
rect 10968 17144 11020 17196
rect 11980 17187 12032 17196
rect 11980 17153 11987 17187
rect 11987 17153 12021 17187
rect 12021 17153 12032 17187
rect 11980 17144 12032 17153
rect 16304 17144 16356 17196
rect 17500 17212 17552 17264
rect 10692 17076 10744 17128
rect 12624 17076 12676 17128
rect 13636 17076 13688 17128
rect 9588 16940 9640 16992
rect 11980 16940 12032 16992
rect 12532 16940 12584 16992
rect 13820 16940 13872 16992
rect 14188 16983 14240 16992
rect 14188 16949 14197 16983
rect 14197 16949 14231 16983
rect 14231 16949 14240 16983
rect 14188 16940 14240 16949
rect 14372 17008 14424 17060
rect 14648 17008 14700 17060
rect 15384 16940 15436 16992
rect 16396 17008 16448 17060
rect 16120 16940 16172 16992
rect 16304 16940 16356 16992
rect 17040 16940 17092 16992
rect 18696 17144 18748 17196
rect 17500 17076 17552 17128
rect 17684 16983 17736 16992
rect 17684 16949 17693 16983
rect 17693 16949 17727 16983
rect 17727 16949 17736 16983
rect 17684 16940 17736 16949
rect 18420 16940 18472 16992
rect 19616 17212 19668 17264
rect 25504 17212 25556 17264
rect 19524 17187 19576 17196
rect 19524 17153 19533 17187
rect 19533 17153 19567 17187
rect 19567 17153 19576 17187
rect 19524 17144 19576 17153
rect 21272 17144 21324 17196
rect 22560 17144 22612 17196
rect 19708 17119 19760 17128
rect 19708 17085 19717 17119
rect 19717 17085 19751 17119
rect 19751 17085 19760 17119
rect 19708 17076 19760 17085
rect 20720 17076 20772 17128
rect 21640 17076 21692 17128
rect 22744 17008 22796 17060
rect 21548 16940 21600 16992
rect 22468 16940 22520 16992
rect 23296 16940 23348 16992
rect 23940 17076 23992 17128
rect 25044 17076 25096 17128
rect 25412 17076 25464 17128
rect 756 16804 808 16856
rect 3917 16838 3969 16890
rect 3981 16838 4033 16890
rect 4045 16838 4097 16890
rect 4109 16838 4161 16890
rect 4173 16838 4225 16890
rect 9851 16838 9903 16890
rect 9915 16838 9967 16890
rect 9979 16838 10031 16890
rect 10043 16838 10095 16890
rect 10107 16838 10159 16890
rect 15785 16838 15837 16890
rect 15849 16838 15901 16890
rect 15913 16838 15965 16890
rect 15977 16838 16029 16890
rect 16041 16838 16093 16890
rect 21719 16838 21771 16890
rect 21783 16838 21835 16890
rect 21847 16838 21899 16890
rect 21911 16838 21963 16890
rect 21975 16838 22027 16890
rect 1308 16736 1360 16788
rect 3516 16736 3568 16788
rect 8392 16736 8444 16788
rect 1676 16668 1728 16720
rect 8300 16668 8352 16720
rect 1584 16575 1636 16584
rect 1584 16541 1593 16575
rect 1593 16541 1627 16575
rect 1627 16541 1636 16575
rect 1584 16532 1636 16541
rect 3700 16600 3752 16652
rect 7196 16643 7248 16652
rect 2044 16532 2096 16584
rect 4252 16532 4304 16584
rect 7196 16609 7205 16643
rect 7205 16609 7239 16643
rect 7239 16609 7248 16643
rect 7196 16600 7248 16609
rect 9772 16600 9824 16652
rect 10324 16600 10376 16652
rect 10692 16600 10744 16652
rect 11704 16736 11756 16788
rect 12072 16736 12124 16788
rect 13452 16736 13504 16788
rect 15660 16736 15712 16788
rect 16120 16736 16172 16788
rect 5356 16532 5408 16584
rect 5448 16464 5500 16516
rect 9588 16464 9640 16516
rect 9772 16464 9824 16516
rect 10232 16464 10284 16516
rect 10876 16464 10928 16516
rect 2504 16396 2556 16448
rect 4988 16396 5040 16448
rect 7932 16396 7984 16448
rect 8392 16396 8444 16448
rect 9404 16396 9456 16448
rect 11796 16396 11848 16448
rect 13360 16600 13412 16652
rect 16028 16600 16080 16652
rect 16672 16736 16724 16788
rect 17316 16779 17368 16788
rect 17316 16745 17325 16779
rect 17325 16745 17359 16779
rect 17359 16745 17368 16779
rect 17316 16736 17368 16745
rect 17684 16736 17736 16788
rect 18328 16668 18380 16720
rect 18696 16668 18748 16720
rect 22652 16736 22704 16788
rect 22744 16736 22796 16788
rect 22376 16668 22428 16720
rect 12532 16532 12584 16584
rect 13452 16532 13504 16584
rect 14372 16575 14424 16584
rect 14372 16541 14379 16575
rect 14379 16541 14413 16575
rect 14413 16541 14424 16575
rect 14372 16532 14424 16541
rect 16396 16575 16448 16584
rect 16396 16541 16405 16575
rect 16405 16541 16439 16575
rect 16439 16541 16448 16575
rect 16396 16532 16448 16541
rect 17316 16532 17368 16584
rect 13452 16396 13504 16448
rect 13544 16396 13596 16448
rect 13636 16439 13688 16448
rect 13636 16405 13645 16439
rect 13645 16405 13679 16439
rect 13679 16405 13688 16439
rect 13636 16396 13688 16405
rect 14556 16396 14608 16448
rect 17500 16464 17552 16516
rect 19248 16532 19300 16584
rect 21272 16575 21324 16584
rect 21272 16541 21306 16575
rect 21306 16541 21324 16575
rect 21272 16532 21324 16541
rect 22468 16575 22520 16584
rect 22468 16541 22477 16575
rect 22477 16541 22511 16575
rect 22511 16541 22520 16575
rect 22468 16532 22520 16541
rect 23112 16532 23164 16584
rect 23296 16575 23348 16584
rect 23296 16541 23305 16575
rect 23305 16541 23339 16575
rect 23339 16541 23348 16575
rect 23296 16532 23348 16541
rect 23940 16643 23992 16652
rect 23940 16609 23949 16643
rect 23949 16609 23983 16643
rect 23983 16609 23992 16643
rect 23940 16600 23992 16609
rect 17868 16396 17920 16448
rect 18052 16396 18104 16448
rect 22560 16439 22612 16448
rect 22560 16405 22569 16439
rect 22569 16405 22603 16439
rect 22603 16405 22612 16439
rect 22560 16396 22612 16405
rect 23388 16396 23440 16448
rect 6884 16294 6936 16346
rect 6948 16294 7000 16346
rect 7012 16294 7064 16346
rect 7076 16294 7128 16346
rect 7140 16294 7192 16346
rect 12818 16294 12870 16346
rect 12882 16294 12934 16346
rect 12946 16294 12998 16346
rect 13010 16294 13062 16346
rect 13074 16294 13126 16346
rect 18752 16294 18804 16346
rect 18816 16294 18868 16346
rect 18880 16294 18932 16346
rect 18944 16294 18996 16346
rect 19008 16294 19060 16346
rect 24686 16294 24738 16346
rect 24750 16294 24802 16346
rect 24814 16294 24866 16346
rect 24878 16294 24930 16346
rect 24942 16294 24994 16346
rect 1584 16192 1636 16244
rect 6736 16192 6788 16244
rect 9588 16192 9640 16244
rect 11428 16192 11480 16244
rect 14096 16192 14148 16244
rect 1492 16167 1544 16176
rect 1492 16133 1501 16167
rect 1501 16133 1535 16167
rect 1535 16133 1544 16167
rect 1492 16124 1544 16133
rect 20 16056 72 16108
rect 480 16056 532 16108
rect 2320 16099 2372 16108
rect 2320 16065 2329 16099
rect 2329 16065 2363 16099
rect 2363 16065 2372 16099
rect 2320 16056 2372 16065
rect 5540 16124 5592 16176
rect 9404 16124 9456 16176
rect 2688 16099 2740 16108
rect 2688 16065 2695 16099
rect 2695 16065 2729 16099
rect 2729 16065 2740 16099
rect 2688 16056 2740 16065
rect 3700 16056 3752 16108
rect 3792 16099 3844 16108
rect 3792 16065 3801 16099
rect 3801 16065 3835 16099
rect 3835 16065 3844 16099
rect 3792 16056 3844 16065
rect 4804 16099 4856 16108
rect 4804 16065 4838 16099
rect 4838 16065 4856 16099
rect 4804 16056 4856 16065
rect 4988 16099 5040 16108
rect 4988 16065 4997 16099
rect 4997 16065 5031 16099
rect 5031 16065 5040 16099
rect 4988 16056 5040 16065
rect 1400 15852 1452 15904
rect 2136 15895 2188 15904
rect 2136 15861 2145 15895
rect 2145 15861 2179 15895
rect 2179 15861 2188 15895
rect 2136 15852 2188 15861
rect 2780 15852 2832 15904
rect 3240 15852 3292 15904
rect 4712 16031 4764 16040
rect 4712 15997 4721 16031
rect 4721 15997 4755 16031
rect 4755 15997 4764 16031
rect 5724 16056 5776 16108
rect 6552 16056 6604 16108
rect 7748 16056 7800 16108
rect 4712 15988 4764 15997
rect 7472 15988 7524 16040
rect 5632 15920 5684 15972
rect 6920 15920 6972 15972
rect 8852 16099 8904 16108
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 8208 15988 8260 16040
rect 8300 16031 8352 16040
rect 8300 15997 8309 16031
rect 8309 15997 8343 16031
rect 8343 15997 8352 16031
rect 8300 15988 8352 15997
rect 8760 15988 8812 16040
rect 4528 15852 4580 15904
rect 7196 15852 7248 15904
rect 7656 15852 7708 15904
rect 7932 15852 7984 15904
rect 8116 15852 8168 15904
rect 13360 16124 13412 16176
rect 14188 16124 14240 16176
rect 10508 16056 10560 16108
rect 11152 16099 11204 16108
rect 11152 16065 11161 16099
rect 11161 16065 11195 16099
rect 11195 16065 11204 16099
rect 11152 16056 11204 16065
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 13544 16056 13596 16108
rect 14556 16124 14608 16176
rect 14740 16167 14792 16176
rect 14740 16133 14749 16167
rect 14749 16133 14783 16167
rect 14783 16133 14792 16167
rect 14740 16124 14792 16133
rect 16948 16124 17000 16176
rect 16212 16056 16264 16108
rect 13636 15988 13688 16040
rect 18236 16192 18288 16244
rect 19800 16192 19852 16244
rect 20076 16192 20128 16244
rect 19340 16167 19392 16176
rect 19340 16133 19374 16167
rect 19374 16133 19392 16167
rect 19340 16124 19392 16133
rect 17960 16099 18012 16108
rect 17960 16065 17969 16099
rect 17969 16065 18003 16099
rect 18003 16065 18012 16099
rect 17960 16056 18012 16065
rect 18420 15988 18472 16040
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 18052 15852 18104 15904
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 20076 15988 20128 16040
rect 22284 16192 22336 16244
rect 23020 16192 23072 16244
rect 24400 16192 24452 16244
rect 23848 16056 23900 16108
rect 21640 15988 21692 16040
rect 23020 15988 23072 16040
rect 24216 15988 24268 16040
rect 19248 15852 19300 15904
rect 19984 15852 20036 15904
rect 20628 15895 20680 15904
rect 20628 15861 20637 15895
rect 20637 15861 20671 15895
rect 20671 15861 20680 15895
rect 20628 15852 20680 15861
rect 20720 15852 20772 15904
rect 21364 15852 21416 15904
rect 23112 15852 23164 15904
rect 23756 15895 23808 15904
rect 23756 15861 23765 15895
rect 23765 15861 23799 15895
rect 23799 15861 23808 15895
rect 23756 15852 23808 15861
rect 3917 15750 3969 15802
rect 3981 15750 4033 15802
rect 4045 15750 4097 15802
rect 4109 15750 4161 15802
rect 4173 15750 4225 15802
rect 9851 15750 9903 15802
rect 9915 15750 9967 15802
rect 9979 15750 10031 15802
rect 10043 15750 10095 15802
rect 10107 15750 10159 15802
rect 15785 15750 15837 15802
rect 15849 15750 15901 15802
rect 15913 15750 15965 15802
rect 15977 15750 16029 15802
rect 16041 15750 16093 15802
rect 21719 15750 21771 15802
rect 21783 15750 21835 15802
rect 21847 15750 21899 15802
rect 21911 15750 21963 15802
rect 21975 15750 22027 15802
rect 2044 15648 2096 15700
rect 4528 15648 4580 15700
rect 4620 15691 4672 15700
rect 4620 15657 4629 15691
rect 4629 15657 4663 15691
rect 4663 15657 4672 15691
rect 4620 15648 4672 15657
rect 1952 15580 2004 15632
rect 2044 15512 2096 15564
rect 2504 15580 2556 15632
rect 3424 15580 3476 15632
rect 2872 15512 2924 15564
rect 3332 15512 3384 15564
rect 5448 15580 5500 15632
rect 1952 15487 2004 15496
rect 1952 15453 1961 15487
rect 1961 15453 1995 15487
rect 1995 15453 2004 15487
rect 1952 15444 2004 15453
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 2596 15308 2648 15360
rect 5816 15512 5868 15564
rect 5264 15444 5316 15496
rect 4620 15376 4672 15428
rect 4712 15376 4764 15428
rect 5908 15487 5960 15496
rect 5908 15453 5917 15487
rect 5917 15453 5951 15487
rect 5951 15453 5960 15487
rect 5908 15444 5960 15453
rect 6000 15444 6052 15496
rect 6276 15419 6328 15428
rect 6276 15385 6285 15419
rect 6285 15385 6319 15419
rect 6319 15385 6328 15419
rect 6276 15376 6328 15385
rect 8116 15648 8168 15700
rect 9220 15648 9272 15700
rect 9588 15648 9640 15700
rect 10600 15648 10652 15700
rect 11152 15648 11204 15700
rect 17500 15648 17552 15700
rect 19340 15648 19392 15700
rect 20536 15648 20588 15700
rect 20628 15648 20680 15700
rect 21364 15648 21416 15700
rect 22560 15648 22612 15700
rect 23388 15648 23440 15700
rect 13360 15580 13412 15632
rect 6828 15512 6880 15564
rect 6920 15512 6972 15564
rect 11244 15512 11296 15564
rect 11428 15512 11480 15564
rect 7196 15444 7248 15496
rect 7380 15444 7432 15496
rect 6644 15351 6696 15360
rect 6644 15317 6653 15351
rect 6653 15317 6687 15351
rect 6687 15317 6696 15351
rect 6644 15308 6696 15317
rect 7932 15376 7984 15428
rect 9588 15487 9640 15496
rect 9588 15453 9597 15487
rect 9597 15453 9631 15487
rect 9631 15453 9640 15487
rect 9588 15444 9640 15453
rect 9772 15444 9824 15496
rect 10416 15487 10468 15496
rect 10416 15453 10450 15487
rect 10450 15453 10468 15487
rect 10416 15444 10468 15453
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 11980 15444 12032 15496
rect 12164 15444 12216 15496
rect 15200 15512 15252 15564
rect 16396 15512 16448 15564
rect 14464 15444 14516 15496
rect 14556 15444 14608 15496
rect 17316 15444 17368 15496
rect 19524 15512 19576 15564
rect 19800 15555 19852 15564
rect 19800 15521 19809 15555
rect 19809 15521 19843 15555
rect 19843 15521 19852 15555
rect 19800 15512 19852 15521
rect 7380 15308 7432 15360
rect 12072 15308 12124 15360
rect 13360 15351 13412 15360
rect 13360 15317 13369 15351
rect 13369 15317 13403 15351
rect 13403 15317 13412 15351
rect 13360 15308 13412 15317
rect 15200 15376 15252 15428
rect 15568 15376 15620 15428
rect 22652 15487 22704 15496
rect 22652 15453 22661 15487
rect 22661 15453 22695 15487
rect 22695 15453 22704 15487
rect 22652 15444 22704 15453
rect 23020 15444 23072 15496
rect 23112 15487 23164 15496
rect 23112 15453 23121 15487
rect 23121 15453 23155 15487
rect 23155 15453 23164 15487
rect 23112 15444 23164 15453
rect 23204 15487 23256 15496
rect 23204 15453 23213 15487
rect 23213 15453 23247 15487
rect 23247 15453 23256 15487
rect 23204 15444 23256 15453
rect 23572 15444 23624 15496
rect 20444 15376 20496 15428
rect 23664 15376 23716 15428
rect 15476 15308 15528 15360
rect 16672 15308 16724 15360
rect 22468 15308 22520 15360
rect 23388 15308 23440 15360
rect 23480 15351 23532 15360
rect 23480 15317 23489 15351
rect 23489 15317 23523 15351
rect 23523 15317 23532 15351
rect 23480 15308 23532 15317
rect 24124 15351 24176 15360
rect 24124 15317 24133 15351
rect 24133 15317 24167 15351
rect 24167 15317 24176 15351
rect 24124 15308 24176 15317
rect 6884 15206 6936 15258
rect 6948 15206 7000 15258
rect 7012 15206 7064 15258
rect 7076 15206 7128 15258
rect 7140 15206 7192 15258
rect 12818 15206 12870 15258
rect 12882 15206 12934 15258
rect 12946 15206 12998 15258
rect 13010 15206 13062 15258
rect 13074 15206 13126 15258
rect 18752 15206 18804 15258
rect 18816 15206 18868 15258
rect 18880 15206 18932 15258
rect 18944 15206 18996 15258
rect 19008 15206 19060 15258
rect 24686 15206 24738 15258
rect 24750 15206 24802 15258
rect 24814 15206 24866 15258
rect 24878 15206 24930 15258
rect 24942 15206 24994 15258
rect 1768 15147 1820 15156
rect 1768 15113 1777 15147
rect 1777 15113 1811 15147
rect 1811 15113 1820 15147
rect 1768 15104 1820 15113
rect 2228 15104 2280 15156
rect 2964 15104 3016 15156
rect 3700 15147 3752 15156
rect 3700 15113 3709 15147
rect 3709 15113 3743 15147
rect 3743 15113 3752 15147
rect 3700 15104 3752 15113
rect 5816 15104 5868 15156
rect 2136 15036 2188 15088
rect 3792 14968 3844 15020
rect 4528 14968 4580 15020
rect 1676 14900 1728 14952
rect 4712 14900 4764 14952
rect 6736 14943 6788 14952
rect 6736 14909 6745 14943
rect 6745 14909 6779 14943
rect 6779 14909 6788 14943
rect 6736 14900 6788 14909
rect 7656 15104 7708 15156
rect 9220 15104 9272 15156
rect 10600 15104 10652 15156
rect 11520 15104 11572 15156
rect 11980 15104 12032 15156
rect 12440 15104 12492 15156
rect 13544 15104 13596 15156
rect 14924 15104 14976 15156
rect 17408 15104 17460 15156
rect 20168 15104 20220 15156
rect 20628 15104 20680 15156
rect 23112 15104 23164 15156
rect 7748 15011 7800 15020
rect 7748 14977 7782 15011
rect 7782 14977 7800 15011
rect 10876 15036 10928 15088
rect 12072 15079 12124 15088
rect 12072 15045 12081 15079
rect 12081 15045 12115 15079
rect 12115 15045 12124 15079
rect 12072 15036 12124 15045
rect 7748 14968 7800 14977
rect 9404 14968 9456 15020
rect 7288 14900 7340 14952
rect 7380 14943 7432 14952
rect 7380 14909 7389 14943
rect 7389 14909 7423 14943
rect 7423 14909 7432 14943
rect 7380 14900 7432 14909
rect 7472 14900 7524 14952
rect 7932 14943 7984 14952
rect 7932 14909 7941 14943
rect 7941 14909 7975 14943
rect 7975 14909 7984 14943
rect 7932 14900 7984 14909
rect 3700 14832 3752 14884
rect 3976 14832 4028 14884
rect 2136 14764 2188 14816
rect 5816 14764 5868 14816
rect 9680 14764 9732 14816
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 14280 15036 14332 15088
rect 16580 15036 16632 15088
rect 11980 14968 12032 14977
rect 13176 14968 13228 15020
rect 11704 14900 11756 14952
rect 14280 14900 14332 14952
rect 14924 14900 14976 14952
rect 15200 14943 15252 14952
rect 15200 14909 15234 14943
rect 15234 14909 15252 14943
rect 15200 14900 15252 14909
rect 16212 14900 16264 14952
rect 17960 14968 18012 15020
rect 22928 15041 22980 15088
rect 18788 14968 18840 15020
rect 19248 14968 19300 15020
rect 22560 15011 22612 15020
rect 22560 14977 22569 15011
rect 22569 14977 22603 15011
rect 22603 14977 22612 15011
rect 22560 14968 22612 14977
rect 22928 15036 22953 15041
rect 22953 15036 22980 15041
rect 23020 15036 23072 15088
rect 23572 15104 23624 15156
rect 23480 15036 23532 15088
rect 21640 14900 21692 14952
rect 14832 14875 14884 14884
rect 14832 14841 14841 14875
rect 14841 14841 14875 14875
rect 14875 14841 14884 14875
rect 14832 14832 14884 14841
rect 10968 14764 11020 14816
rect 14648 14764 14700 14816
rect 14924 14764 14976 14816
rect 15200 14764 15252 14816
rect 19616 14807 19668 14816
rect 19616 14773 19625 14807
rect 19625 14773 19659 14807
rect 19659 14773 19668 14807
rect 19616 14764 19668 14773
rect 24400 14807 24452 14816
rect 24400 14773 24409 14807
rect 24409 14773 24443 14807
rect 24443 14773 24452 14807
rect 24400 14764 24452 14773
rect 3917 14662 3969 14714
rect 3981 14662 4033 14714
rect 4045 14662 4097 14714
rect 4109 14662 4161 14714
rect 4173 14662 4225 14714
rect 9851 14662 9903 14714
rect 9915 14662 9967 14714
rect 9979 14662 10031 14714
rect 10043 14662 10095 14714
rect 10107 14662 10159 14714
rect 15785 14662 15837 14714
rect 15849 14662 15901 14714
rect 15913 14662 15965 14714
rect 15977 14662 16029 14714
rect 16041 14662 16093 14714
rect 21719 14662 21771 14714
rect 21783 14662 21835 14714
rect 21847 14662 21899 14714
rect 21911 14662 21963 14714
rect 21975 14662 22027 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 1308 14492 1360 14544
rect 3424 14424 3476 14476
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 2228 14356 2280 14365
rect 1308 14288 1360 14340
rect 2504 14356 2556 14408
rect 5816 14560 5868 14612
rect 5908 14560 5960 14612
rect 7932 14560 7984 14612
rect 11704 14560 11756 14612
rect 4160 14535 4212 14544
rect 4160 14501 4169 14535
rect 4169 14501 4203 14535
rect 4203 14501 4212 14535
rect 4160 14492 4212 14501
rect 8392 14492 8444 14544
rect 10140 14492 10192 14544
rect 4712 14424 4764 14476
rect 5540 14467 5592 14476
rect 5540 14433 5549 14467
rect 5549 14433 5583 14467
rect 5583 14433 5592 14467
rect 5540 14424 5592 14433
rect 6644 14424 6696 14476
rect 6828 14424 6880 14476
rect 12716 14424 12768 14476
rect 14832 14560 14884 14612
rect 16212 14560 16264 14612
rect 18236 14560 18288 14612
rect 3792 14356 3844 14408
rect 11060 14399 11112 14408
rect 11060 14365 11067 14399
rect 11067 14365 11101 14399
rect 11101 14365 11112 14399
rect 11060 14356 11112 14365
rect 11796 14356 11848 14408
rect 2044 14263 2096 14272
rect 2044 14229 2053 14263
rect 2053 14229 2087 14263
rect 2087 14229 2096 14263
rect 2044 14220 2096 14229
rect 2964 14331 3016 14340
rect 2964 14297 2973 14331
rect 2973 14297 3007 14331
rect 3007 14297 3016 14331
rect 2964 14288 3016 14297
rect 2780 14220 2832 14272
rect 3516 14220 3568 14272
rect 4712 14288 4764 14340
rect 7840 14288 7892 14340
rect 10876 14288 10928 14340
rect 17040 14356 17092 14408
rect 19340 14492 19392 14544
rect 19800 14492 19852 14544
rect 18788 14424 18840 14476
rect 19248 14424 19300 14476
rect 20720 14467 20772 14476
rect 20720 14433 20729 14467
rect 20729 14433 20763 14467
rect 20763 14433 20772 14467
rect 20720 14424 20772 14433
rect 22560 14560 22612 14612
rect 19616 14356 19668 14408
rect 22192 14399 22244 14408
rect 22192 14365 22201 14399
rect 22201 14365 22235 14399
rect 22235 14365 22244 14399
rect 22192 14356 22244 14365
rect 5540 14220 5592 14272
rect 10232 14220 10284 14272
rect 11152 14220 11204 14272
rect 13820 14220 13872 14272
rect 14188 14220 14240 14272
rect 15844 14220 15896 14272
rect 19524 14288 19576 14340
rect 19708 14220 19760 14272
rect 20260 14220 20312 14272
rect 20904 14288 20956 14340
rect 23112 14331 23164 14340
rect 21364 14220 21416 14272
rect 23112 14297 23146 14331
rect 23146 14297 23164 14331
rect 23112 14288 23164 14297
rect 22284 14263 22336 14272
rect 22284 14229 22293 14263
rect 22293 14229 22327 14263
rect 22327 14229 22336 14263
rect 22284 14220 22336 14229
rect 23204 14220 23256 14272
rect 6884 14118 6936 14170
rect 6948 14118 7000 14170
rect 7012 14118 7064 14170
rect 7076 14118 7128 14170
rect 7140 14118 7192 14170
rect 12818 14118 12870 14170
rect 12882 14118 12934 14170
rect 12946 14118 12998 14170
rect 13010 14118 13062 14170
rect 13074 14118 13126 14170
rect 18752 14118 18804 14170
rect 18816 14118 18868 14170
rect 18880 14118 18932 14170
rect 18944 14118 18996 14170
rect 19008 14118 19060 14170
rect 24686 14118 24738 14170
rect 24750 14118 24802 14170
rect 24814 14118 24866 14170
rect 24878 14118 24930 14170
rect 24942 14118 24994 14170
rect 1400 14016 1452 14068
rect 2688 14016 2740 14068
rect 3700 14016 3752 14068
rect 1400 13880 1452 13932
rect 1860 13948 1912 14000
rect 3056 13880 3108 13932
rect 9220 14016 9272 14068
rect 9680 14016 9732 14068
rect 7380 13948 7432 14000
rect 10784 14016 10836 14068
rect 13544 14016 13596 14068
rect 6644 13880 6696 13932
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 8668 13923 8720 13932
rect 8668 13889 8675 13923
rect 8675 13889 8709 13923
rect 8709 13889 8720 13923
rect 8668 13880 8720 13889
rect 9496 13880 9548 13932
rect 10784 13880 10836 13932
rect 3792 13812 3844 13864
rect 9220 13812 9272 13864
rect 12716 13855 12768 13864
rect 12716 13821 12725 13855
rect 12725 13821 12759 13855
rect 12759 13821 12768 13855
rect 12716 13812 12768 13821
rect 1400 13676 1452 13728
rect 2320 13719 2372 13728
rect 2320 13685 2329 13719
rect 2329 13685 2363 13719
rect 2363 13685 2372 13719
rect 2320 13676 2372 13685
rect 2964 13676 3016 13728
rect 3056 13676 3108 13728
rect 3700 13719 3752 13728
rect 3700 13685 3709 13719
rect 3709 13685 3743 13719
rect 3743 13685 3752 13719
rect 3700 13676 3752 13685
rect 4988 13676 5040 13728
rect 6552 13676 6604 13728
rect 6736 13676 6788 13728
rect 13728 13719 13780 13728
rect 13728 13685 13737 13719
rect 13737 13685 13771 13719
rect 13771 13685 13780 13719
rect 13728 13676 13780 13685
rect 14372 13744 14424 13796
rect 16304 14016 16356 14068
rect 19892 14016 19944 14068
rect 22192 14016 22244 14068
rect 23480 14016 23532 14068
rect 15292 13948 15344 14000
rect 23020 13948 23072 14000
rect 15844 13880 15896 13932
rect 16304 13880 16356 13932
rect 17316 13880 17368 13932
rect 17592 13880 17644 13932
rect 18236 13880 18288 13932
rect 18696 13880 18748 13932
rect 19340 13880 19392 13932
rect 19800 13880 19852 13932
rect 19432 13855 19484 13864
rect 19432 13821 19441 13855
rect 19441 13821 19475 13855
rect 19475 13821 19484 13855
rect 19432 13812 19484 13821
rect 20904 13880 20956 13932
rect 22192 13880 22244 13932
rect 22468 13880 22520 13932
rect 23296 13880 23348 13932
rect 23572 13880 23624 13932
rect 23664 13923 23716 13932
rect 23664 13889 23673 13923
rect 23673 13889 23707 13923
rect 23707 13889 23716 13923
rect 23664 13880 23716 13889
rect 21640 13812 21692 13864
rect 15200 13744 15252 13796
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 17684 13719 17736 13728
rect 17684 13685 17693 13719
rect 17693 13685 17727 13719
rect 17727 13685 17736 13719
rect 17684 13676 17736 13685
rect 19064 13719 19116 13728
rect 19064 13685 19073 13719
rect 19073 13685 19107 13719
rect 19107 13685 19116 13719
rect 19064 13676 19116 13685
rect 20168 13676 20220 13728
rect 22928 13676 22980 13728
rect 3917 13574 3969 13626
rect 3981 13574 4033 13626
rect 4045 13574 4097 13626
rect 4109 13574 4161 13626
rect 4173 13574 4225 13626
rect 9851 13574 9903 13626
rect 9915 13574 9967 13626
rect 9979 13574 10031 13626
rect 10043 13574 10095 13626
rect 10107 13574 10159 13626
rect 15785 13574 15837 13626
rect 15849 13574 15901 13626
rect 15913 13574 15965 13626
rect 15977 13574 16029 13626
rect 16041 13574 16093 13626
rect 21719 13574 21771 13626
rect 21783 13574 21835 13626
rect 21847 13574 21899 13626
rect 21911 13574 21963 13626
rect 21975 13574 22027 13626
rect 1768 13515 1820 13524
rect 1768 13481 1777 13515
rect 1777 13481 1811 13515
rect 1811 13481 1820 13515
rect 1768 13472 1820 13481
rect 2228 13472 2280 13524
rect 1584 13336 1636 13388
rect 3240 13336 3292 13388
rect 3516 13472 3568 13524
rect 3700 13404 3752 13456
rect 4528 13336 4580 13388
rect 4712 13379 4764 13388
rect 4712 13345 4721 13379
rect 4721 13345 4755 13379
rect 4755 13345 4764 13379
rect 4712 13336 4764 13345
rect 4804 13379 4856 13388
rect 4804 13345 4838 13379
rect 4838 13345 4856 13379
rect 4804 13336 4856 13345
rect 4988 13379 5040 13388
rect 4988 13345 4997 13379
rect 4997 13345 5031 13379
rect 5031 13345 5040 13379
rect 4988 13336 5040 13345
rect 6644 13336 6696 13388
rect 2044 13268 2096 13320
rect 3056 13268 3108 13320
rect 3700 13268 3752 13320
rect 7380 13268 7432 13320
rect 8944 13472 8996 13524
rect 9680 13472 9732 13524
rect 10140 13472 10192 13524
rect 10232 13472 10284 13524
rect 10784 13515 10836 13524
rect 10784 13481 10793 13515
rect 10793 13481 10827 13515
rect 10827 13481 10836 13515
rect 10784 13472 10836 13481
rect 8576 13336 8628 13388
rect 9496 13336 9548 13388
rect 9680 13336 9732 13388
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 10784 13336 10836 13388
rect 10876 13379 10928 13388
rect 10876 13345 10885 13379
rect 10885 13345 10919 13379
rect 10919 13345 10928 13379
rect 10876 13336 10928 13345
rect 12716 13472 12768 13524
rect 15292 13472 15344 13524
rect 15568 13472 15620 13524
rect 15476 13404 15528 13456
rect 16212 13404 16264 13456
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 16580 13472 16632 13524
rect 16856 13472 16908 13524
rect 17500 13515 17552 13524
rect 17500 13481 17509 13515
rect 17509 13481 17543 13515
rect 17543 13481 17552 13515
rect 17500 13472 17552 13481
rect 17868 13472 17920 13524
rect 18236 13472 18288 13524
rect 19708 13472 19760 13524
rect 22284 13515 22336 13524
rect 22284 13481 22293 13515
rect 22293 13481 22327 13515
rect 22327 13481 22336 13515
rect 22284 13472 22336 13481
rect 17684 13336 17736 13388
rect 19064 13404 19116 13456
rect 1768 13132 1820 13184
rect 3240 13175 3292 13184
rect 3240 13141 3249 13175
rect 3249 13141 3283 13175
rect 3283 13141 3292 13175
rect 3240 13132 3292 13141
rect 7932 13200 7984 13252
rect 9864 13311 9916 13320
rect 9864 13277 9873 13311
rect 9873 13277 9907 13311
rect 9907 13277 9916 13311
rect 9864 13268 9916 13277
rect 11520 13268 11572 13320
rect 12532 13311 12584 13320
rect 12532 13277 12539 13311
rect 12539 13277 12573 13311
rect 12573 13277 12584 13311
rect 12532 13268 12584 13277
rect 9496 13132 9548 13184
rect 9864 13132 9916 13184
rect 11796 13132 11848 13184
rect 11888 13175 11940 13184
rect 11888 13141 11897 13175
rect 11897 13141 11931 13175
rect 11931 13141 11940 13175
rect 11888 13132 11940 13141
rect 12256 13200 12308 13252
rect 12624 13132 12676 13184
rect 13268 13175 13320 13184
rect 13268 13141 13277 13175
rect 13277 13141 13311 13175
rect 13311 13141 13320 13175
rect 13268 13132 13320 13141
rect 15384 13132 15436 13184
rect 16580 13311 16632 13320
rect 16580 13277 16589 13311
rect 16589 13277 16623 13311
rect 16623 13277 16632 13311
rect 16580 13268 16632 13277
rect 23204 13472 23256 13524
rect 18604 13311 18656 13320
rect 18604 13277 18613 13311
rect 18613 13277 18647 13311
rect 18647 13277 18656 13311
rect 18604 13268 18656 13277
rect 19432 13268 19484 13320
rect 20076 13311 20128 13320
rect 18420 13243 18472 13252
rect 18420 13209 18429 13243
rect 18429 13209 18463 13243
rect 18463 13209 18472 13243
rect 18420 13200 18472 13209
rect 20076 13277 20085 13311
rect 20085 13277 20119 13311
rect 20119 13277 20128 13311
rect 20076 13268 20128 13277
rect 20260 13311 20312 13320
rect 20260 13277 20269 13311
rect 20269 13277 20303 13311
rect 20303 13277 20312 13311
rect 20260 13268 20312 13277
rect 22928 13404 22980 13456
rect 22652 13336 22704 13388
rect 16396 13132 16448 13184
rect 20168 13132 20220 13184
rect 20536 13132 20588 13184
rect 22376 13132 22428 13184
rect 22468 13175 22520 13184
rect 22468 13141 22477 13175
rect 22477 13141 22511 13175
rect 22511 13141 22520 13175
rect 22468 13132 22520 13141
rect 24676 13404 24728 13456
rect 23296 13268 23348 13320
rect 25688 13268 25740 13320
rect 24032 13243 24084 13252
rect 24032 13209 24041 13243
rect 24041 13209 24075 13243
rect 24075 13209 24084 13243
rect 24032 13200 24084 13209
rect 23112 13132 23164 13184
rect 6884 13030 6936 13082
rect 6948 13030 7000 13082
rect 7012 13030 7064 13082
rect 7076 13030 7128 13082
rect 7140 13030 7192 13082
rect 12818 13030 12870 13082
rect 12882 13030 12934 13082
rect 12946 13030 12998 13082
rect 13010 13030 13062 13082
rect 13074 13030 13126 13082
rect 18752 13030 18804 13082
rect 18816 13030 18868 13082
rect 18880 13030 18932 13082
rect 18944 13030 18996 13082
rect 19008 13030 19060 13082
rect 24686 13030 24738 13082
rect 24750 13030 24802 13082
rect 24814 13030 24866 13082
rect 24878 13030 24930 13082
rect 24942 13030 24994 13082
rect 1676 12971 1728 12980
rect 1676 12937 1685 12971
rect 1685 12937 1719 12971
rect 1719 12937 1728 12971
rect 1676 12928 1728 12937
rect 2044 12928 2096 12980
rect 2688 12928 2740 12980
rect 3056 12928 3108 12980
rect 3332 12928 3384 12980
rect 3516 12928 3568 12980
rect 4528 12928 4580 12980
rect 18420 12928 18472 12980
rect 18604 12928 18656 12980
rect 19432 12971 19484 12980
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 19984 12928 20036 12980
rect 20444 12928 20496 12980
rect 22468 12928 22520 12980
rect 24492 12928 24544 12980
rect 3884 12860 3936 12912
rect 1952 12724 2004 12776
rect 2136 12724 2188 12776
rect 3056 12835 3108 12844
rect 3056 12801 3090 12835
rect 3090 12801 3108 12835
rect 3056 12792 3108 12801
rect 3976 12792 4028 12844
rect 2780 12724 2832 12776
rect 2964 12767 3016 12776
rect 2964 12733 2973 12767
rect 2973 12733 3007 12767
rect 3007 12733 3016 12767
rect 2964 12724 3016 12733
rect 2412 12656 2464 12708
rect 2688 12699 2740 12708
rect 2688 12665 2697 12699
rect 2697 12665 2731 12699
rect 2731 12665 2740 12699
rect 2688 12656 2740 12665
rect 6552 12860 6604 12912
rect 14464 12903 14516 12912
rect 14464 12869 14473 12903
rect 14473 12869 14507 12903
rect 14507 12869 14516 12903
rect 14464 12860 14516 12869
rect 14648 12860 14700 12912
rect 15384 12860 15436 12912
rect 16580 12860 16632 12912
rect 4620 12792 4672 12844
rect 9588 12835 9640 12844
rect 9588 12801 9597 12835
rect 9597 12801 9631 12835
rect 9631 12801 9640 12835
rect 9588 12792 9640 12801
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 13636 12835 13688 12844
rect 13636 12801 13670 12835
rect 13670 12801 13688 12835
rect 13636 12792 13688 12801
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 1952 12588 2004 12640
rect 3700 12588 3752 12640
rect 9496 12724 9548 12776
rect 5908 12631 5960 12640
rect 5908 12597 5917 12631
rect 5917 12597 5951 12631
rect 5951 12597 5960 12631
rect 5908 12588 5960 12597
rect 10048 12699 10100 12708
rect 10048 12665 10057 12699
rect 10057 12665 10091 12699
rect 10091 12665 10100 12699
rect 10048 12656 10100 12665
rect 6644 12588 6696 12640
rect 7104 12588 7156 12640
rect 9220 12588 9272 12640
rect 9404 12588 9456 12640
rect 10416 12767 10468 12776
rect 10416 12733 10450 12767
rect 10450 12733 10468 12767
rect 10416 12724 10468 12733
rect 10600 12767 10652 12776
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 11520 12656 11572 12708
rect 13084 12656 13136 12708
rect 11612 12588 11664 12640
rect 13268 12767 13320 12776
rect 13268 12733 13277 12767
rect 13277 12733 13311 12767
rect 13311 12733 13320 12767
rect 13268 12724 13320 12733
rect 14004 12724 14056 12776
rect 17960 12767 18012 12776
rect 17960 12733 17969 12767
rect 17969 12733 18003 12767
rect 18003 12733 18012 12767
rect 17960 12724 18012 12733
rect 20536 12792 20588 12844
rect 21180 12835 21232 12844
rect 21180 12801 21189 12835
rect 21189 12801 21223 12835
rect 21223 12801 21232 12835
rect 21180 12792 21232 12801
rect 21364 12835 21416 12844
rect 21364 12801 21373 12835
rect 21373 12801 21407 12835
rect 21407 12801 21416 12835
rect 21364 12792 21416 12801
rect 21456 12792 21508 12844
rect 22376 12792 22428 12844
rect 23480 12792 23532 12844
rect 25320 12792 25372 12844
rect 25320 12656 25372 12708
rect 25688 12656 25740 12708
rect 14556 12588 14608 12640
rect 15568 12631 15620 12640
rect 15568 12597 15577 12631
rect 15577 12597 15611 12631
rect 15611 12597 15620 12631
rect 15568 12588 15620 12597
rect 15660 12588 15712 12640
rect 17500 12588 17552 12640
rect 20996 12631 21048 12640
rect 20996 12597 21005 12631
rect 21005 12597 21039 12631
rect 21039 12597 21048 12631
rect 20996 12588 21048 12597
rect 21272 12631 21324 12640
rect 21272 12597 21281 12631
rect 21281 12597 21315 12631
rect 21315 12597 21324 12631
rect 21272 12588 21324 12597
rect 23848 12631 23900 12640
rect 23848 12597 23857 12631
rect 23857 12597 23891 12631
rect 23891 12597 23900 12631
rect 23848 12588 23900 12597
rect 3917 12486 3969 12538
rect 3981 12486 4033 12538
rect 4045 12486 4097 12538
rect 4109 12486 4161 12538
rect 4173 12486 4225 12538
rect 9851 12486 9903 12538
rect 9915 12486 9967 12538
rect 9979 12486 10031 12538
rect 10043 12486 10095 12538
rect 10107 12486 10159 12538
rect 15785 12486 15837 12538
rect 15849 12486 15901 12538
rect 15913 12486 15965 12538
rect 15977 12486 16029 12538
rect 16041 12486 16093 12538
rect 21719 12486 21771 12538
rect 21783 12486 21835 12538
rect 21847 12486 21899 12538
rect 21911 12486 21963 12538
rect 21975 12486 22027 12538
rect 1400 12427 1452 12436
rect 1400 12393 1409 12427
rect 1409 12393 1443 12427
rect 1443 12393 1452 12427
rect 1400 12384 1452 12393
rect 2688 12427 2740 12436
rect 2688 12393 2697 12427
rect 2697 12393 2731 12427
rect 2731 12393 2740 12427
rect 2688 12384 2740 12393
rect 4528 12384 4580 12436
rect 5172 12384 5224 12436
rect 5540 12384 5592 12436
rect 3608 12316 3660 12368
rect 5356 12316 5408 12368
rect 1492 12248 1544 12300
rect 2412 12248 2464 12300
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 5908 12384 5960 12436
rect 6000 12384 6052 12436
rect 6644 12316 6696 12368
rect 7012 12248 7064 12300
rect 7564 12359 7616 12368
rect 7564 12325 7573 12359
rect 7573 12325 7607 12359
rect 7607 12325 7616 12359
rect 7564 12316 7616 12325
rect 7472 12248 7524 12300
rect 1308 12112 1360 12164
rect 2320 12180 2372 12232
rect 3148 12155 3200 12164
rect 3148 12121 3157 12155
rect 3157 12121 3191 12155
rect 3191 12121 3200 12155
rect 3148 12112 3200 12121
rect 4620 12180 4672 12232
rect 5080 12180 5132 12232
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 5908 12180 5960 12189
rect 4712 12112 4764 12164
rect 3976 12087 4028 12096
rect 3976 12053 3985 12087
rect 3985 12053 4019 12087
rect 4019 12053 4028 12087
rect 3976 12044 4028 12053
rect 5172 12044 5224 12096
rect 7840 12223 7892 12232
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 9312 12248 9364 12300
rect 9496 12248 9548 12300
rect 10876 12384 10928 12436
rect 12624 12384 12676 12436
rect 13268 12384 13320 12436
rect 15660 12384 15712 12436
rect 16304 12384 16356 12436
rect 16856 12384 16908 12436
rect 17040 12359 17092 12368
rect 17040 12325 17049 12359
rect 17049 12325 17083 12359
rect 17083 12325 17092 12359
rect 17040 12316 17092 12325
rect 13084 12248 13136 12300
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 10048 12223 10100 12232
rect 10048 12189 10055 12223
rect 10055 12189 10089 12223
rect 10089 12189 10100 12223
rect 10048 12180 10100 12189
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 11980 12180 12032 12232
rect 12716 12180 12768 12232
rect 13176 12180 13228 12232
rect 9680 12112 9732 12164
rect 8208 12044 8260 12096
rect 8760 12044 8812 12096
rect 11336 12087 11388 12096
rect 11336 12053 11345 12087
rect 11345 12053 11379 12087
rect 11379 12053 11388 12087
rect 11336 12044 11388 12053
rect 14280 12248 14332 12300
rect 15384 12248 15436 12300
rect 16304 12248 16356 12300
rect 17316 12384 17368 12436
rect 18328 12316 18380 12368
rect 19248 12316 19300 12368
rect 15568 12180 15620 12232
rect 12440 12087 12492 12096
rect 12440 12053 12449 12087
rect 12449 12053 12483 12087
rect 12483 12053 12492 12087
rect 12440 12044 12492 12053
rect 13912 12112 13964 12164
rect 14464 12112 14516 12164
rect 15200 12112 15252 12164
rect 13820 12044 13872 12096
rect 14096 12044 14148 12096
rect 14648 12044 14700 12096
rect 14740 12044 14792 12096
rect 14924 12044 14976 12096
rect 18144 12248 18196 12300
rect 17500 12180 17552 12232
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 20168 12180 20220 12232
rect 20720 12384 20772 12436
rect 21180 12384 21232 12436
rect 21548 12384 21600 12436
rect 22652 12427 22704 12436
rect 22652 12393 22661 12427
rect 22661 12393 22695 12427
rect 22695 12393 22704 12427
rect 22652 12384 22704 12393
rect 20812 12291 20864 12300
rect 20812 12257 20821 12291
rect 20821 12257 20855 12291
rect 20855 12257 20864 12291
rect 20812 12248 20864 12257
rect 22008 12248 22060 12300
rect 22652 12180 22704 12232
rect 21088 12155 21140 12164
rect 21088 12121 21122 12155
rect 21122 12121 21140 12155
rect 21088 12112 21140 12121
rect 21456 12112 21508 12164
rect 21548 12112 21600 12164
rect 22928 12112 22980 12164
rect 18052 12044 18104 12096
rect 18236 12087 18288 12096
rect 18236 12053 18245 12087
rect 18245 12053 18279 12087
rect 18279 12053 18288 12087
rect 18236 12044 18288 12053
rect 22192 12087 22244 12096
rect 22192 12053 22201 12087
rect 22201 12053 22235 12087
rect 22235 12053 22244 12087
rect 22192 12044 22244 12053
rect 22468 12044 22520 12096
rect 23848 12087 23900 12096
rect 23848 12053 23857 12087
rect 23857 12053 23891 12087
rect 23891 12053 23900 12087
rect 23848 12044 23900 12053
rect 25688 12044 25740 12096
rect 6884 11942 6936 11994
rect 6948 11942 7000 11994
rect 7012 11942 7064 11994
rect 7076 11942 7128 11994
rect 7140 11942 7192 11994
rect 12818 11942 12870 11994
rect 12882 11942 12934 11994
rect 12946 11942 12998 11994
rect 13010 11942 13062 11994
rect 13074 11942 13126 11994
rect 18752 11942 18804 11994
rect 18816 11942 18868 11994
rect 18880 11942 18932 11994
rect 18944 11942 18996 11994
rect 19008 11942 19060 11994
rect 24686 11942 24738 11994
rect 24750 11942 24802 11994
rect 24814 11942 24866 11994
rect 24878 11942 24930 11994
rect 24942 11942 24994 11994
rect 1492 11840 1544 11892
rect 2136 11772 2188 11824
rect 112 11636 164 11688
rect 2872 11704 2924 11756
rect 1860 11636 1912 11688
rect 3148 11840 3200 11892
rect 5172 11840 5224 11892
rect 5264 11840 5316 11892
rect 6000 11840 6052 11892
rect 6552 11840 6604 11892
rect 4068 11704 4120 11756
rect 4344 11704 4396 11756
rect 5448 11704 5500 11756
rect 7380 11772 7432 11824
rect 7564 11840 7616 11892
rect 8116 11840 8168 11892
rect 10048 11840 10100 11892
rect 10324 11840 10376 11892
rect 10600 11840 10652 11892
rect 8760 11772 8812 11824
rect 12348 11772 12400 11824
rect 12440 11772 12492 11824
rect 13176 11772 13228 11824
rect 10968 11704 11020 11756
rect 13636 11747 13688 11756
rect 13636 11713 13643 11747
rect 13643 11713 13677 11747
rect 13677 11713 13688 11747
rect 13636 11704 13688 11713
rect 14004 11704 14056 11756
rect 2412 11500 2464 11552
rect 3056 11543 3108 11552
rect 3056 11509 3065 11543
rect 3065 11509 3099 11543
rect 3099 11509 3108 11543
rect 3056 11500 3108 11509
rect 4620 11636 4672 11688
rect 5540 11636 5592 11688
rect 4804 11568 4856 11620
rect 5080 11568 5132 11620
rect 4160 11500 4212 11552
rect 4620 11500 4672 11552
rect 9588 11636 9640 11688
rect 8944 11568 8996 11620
rect 10784 11636 10836 11688
rect 9220 11500 9272 11552
rect 13084 11568 13136 11620
rect 10784 11500 10836 11552
rect 13452 11500 13504 11552
rect 14280 11840 14332 11892
rect 16948 11840 17000 11892
rect 14464 11772 14516 11824
rect 17316 11772 17368 11824
rect 18144 11840 18196 11892
rect 18328 11840 18380 11892
rect 21364 11840 21416 11892
rect 22192 11840 22244 11892
rect 23756 11840 23808 11892
rect 23848 11840 23900 11892
rect 24400 11883 24452 11892
rect 24400 11849 24409 11883
rect 24409 11849 24443 11883
rect 24443 11849 24452 11883
rect 24400 11840 24452 11849
rect 14280 11704 14332 11756
rect 16488 11704 16540 11756
rect 17040 11704 17092 11756
rect 14648 11636 14700 11688
rect 16672 11679 16724 11688
rect 16672 11645 16681 11679
rect 16681 11645 16715 11679
rect 16715 11645 16724 11679
rect 16672 11636 16724 11645
rect 17684 11704 17736 11756
rect 21916 11772 21968 11824
rect 17500 11636 17552 11688
rect 20720 11747 20772 11756
rect 20720 11713 20729 11747
rect 20729 11713 20763 11747
rect 20763 11713 20772 11747
rect 20720 11704 20772 11713
rect 20996 11747 21048 11756
rect 20996 11713 21005 11747
rect 21005 11713 21039 11747
rect 21039 11713 21048 11747
rect 20996 11704 21048 11713
rect 21364 11747 21416 11756
rect 21364 11713 21373 11747
rect 21373 11713 21407 11747
rect 21407 11713 21416 11747
rect 21364 11704 21416 11713
rect 22836 11704 22888 11756
rect 23480 11704 23532 11756
rect 19248 11636 19300 11688
rect 22468 11636 22520 11688
rect 22652 11679 22704 11688
rect 22652 11645 22661 11679
rect 22661 11645 22695 11679
rect 22695 11645 22704 11679
rect 22652 11636 22704 11645
rect 22468 11500 22520 11552
rect 23480 11500 23532 11552
rect 23664 11543 23716 11552
rect 23664 11509 23673 11543
rect 23673 11509 23707 11543
rect 23707 11509 23716 11543
rect 23664 11500 23716 11509
rect 3917 11398 3969 11450
rect 3981 11398 4033 11450
rect 4045 11398 4097 11450
rect 4109 11398 4161 11450
rect 4173 11398 4225 11450
rect 9851 11398 9903 11450
rect 9915 11398 9967 11450
rect 9979 11398 10031 11450
rect 10043 11398 10095 11450
rect 10107 11398 10159 11450
rect 15785 11398 15837 11450
rect 15849 11398 15901 11450
rect 15913 11398 15965 11450
rect 15977 11398 16029 11450
rect 16041 11398 16093 11450
rect 21719 11398 21771 11450
rect 21783 11398 21835 11450
rect 21847 11398 21899 11450
rect 21911 11398 21963 11450
rect 21975 11398 22027 11450
rect 1768 11296 1820 11348
rect 1860 11296 1912 11348
rect 2228 11296 2280 11348
rect 756 11160 808 11212
rect 3056 11296 3108 11348
rect 4620 11296 4672 11348
rect 5816 11296 5868 11348
rect 7380 11228 7432 11280
rect 8300 11228 8352 11280
rect 10232 11296 10284 11348
rect 12440 11228 12492 11280
rect 14280 11228 14332 11280
rect 3332 11160 3384 11212
rect 4252 11160 4304 11212
rect 4804 11203 4856 11212
rect 4804 11169 4813 11203
rect 4813 11169 4847 11203
rect 4847 11169 4856 11203
rect 4804 11160 4856 11169
rect 4988 11160 5040 11212
rect 5632 11160 5684 11212
rect 6000 11160 6052 11212
rect 6644 11160 6696 11212
rect 7472 11160 7524 11212
rect 8760 11160 8812 11212
rect 10140 11160 10192 11212
rect 11152 11160 11204 11212
rect 13084 11160 13136 11212
rect 14648 11160 14700 11212
rect 15292 11160 15344 11212
rect 15844 11203 15896 11212
rect 15844 11169 15853 11203
rect 15853 11169 15887 11203
rect 15887 11169 15896 11203
rect 15844 11160 15896 11169
rect 1860 11092 1912 11144
rect 2688 11135 2740 11144
rect 2688 11101 2697 11135
rect 2697 11101 2731 11135
rect 2731 11101 2740 11135
rect 2688 11092 2740 11101
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 3884 11135 3936 11144
rect 3884 11101 3893 11135
rect 3893 11101 3927 11135
rect 3927 11101 3936 11135
rect 3884 11092 3936 11101
rect 3976 11092 4028 11144
rect 5080 11135 5132 11144
rect 5080 11101 5089 11135
rect 5089 11101 5123 11135
rect 5123 11101 5132 11135
rect 5080 11092 5132 11101
rect 6368 11092 6420 11144
rect 7656 11092 7708 11144
rect 8024 11092 8076 11144
rect 8944 11092 8996 11144
rect 1400 10999 1452 11008
rect 1400 10965 1409 10999
rect 1409 10965 1443 10999
rect 1443 10965 1452 10999
rect 1400 10956 1452 10965
rect 5632 11024 5684 11076
rect 6552 11024 6604 11076
rect 7564 11024 7616 11076
rect 15016 11092 15068 11144
rect 15200 11135 15252 11144
rect 15200 11101 15209 11135
rect 15209 11101 15243 11135
rect 15243 11101 15252 11135
rect 15200 11092 15252 11101
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 16120 11135 16172 11144
rect 16120 11101 16129 11135
rect 16129 11101 16163 11135
rect 16163 11101 16172 11135
rect 16120 11092 16172 11101
rect 22468 11296 22520 11348
rect 9496 11024 9548 11076
rect 10508 11024 10560 11076
rect 4988 10956 5040 11008
rect 12072 10956 12124 11008
rect 16948 11024 17000 11076
rect 17224 11024 17276 11076
rect 17776 11092 17828 11144
rect 18236 11024 18288 11076
rect 19248 11135 19300 11144
rect 19248 11101 19257 11135
rect 19257 11101 19291 11135
rect 19291 11101 19300 11135
rect 19248 11092 19300 11101
rect 22100 11092 22152 11144
rect 23664 11296 23716 11348
rect 22928 11092 22980 11144
rect 23020 11135 23072 11144
rect 23020 11101 23027 11135
rect 23027 11101 23061 11135
rect 23061 11101 23072 11135
rect 23020 11092 23072 11101
rect 19340 10956 19392 11008
rect 23664 10956 23716 11008
rect 6884 10854 6936 10906
rect 6948 10854 7000 10906
rect 7012 10854 7064 10906
rect 7076 10854 7128 10906
rect 7140 10854 7192 10906
rect 12818 10854 12870 10906
rect 12882 10854 12934 10906
rect 12946 10854 12998 10906
rect 13010 10854 13062 10906
rect 13074 10854 13126 10906
rect 18752 10854 18804 10906
rect 18816 10854 18868 10906
rect 18880 10854 18932 10906
rect 18944 10854 18996 10906
rect 19008 10854 19060 10906
rect 24686 10854 24738 10906
rect 24750 10854 24802 10906
rect 24814 10854 24866 10906
rect 24878 10854 24930 10906
rect 24942 10854 24994 10906
rect 2964 10752 3016 10804
rect 4988 10752 5040 10804
rect 5080 10752 5132 10804
rect 5540 10752 5592 10804
rect 5908 10752 5960 10804
rect 11796 10752 11848 10804
rect 12256 10752 12308 10804
rect 13544 10752 13596 10804
rect 2596 10616 2648 10668
rect 3976 10659 4028 10668
rect 3976 10625 3985 10659
rect 3985 10625 4019 10659
rect 4019 10625 4028 10659
rect 3976 10616 4028 10625
rect 4160 10616 4212 10668
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 6736 10616 6788 10668
rect 2412 10591 2464 10600
rect 2412 10557 2421 10591
rect 2421 10557 2455 10591
rect 2455 10557 2464 10591
rect 2412 10548 2464 10557
rect 3700 10548 3752 10600
rect 4068 10548 4120 10600
rect 6552 10591 6604 10600
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 7288 10591 7340 10600
rect 7288 10557 7297 10591
rect 7297 10557 7331 10591
rect 7331 10557 7340 10591
rect 7288 10548 7340 10557
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 10140 10684 10192 10736
rect 11336 10684 11388 10736
rect 11612 10684 11664 10736
rect 11980 10727 12032 10736
rect 11980 10693 11989 10727
rect 11989 10693 12023 10727
rect 12023 10693 12032 10727
rect 11980 10684 12032 10693
rect 12072 10727 12124 10736
rect 12072 10693 12081 10727
rect 12081 10693 12115 10727
rect 12115 10693 12124 10727
rect 12072 10684 12124 10693
rect 12716 10684 12768 10736
rect 13176 10684 13228 10736
rect 13728 10727 13780 10736
rect 13728 10693 13737 10727
rect 13737 10693 13771 10727
rect 13771 10693 13780 10727
rect 13728 10684 13780 10693
rect 14188 10752 14240 10804
rect 13912 10684 13964 10736
rect 14832 10727 14884 10736
rect 14832 10693 14841 10727
rect 14841 10693 14875 10727
rect 14875 10693 14884 10727
rect 14832 10684 14884 10693
rect 15292 10752 15344 10804
rect 15844 10752 15896 10804
rect 16672 10752 16724 10804
rect 16948 10752 17000 10804
rect 17040 10752 17092 10804
rect 14096 10659 14148 10668
rect 14096 10625 14105 10659
rect 14105 10625 14139 10659
rect 14139 10625 14148 10659
rect 14096 10616 14148 10625
rect 14464 10659 14516 10668
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 14648 10616 14700 10668
rect 17500 10684 17552 10736
rect 18052 10684 18104 10736
rect 19708 10684 19760 10736
rect 19892 10689 19944 10736
rect 15568 10616 15620 10668
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 19340 10659 19392 10668
rect 19340 10625 19349 10659
rect 19349 10625 19383 10659
rect 19383 10625 19392 10659
rect 19340 10616 19392 10625
rect 19524 10659 19576 10668
rect 19524 10625 19533 10659
rect 19533 10625 19567 10659
rect 19567 10625 19576 10659
rect 19524 10616 19576 10625
rect 19892 10684 19917 10689
rect 19917 10684 19944 10689
rect 20168 10752 20220 10804
rect 22376 10659 22428 10668
rect 22376 10625 22385 10659
rect 22385 10625 22419 10659
rect 22419 10625 22428 10659
rect 22376 10616 22428 10625
rect 22652 10659 22704 10668
rect 22652 10625 22661 10659
rect 22661 10625 22695 10659
rect 22695 10625 22704 10659
rect 22652 10616 22704 10625
rect 8116 10548 8168 10600
rect 3424 10480 3476 10532
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 2872 10412 2924 10464
rect 5540 10480 5592 10532
rect 13636 10548 13688 10600
rect 14832 10548 14884 10600
rect 22100 10548 22152 10600
rect 15292 10412 15344 10464
rect 23204 10659 23256 10668
rect 23204 10625 23213 10659
rect 23213 10625 23247 10659
rect 23247 10625 23256 10659
rect 23204 10616 23256 10625
rect 23480 10684 23532 10736
rect 23664 10684 23716 10736
rect 24492 10659 24544 10668
rect 24492 10625 24501 10659
rect 24501 10625 24535 10659
rect 24535 10625 24544 10659
rect 24492 10616 24544 10625
rect 25596 10548 25648 10600
rect 25412 10480 25464 10532
rect 20904 10412 20956 10464
rect 22836 10412 22888 10464
rect 23848 10455 23900 10464
rect 23848 10421 23857 10455
rect 23857 10421 23891 10455
rect 23891 10421 23900 10455
rect 23848 10412 23900 10421
rect 3917 10310 3969 10362
rect 3981 10310 4033 10362
rect 4045 10310 4097 10362
rect 4109 10310 4161 10362
rect 4173 10310 4225 10362
rect 9851 10310 9903 10362
rect 9915 10310 9967 10362
rect 9979 10310 10031 10362
rect 10043 10310 10095 10362
rect 10107 10310 10159 10362
rect 15785 10310 15837 10362
rect 15849 10310 15901 10362
rect 15913 10310 15965 10362
rect 15977 10310 16029 10362
rect 16041 10310 16093 10362
rect 21719 10310 21771 10362
rect 21783 10310 21835 10362
rect 21847 10310 21899 10362
rect 21911 10310 21963 10362
rect 21975 10310 22027 10362
rect 3240 10251 3292 10260
rect 3240 10217 3249 10251
rect 3249 10217 3283 10251
rect 3283 10217 3292 10251
rect 3240 10208 3292 10217
rect 1676 10183 1728 10192
rect 1676 10149 1685 10183
rect 1685 10149 1719 10183
rect 1719 10149 1728 10183
rect 1676 10140 1728 10149
rect 2780 10072 2832 10124
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 5908 10208 5960 10260
rect 6828 10208 6880 10260
rect 6920 10251 6972 10260
rect 6920 10217 6929 10251
rect 6929 10217 6963 10251
rect 6963 10217 6972 10251
rect 6920 10208 6972 10217
rect 1400 10004 1452 10056
rect 4344 10072 4396 10124
rect 2688 9936 2740 9988
rect 2964 9936 3016 9988
rect 3884 9979 3936 9988
rect 3884 9945 3893 9979
rect 3893 9945 3927 9979
rect 3927 9945 3936 9979
rect 3884 9936 3936 9945
rect 4804 10047 4856 10056
rect 4804 10013 4811 10047
rect 4811 10013 4845 10047
rect 4845 10013 4856 10047
rect 4804 10004 4856 10013
rect 5816 9936 5868 9988
rect 6276 9936 6328 9988
rect 2872 9911 2924 9920
rect 2872 9877 2881 9911
rect 2881 9877 2915 9911
rect 2915 9877 2924 9911
rect 2872 9868 2924 9877
rect 3332 9868 3384 9920
rect 5448 9868 5500 9920
rect 9128 10115 9180 10124
rect 9128 10081 9137 10115
rect 9137 10081 9171 10115
rect 9171 10081 9180 10115
rect 9128 10072 9180 10081
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 9864 10115 9916 10124
rect 9864 10081 9873 10115
rect 9873 10081 9907 10115
rect 9907 10081 9916 10115
rect 9864 10072 9916 10081
rect 12256 10208 12308 10260
rect 12440 10208 12492 10260
rect 8300 10004 8352 10056
rect 8760 10004 8812 10056
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 10876 10004 10928 10056
rect 10416 9868 10468 9920
rect 12348 10004 12400 10056
rect 13636 10251 13688 10260
rect 13636 10217 13645 10251
rect 13645 10217 13679 10251
rect 13679 10217 13688 10251
rect 13636 10208 13688 10217
rect 14096 10208 14148 10260
rect 18880 10208 18932 10260
rect 19524 10251 19576 10260
rect 19524 10217 19533 10251
rect 19533 10217 19567 10251
rect 19567 10217 19576 10251
rect 19524 10208 19576 10217
rect 22376 10251 22428 10260
rect 22376 10217 22385 10251
rect 22385 10217 22419 10251
rect 22419 10217 22428 10251
rect 22376 10208 22428 10217
rect 22652 10251 22704 10260
rect 22652 10217 22661 10251
rect 22661 10217 22695 10251
rect 22695 10217 22704 10251
rect 22652 10208 22704 10217
rect 22836 10208 22888 10260
rect 14004 10072 14056 10124
rect 14372 10047 14424 10056
rect 14372 10013 14397 10047
rect 14397 10013 14424 10047
rect 14372 10004 14424 10013
rect 16856 10004 16908 10056
rect 17408 10004 17460 10056
rect 22100 10140 22152 10192
rect 11336 9936 11388 9988
rect 11888 9868 11940 9920
rect 12072 9868 12124 9920
rect 17684 9936 17736 9988
rect 19340 9936 19392 9988
rect 19708 10047 19760 10056
rect 19708 10013 19717 10047
rect 19717 10013 19751 10047
rect 19751 10013 19760 10047
rect 19708 10004 19760 10013
rect 21180 10047 21232 10056
rect 21180 10013 21189 10047
rect 21189 10013 21232 10047
rect 21180 10004 21232 10013
rect 21732 10004 21784 10056
rect 19984 9936 20036 9988
rect 20996 9936 21048 9988
rect 21548 9936 21600 9988
rect 22928 9936 22980 9988
rect 17316 9868 17368 9920
rect 24124 9868 24176 9920
rect 6884 9766 6936 9818
rect 6948 9766 7000 9818
rect 7012 9766 7064 9818
rect 7076 9766 7128 9818
rect 7140 9766 7192 9818
rect 12818 9766 12870 9818
rect 12882 9766 12934 9818
rect 12946 9766 12998 9818
rect 13010 9766 13062 9818
rect 13074 9766 13126 9818
rect 18752 9766 18804 9818
rect 18816 9766 18868 9818
rect 18880 9766 18932 9818
rect 18944 9766 18996 9818
rect 19008 9766 19060 9818
rect 24686 9766 24738 9818
rect 24750 9766 24802 9818
rect 24814 9766 24866 9818
rect 24878 9766 24930 9818
rect 24942 9766 24994 9818
rect 1768 9707 1820 9716
rect 1768 9673 1777 9707
rect 1777 9673 1811 9707
rect 1811 9673 1820 9707
rect 1768 9664 1820 9673
rect 2320 9707 2372 9716
rect 2320 9673 2329 9707
rect 2329 9673 2363 9707
rect 2363 9673 2372 9707
rect 2320 9664 2372 9673
rect 3884 9664 3936 9716
rect 5724 9664 5776 9716
rect 6552 9664 6604 9716
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 2596 9528 2648 9580
rect 2964 9528 3016 9580
rect 3148 9639 3200 9648
rect 3148 9605 3157 9639
rect 3157 9605 3191 9639
rect 3191 9605 3200 9639
rect 3148 9596 3200 9605
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 4344 9528 4396 9580
rect 4528 9528 4580 9580
rect 6092 9596 6144 9648
rect 5172 9528 5224 9580
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 5908 9571 5960 9580
rect 5908 9537 5917 9571
rect 5917 9537 5951 9571
rect 5951 9537 5960 9571
rect 5908 9528 5960 9537
rect 9588 9664 9640 9716
rect 10140 9664 10192 9716
rect 9036 9596 9088 9648
rect 11060 9596 11112 9648
rect 11612 9596 11664 9648
rect 11980 9639 12032 9648
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 3424 9392 3476 9444
rect 7196 9460 7248 9512
rect 5816 9392 5868 9444
rect 6736 9392 6788 9444
rect 4528 9367 4580 9376
rect 4528 9333 4537 9367
rect 4537 9333 4571 9367
rect 4571 9333 4580 9367
rect 4528 9324 4580 9333
rect 4620 9324 4672 9376
rect 5724 9367 5776 9376
rect 5724 9333 5733 9367
rect 5733 9333 5767 9367
rect 5767 9333 5776 9367
rect 5724 9324 5776 9333
rect 8944 9324 8996 9376
rect 10968 9528 11020 9580
rect 11796 9528 11848 9580
rect 12256 9528 12308 9580
rect 12348 9528 12400 9580
rect 12532 9528 12584 9580
rect 12808 9639 12860 9648
rect 12808 9605 12817 9639
rect 12817 9605 12851 9639
rect 12851 9605 12860 9639
rect 12808 9596 12860 9605
rect 16672 9596 16724 9648
rect 17224 9596 17276 9648
rect 19248 9596 19300 9648
rect 19708 9664 19760 9716
rect 21272 9664 21324 9716
rect 21732 9664 21784 9716
rect 22376 9664 22428 9716
rect 23112 9664 23164 9716
rect 23204 9707 23256 9716
rect 23204 9673 23213 9707
rect 23213 9673 23247 9707
rect 23247 9673 23256 9707
rect 23204 9664 23256 9673
rect 24216 9664 24268 9716
rect 24952 9664 25004 9716
rect 23756 9596 23808 9648
rect 25044 9596 25096 9648
rect 11336 9460 11388 9512
rect 11888 9460 11940 9512
rect 17040 9528 17092 9580
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 19432 9392 19484 9444
rect 20812 9460 20864 9512
rect 21548 9460 21600 9512
rect 23572 9571 23624 9580
rect 23572 9537 23581 9571
rect 23581 9537 23615 9571
rect 23615 9537 23624 9571
rect 23572 9528 23624 9537
rect 23940 9571 23992 9580
rect 23940 9537 23949 9571
rect 23949 9537 23983 9571
rect 23983 9537 23992 9571
rect 23940 9528 23992 9537
rect 24216 9528 24268 9580
rect 17132 9324 17184 9376
rect 17684 9367 17736 9376
rect 17684 9333 17693 9367
rect 17693 9333 17727 9367
rect 17727 9333 17736 9367
rect 17684 9324 17736 9333
rect 20996 9392 21048 9444
rect 20444 9324 20496 9376
rect 21364 9324 21416 9376
rect 23112 9324 23164 9376
rect 3917 9222 3969 9274
rect 3981 9222 4033 9274
rect 4045 9222 4097 9274
rect 4109 9222 4161 9274
rect 4173 9222 4225 9274
rect 9851 9222 9903 9274
rect 9915 9222 9967 9274
rect 9979 9222 10031 9274
rect 10043 9222 10095 9274
rect 10107 9222 10159 9274
rect 15785 9222 15837 9274
rect 15849 9222 15901 9274
rect 15913 9222 15965 9274
rect 15977 9222 16029 9274
rect 16041 9222 16093 9274
rect 21719 9222 21771 9274
rect 21783 9222 21835 9274
rect 21847 9222 21899 9274
rect 21911 9222 21963 9274
rect 21975 9222 22027 9274
rect 1308 9120 1360 9172
rect 2228 9120 2280 9172
rect 2964 9120 3016 9172
rect 4344 9120 4396 9172
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 2596 9052 2648 9104
rect 3424 9052 3476 9104
rect 4160 9052 4212 9104
rect 4528 9120 4580 9172
rect 4712 9120 4764 9172
rect 7196 9120 7248 9172
rect 12164 9120 12216 9172
rect 12256 9120 12308 9172
rect 17132 9120 17184 9172
rect 7362 9095 7414 9104
rect 7362 9061 7389 9095
rect 7389 9061 7414 9095
rect 7362 9052 7414 9061
rect 8392 9052 8444 9104
rect 2596 8916 2648 8968
rect 4528 8984 4580 9036
rect 4896 8984 4948 9036
rect 6920 9027 6972 9036
rect 6920 8993 6929 9027
rect 6929 8993 6963 9027
rect 6963 8993 6972 9027
rect 6920 8984 6972 8993
rect 7656 9027 7708 9036
rect 1308 8848 1360 8900
rect 3608 8916 3660 8968
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 4988 8959 5040 8968
rect 4988 8925 4997 8959
rect 4997 8925 5031 8959
rect 5031 8925 5040 8959
rect 4988 8916 5040 8925
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 8116 8984 8168 9036
rect 8484 8984 8536 9036
rect 9772 9052 9824 9104
rect 16488 9052 16540 9104
rect 18144 9052 18196 9104
rect 17132 9027 17184 9036
rect 17132 8993 17141 9027
rect 17141 8993 17175 9027
rect 17175 8993 17184 9027
rect 17132 8984 17184 8993
rect 18328 9027 18380 9036
rect 18328 8993 18337 9027
rect 18337 8993 18371 9027
rect 18371 8993 18380 9027
rect 18328 8984 18380 8993
rect 2780 8823 2832 8832
rect 2780 8789 2789 8823
rect 2789 8789 2823 8823
rect 2823 8789 2832 8823
rect 2780 8780 2832 8789
rect 5540 8848 5592 8900
rect 6184 8848 6236 8900
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 9128 8916 9180 8968
rect 10416 8916 10468 8968
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 11888 8959 11940 8968
rect 11888 8925 11897 8959
rect 11897 8925 11931 8959
rect 11931 8925 11940 8959
rect 11888 8916 11940 8925
rect 12072 8916 12124 8968
rect 14832 8916 14884 8968
rect 15476 8916 15528 8968
rect 17408 8959 17460 8968
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 17500 8959 17552 8968
rect 17500 8925 17534 8959
rect 17534 8925 17552 8959
rect 17500 8916 17552 8925
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 3424 8780 3476 8832
rect 4712 8780 4764 8832
rect 5080 8780 5132 8832
rect 6460 8780 6512 8832
rect 7472 8780 7524 8832
rect 10232 8780 10284 8832
rect 15568 8848 15620 8900
rect 11152 8823 11204 8832
rect 11152 8789 11161 8823
rect 11161 8789 11195 8823
rect 11195 8789 11204 8823
rect 11152 8780 11204 8789
rect 12440 8780 12492 8832
rect 14096 8780 14148 8832
rect 15016 8780 15068 8832
rect 16120 8823 16172 8832
rect 16120 8789 16129 8823
rect 16129 8789 16163 8823
rect 16163 8789 16172 8823
rect 16120 8780 16172 8789
rect 20444 8916 20496 8968
rect 21640 8984 21692 9036
rect 25504 8984 25556 9036
rect 20812 8780 20864 8832
rect 21824 8959 21876 8968
rect 21824 8925 21833 8959
rect 21833 8925 21867 8959
rect 21867 8925 21876 8959
rect 21824 8916 21876 8925
rect 23296 8959 23348 8968
rect 23296 8925 23305 8959
rect 23305 8925 23339 8959
rect 23339 8925 23348 8959
rect 23296 8916 23348 8925
rect 23480 8959 23532 8968
rect 23480 8925 23489 8959
rect 23489 8925 23523 8959
rect 23523 8925 23532 8959
rect 23480 8916 23532 8925
rect 24032 8959 24084 8968
rect 24032 8925 24041 8959
rect 24041 8925 24075 8959
rect 24075 8925 24084 8959
rect 24032 8916 24084 8925
rect 23940 8848 23992 8900
rect 23204 8780 23256 8832
rect 6884 8678 6936 8730
rect 6948 8678 7000 8730
rect 7012 8678 7064 8730
rect 7076 8678 7128 8730
rect 7140 8678 7192 8730
rect 12818 8678 12870 8730
rect 12882 8678 12934 8730
rect 12946 8678 12998 8730
rect 13010 8678 13062 8730
rect 13074 8678 13126 8730
rect 18752 8678 18804 8730
rect 18816 8678 18868 8730
rect 18880 8678 18932 8730
rect 18944 8678 18996 8730
rect 19008 8678 19060 8730
rect 24686 8678 24738 8730
rect 24750 8678 24802 8730
rect 24814 8678 24866 8730
rect 24878 8678 24930 8730
rect 24942 8678 24994 8730
rect 1676 8576 1728 8628
rect 4988 8576 5040 8628
rect 5264 8576 5316 8628
rect 5540 8576 5592 8628
rect 5724 8576 5776 8628
rect 6736 8576 6788 8628
rect 7196 8576 7248 8628
rect 7288 8576 7340 8628
rect 7564 8576 7616 8628
rect 7932 8576 7984 8628
rect 10508 8619 10560 8628
rect 10508 8585 10517 8619
rect 10517 8585 10551 8619
rect 10551 8585 10560 8619
rect 10508 8576 10560 8585
rect 10600 8576 10652 8628
rect 10876 8576 10928 8628
rect 11888 8576 11940 8628
rect 1400 8508 1452 8560
rect 1676 8372 1728 8424
rect 2320 8372 2372 8424
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 2596 8372 2648 8424
rect 2780 8372 2832 8424
rect 2964 8415 3016 8424
rect 2964 8381 2973 8415
rect 2973 8381 3007 8415
rect 3007 8381 3016 8415
rect 2964 8372 3016 8381
rect 3424 8372 3476 8424
rect 6552 8440 6604 8492
rect 7656 8508 7708 8560
rect 12256 8508 12308 8560
rect 12440 8551 12492 8560
rect 12440 8517 12449 8551
rect 12449 8517 12483 8551
rect 12483 8517 12492 8551
rect 12440 8508 12492 8517
rect 7932 8440 7984 8492
rect 12348 8440 12400 8492
rect 14464 8576 14516 8628
rect 13176 8508 13228 8560
rect 13636 8508 13688 8560
rect 16580 8576 16632 8628
rect 16764 8576 16816 8628
rect 17040 8576 17092 8628
rect 17132 8576 17184 8628
rect 21824 8576 21876 8628
rect 23480 8576 23532 8628
rect 3976 8372 4028 8424
rect 4160 8236 4212 8288
rect 6644 8372 6696 8424
rect 9312 8372 9364 8424
rect 12992 8372 13044 8424
rect 14004 8440 14056 8492
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 14924 8551 14976 8560
rect 14924 8517 14933 8551
rect 14933 8517 14967 8551
rect 14967 8517 14976 8551
rect 14924 8508 14976 8517
rect 16672 8483 16724 8492
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 19432 8508 19484 8560
rect 18052 8440 18104 8492
rect 19248 8440 19300 8492
rect 21088 8440 21140 8492
rect 23664 8508 23716 8560
rect 23204 8440 23256 8492
rect 23756 8440 23808 8492
rect 5172 8304 5224 8356
rect 6092 8304 6144 8356
rect 6828 8236 6880 8288
rect 9220 8236 9272 8288
rect 9496 8236 9548 8288
rect 11060 8236 11112 8288
rect 13452 8347 13504 8356
rect 13452 8313 13461 8347
rect 13461 8313 13495 8347
rect 13495 8313 13504 8347
rect 13452 8304 13504 8313
rect 21548 8372 21600 8424
rect 16396 8304 16448 8356
rect 13636 8236 13688 8288
rect 13820 8236 13872 8288
rect 15016 8236 15068 8288
rect 21640 8304 21692 8356
rect 22100 8236 22152 8288
rect 3917 8134 3969 8186
rect 3981 8134 4033 8186
rect 4045 8134 4097 8186
rect 4109 8134 4161 8186
rect 4173 8134 4225 8186
rect 9851 8134 9903 8186
rect 9915 8134 9967 8186
rect 9979 8134 10031 8186
rect 10043 8134 10095 8186
rect 10107 8134 10159 8186
rect 15785 8134 15837 8186
rect 15849 8134 15901 8186
rect 15913 8134 15965 8186
rect 15977 8134 16029 8186
rect 16041 8134 16093 8186
rect 21719 8134 21771 8186
rect 21783 8134 21835 8186
rect 21847 8134 21899 8186
rect 21911 8134 21963 8186
rect 21975 8134 22027 8186
rect 1492 8032 1544 8084
rect 1952 8075 2004 8084
rect 1952 8041 1961 8075
rect 1961 8041 1995 8075
rect 1995 8041 2004 8075
rect 1952 8032 2004 8041
rect 2504 8032 2556 8084
rect 3240 8075 3292 8084
rect 3240 8041 3249 8075
rect 3249 8041 3283 8075
rect 3283 8041 3292 8075
rect 3240 8032 3292 8041
rect 4344 8032 4396 8084
rect 6828 8032 6880 8084
rect 7288 8007 7340 8016
rect 7288 7973 7297 8007
rect 7297 7973 7331 8007
rect 7331 7973 7340 8007
rect 7288 7964 7340 7973
rect 1216 7896 1268 7948
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 1492 7803 1544 7812
rect 1492 7769 1501 7803
rect 1501 7769 1535 7803
rect 1535 7769 1544 7803
rect 1492 7760 1544 7769
rect 3332 7828 3384 7880
rect 6000 7896 6052 7948
rect 6184 7896 6236 7948
rect 6460 7939 6512 7948
rect 6460 7905 6494 7939
rect 6494 7905 6512 7939
rect 6460 7896 6512 7905
rect 8668 7964 8720 8016
rect 9772 8032 9824 8084
rect 13452 7964 13504 8016
rect 8392 7896 8444 7948
rect 11796 7896 11848 7948
rect 16488 8032 16540 8084
rect 16120 7964 16172 8016
rect 20628 8032 20680 8084
rect 16304 7939 16356 7948
rect 16304 7905 16313 7939
rect 16313 7905 16347 7939
rect 16347 7905 16356 7939
rect 16304 7896 16356 7905
rect 16396 7939 16448 7948
rect 16396 7905 16430 7939
rect 16430 7905 16448 7939
rect 16396 7896 16448 7905
rect 5540 7828 5592 7880
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 7564 7828 7616 7880
rect 7196 7760 7248 7812
rect 9220 7871 9272 7880
rect 9220 7837 9227 7871
rect 9227 7837 9261 7871
rect 9261 7837 9272 7871
rect 9220 7828 9272 7837
rect 9312 7760 9364 7812
rect 9864 7760 9916 7812
rect 11704 7828 11756 7880
rect 15200 7828 15252 7880
rect 15476 7828 15528 7880
rect 16580 7871 16632 7880
rect 16580 7837 16589 7871
rect 16589 7837 16623 7871
rect 16623 7837 16632 7871
rect 16580 7828 16632 7837
rect 11704 7692 11756 7744
rect 12992 7760 13044 7812
rect 13912 7760 13964 7812
rect 19708 7871 19760 7880
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 19708 7828 19760 7837
rect 20168 7760 20220 7812
rect 20720 7871 20772 7880
rect 20720 7837 20729 7871
rect 20729 7837 20763 7871
rect 20763 7837 20772 7871
rect 20720 7828 20772 7837
rect 20996 8032 21048 8084
rect 23296 8075 23348 8084
rect 23296 8041 23305 8075
rect 23305 8041 23339 8075
rect 23339 8041 23348 8075
rect 23296 8032 23348 8041
rect 23480 8032 23532 8084
rect 23572 8032 23624 8084
rect 24216 7964 24268 8016
rect 22192 7828 22244 7880
rect 22560 7871 22612 7880
rect 22560 7837 22567 7871
rect 22567 7837 22601 7871
rect 22601 7837 22612 7871
rect 22560 7828 22612 7837
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 24124 7871 24176 7880
rect 24124 7837 24133 7871
rect 24133 7837 24167 7871
rect 24167 7837 24176 7871
rect 24124 7828 24176 7837
rect 24216 7760 24268 7812
rect 20536 7692 20588 7744
rect 22100 7692 22152 7744
rect 22192 7692 22244 7744
rect 22560 7692 22612 7744
rect 6884 7590 6936 7642
rect 6948 7590 7000 7642
rect 7012 7590 7064 7642
rect 7076 7590 7128 7642
rect 7140 7590 7192 7642
rect 12818 7590 12870 7642
rect 12882 7590 12934 7642
rect 12946 7590 12998 7642
rect 13010 7590 13062 7642
rect 13074 7590 13126 7642
rect 18752 7590 18804 7642
rect 18816 7590 18868 7642
rect 18880 7590 18932 7642
rect 18944 7590 18996 7642
rect 19008 7590 19060 7642
rect 24686 7590 24738 7642
rect 24750 7590 24802 7642
rect 24814 7590 24866 7642
rect 24878 7590 24930 7642
rect 24942 7590 24994 7642
rect 1308 7488 1360 7540
rect 1860 7463 1912 7472
rect 1860 7429 1869 7463
rect 1869 7429 1903 7463
rect 1903 7429 1912 7463
rect 1860 7420 1912 7429
rect 2872 7420 2924 7472
rect 4252 7488 4304 7540
rect 7288 7488 7340 7540
rect 7380 7488 7432 7540
rect 7656 7488 7708 7540
rect 9404 7531 9456 7540
rect 9404 7497 9413 7531
rect 9413 7497 9447 7531
rect 9447 7497 9456 7531
rect 9404 7488 9456 7497
rect 1952 7352 2004 7404
rect 2504 7352 2556 7404
rect 3700 7352 3752 7404
rect 7932 7420 7984 7472
rect 9864 7420 9916 7472
rect 6000 7352 6052 7404
rect 6828 7352 6880 7404
rect 7288 7352 7340 7404
rect 9680 7352 9732 7404
rect 1308 7216 1360 7268
rect 2964 7216 3016 7268
rect 3700 7216 3752 7268
rect 6092 7284 6144 7336
rect 6184 7216 6236 7268
rect 9220 7216 9272 7268
rect 10968 7352 11020 7404
rect 12532 7420 12584 7472
rect 13820 7488 13872 7540
rect 14188 7488 14240 7540
rect 16580 7488 16632 7540
rect 11888 7352 11940 7404
rect 13268 7420 13320 7472
rect 19708 7488 19760 7540
rect 20536 7488 20588 7540
rect 13452 7352 13504 7404
rect 16396 7352 16448 7404
rect 18236 7395 18288 7404
rect 18236 7361 18245 7395
rect 18245 7361 18279 7395
rect 18279 7361 18288 7395
rect 18236 7352 18288 7361
rect 18788 7352 18840 7404
rect 5080 7148 5132 7200
rect 11060 7148 11112 7200
rect 14832 7284 14884 7336
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 18328 7327 18380 7336
rect 18328 7293 18337 7327
rect 18337 7293 18371 7327
rect 18371 7293 18380 7327
rect 18328 7284 18380 7293
rect 20720 7488 20772 7540
rect 21456 7488 21508 7540
rect 23664 7531 23716 7540
rect 23664 7497 23673 7531
rect 23673 7497 23707 7531
rect 23707 7497 23716 7531
rect 23664 7488 23716 7497
rect 24032 7531 24084 7540
rect 24032 7497 24041 7531
rect 24041 7497 24075 7531
rect 24075 7497 24084 7531
rect 24032 7488 24084 7497
rect 24216 7488 24268 7540
rect 19248 7395 19300 7404
rect 19248 7361 19257 7395
rect 19257 7361 19291 7395
rect 19291 7361 19300 7395
rect 19248 7352 19300 7361
rect 22008 7420 22060 7472
rect 21088 7284 21140 7336
rect 21272 7284 21324 7336
rect 22100 7352 22152 7404
rect 14188 7148 14240 7200
rect 15292 7148 15344 7200
rect 15568 7148 15620 7200
rect 18420 7148 18472 7200
rect 22744 7395 22796 7404
rect 22744 7361 22753 7395
rect 22753 7361 22787 7395
rect 22787 7361 22796 7395
rect 22744 7352 22796 7361
rect 23204 7395 23256 7404
rect 23204 7361 23213 7395
rect 23213 7361 23247 7395
rect 23247 7361 23256 7395
rect 23204 7352 23256 7361
rect 23480 7395 23532 7404
rect 23480 7361 23489 7395
rect 23489 7361 23523 7395
rect 23523 7361 23532 7395
rect 23480 7352 23532 7361
rect 23572 7352 23624 7404
rect 23756 7352 23808 7404
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 20812 7148 20864 7200
rect 21088 7148 21140 7200
rect 22192 7148 22244 7200
rect 22284 7191 22336 7200
rect 22284 7157 22293 7191
rect 22293 7157 22327 7191
rect 22327 7157 22336 7191
rect 22284 7148 22336 7157
rect 23020 7191 23072 7200
rect 23020 7157 23029 7191
rect 23029 7157 23063 7191
rect 23063 7157 23072 7191
rect 23020 7148 23072 7157
rect 3917 7046 3969 7098
rect 3981 7046 4033 7098
rect 4045 7046 4097 7098
rect 4109 7046 4161 7098
rect 4173 7046 4225 7098
rect 9851 7046 9903 7098
rect 9915 7046 9967 7098
rect 9979 7046 10031 7098
rect 10043 7046 10095 7098
rect 10107 7046 10159 7098
rect 15785 7046 15837 7098
rect 15849 7046 15901 7098
rect 15913 7046 15965 7098
rect 15977 7046 16029 7098
rect 16041 7046 16093 7098
rect 21719 7046 21771 7098
rect 21783 7046 21835 7098
rect 21847 7046 21899 7098
rect 21911 7046 21963 7098
rect 21975 7046 22027 7098
rect 1768 6987 1820 6996
rect 1768 6953 1777 6987
rect 1777 6953 1811 6987
rect 1811 6953 1820 6987
rect 1768 6944 1820 6953
rect 1952 6944 2004 6996
rect 4712 6944 4764 6996
rect 2964 6876 3016 6928
rect 11152 6944 11204 6996
rect 6092 6876 6144 6928
rect 6644 6876 6696 6928
rect 1216 6808 1268 6860
rect 3056 6851 3108 6860
rect 3056 6817 3065 6851
rect 3065 6817 3099 6851
rect 3099 6817 3108 6851
rect 3056 6808 3108 6817
rect 3332 6808 3384 6860
rect 2136 6740 2188 6792
rect 1952 6672 2004 6724
rect 2228 6715 2280 6724
rect 2228 6681 2237 6715
rect 2237 6681 2271 6715
rect 2271 6681 2280 6715
rect 2228 6672 2280 6681
rect 2504 6672 2556 6724
rect 2780 6715 2832 6724
rect 2780 6681 2789 6715
rect 2789 6681 2823 6715
rect 2823 6681 2832 6715
rect 2780 6672 2832 6681
rect 3700 6740 3752 6792
rect 4988 6808 5040 6860
rect 6368 6808 6420 6860
rect 11060 6876 11112 6928
rect 6644 6740 6696 6792
rect 8024 6808 8076 6860
rect 10416 6808 10468 6860
rect 12532 6876 12584 6928
rect 18236 6944 18288 6996
rect 18788 6944 18840 6996
rect 19616 6944 19668 6996
rect 20168 6944 20220 6996
rect 21272 6987 21324 6996
rect 21272 6953 21281 6987
rect 21281 6953 21315 6987
rect 21315 6953 21324 6987
rect 21272 6944 21324 6953
rect 21456 6944 21508 6996
rect 21916 6944 21968 6996
rect 22468 6944 22520 6996
rect 22744 6944 22796 6996
rect 7380 6740 7432 6792
rect 7564 6740 7616 6792
rect 2044 6604 2096 6656
rect 3332 6604 3384 6656
rect 3700 6604 3752 6656
rect 4344 6647 4396 6656
rect 4344 6613 4353 6647
rect 4353 6613 4387 6647
rect 4387 6613 4396 6647
rect 4344 6604 4396 6613
rect 4620 6647 4672 6656
rect 4620 6613 4629 6647
rect 4629 6613 4663 6647
rect 4663 6613 4672 6647
rect 4620 6604 4672 6613
rect 8576 6672 8628 6724
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 11520 6783 11572 6792
rect 11520 6749 11554 6783
rect 11554 6749 11572 6783
rect 11520 6740 11572 6749
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 9404 6672 9456 6724
rect 12348 6740 12400 6792
rect 15292 6740 15344 6792
rect 15660 6740 15712 6792
rect 17868 6740 17920 6792
rect 18604 6783 18656 6792
rect 18604 6749 18613 6783
rect 18613 6749 18647 6783
rect 18647 6749 18656 6783
rect 18604 6740 18656 6749
rect 12532 6672 12584 6724
rect 13452 6672 13504 6724
rect 19156 6740 19208 6792
rect 19432 6740 19484 6792
rect 19984 6740 20036 6792
rect 24492 6876 24544 6928
rect 21548 6851 21600 6860
rect 21548 6817 21557 6851
rect 21557 6817 21591 6851
rect 21591 6817 21600 6851
rect 21548 6808 21600 6817
rect 20720 6672 20772 6724
rect 22744 6740 22796 6792
rect 21640 6672 21692 6724
rect 7380 6604 7432 6656
rect 7472 6604 7524 6656
rect 8024 6604 8076 6656
rect 8208 6647 8260 6656
rect 8208 6613 8217 6647
rect 8217 6613 8251 6647
rect 8251 6613 8260 6647
rect 8208 6604 8260 6613
rect 9036 6604 9088 6656
rect 11244 6604 11296 6656
rect 12256 6604 12308 6656
rect 12348 6647 12400 6656
rect 12348 6613 12357 6647
rect 12357 6613 12391 6647
rect 12391 6613 12400 6647
rect 12348 6604 12400 6613
rect 12440 6604 12492 6656
rect 17500 6604 17552 6656
rect 18328 6604 18380 6656
rect 21364 6604 21416 6656
rect 23572 6740 23624 6792
rect 6884 6502 6936 6554
rect 6948 6502 7000 6554
rect 7012 6502 7064 6554
rect 7076 6502 7128 6554
rect 7140 6502 7192 6554
rect 12818 6502 12870 6554
rect 12882 6502 12934 6554
rect 12946 6502 12998 6554
rect 13010 6502 13062 6554
rect 13074 6502 13126 6554
rect 18752 6502 18804 6554
rect 18816 6502 18868 6554
rect 18880 6502 18932 6554
rect 18944 6502 18996 6554
rect 19008 6502 19060 6554
rect 24686 6502 24738 6554
rect 24750 6502 24802 6554
rect 24814 6502 24866 6554
rect 24878 6502 24930 6554
rect 24942 6502 24994 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 2780 6400 2832 6452
rect 4344 6400 4396 6452
rect 5356 6400 5408 6452
rect 8944 6400 8996 6452
rect 9680 6443 9732 6452
rect 9680 6409 9689 6443
rect 9689 6409 9723 6443
rect 9723 6409 9732 6443
rect 9680 6400 9732 6409
rect 10508 6400 10560 6452
rect 1308 6264 1360 6316
rect 1860 6264 1912 6316
rect 3608 6307 3660 6316
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 3700 6264 3752 6273
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 4896 6307 4948 6316
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 8208 6264 8260 6316
rect 8852 6264 8904 6316
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 10416 6264 10468 6316
rect 15568 6400 15620 6452
rect 18604 6400 18656 6452
rect 19156 6400 19208 6452
rect 20628 6400 20680 6452
rect 21364 6400 21416 6452
rect 21456 6400 21508 6452
rect 23020 6400 23072 6452
rect 11060 6332 11112 6384
rect 11612 6264 11664 6316
rect 3516 6196 3568 6248
rect 4436 6196 4488 6248
rect 5448 6196 5500 6248
rect 7840 6239 7892 6248
rect 7840 6205 7849 6239
rect 7849 6205 7883 6239
rect 7883 6205 7892 6239
rect 7840 6196 7892 6205
rect 1860 6128 1912 6180
rect 2412 6060 2464 6112
rect 2964 6060 3016 6112
rect 4344 6171 4396 6180
rect 4344 6137 4353 6171
rect 4353 6137 4387 6171
rect 4387 6137 4396 6171
rect 4344 6128 4396 6137
rect 8300 6128 8352 6180
rect 11796 6196 11848 6248
rect 12440 6307 12492 6316
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 15292 6332 15344 6384
rect 19340 6332 19392 6384
rect 12716 6239 12768 6248
rect 12716 6205 12725 6239
rect 12725 6205 12759 6239
rect 12759 6205 12768 6239
rect 12716 6196 12768 6205
rect 11060 6128 11112 6180
rect 11152 6128 11204 6180
rect 6092 6060 6144 6112
rect 6184 6060 6236 6112
rect 6368 6060 6420 6112
rect 6644 6060 6696 6112
rect 13820 6060 13872 6112
rect 17224 6196 17276 6248
rect 16120 6128 16172 6180
rect 15660 6060 15712 6112
rect 16488 6060 16540 6112
rect 17500 6060 17552 6112
rect 20628 6307 20680 6316
rect 20628 6273 20637 6307
rect 20637 6273 20671 6307
rect 20671 6273 20680 6307
rect 20628 6264 20680 6273
rect 19064 6128 19116 6180
rect 21272 6264 21324 6316
rect 21364 6264 21416 6316
rect 22100 6264 22152 6316
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 22192 6264 22244 6273
rect 22284 6264 22336 6316
rect 23020 6264 23072 6316
rect 21548 6196 21600 6248
rect 21916 6128 21968 6180
rect 22192 6128 22244 6180
rect 22652 6171 22704 6180
rect 22652 6137 22661 6171
rect 22661 6137 22695 6171
rect 22695 6137 22704 6171
rect 22652 6128 22704 6137
rect 20720 6060 20772 6112
rect 21180 6060 21232 6112
rect 21548 6060 21600 6112
rect 23756 6060 23808 6112
rect 3917 5958 3969 6010
rect 3981 5958 4033 6010
rect 4045 5958 4097 6010
rect 4109 5958 4161 6010
rect 4173 5958 4225 6010
rect 9851 5958 9903 6010
rect 9915 5958 9967 6010
rect 9979 5958 10031 6010
rect 10043 5958 10095 6010
rect 10107 5958 10159 6010
rect 15785 5958 15837 6010
rect 15849 5958 15901 6010
rect 15913 5958 15965 6010
rect 15977 5958 16029 6010
rect 16041 5958 16093 6010
rect 21719 5958 21771 6010
rect 21783 5958 21835 6010
rect 21847 5958 21899 6010
rect 21911 5958 21963 6010
rect 21975 5958 22027 6010
rect 2228 5856 2280 5908
rect 1768 5763 1820 5772
rect 1768 5729 1777 5763
rect 1777 5729 1811 5763
rect 1811 5729 1820 5763
rect 1768 5720 1820 5729
rect 2320 5720 2372 5772
rect 2412 5763 2464 5772
rect 2412 5729 2421 5763
rect 2421 5729 2455 5763
rect 2455 5729 2464 5763
rect 2412 5720 2464 5729
rect 2780 5856 2832 5908
rect 2872 5856 2924 5908
rect 3424 5856 3476 5908
rect 3608 5899 3660 5908
rect 3608 5865 3617 5899
rect 3617 5865 3651 5899
rect 3651 5865 3660 5899
rect 3608 5856 3660 5865
rect 4896 5856 4948 5908
rect 2872 5720 2924 5772
rect 2964 5763 3016 5772
rect 2964 5729 2973 5763
rect 2973 5729 3007 5763
rect 3007 5729 3016 5763
rect 2964 5720 3016 5729
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 3700 5652 3752 5704
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 5356 5652 5408 5704
rect 3516 5584 3568 5636
rect 6092 5856 6144 5908
rect 5632 5788 5684 5840
rect 7380 5899 7432 5908
rect 7380 5865 7389 5899
rect 7389 5865 7423 5899
rect 7423 5865 7432 5899
rect 7380 5856 7432 5865
rect 7840 5856 7892 5908
rect 8852 5856 8904 5908
rect 11244 5856 11296 5908
rect 12716 5856 12768 5908
rect 13912 5856 13964 5908
rect 15660 5856 15712 5908
rect 15752 5856 15804 5908
rect 16304 5856 16356 5908
rect 6184 5763 6236 5772
rect 6184 5729 6193 5763
rect 6193 5729 6227 5763
rect 6227 5729 6236 5763
rect 6184 5720 6236 5729
rect 6552 5763 6604 5772
rect 6552 5729 6586 5763
rect 6586 5729 6604 5763
rect 6552 5720 6604 5729
rect 7380 5720 7432 5772
rect 10876 5763 10928 5772
rect 10876 5729 10885 5763
rect 10885 5729 10919 5763
rect 10919 5729 10928 5763
rect 10876 5720 10928 5729
rect 5540 5695 5592 5704
rect 5540 5661 5549 5695
rect 5549 5661 5583 5695
rect 5583 5661 5592 5695
rect 5540 5652 5592 5661
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 2320 5516 2372 5568
rect 4528 5516 4580 5568
rect 5172 5516 5224 5568
rect 8760 5652 8812 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 9312 5652 9364 5704
rect 10232 5652 10284 5704
rect 7564 5584 7616 5636
rect 10508 5584 10560 5636
rect 10140 5559 10192 5568
rect 10140 5525 10149 5559
rect 10149 5525 10183 5559
rect 10183 5525 10192 5559
rect 10140 5516 10192 5525
rect 10232 5516 10284 5568
rect 12072 5788 12124 5840
rect 12256 5763 12308 5772
rect 12256 5729 12265 5763
rect 12265 5729 12299 5763
rect 12299 5729 12308 5763
rect 12256 5720 12308 5729
rect 16304 5720 16356 5772
rect 20628 5856 20680 5908
rect 21180 5899 21232 5908
rect 21180 5865 21189 5899
rect 21189 5865 21223 5899
rect 21223 5865 21232 5899
rect 21180 5856 21232 5865
rect 21548 5899 21600 5908
rect 21548 5865 21557 5899
rect 21557 5865 21591 5899
rect 21591 5865 21600 5899
rect 21548 5856 21600 5865
rect 21640 5856 21692 5908
rect 17132 5763 17184 5772
rect 17132 5729 17141 5763
rect 17141 5729 17175 5763
rect 17175 5729 17184 5763
rect 17132 5720 17184 5729
rect 11612 5652 11664 5704
rect 11888 5652 11940 5704
rect 11060 5584 11112 5636
rect 13268 5652 13320 5704
rect 15200 5695 15252 5704
rect 15200 5661 15209 5695
rect 15209 5661 15243 5695
rect 15243 5661 15252 5695
rect 15200 5652 15252 5661
rect 15292 5652 15344 5704
rect 15568 5652 15620 5704
rect 17408 5695 17460 5704
rect 17408 5661 17415 5695
rect 17415 5661 17449 5695
rect 17449 5661 17460 5695
rect 17408 5652 17460 5661
rect 17500 5652 17552 5704
rect 21456 5788 21508 5840
rect 21732 5788 21784 5840
rect 20904 5763 20956 5772
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 20996 5720 21048 5772
rect 24216 5899 24268 5908
rect 24216 5865 24225 5899
rect 24225 5865 24259 5899
rect 24259 5865 24268 5899
rect 24216 5856 24268 5865
rect 21272 5652 21324 5704
rect 18052 5516 18104 5568
rect 19064 5516 19116 5568
rect 20812 5516 20864 5568
rect 21640 5695 21692 5704
rect 21640 5661 21649 5695
rect 21649 5661 21683 5695
rect 21683 5661 21692 5695
rect 21640 5652 21692 5661
rect 21916 5652 21968 5704
rect 22100 5695 22152 5704
rect 22100 5661 22109 5695
rect 22109 5661 22143 5695
rect 22143 5661 22152 5695
rect 22100 5652 22152 5661
rect 22560 5652 22612 5704
rect 25872 5720 25924 5772
rect 23940 5695 23992 5704
rect 23940 5661 23949 5695
rect 23949 5661 23983 5695
rect 23983 5661 23992 5695
rect 23940 5652 23992 5661
rect 25320 5652 25372 5704
rect 22928 5584 22980 5636
rect 22744 5516 22796 5568
rect 6884 5414 6936 5466
rect 6948 5414 7000 5466
rect 7012 5414 7064 5466
rect 7076 5414 7128 5466
rect 7140 5414 7192 5466
rect 12818 5414 12870 5466
rect 12882 5414 12934 5466
rect 12946 5414 12998 5466
rect 13010 5414 13062 5466
rect 13074 5414 13126 5466
rect 18752 5414 18804 5466
rect 18816 5414 18868 5466
rect 18880 5414 18932 5466
rect 18944 5414 18996 5466
rect 19008 5414 19060 5466
rect 24686 5414 24738 5466
rect 24750 5414 24802 5466
rect 24814 5414 24866 5466
rect 24878 5414 24930 5466
rect 24942 5414 24994 5466
rect 1400 5312 1452 5364
rect 2136 5355 2188 5364
rect 2136 5321 2145 5355
rect 2145 5321 2179 5355
rect 2179 5321 2188 5355
rect 2136 5312 2188 5321
rect 2596 5312 2648 5364
rect 2780 5312 2832 5364
rect 2044 5287 2096 5296
rect 2044 5253 2053 5287
rect 2053 5253 2087 5287
rect 2087 5253 2096 5287
rect 2044 5244 2096 5253
rect 4068 5312 4120 5364
rect 4344 5355 4396 5364
rect 4344 5321 4353 5355
rect 4353 5321 4387 5355
rect 4387 5321 4396 5355
rect 4344 5312 4396 5321
rect 6184 5312 6236 5364
rect 7380 5355 7432 5364
rect 7380 5321 7389 5355
rect 7389 5321 7423 5355
rect 7423 5321 7432 5355
rect 7380 5312 7432 5321
rect 7472 5312 7524 5364
rect 9588 5312 9640 5364
rect 2596 5219 2648 5228
rect 2596 5185 2605 5219
rect 2605 5185 2639 5219
rect 2639 5185 2648 5219
rect 2596 5176 2648 5185
rect 4528 5176 4580 5228
rect 4804 5176 4856 5228
rect 6276 5176 6328 5228
rect 7288 5176 7340 5228
rect 8484 5176 8536 5228
rect 9128 5176 9180 5228
rect 9496 5219 9548 5228
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 10600 5176 10652 5228
rect 4068 5108 4120 5160
rect 3056 5015 3108 5024
rect 3056 4981 3065 5015
rect 3065 4981 3099 5015
rect 3099 4981 3108 5015
rect 3056 4972 3108 4981
rect 3332 4972 3384 5024
rect 9680 5151 9732 5160
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 9680 5108 9732 5117
rect 10140 5151 10192 5160
rect 10140 5117 10149 5151
rect 10149 5117 10183 5151
rect 10183 5117 10192 5151
rect 10140 5108 10192 5117
rect 10416 5151 10468 5160
rect 8300 5040 8352 5092
rect 8668 5040 8720 5092
rect 10416 5117 10425 5151
rect 10425 5117 10459 5151
rect 10459 5117 10468 5151
rect 10416 5108 10468 5117
rect 11244 5108 11296 5160
rect 7380 4972 7432 5024
rect 13544 5312 13596 5364
rect 14556 5312 14608 5364
rect 15292 5312 15344 5364
rect 16580 5312 16632 5364
rect 20720 5312 20772 5364
rect 20904 5312 20956 5364
rect 21180 5312 21232 5364
rect 21272 5312 21324 5364
rect 12532 5249 12584 5296
rect 12532 5244 12557 5249
rect 12557 5244 12584 5249
rect 13636 5219 13688 5228
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 14832 5219 14884 5228
rect 14832 5185 14841 5219
rect 14841 5185 14875 5219
rect 14875 5185 14884 5219
rect 14832 5176 14884 5185
rect 12256 5151 12308 5160
rect 12256 5117 12265 5151
rect 12265 5117 12299 5151
rect 12299 5117 12308 5151
rect 12256 5108 12308 5117
rect 14004 5108 14056 5160
rect 14556 5151 14608 5160
rect 14556 5117 14565 5151
rect 14565 5117 14599 5151
rect 14599 5117 14608 5151
rect 14556 5108 14608 5117
rect 14648 5108 14700 5160
rect 18144 5244 18196 5296
rect 18696 5244 18748 5296
rect 17408 5176 17460 5228
rect 19800 5176 19852 5228
rect 17224 5108 17276 5160
rect 17868 5108 17920 5160
rect 19984 5040 20036 5092
rect 16948 4972 17000 5024
rect 20720 5219 20772 5228
rect 20720 5185 20729 5219
rect 20729 5185 20763 5219
rect 20763 5185 20772 5219
rect 20720 5176 20772 5185
rect 22284 5355 22336 5364
rect 22284 5321 22293 5355
rect 22293 5321 22327 5355
rect 22327 5321 22336 5355
rect 22284 5312 22336 5321
rect 22560 5355 22612 5364
rect 22560 5321 22569 5355
rect 22569 5321 22603 5355
rect 22603 5321 22612 5355
rect 22560 5312 22612 5321
rect 23664 5312 23716 5364
rect 24400 5355 24452 5364
rect 24400 5321 24409 5355
rect 24409 5321 24443 5355
rect 24443 5321 24452 5355
rect 24400 5312 24452 5321
rect 20812 5108 20864 5160
rect 21548 5108 21600 5160
rect 22284 5176 22336 5228
rect 22468 5176 22520 5228
rect 22928 5176 22980 5228
rect 23112 5219 23164 5228
rect 23112 5185 23121 5219
rect 23121 5185 23155 5219
rect 23155 5185 23164 5219
rect 23112 5176 23164 5185
rect 23756 5287 23808 5296
rect 23756 5253 23765 5287
rect 23765 5253 23799 5287
rect 23799 5253 23808 5287
rect 23756 5244 23808 5253
rect 24032 5219 24084 5228
rect 24032 5185 24041 5219
rect 24041 5185 24075 5219
rect 24075 5185 24084 5219
rect 24032 5176 24084 5185
rect 25044 5176 25096 5228
rect 24216 5108 24268 5160
rect 23388 5040 23440 5092
rect 23480 5083 23532 5092
rect 23480 5049 23489 5083
rect 23489 5049 23523 5083
rect 23523 5049 23532 5083
rect 23480 5040 23532 5049
rect 22928 5015 22980 5024
rect 22928 4981 22937 5015
rect 22937 4981 22971 5015
rect 22971 4981 22980 5015
rect 22928 4972 22980 4981
rect 24124 4972 24176 5024
rect 3917 4870 3969 4922
rect 3981 4870 4033 4922
rect 4045 4870 4097 4922
rect 4109 4870 4161 4922
rect 4173 4870 4225 4922
rect 9851 4870 9903 4922
rect 9915 4870 9967 4922
rect 9979 4870 10031 4922
rect 10043 4870 10095 4922
rect 10107 4870 10159 4922
rect 15785 4870 15837 4922
rect 15849 4870 15901 4922
rect 15913 4870 15965 4922
rect 15977 4870 16029 4922
rect 16041 4870 16093 4922
rect 21719 4870 21771 4922
rect 21783 4870 21835 4922
rect 21847 4870 21899 4922
rect 21911 4870 21963 4922
rect 21975 4870 22027 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 2596 4768 2648 4820
rect 2688 4768 2740 4820
rect 3056 4768 3108 4820
rect 4712 4811 4764 4820
rect 4712 4777 4721 4811
rect 4721 4777 4755 4811
rect 4755 4777 4764 4811
rect 4712 4768 4764 4777
rect 8300 4768 8352 4820
rect 9680 4768 9732 4820
rect 1952 4632 2004 4684
rect 9128 4700 9180 4752
rect 10048 4700 10100 4752
rect 11152 4811 11204 4820
rect 11152 4777 11161 4811
rect 11161 4777 11195 4811
rect 11195 4777 11204 4811
rect 11152 4768 11204 4777
rect 12716 4768 12768 4820
rect 12348 4700 12400 4752
rect 14832 4768 14884 4820
rect 2320 4564 2372 4616
rect 2872 4564 2924 4616
rect 3424 4564 3476 4616
rect 7380 4632 7432 4684
rect 8484 4632 8536 4684
rect 10140 4675 10192 4684
rect 10140 4641 10149 4675
rect 10149 4641 10183 4675
rect 10183 4641 10192 4675
rect 10140 4632 10192 4641
rect 11612 4675 11664 4684
rect 11612 4641 11621 4675
rect 11621 4641 11655 4675
rect 11655 4641 11664 4675
rect 11612 4632 11664 4641
rect 16948 4700 17000 4752
rect 14832 4632 14884 4684
rect 5172 4564 5224 4616
rect 7288 4564 7340 4616
rect 1124 4428 1176 4480
rect 3332 4471 3384 4480
rect 3332 4437 3341 4471
rect 3341 4437 3375 4471
rect 3375 4437 3384 4471
rect 3332 4428 3384 4437
rect 4068 4428 4120 4480
rect 7472 4428 7524 4480
rect 9772 4564 9824 4616
rect 10324 4564 10376 4616
rect 10508 4564 10560 4616
rect 12532 4564 12584 4616
rect 14372 4607 14424 4616
rect 14372 4573 14379 4607
rect 14379 4573 14413 4607
rect 14413 4573 14424 4607
rect 14372 4564 14424 4573
rect 17224 4607 17276 4616
rect 17224 4573 17233 4607
rect 17233 4573 17267 4607
rect 17267 4573 17276 4607
rect 17224 4564 17276 4573
rect 8760 4428 8812 4480
rect 8852 4428 8904 4480
rect 12348 4428 12400 4480
rect 12716 4428 12768 4480
rect 17316 4428 17368 4480
rect 18236 4471 18288 4480
rect 18236 4437 18245 4471
rect 18245 4437 18279 4471
rect 18279 4437 18288 4471
rect 18236 4428 18288 4437
rect 18696 4811 18748 4820
rect 18696 4777 18705 4811
rect 18705 4777 18739 4811
rect 18739 4777 18748 4811
rect 18696 4768 18748 4777
rect 19708 4768 19760 4820
rect 19800 4811 19852 4820
rect 19800 4777 19809 4811
rect 19809 4777 19843 4811
rect 19843 4777 19852 4811
rect 19800 4768 19852 4777
rect 20720 4768 20772 4820
rect 21548 4768 21600 4820
rect 22376 4768 22428 4820
rect 25412 4768 25464 4820
rect 20168 4700 20220 4752
rect 20536 4675 20588 4684
rect 20536 4641 20545 4675
rect 20545 4641 20579 4675
rect 20579 4641 20588 4675
rect 20536 4632 20588 4641
rect 18696 4564 18748 4616
rect 19340 4564 19392 4616
rect 19616 4607 19668 4616
rect 19616 4573 19625 4607
rect 19625 4573 19659 4607
rect 19659 4573 19668 4607
rect 19616 4564 19668 4573
rect 19524 4496 19576 4548
rect 19984 4607 20036 4616
rect 19984 4573 19993 4607
rect 19993 4573 20027 4607
rect 20027 4573 20036 4607
rect 19984 4564 20036 4573
rect 20168 4607 20220 4616
rect 20168 4573 20177 4607
rect 20177 4573 20211 4607
rect 20211 4573 20220 4607
rect 20168 4564 20220 4573
rect 20444 4607 20496 4616
rect 20444 4573 20453 4607
rect 20453 4573 20487 4607
rect 20487 4573 20496 4607
rect 22928 4632 22980 4684
rect 23204 4675 23256 4684
rect 23204 4641 23213 4675
rect 23213 4641 23247 4675
rect 23247 4641 23256 4675
rect 23204 4632 23256 4641
rect 20444 4564 20496 4573
rect 20168 4428 20220 4480
rect 20996 4496 21048 4548
rect 21088 4496 21140 4548
rect 22560 4564 22612 4616
rect 22652 4607 22704 4616
rect 22652 4573 22661 4607
rect 22661 4573 22695 4607
rect 22695 4573 22704 4607
rect 22652 4564 22704 4573
rect 23664 4496 23716 4548
rect 20536 4428 20588 4480
rect 6884 4326 6936 4378
rect 6948 4326 7000 4378
rect 7012 4326 7064 4378
rect 7076 4326 7128 4378
rect 7140 4326 7192 4378
rect 12818 4326 12870 4378
rect 12882 4326 12934 4378
rect 12946 4326 12998 4378
rect 13010 4326 13062 4378
rect 13074 4326 13126 4378
rect 18752 4326 18804 4378
rect 18816 4326 18868 4378
rect 18880 4326 18932 4378
rect 18944 4326 18996 4378
rect 19008 4326 19060 4378
rect 24686 4326 24738 4378
rect 24750 4326 24802 4378
rect 24814 4326 24866 4378
rect 24878 4326 24930 4378
rect 24942 4326 24994 4378
rect 1584 4267 1636 4276
rect 1584 4233 1593 4267
rect 1593 4233 1627 4267
rect 1627 4233 1636 4267
rect 1584 4224 1636 4233
rect 3332 4224 3384 4276
rect 3700 4224 3752 4276
rect 5172 4267 5224 4276
rect 5172 4233 5181 4267
rect 5181 4233 5215 4267
rect 5215 4233 5224 4267
rect 5172 4224 5224 4233
rect 9404 4267 9456 4276
rect 9404 4233 9413 4267
rect 9413 4233 9447 4267
rect 9447 4233 9456 4267
rect 9404 4224 9456 4233
rect 1860 4088 1912 4140
rect 2596 4088 2648 4140
rect 3240 4088 3292 4140
rect 3516 4131 3568 4140
rect 3516 4097 3525 4131
rect 3525 4097 3559 4131
rect 3559 4097 3568 4131
rect 3516 4088 3568 4097
rect 4436 4088 4488 4140
rect 8760 4131 8812 4140
rect 8760 4097 8769 4131
rect 8769 4097 8803 4131
rect 8803 4097 8812 4131
rect 8760 4088 8812 4097
rect 12164 4267 12216 4276
rect 12164 4233 12173 4267
rect 12173 4233 12207 4267
rect 12207 4233 12216 4267
rect 12164 4224 12216 4233
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 12532 4199 12584 4208
rect 12532 4165 12541 4199
rect 12541 4165 12575 4199
rect 12575 4165 12584 4199
rect 12532 4156 12584 4165
rect 13636 4156 13688 4208
rect 12624 4088 12676 4140
rect 15200 4224 15252 4276
rect 15016 4088 15068 4140
rect 15660 4131 15712 4140
rect 15660 4097 15694 4131
rect 15694 4097 15712 4131
rect 15660 4088 15712 4097
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 5540 3995 5592 4004
rect 5540 3961 5549 3995
rect 5549 3961 5583 3995
rect 5583 3961 5592 3995
rect 5540 3952 5592 3961
rect 7840 4020 7892 4072
rect 8116 3952 8168 4004
rect 8208 3995 8260 4004
rect 8208 3961 8217 3995
rect 8217 3961 8251 3995
rect 8251 3961 8260 3995
rect 8208 3952 8260 3961
rect 5264 3884 5316 3936
rect 6644 3884 6696 3936
rect 8668 4020 8720 4072
rect 10968 4020 11020 4072
rect 12348 4020 12400 4072
rect 14556 4020 14608 4072
rect 9772 3952 9824 4004
rect 11612 3952 11664 4004
rect 13912 3995 13964 4004
rect 13912 3961 13921 3995
rect 13921 3961 13955 3995
rect 13955 3961 13964 3995
rect 15568 4063 15620 4072
rect 15568 4029 15577 4063
rect 15577 4029 15611 4063
rect 15611 4029 15620 4063
rect 15568 4020 15620 4029
rect 17040 4020 17092 4072
rect 18236 4156 18288 4208
rect 13912 3952 13964 3961
rect 15384 3952 15436 4004
rect 18144 4020 18196 4072
rect 18512 4131 18564 4140
rect 18512 4097 18521 4131
rect 18521 4097 18555 4131
rect 18555 4097 18564 4131
rect 19340 4224 19392 4276
rect 19616 4224 19668 4276
rect 20444 4156 20496 4208
rect 24400 4224 24452 4276
rect 18512 4088 18564 4097
rect 19800 4088 19852 4140
rect 21548 4088 21600 4140
rect 20444 4020 20496 4072
rect 22100 4131 22152 4140
rect 22100 4097 22107 4131
rect 22107 4097 22141 4131
rect 22141 4097 22152 4131
rect 22100 4088 22152 4097
rect 25688 4088 25740 4140
rect 24216 4020 24268 4072
rect 20168 3952 20220 4004
rect 8576 3884 8628 3936
rect 9496 3884 9548 3936
rect 12072 3884 12124 3936
rect 14464 3884 14516 3936
rect 18328 3884 18380 3936
rect 18880 3927 18932 3936
rect 18880 3893 18889 3927
rect 18889 3893 18923 3927
rect 18923 3893 18932 3927
rect 18880 3884 18932 3893
rect 19156 3884 19208 3936
rect 20996 3884 21048 3936
rect 21180 3884 21232 3936
rect 21456 3884 21508 3936
rect 22284 3884 22336 3936
rect 3917 3782 3969 3834
rect 3981 3782 4033 3834
rect 4045 3782 4097 3834
rect 4109 3782 4161 3834
rect 4173 3782 4225 3834
rect 9851 3782 9903 3834
rect 9915 3782 9967 3834
rect 9979 3782 10031 3834
rect 10043 3782 10095 3834
rect 10107 3782 10159 3834
rect 15785 3782 15837 3834
rect 15849 3782 15901 3834
rect 15913 3782 15965 3834
rect 15977 3782 16029 3834
rect 16041 3782 16093 3834
rect 21719 3782 21771 3834
rect 21783 3782 21835 3834
rect 21847 3782 21899 3834
rect 21911 3782 21963 3834
rect 21975 3782 22027 3834
rect 1492 3680 1544 3732
rect 2412 3680 2464 3732
rect 4528 3680 4580 3732
rect 5172 3680 5224 3732
rect 5908 3680 5960 3732
rect 8208 3680 8260 3732
rect 8300 3680 8352 3732
rect 14464 3680 14516 3732
rect 7288 3544 7340 3596
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 1860 3476 1912 3528
rect 2964 3476 3016 3528
rect 6736 3476 6788 3528
rect 9772 3587 9824 3596
rect 9772 3553 9781 3587
rect 9781 3553 9815 3587
rect 9815 3553 9824 3587
rect 9772 3544 9824 3553
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 9496 3476 9548 3528
rect 11060 3476 11112 3528
rect 11152 3476 11204 3528
rect 13268 3612 13320 3664
rect 13912 3612 13964 3664
rect 12716 3544 12768 3596
rect 11980 3476 12032 3528
rect 15384 3680 15436 3732
rect 16120 3680 16172 3732
rect 17040 3723 17092 3732
rect 17040 3689 17049 3723
rect 17049 3689 17083 3723
rect 17083 3689 17092 3723
rect 17040 3680 17092 3689
rect 18328 3723 18380 3732
rect 18328 3689 18337 3723
rect 18337 3689 18371 3723
rect 18371 3689 18380 3723
rect 18328 3680 18380 3689
rect 14924 3519 14976 3528
rect 14924 3485 14931 3519
rect 14931 3485 14965 3519
rect 14965 3485 14976 3519
rect 14924 3476 14976 3485
rect 8392 3408 8444 3460
rect 8576 3408 8628 3460
rect 8760 3340 8812 3392
rect 8944 3383 8996 3392
rect 8944 3349 8953 3383
rect 8953 3349 8987 3383
rect 8987 3349 8996 3383
rect 8944 3340 8996 3349
rect 10232 3340 10284 3392
rect 11520 3383 11572 3392
rect 11520 3349 11529 3383
rect 11529 3349 11563 3383
rect 11563 3349 11572 3383
rect 11520 3340 11572 3349
rect 11796 3408 11848 3460
rect 15568 3408 15620 3460
rect 13452 3340 13504 3392
rect 13820 3340 13872 3392
rect 13912 3340 13964 3392
rect 16396 3476 16448 3528
rect 17592 3476 17644 3528
rect 18144 3544 18196 3596
rect 18880 3544 18932 3596
rect 17132 3408 17184 3460
rect 17500 3383 17552 3392
rect 17500 3349 17509 3383
rect 17509 3349 17543 3383
rect 17543 3349 17552 3383
rect 17500 3340 17552 3349
rect 17868 3451 17920 3460
rect 17868 3417 17877 3451
rect 17877 3417 17911 3451
rect 17911 3417 17920 3451
rect 17868 3408 17920 3417
rect 18236 3519 18288 3528
rect 18236 3485 18245 3519
rect 18245 3485 18279 3519
rect 18279 3485 18288 3519
rect 18236 3476 18288 3485
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 19248 3476 19300 3528
rect 19892 3544 19944 3596
rect 20168 3544 20220 3596
rect 22468 3680 22520 3732
rect 25596 3680 25648 3732
rect 21364 3612 21416 3664
rect 22652 3612 22704 3664
rect 23572 3612 23624 3664
rect 20720 3544 20772 3596
rect 22284 3544 22336 3596
rect 23020 3587 23072 3596
rect 23020 3553 23029 3587
rect 23029 3553 23063 3587
rect 23063 3553 23072 3587
rect 23020 3544 23072 3553
rect 19708 3451 19760 3460
rect 19708 3417 19717 3451
rect 19717 3417 19751 3451
rect 19751 3417 19760 3451
rect 19708 3408 19760 3417
rect 19892 3408 19944 3460
rect 18604 3340 18656 3392
rect 19248 3383 19300 3392
rect 19248 3349 19257 3383
rect 19257 3349 19291 3383
rect 19291 3349 19300 3383
rect 19248 3340 19300 3349
rect 19524 3340 19576 3392
rect 20168 3340 20220 3392
rect 20996 3408 21048 3460
rect 21640 3519 21692 3528
rect 21640 3485 21649 3519
rect 21649 3485 21683 3519
rect 21683 3485 21692 3519
rect 21640 3476 21692 3485
rect 22100 3519 22152 3528
rect 22100 3485 22109 3519
rect 22109 3485 22143 3519
rect 22143 3485 22152 3519
rect 22100 3476 22152 3485
rect 22652 3519 22704 3528
rect 22652 3485 22661 3519
rect 22661 3485 22695 3519
rect 22695 3485 22704 3519
rect 22652 3476 22704 3485
rect 23112 3476 23164 3528
rect 6884 3238 6936 3290
rect 6948 3238 7000 3290
rect 7012 3238 7064 3290
rect 7076 3238 7128 3290
rect 7140 3238 7192 3290
rect 12818 3238 12870 3290
rect 12882 3238 12934 3290
rect 12946 3238 12998 3290
rect 13010 3238 13062 3290
rect 13074 3238 13126 3290
rect 18752 3238 18804 3290
rect 18816 3238 18868 3290
rect 18880 3238 18932 3290
rect 18944 3238 18996 3290
rect 19008 3238 19060 3290
rect 24686 3238 24738 3290
rect 24750 3238 24802 3290
rect 24814 3238 24866 3290
rect 24878 3238 24930 3290
rect 24942 3238 24994 3290
rect 1584 3136 1636 3188
rect 11152 3136 11204 3188
rect 11520 3136 11572 3188
rect 12532 3136 12584 3188
rect 14372 3136 14424 3188
rect 1952 3068 2004 3120
rect 4344 3068 4396 3120
rect 4436 3111 4488 3120
rect 4436 3077 4445 3111
rect 4445 3077 4479 3111
rect 4479 3077 4488 3111
rect 4436 3068 4488 3077
rect 6184 3068 6236 3120
rect 572 2932 624 2984
rect 4620 2975 4672 2984
rect 4620 2941 4629 2975
rect 4629 2941 4663 2975
rect 4663 2941 4672 2975
rect 4620 2932 4672 2941
rect 4896 2975 4948 2984
rect 4896 2941 4905 2975
rect 4905 2941 4939 2975
rect 4939 2941 4948 2975
rect 4896 2932 4948 2941
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 10140 3111 10192 3120
rect 10140 3077 10149 3111
rect 10149 3077 10183 3111
rect 10183 3077 10192 3111
rect 10140 3068 10192 3077
rect 10232 3111 10284 3120
rect 10232 3077 10241 3111
rect 10241 3077 10275 3111
rect 10275 3077 10284 3111
rect 10232 3068 10284 3077
rect 10416 3068 10468 3120
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 8668 3000 8720 3052
rect 8760 3043 8812 3052
rect 8760 3009 8769 3043
rect 8769 3009 8803 3043
rect 8803 3009 8812 3043
rect 8760 3000 8812 3009
rect 9404 3000 9456 3052
rect 11612 3068 11664 3120
rect 6552 2864 6604 2916
rect 5356 2796 5408 2848
rect 6460 2839 6512 2848
rect 6460 2805 6469 2839
rect 6469 2805 6503 2839
rect 6503 2805 6512 2839
rect 6460 2796 6512 2805
rect 6736 2839 6788 2848
rect 6736 2805 6745 2839
rect 6745 2805 6779 2839
rect 6779 2805 6788 2839
rect 6736 2796 6788 2805
rect 7288 2839 7340 2848
rect 7288 2805 7297 2839
rect 7297 2805 7331 2839
rect 7331 2805 7340 2839
rect 7288 2796 7340 2805
rect 7656 2932 7708 2984
rect 7840 2932 7892 2984
rect 8116 2932 8168 2984
rect 10232 2932 10284 2984
rect 10968 2932 11020 2984
rect 12072 3068 12124 3120
rect 12164 3043 12216 3052
rect 12164 3009 12173 3043
rect 12173 3009 12207 3043
rect 12207 3009 12216 3043
rect 12164 3000 12216 3009
rect 12900 3000 12952 3052
rect 13728 3000 13780 3052
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 17040 3068 17092 3120
rect 18512 3136 18564 3188
rect 19340 3136 19392 3188
rect 19432 3179 19484 3188
rect 19432 3145 19441 3179
rect 19441 3145 19475 3179
rect 19475 3145 19484 3179
rect 19432 3136 19484 3145
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 18236 3068 18288 3120
rect 8208 2907 8260 2916
rect 8208 2873 8217 2907
rect 8217 2873 8251 2907
rect 8251 2873 8260 2907
rect 8208 2864 8260 2873
rect 9312 2864 9364 2916
rect 11060 2864 11112 2916
rect 17684 3043 17736 3052
rect 17684 3009 17693 3043
rect 17693 3009 17727 3043
rect 17727 3009 17736 3043
rect 17684 3000 17736 3009
rect 17868 3000 17920 3052
rect 19340 3000 19392 3052
rect 11796 2796 11848 2848
rect 19616 3111 19668 3120
rect 19616 3077 19625 3111
rect 19625 3077 19659 3111
rect 19659 3077 19668 3111
rect 19616 3068 19668 3077
rect 22744 3068 22796 3120
rect 22836 3111 22888 3120
rect 22836 3077 22845 3111
rect 22845 3077 22879 3111
rect 22879 3077 22888 3111
rect 22836 3068 22888 3077
rect 23020 3068 23072 3120
rect 24124 3068 24176 3120
rect 21640 3000 21692 3052
rect 22284 3000 22336 3052
rect 14372 2796 14424 2848
rect 16580 2796 16632 2848
rect 16856 2796 16908 2848
rect 17316 2864 17368 2916
rect 17960 2864 18012 2916
rect 17224 2839 17276 2848
rect 17224 2805 17233 2839
rect 17233 2805 17267 2839
rect 17267 2805 17276 2839
rect 17224 2796 17276 2805
rect 17684 2796 17736 2848
rect 19156 2864 19208 2916
rect 19708 2932 19760 2984
rect 20904 2932 20956 2984
rect 19984 2864 20036 2916
rect 18236 2796 18288 2848
rect 18420 2796 18472 2848
rect 19524 2796 19576 2848
rect 19800 2796 19852 2848
rect 20720 2864 20772 2916
rect 22468 2932 22520 2984
rect 21272 2796 21324 2848
rect 21548 2796 21600 2848
rect 24216 2796 24268 2848
rect 24492 2839 24544 2848
rect 24492 2805 24501 2839
rect 24501 2805 24535 2839
rect 24535 2805 24544 2839
rect 24492 2796 24544 2805
rect 3917 2694 3969 2746
rect 3981 2694 4033 2746
rect 4045 2694 4097 2746
rect 4109 2694 4161 2746
rect 4173 2694 4225 2746
rect 9851 2694 9903 2746
rect 9915 2694 9967 2746
rect 9979 2694 10031 2746
rect 10043 2694 10095 2746
rect 10107 2694 10159 2746
rect 15785 2694 15837 2746
rect 15849 2694 15901 2746
rect 15913 2694 15965 2746
rect 15977 2694 16029 2746
rect 16041 2694 16093 2746
rect 21719 2694 21771 2746
rect 21783 2694 21835 2746
rect 21847 2694 21899 2746
rect 21911 2694 21963 2746
rect 21975 2694 22027 2746
rect 1952 2635 2004 2644
rect 1952 2601 1961 2635
rect 1961 2601 1995 2635
rect 1995 2601 2004 2635
rect 1952 2592 2004 2601
rect 4436 2592 4488 2644
rect 4988 2592 5040 2644
rect 5172 2635 5224 2644
rect 5172 2601 5181 2635
rect 5181 2601 5215 2635
rect 5215 2601 5224 2635
rect 5172 2592 5224 2601
rect 6828 2592 6880 2644
rect 8208 2592 8260 2644
rect 8392 2592 8444 2644
rect 9404 2635 9456 2644
rect 9404 2601 9413 2635
rect 9413 2601 9447 2635
rect 9447 2601 9456 2635
rect 9404 2592 9456 2601
rect 940 2388 992 2440
rect 1492 2388 1544 2440
rect 2504 2431 2556 2440
rect 2504 2397 2513 2431
rect 2513 2397 2547 2431
rect 2547 2397 2556 2431
rect 2504 2388 2556 2397
rect 9680 2524 9732 2576
rect 5356 2456 5408 2508
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 756 2320 808 2372
rect 4528 2320 4580 2372
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 5908 2388 5960 2440
rect 5264 2320 5316 2372
rect 4068 2252 4120 2304
rect 5540 2252 5592 2304
rect 5816 2363 5868 2372
rect 5816 2329 5825 2363
rect 5825 2329 5859 2363
rect 5859 2329 5868 2363
rect 5816 2320 5868 2329
rect 7104 2388 7156 2440
rect 7564 2388 7616 2440
rect 6368 2252 6420 2304
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 11060 2592 11112 2644
rect 11244 2635 11296 2644
rect 11244 2601 11253 2635
rect 11253 2601 11287 2635
rect 11287 2601 11296 2635
rect 11244 2592 11296 2601
rect 14004 2592 14056 2644
rect 16764 2592 16816 2644
rect 17408 2592 17460 2644
rect 19064 2592 19116 2644
rect 11336 2456 11388 2508
rect 13912 2524 13964 2576
rect 20076 2592 20128 2644
rect 21916 2635 21968 2644
rect 21916 2601 21925 2635
rect 21925 2601 21959 2635
rect 21959 2601 21968 2635
rect 21916 2592 21968 2601
rect 24584 2592 24636 2644
rect 8668 2320 8720 2372
rect 11520 2320 11572 2372
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 7932 2252 7984 2304
rect 8576 2295 8628 2304
rect 8576 2261 8585 2295
rect 8585 2261 8619 2295
rect 8619 2261 8628 2295
rect 8576 2252 8628 2261
rect 9588 2295 9640 2304
rect 9588 2261 9597 2295
rect 9597 2261 9631 2295
rect 9631 2261 9640 2295
rect 9588 2252 9640 2261
rect 10784 2252 10836 2304
rect 11704 2252 11756 2304
rect 11796 2295 11848 2304
rect 11796 2261 11805 2295
rect 11805 2261 11839 2295
rect 11839 2261 11848 2295
rect 11796 2252 11848 2261
rect 12072 2295 12124 2304
rect 12072 2261 12081 2295
rect 12081 2261 12115 2295
rect 12115 2261 12124 2295
rect 12072 2252 12124 2261
rect 12440 2388 12492 2440
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 13544 2431 13596 2440
rect 13544 2397 13553 2431
rect 13553 2397 13587 2431
rect 13587 2397 13596 2431
rect 13544 2388 13596 2397
rect 14740 2388 14792 2440
rect 14832 2431 14884 2440
rect 14832 2397 14841 2431
rect 14841 2397 14875 2431
rect 14875 2397 14884 2431
rect 14832 2388 14884 2397
rect 15108 2431 15160 2440
rect 15108 2397 15117 2431
rect 15117 2397 15151 2431
rect 15151 2397 15160 2431
rect 15108 2388 15160 2397
rect 15476 2431 15528 2440
rect 15476 2397 15485 2431
rect 15485 2397 15519 2431
rect 15519 2397 15528 2431
rect 15476 2388 15528 2397
rect 16948 2456 17000 2508
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 18328 2456 18380 2508
rect 18604 2456 18656 2508
rect 17316 2388 17368 2440
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 12440 2252 12492 2304
rect 13176 2252 13228 2304
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13360 2252 13412 2261
rect 13636 2295 13688 2304
rect 13636 2261 13645 2295
rect 13645 2261 13679 2295
rect 13679 2261 13688 2295
rect 13636 2252 13688 2261
rect 14556 2252 14608 2304
rect 14924 2295 14976 2304
rect 14924 2261 14933 2295
rect 14933 2261 14967 2295
rect 14967 2261 14976 2295
rect 14924 2252 14976 2261
rect 15844 2295 15896 2304
rect 15844 2261 15853 2295
rect 15853 2261 15887 2295
rect 15887 2261 15896 2295
rect 15844 2252 15896 2261
rect 16672 2295 16724 2304
rect 16672 2261 16681 2295
rect 16681 2261 16715 2295
rect 16715 2261 16724 2295
rect 16672 2252 16724 2261
rect 19340 2320 19392 2372
rect 17132 2252 17184 2304
rect 17316 2295 17368 2304
rect 17316 2261 17325 2295
rect 17325 2261 17359 2295
rect 17359 2261 17368 2295
rect 17316 2252 17368 2261
rect 17776 2295 17828 2304
rect 17776 2261 17785 2295
rect 17785 2261 17819 2295
rect 17819 2261 17828 2295
rect 17776 2252 17828 2261
rect 18604 2252 18656 2304
rect 20812 2456 20864 2508
rect 22468 2499 22520 2508
rect 22468 2465 22477 2499
rect 22477 2465 22511 2499
rect 22511 2465 22520 2499
rect 22468 2456 22520 2465
rect 23756 2388 23808 2440
rect 23848 2388 23900 2440
rect 19800 2252 19852 2304
rect 20628 2363 20680 2372
rect 20628 2329 20637 2363
rect 20637 2329 20671 2363
rect 20671 2329 20680 2363
rect 20628 2320 20680 2329
rect 21456 2320 21508 2372
rect 21732 2320 21784 2372
rect 23480 2320 23532 2372
rect 25136 2320 25188 2372
rect 6884 2150 6936 2202
rect 6948 2150 7000 2202
rect 7012 2150 7064 2202
rect 7076 2150 7128 2202
rect 7140 2150 7192 2202
rect 12818 2150 12870 2202
rect 12882 2150 12934 2202
rect 12946 2150 12998 2202
rect 13010 2150 13062 2202
rect 13074 2150 13126 2202
rect 18752 2150 18804 2202
rect 18816 2150 18868 2202
rect 18880 2150 18932 2202
rect 18944 2150 18996 2202
rect 19008 2150 19060 2202
rect 24686 2150 24738 2202
rect 24750 2150 24802 2202
rect 24814 2150 24866 2202
rect 24878 2150 24930 2202
rect 24942 2150 24994 2202
rect 3056 2048 3108 2100
rect 3608 2048 3660 2100
rect 3976 2048 4028 2100
rect 4068 2091 4120 2100
rect 4068 2057 4077 2091
rect 4077 2057 4111 2091
rect 4111 2057 4120 2091
rect 4068 2048 4120 2057
rect 4252 2048 4304 2100
rect 4436 2091 4488 2100
rect 4436 2057 4445 2091
rect 4445 2057 4479 2091
rect 4479 2057 4488 2091
rect 4436 2048 4488 2057
rect 5080 2048 5132 2100
rect 5172 2048 5224 2100
rect 2872 1980 2924 2032
rect 204 1912 256 1964
rect 848 1844 900 1896
rect 1032 1776 1084 1828
rect 2780 1955 2832 1964
rect 2780 1921 2789 1955
rect 2789 1921 2823 1955
rect 2823 1921 2832 1955
rect 2780 1912 2832 1921
rect 3056 1955 3108 1964
rect 3056 1921 3065 1955
rect 3065 1921 3099 1955
rect 3099 1921 3108 1955
rect 3056 1912 3108 1921
rect 3516 1955 3568 1964
rect 3516 1921 3525 1955
rect 3525 1921 3559 1955
rect 3559 1921 3568 1955
rect 3516 1912 3568 1921
rect 3700 1912 3752 1964
rect 5632 1980 5684 2032
rect 5816 2048 5868 2100
rect 6000 2048 6052 2100
rect 7012 2091 7064 2100
rect 7012 2057 7021 2091
rect 7021 2057 7055 2091
rect 7055 2057 7064 2091
rect 7012 2048 7064 2057
rect 7748 2091 7800 2100
rect 7748 2057 7757 2091
rect 7757 2057 7791 2091
rect 7791 2057 7800 2091
rect 7748 2048 7800 2057
rect 7932 2048 7984 2100
rect 8116 2091 8168 2100
rect 8116 2057 8125 2091
rect 8125 2057 8159 2091
rect 8159 2057 8168 2091
rect 8116 2048 8168 2057
rect 8484 2091 8536 2100
rect 8484 2057 8493 2091
rect 8493 2057 8527 2091
rect 8527 2057 8536 2091
rect 8484 2048 8536 2057
rect 8576 2048 8628 2100
rect 8852 2091 8904 2100
rect 8852 2057 8861 2091
rect 8861 2057 8895 2091
rect 8895 2057 8904 2091
rect 8852 2048 8904 2057
rect 4068 1844 4120 1896
rect 5080 1912 5132 1964
rect 6368 1912 6420 1964
rect 5724 1844 5776 1896
rect 6552 2023 6604 2032
rect 6552 1989 6561 2023
rect 6561 1989 6595 2023
rect 6595 1989 6604 2023
rect 6552 1980 6604 1989
rect 7288 1980 7340 2032
rect 8944 1980 8996 2032
rect 7472 1912 7524 1964
rect 8024 1844 8076 1896
rect 8300 1912 8352 1964
rect 9864 2048 9916 2100
rect 10232 2048 10284 2100
rect 10324 1980 10376 2032
rect 9404 1912 9456 1964
rect 10416 1912 10468 1964
rect 13360 2048 13412 2100
rect 13636 2048 13688 2100
rect 14924 2048 14976 2100
rect 15844 2048 15896 2100
rect 17316 2048 17368 2100
rect 18604 2048 18656 2100
rect 19340 2048 19392 2100
rect 19800 2048 19852 2100
rect 20352 2048 20404 2100
rect 21732 2048 21784 2100
rect 23480 2048 23532 2100
rect 23940 2048 23992 2100
rect 24492 2048 24544 2100
rect 11704 1980 11756 2032
rect 12348 1955 12400 1964
rect 12348 1921 12357 1955
rect 12357 1921 12391 1955
rect 12391 1921 12400 1955
rect 12348 1912 12400 1921
rect 13728 1912 13780 1964
rect 13820 1955 13872 1964
rect 13820 1921 13829 1955
rect 13829 1921 13863 1955
rect 13863 1921 13872 1955
rect 13820 1912 13872 1921
rect 14280 1955 14332 1964
rect 14280 1921 14289 1955
rect 14289 1921 14323 1955
rect 14323 1921 14332 1955
rect 14280 1912 14332 1921
rect 17592 1980 17644 2032
rect 18512 1980 18564 2032
rect 3332 1751 3384 1760
rect 3332 1717 3341 1751
rect 3341 1717 3375 1751
rect 3375 1717 3384 1751
rect 3332 1708 3384 1717
rect 4804 1708 4856 1760
rect 5356 1708 5408 1760
rect 11704 1844 11756 1896
rect 16120 1955 16172 1964
rect 16120 1921 16129 1955
rect 16129 1921 16163 1955
rect 16163 1921 16172 1955
rect 16120 1912 16172 1921
rect 16856 1912 16908 1964
rect 18604 1912 18656 1964
rect 19524 1912 19576 1964
rect 20260 1912 20312 1964
rect 20720 1955 20772 1964
rect 20720 1921 20729 1955
rect 20729 1921 20763 1955
rect 20763 1921 20772 1955
rect 20720 1912 20772 1921
rect 21364 1912 21416 1964
rect 24308 1955 24360 1964
rect 24308 1921 24317 1955
rect 24317 1921 24351 1955
rect 24351 1921 24360 1955
rect 24308 1912 24360 1921
rect 11152 1819 11204 1828
rect 11152 1785 11161 1819
rect 11161 1785 11195 1819
rect 11195 1785 11204 1819
rect 11152 1776 11204 1785
rect 11888 1776 11940 1828
rect 15384 1776 15436 1828
rect 12256 1708 12308 1760
rect 12624 1751 12676 1760
rect 12624 1717 12633 1751
rect 12633 1717 12667 1751
rect 12667 1717 12676 1751
rect 12624 1708 12676 1717
rect 13360 1751 13412 1760
rect 13360 1717 13369 1751
rect 13369 1717 13403 1751
rect 13403 1717 13412 1751
rect 13360 1708 13412 1717
rect 13636 1751 13688 1760
rect 13636 1717 13645 1751
rect 13645 1717 13679 1751
rect 13679 1717 13688 1751
rect 13636 1708 13688 1717
rect 14096 1751 14148 1760
rect 14096 1717 14105 1751
rect 14105 1717 14139 1751
rect 14139 1717 14148 1751
rect 14096 1708 14148 1717
rect 14280 1708 14332 1760
rect 14740 1708 14792 1760
rect 15752 1751 15804 1760
rect 15752 1717 15761 1751
rect 15761 1717 15795 1751
rect 15795 1717 15804 1751
rect 15752 1708 15804 1717
rect 17132 1776 17184 1828
rect 19800 1844 19852 1896
rect 25320 1844 25372 1896
rect 16856 1751 16908 1760
rect 16856 1717 16865 1751
rect 16865 1717 16899 1751
rect 16899 1717 16908 1751
rect 16856 1708 16908 1717
rect 17960 1751 18012 1760
rect 17960 1717 17969 1751
rect 17969 1717 18003 1751
rect 18003 1717 18012 1751
rect 17960 1708 18012 1717
rect 18144 1708 18196 1760
rect 22744 1776 22796 1828
rect 19524 1708 19576 1760
rect 20168 1708 20220 1760
rect 3917 1606 3969 1658
rect 3981 1606 4033 1658
rect 4045 1606 4097 1658
rect 4109 1606 4161 1658
rect 4173 1606 4225 1658
rect 9851 1606 9903 1658
rect 9915 1606 9967 1658
rect 9979 1606 10031 1658
rect 10043 1606 10095 1658
rect 10107 1606 10159 1658
rect 15785 1606 15837 1658
rect 15849 1606 15901 1658
rect 15913 1606 15965 1658
rect 15977 1606 16029 1658
rect 16041 1606 16093 1658
rect 21719 1606 21771 1658
rect 21783 1606 21835 1658
rect 21847 1606 21899 1658
rect 21911 1606 21963 1658
rect 21975 1606 22027 1658
rect 3332 1504 3384 1556
rect 4436 1504 4488 1556
rect 4528 1504 4580 1556
rect 9036 1504 9088 1556
rect 10416 1504 10468 1556
rect 10968 1504 11020 1556
rect 1676 1300 1728 1352
rect 2044 1300 2096 1352
rect 2228 1343 2280 1352
rect 2228 1309 2237 1343
rect 2237 1309 2271 1343
rect 2271 1309 2280 1343
rect 2228 1300 2280 1309
rect 2596 1300 2648 1352
rect 3792 1300 3844 1352
rect 7748 1436 7800 1488
rect 6460 1368 6512 1420
rect 1584 1275 1636 1284
rect 1584 1241 1593 1275
rect 1593 1241 1627 1275
rect 1627 1241 1636 1275
rect 1584 1232 1636 1241
rect 1952 1275 2004 1284
rect 1952 1241 1961 1275
rect 1961 1241 1995 1275
rect 1995 1241 2004 1275
rect 1952 1232 2004 1241
rect 2964 1232 3016 1284
rect 3884 1207 3936 1216
rect 3884 1173 3893 1207
rect 3893 1173 3927 1207
rect 3927 1173 3936 1207
rect 3884 1164 3936 1173
rect 4068 1164 4120 1216
rect 4436 1343 4488 1352
rect 4436 1309 4445 1343
rect 4445 1309 4479 1343
rect 4479 1309 4488 1343
rect 4436 1300 4488 1309
rect 5816 1300 5868 1352
rect 6276 1300 6328 1352
rect 6368 1300 6420 1352
rect 6736 1343 6788 1352
rect 6736 1309 6745 1343
rect 6745 1309 6779 1343
rect 6779 1309 6788 1343
rect 6736 1300 6788 1309
rect 6920 1368 6972 1420
rect 8208 1300 8260 1352
rect 9036 1300 9088 1352
rect 10232 1368 10284 1420
rect 9588 1343 9640 1352
rect 9588 1309 9597 1343
rect 9597 1309 9631 1343
rect 9631 1309 9640 1343
rect 9588 1300 9640 1309
rect 9680 1300 9732 1352
rect 6000 1232 6052 1284
rect 5080 1207 5132 1216
rect 5080 1173 5089 1207
rect 5089 1173 5123 1207
rect 5123 1173 5132 1207
rect 5080 1164 5132 1173
rect 5540 1207 5592 1216
rect 5540 1173 5549 1207
rect 5549 1173 5583 1207
rect 5583 1173 5592 1207
rect 5540 1164 5592 1173
rect 6092 1207 6144 1216
rect 6092 1173 6101 1207
rect 6101 1173 6135 1207
rect 6135 1173 6144 1207
rect 6092 1164 6144 1173
rect 6460 1164 6512 1216
rect 6552 1164 6604 1216
rect 6736 1164 6788 1216
rect 6920 1164 6972 1216
rect 7564 1207 7616 1216
rect 7564 1173 7573 1207
rect 7573 1173 7607 1207
rect 7607 1173 7616 1207
rect 7564 1164 7616 1173
rect 7932 1207 7984 1216
rect 7932 1173 7941 1207
rect 7941 1173 7975 1207
rect 7975 1173 7984 1207
rect 7932 1164 7984 1173
rect 8944 1207 8996 1216
rect 8944 1173 8953 1207
rect 8953 1173 8987 1207
rect 8987 1173 8996 1207
rect 8944 1164 8996 1173
rect 9772 1207 9824 1216
rect 9772 1173 9781 1207
rect 9781 1173 9815 1207
rect 9815 1173 9824 1207
rect 9772 1164 9824 1173
rect 10784 1232 10836 1284
rect 12440 1504 12492 1556
rect 12532 1504 12584 1556
rect 13360 1504 13412 1556
rect 13728 1504 13780 1556
rect 14924 1504 14976 1556
rect 11704 1436 11756 1488
rect 11980 1436 12032 1488
rect 12072 1436 12124 1488
rect 11336 1368 11388 1420
rect 12256 1368 12308 1420
rect 11796 1300 11848 1352
rect 14096 1436 14148 1488
rect 14188 1436 14240 1488
rect 15200 1436 15252 1488
rect 16120 1504 16172 1556
rect 16028 1436 16080 1488
rect 11152 1232 11204 1284
rect 13176 1300 13228 1352
rect 13636 1343 13688 1352
rect 13636 1309 13645 1343
rect 13645 1309 13679 1343
rect 13679 1309 13688 1343
rect 13636 1300 13688 1309
rect 10600 1164 10652 1216
rect 11244 1207 11296 1216
rect 11244 1173 11253 1207
rect 11253 1173 11287 1207
rect 11287 1173 11296 1207
rect 11244 1164 11296 1173
rect 11520 1164 11572 1216
rect 11704 1207 11756 1216
rect 11704 1173 11713 1207
rect 11713 1173 11747 1207
rect 11747 1173 11756 1207
rect 11704 1164 11756 1173
rect 14556 1232 14608 1284
rect 16212 1368 16264 1420
rect 18328 1504 18380 1556
rect 24492 1504 24544 1556
rect 21272 1436 21324 1488
rect 16488 1343 16540 1352
rect 16488 1309 16497 1343
rect 16497 1309 16531 1343
rect 16531 1309 16540 1343
rect 16488 1300 16540 1309
rect 16672 1300 16724 1352
rect 17224 1300 17276 1352
rect 19800 1368 19852 1420
rect 17684 1300 17736 1352
rect 18512 1343 18564 1352
rect 18512 1309 18521 1343
rect 18521 1309 18555 1343
rect 18555 1309 18564 1343
rect 18512 1300 18564 1309
rect 19432 1343 19484 1352
rect 19432 1309 19441 1343
rect 19441 1309 19475 1343
rect 19475 1309 19484 1343
rect 19432 1300 19484 1309
rect 20352 1300 20404 1352
rect 20444 1343 20496 1352
rect 20444 1309 20453 1343
rect 20453 1309 20487 1343
rect 20487 1309 20496 1343
rect 20444 1300 20496 1309
rect 20996 1300 21048 1352
rect 23020 1300 23072 1352
rect 13452 1207 13504 1216
rect 13452 1173 13461 1207
rect 13461 1173 13495 1207
rect 13495 1173 13504 1207
rect 13452 1164 13504 1173
rect 13636 1164 13688 1216
rect 14004 1164 14056 1216
rect 16488 1164 16540 1216
rect 19616 1232 19668 1284
rect 21272 1275 21324 1284
rect 21272 1241 21281 1275
rect 21281 1241 21315 1275
rect 21315 1241 21324 1275
rect 21272 1232 21324 1241
rect 22192 1232 22244 1284
rect 22468 1275 22520 1284
rect 22468 1241 22477 1275
rect 22477 1241 22511 1275
rect 22511 1241 22520 1275
rect 22468 1232 22520 1241
rect 20904 1164 20956 1216
rect 6884 1062 6936 1114
rect 6948 1062 7000 1114
rect 7012 1062 7064 1114
rect 7076 1062 7128 1114
rect 7140 1062 7192 1114
rect 12818 1062 12870 1114
rect 12882 1062 12934 1114
rect 12946 1062 12998 1114
rect 13010 1062 13062 1114
rect 13074 1062 13126 1114
rect 18752 1062 18804 1114
rect 18816 1062 18868 1114
rect 18880 1062 18932 1114
rect 18944 1062 18996 1114
rect 19008 1062 19060 1114
rect 24686 1062 24738 1114
rect 24750 1062 24802 1114
rect 24814 1062 24866 1114
rect 24878 1062 24930 1114
rect 24942 1062 24994 1114
rect 5080 960 5132 1012
rect 8300 960 8352 1012
rect 8668 960 8720 1012
rect 11244 960 11296 1012
rect 12900 960 12952 1012
rect 14372 960 14424 1012
rect 21272 960 21324 1012
rect 3884 892 3936 944
rect 7472 892 7524 944
rect 6460 824 6512 876
rect 8944 892 8996 944
rect 11336 892 11388 944
rect 19432 892 19484 944
rect 22836 892 22888 944
rect 572 756 624 808
rect 11520 756 11572 808
rect 6184 688 6236 740
rect 7104 688 7156 740
rect 7564 688 7616 740
rect 9036 688 9088 740
rect 9680 688 9732 740
rect 12716 620 12768 672
rect 21272 620 21324 672
rect 22468 620 22520 672
rect 6368 552 6420 604
rect 9588 552 9640 604
rect 5816 484 5868 536
rect 9036 484 9088 536
rect 6736 348 6788 400
rect 11428 348 11480 400
<< metal2 >>
rect 202 44840 258 45000
rect 478 44840 534 45000
rect 754 44840 810 45000
rect 1030 44840 1086 45000
rect 1306 44840 1362 45000
rect 1582 44840 1638 45000
rect 1858 44962 1914 45000
rect 1858 44934 2084 44962
rect 1858 44840 1914 44934
rect 216 41274 244 44840
rect 492 42090 520 44840
rect 480 42084 532 42090
rect 480 42026 532 42032
rect 768 41614 796 44840
rect 1044 42362 1072 44840
rect 1032 42356 1084 42362
rect 1032 42298 1084 42304
rect 1320 42022 1348 44840
rect 1400 42628 1452 42634
rect 1452 42588 1532 42616
rect 1400 42570 1452 42576
rect 1400 42220 1452 42226
rect 1400 42162 1452 42168
rect 1308 42016 1360 42022
rect 1308 41958 1360 41964
rect 1030 41712 1086 41721
rect 1030 41647 1086 41656
rect 756 41608 808 41614
rect 756 41550 808 41556
rect 204 41268 256 41274
rect 204 41210 256 41216
rect 662 40216 718 40225
rect 662 40151 718 40160
rect 572 39636 624 39642
rect 572 39578 624 39584
rect 20 36712 72 36718
rect 20 36654 72 36660
rect 32 33726 60 36654
rect 478 36136 534 36145
rect 478 36071 534 36080
rect 20 33720 72 33726
rect 20 33662 72 33668
rect 32 26738 60 33662
rect 112 33584 164 33590
rect 112 33526 164 33532
rect 124 27010 152 33526
rect 492 31686 520 36071
rect 480 31680 532 31686
rect 480 31622 532 31628
rect 480 30864 532 30870
rect 480 30806 532 30812
rect 124 26982 428 27010
rect 492 26994 520 30806
rect 296 26920 348 26926
rect 296 26862 348 26868
rect 32 26710 244 26738
rect 20 26648 72 26654
rect 20 26590 72 26596
rect 32 22234 60 26590
rect 112 26512 164 26518
rect 112 26454 164 26460
rect 124 24886 152 26454
rect 112 24880 164 24886
rect 112 24822 164 24828
rect 20 22228 72 22234
rect 20 22170 72 22176
rect 20 16108 72 16114
rect 20 16050 72 16056
rect 32 1873 60 16050
rect 124 11694 152 24822
rect 216 19718 244 26710
rect 308 25022 336 26862
rect 296 25016 348 25022
rect 296 24958 348 24964
rect 400 24546 428 26982
rect 480 26988 532 26994
rect 480 26930 532 26936
rect 478 26888 534 26897
rect 478 26823 534 26832
rect 388 24540 440 24546
rect 388 24482 440 24488
rect 492 24426 520 26823
rect 308 24398 520 24426
rect 204 19712 256 19718
rect 204 19654 256 19660
rect 308 17134 336 24398
rect 388 24336 440 24342
rect 388 24278 440 24284
rect 296 17128 348 17134
rect 296 17070 348 17076
rect 400 16130 428 24278
rect 478 19816 534 19825
rect 478 19751 534 19760
rect 308 16102 428 16130
rect 492 16114 520 19751
rect 480 16108 532 16114
rect 308 15858 336 16102
rect 480 16050 532 16056
rect 308 15830 428 15858
rect 112 11688 164 11694
rect 112 11630 164 11636
rect 204 1964 256 1970
rect 204 1906 256 1912
rect 18 1864 74 1873
rect 18 1799 74 1808
rect 216 160 244 1906
rect 400 1465 428 15830
rect 584 2990 612 39578
rect 676 31754 704 40151
rect 938 40080 994 40089
rect 860 40038 938 40066
rect 860 33522 888 40038
rect 938 40015 994 40024
rect 940 39296 992 39302
rect 940 39238 992 39244
rect 848 33516 900 33522
rect 848 33458 900 33464
rect 676 31726 888 31754
rect 664 31680 716 31686
rect 664 31622 716 31628
rect 676 26081 704 31622
rect 756 28484 808 28490
rect 756 28426 808 28432
rect 768 28121 796 28426
rect 754 28112 810 28121
rect 754 28047 810 28056
rect 860 27962 888 31726
rect 768 27934 888 27962
rect 662 26072 718 26081
rect 662 26007 718 26016
rect 664 25016 716 25022
rect 664 24958 716 24964
rect 768 24970 796 27934
rect 952 27010 980 39238
rect 860 26982 980 27010
rect 860 26654 888 26982
rect 848 26648 900 26654
rect 848 26590 900 26596
rect 940 26036 992 26042
rect 940 25978 992 25984
rect 848 25968 900 25974
rect 848 25910 900 25916
rect 860 25129 888 25910
rect 952 25401 980 25978
rect 938 25392 994 25401
rect 938 25327 994 25336
rect 940 25152 992 25158
rect 846 25120 902 25129
rect 940 25094 992 25100
rect 846 25055 902 25064
rect 676 24834 704 24958
rect 768 24942 888 24970
rect 676 24806 796 24834
rect 662 22808 718 22817
rect 662 22743 718 22752
rect 676 17218 704 22743
rect 768 19666 796 24806
rect 860 24721 888 24942
rect 846 24712 902 24721
rect 846 24647 902 24656
rect 952 23905 980 25094
rect 938 23896 994 23905
rect 938 23831 994 23840
rect 1044 22094 1072 41647
rect 1412 39545 1440 42162
rect 1398 39536 1454 39545
rect 1398 39471 1454 39480
rect 1504 39137 1532 42588
rect 1596 42294 1624 44840
rect 1768 43648 1820 43654
rect 1768 43590 1820 43596
rect 1780 43314 1808 43590
rect 2056 43330 2084 44934
rect 2134 44840 2190 45000
rect 2410 44840 2466 45000
rect 2686 44840 2742 45000
rect 2962 44840 3018 45000
rect 3238 44962 3294 45000
rect 3514 44962 3570 45000
rect 3238 44934 3372 44962
rect 3238 44840 3294 44934
rect 2148 43450 2176 44840
rect 2424 43450 2452 44840
rect 2136 43444 2188 43450
rect 2136 43386 2188 43392
rect 2412 43444 2464 43450
rect 2412 43386 2464 43392
rect 1676 43308 1728 43314
rect 1676 43250 1728 43256
rect 1768 43308 1820 43314
rect 2056 43302 2176 43330
rect 1768 43250 1820 43256
rect 1584 42288 1636 42294
rect 1584 42230 1636 42236
rect 1688 41414 1716 43250
rect 2044 42628 2096 42634
rect 2044 42570 2096 42576
rect 1688 41386 1808 41414
rect 1674 41032 1730 41041
rect 1674 40967 1676 40976
rect 1728 40967 1730 40976
rect 1676 40938 1728 40944
rect 1676 40520 1728 40526
rect 1676 40462 1728 40468
rect 1584 39432 1636 39438
rect 1584 39374 1636 39380
rect 1490 39128 1546 39137
rect 1490 39063 1546 39072
rect 1400 38956 1452 38962
rect 1452 38916 1532 38944
rect 1400 38898 1452 38904
rect 1398 38720 1454 38729
rect 1398 38655 1454 38664
rect 1412 38350 1440 38655
rect 1504 38457 1532 38916
rect 1490 38448 1546 38457
rect 1490 38383 1546 38392
rect 1400 38344 1452 38350
rect 1400 38286 1452 38292
rect 1216 38208 1268 38214
rect 1216 38150 1268 38156
rect 1306 38176 1362 38185
rect 1228 37641 1256 38150
rect 1306 38111 1362 38120
rect 1320 38010 1348 38111
rect 1308 38004 1360 38010
rect 1308 37946 1360 37952
rect 1214 37632 1270 37641
rect 1214 37567 1270 37576
rect 1308 37120 1360 37126
rect 1596 37097 1624 39374
rect 1688 38321 1716 40462
rect 1674 38312 1730 38321
rect 1674 38247 1730 38256
rect 1780 37890 1808 41386
rect 2056 40361 2084 42570
rect 2148 41138 2176 43302
rect 2700 42770 2728 44840
rect 2976 43450 3004 44840
rect 2964 43444 3016 43450
rect 2964 43386 3016 43392
rect 2872 43308 2924 43314
rect 2872 43250 2924 43256
rect 2688 42764 2740 42770
rect 2688 42706 2740 42712
rect 2502 42256 2558 42265
rect 2502 42191 2504 42200
rect 2556 42191 2558 42200
rect 2504 42162 2556 42168
rect 2228 42152 2280 42158
rect 2226 42120 2228 42129
rect 2280 42120 2282 42129
rect 2226 42055 2282 42064
rect 2412 41540 2464 41546
rect 2412 41482 2464 41488
rect 2136 41132 2188 41138
rect 2136 41074 2188 41080
rect 2320 41132 2372 41138
rect 2320 41074 2372 41080
rect 2226 40624 2282 40633
rect 2226 40559 2282 40568
rect 2042 40352 2098 40361
rect 2042 40287 2098 40296
rect 1860 39840 1912 39846
rect 1860 39782 1912 39788
rect 1872 39574 1900 39782
rect 1860 39568 1912 39574
rect 1860 39510 1912 39516
rect 1872 39098 1900 39510
rect 1952 39432 2004 39438
rect 1952 39374 2004 39380
rect 1860 39092 1912 39098
rect 1860 39034 1912 39040
rect 1860 38956 1912 38962
rect 1860 38898 1912 38904
rect 1688 37862 1808 37890
rect 1308 37062 1360 37068
rect 1582 37088 1638 37097
rect 1216 36780 1268 36786
rect 1216 36722 1268 36728
rect 1124 36032 1176 36038
rect 1124 35974 1176 35980
rect 1136 34388 1164 35974
rect 1228 34513 1256 36722
rect 1320 36009 1348 37062
rect 1582 37023 1638 37032
rect 1688 36689 1716 37862
rect 1872 37856 1900 38898
rect 1964 38729 1992 39374
rect 2044 39364 2096 39370
rect 2044 39306 2096 39312
rect 2056 38962 2084 39306
rect 2044 38956 2096 38962
rect 2044 38898 2096 38904
rect 2240 38894 2268 40559
rect 2332 39273 2360 41074
rect 2424 39817 2452 41482
rect 2780 41472 2832 41478
rect 2780 41414 2832 41420
rect 2688 41132 2740 41138
rect 2688 41074 2740 41080
rect 2594 40624 2650 40633
rect 2594 40559 2650 40568
rect 2608 40526 2636 40559
rect 2596 40520 2648 40526
rect 2700 40497 2728 41074
rect 2596 40462 2648 40468
rect 2686 40488 2742 40497
rect 2686 40423 2742 40432
rect 2504 40044 2556 40050
rect 2504 39986 2556 39992
rect 2410 39808 2466 39817
rect 2410 39743 2466 39752
rect 2516 39545 2544 39986
rect 2596 39840 2648 39846
rect 2596 39782 2648 39788
rect 2502 39536 2558 39545
rect 2502 39471 2558 39480
rect 2318 39264 2374 39273
rect 2318 39199 2374 39208
rect 2228 38888 2280 38894
rect 2228 38830 2280 38836
rect 2044 38820 2096 38826
rect 2044 38762 2096 38768
rect 1950 38720 2006 38729
rect 1950 38655 2006 38664
rect 1872 37828 1992 37856
rect 1768 37800 1820 37806
rect 1768 37742 1820 37748
rect 1780 37466 1808 37742
rect 1860 37732 1912 37738
rect 1860 37674 1912 37680
rect 1768 37460 1820 37466
rect 1768 37402 1820 37408
rect 1768 36712 1820 36718
rect 1674 36680 1730 36689
rect 1768 36654 1820 36660
rect 1674 36615 1730 36624
rect 1400 36168 1452 36174
rect 1400 36110 1452 36116
rect 1306 36000 1362 36009
rect 1306 35935 1362 35944
rect 1308 35760 1360 35766
rect 1308 35702 1360 35708
rect 1320 34921 1348 35702
rect 1306 34912 1362 34921
rect 1306 34847 1362 34856
rect 1214 34504 1270 34513
rect 1214 34439 1270 34448
rect 1136 34360 1256 34388
rect 1124 33516 1176 33522
rect 1124 33458 1176 33464
rect 1136 31754 1164 33458
rect 1228 32570 1256 34360
rect 1412 34105 1440 36110
rect 1492 35692 1544 35698
rect 1492 35634 1544 35640
rect 1504 34626 1532 35634
rect 1676 35624 1728 35630
rect 1674 35592 1676 35601
rect 1728 35592 1730 35601
rect 1674 35527 1730 35536
rect 1676 35148 1728 35154
rect 1676 35090 1728 35096
rect 1504 34598 1624 34626
rect 1492 34536 1544 34542
rect 1492 34478 1544 34484
rect 1398 34096 1454 34105
rect 1398 34031 1454 34040
rect 1504 33862 1532 34478
rect 1492 33856 1544 33862
rect 1492 33798 1544 33804
rect 1400 33516 1452 33522
rect 1400 33458 1452 33464
rect 1308 32836 1360 32842
rect 1308 32778 1360 32784
rect 1216 32564 1268 32570
rect 1216 32506 1268 32512
rect 1228 32230 1256 32506
rect 1320 32473 1348 32778
rect 1306 32464 1362 32473
rect 1306 32399 1362 32408
rect 1216 32224 1268 32230
rect 1216 32166 1268 32172
rect 1412 32065 1440 33458
rect 1504 32892 1532 33798
rect 1596 33561 1624 34598
rect 1688 34388 1716 35090
rect 1780 34746 1808 36654
rect 1768 34740 1820 34746
rect 1768 34682 1820 34688
rect 1768 34400 1820 34406
rect 1688 34360 1768 34388
rect 1768 34342 1820 34348
rect 1674 33688 1730 33697
rect 1674 33623 1730 33632
rect 1582 33552 1638 33561
rect 1688 33522 1716 33623
rect 1582 33487 1638 33496
rect 1676 33516 1728 33522
rect 1676 33458 1728 33464
rect 1872 33114 1900 37674
rect 1964 33862 1992 37828
rect 1952 33856 2004 33862
rect 1952 33798 2004 33804
rect 1952 33516 2004 33522
rect 1952 33458 2004 33464
rect 1860 33108 1912 33114
rect 1860 33050 1912 33056
rect 1584 32904 1636 32910
rect 1504 32864 1584 32892
rect 1584 32846 1636 32852
rect 1676 32904 1728 32910
rect 1676 32846 1728 32852
rect 1492 32768 1544 32774
rect 1492 32710 1544 32716
rect 1504 32366 1532 32710
rect 1492 32360 1544 32366
rect 1492 32302 1544 32308
rect 1398 32056 1454 32065
rect 1398 31991 1454 32000
rect 1136 31726 1256 31754
rect 1124 31408 1176 31414
rect 1124 31350 1176 31356
rect 1136 30841 1164 31350
rect 1122 30832 1178 30841
rect 1122 30767 1178 30776
rect 1122 29744 1178 29753
rect 1122 29679 1178 29688
rect 1136 29306 1164 29679
rect 1124 29300 1176 29306
rect 1124 29242 1176 29248
rect 1228 29186 1256 31726
rect 1596 31686 1624 32846
rect 1688 32473 1716 32846
rect 1674 32464 1730 32473
rect 1674 32399 1730 32408
rect 1676 32360 1728 32366
rect 1728 32308 1808 32314
rect 1676 32302 1808 32308
rect 1688 32286 1808 32302
rect 1676 32224 1728 32230
rect 1676 32166 1728 32172
rect 1584 31680 1636 31686
rect 1584 31622 1636 31628
rect 1490 31512 1546 31521
rect 1490 31447 1546 31456
rect 1400 30728 1452 30734
rect 1400 30670 1452 30676
rect 1306 30560 1362 30569
rect 1306 30495 1362 30504
rect 1320 30394 1348 30495
rect 1308 30388 1360 30394
rect 1308 30330 1360 30336
rect 1412 30297 1440 30670
rect 1398 30288 1454 30297
rect 1504 30258 1532 31447
rect 1584 31340 1636 31346
rect 1584 31282 1636 31288
rect 1596 30297 1624 31282
rect 1688 30580 1716 32166
rect 1780 31822 1808 32286
rect 1860 32292 1912 32298
rect 1860 32234 1912 32240
rect 1768 31816 1820 31822
rect 1768 31758 1820 31764
rect 1768 31680 1820 31686
rect 1768 31622 1820 31628
rect 1780 31278 1808 31622
rect 1768 31272 1820 31278
rect 1768 31214 1820 31220
rect 1780 30734 1808 31214
rect 1768 30728 1820 30734
rect 1768 30670 1820 30676
rect 1688 30552 1808 30580
rect 1582 30288 1638 30297
rect 1398 30223 1454 30232
rect 1492 30252 1544 30258
rect 1582 30223 1638 30232
rect 1676 30252 1728 30258
rect 1492 30194 1544 30200
rect 1676 30194 1728 30200
rect 1584 30184 1636 30190
rect 1584 30126 1636 30132
rect 1492 30116 1544 30122
rect 1492 30058 1544 30064
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1308 29572 1360 29578
rect 1308 29514 1360 29520
rect 1320 29481 1348 29514
rect 1306 29472 1362 29481
rect 1306 29407 1362 29416
rect 1412 29322 1440 29582
rect 1136 29158 1256 29186
rect 1320 29294 1440 29322
rect 1136 23089 1164 29158
rect 1214 28656 1270 28665
rect 1214 28591 1270 28600
rect 1228 28558 1256 28591
rect 1216 28552 1268 28558
rect 1216 28494 1268 28500
rect 1320 27996 1348 29294
rect 1400 29096 1452 29102
rect 1400 29038 1452 29044
rect 1412 28121 1440 29038
rect 1398 28112 1454 28121
rect 1398 28047 1454 28056
rect 1400 28008 1452 28014
rect 1320 27968 1400 27996
rect 1400 27950 1452 27956
rect 1412 27470 1440 27950
rect 1400 27464 1452 27470
rect 1214 27432 1270 27441
rect 1400 27406 1452 27412
rect 1214 27367 1270 27376
rect 1228 27033 1256 27367
rect 1308 27056 1360 27062
rect 1214 27024 1270 27033
rect 1308 26998 1360 27004
rect 1214 26959 1270 26968
rect 1320 26761 1348 26998
rect 1306 26752 1362 26761
rect 1306 26687 1362 26696
rect 1412 26586 1440 27406
rect 1400 26580 1452 26586
rect 1400 26522 1452 26528
rect 1504 26466 1532 30058
rect 1596 28966 1624 30126
rect 1584 28960 1636 28966
rect 1688 28937 1716 30194
rect 1584 28902 1636 28908
rect 1674 28928 1730 28937
rect 1674 28863 1730 28872
rect 1780 28082 1808 30552
rect 1872 29186 1900 32234
rect 1964 32201 1992 33458
rect 1950 32192 2006 32201
rect 1950 32127 2006 32136
rect 2056 31346 2084 38762
rect 2136 37732 2188 37738
rect 2136 37674 2188 37680
rect 2148 37466 2176 37674
rect 2136 37460 2188 37466
rect 2136 37402 2188 37408
rect 2136 37256 2188 37262
rect 2240 37244 2268 38830
rect 2516 38418 2544 39471
rect 2504 38412 2556 38418
rect 2504 38354 2556 38360
rect 2608 37874 2636 39782
rect 2792 39114 2820 41414
rect 2884 40186 2912 43250
rect 3344 42906 3372 44934
rect 3514 44934 3740 44962
rect 3514 44840 3570 44934
rect 3516 44056 3568 44062
rect 3516 43998 3568 44004
rect 3424 43716 3476 43722
rect 3424 43658 3476 43664
rect 3332 42900 3384 42906
rect 3332 42842 3384 42848
rect 3056 42628 3108 42634
rect 3056 42570 3108 42576
rect 3240 42628 3292 42634
rect 3240 42570 3292 42576
rect 2964 41064 3016 41070
rect 2964 41006 3016 41012
rect 2976 40186 3004 41006
rect 2872 40180 2924 40186
rect 2872 40122 2924 40128
rect 2964 40180 3016 40186
rect 2964 40122 3016 40128
rect 2964 40044 3016 40050
rect 2964 39986 3016 39992
rect 2792 39086 2912 39114
rect 2780 38956 2832 38962
rect 2780 38898 2832 38904
rect 2688 38276 2740 38282
rect 2688 38218 2740 38224
rect 2596 37868 2648 37874
rect 2596 37810 2648 37816
rect 2320 37800 2372 37806
rect 2320 37742 2372 37748
rect 2188 37216 2268 37244
rect 2136 37198 2188 37204
rect 2148 33946 2176 37198
rect 2332 36718 2360 37742
rect 2504 37664 2556 37670
rect 2504 37606 2556 37612
rect 2320 36712 2372 36718
rect 2320 36654 2372 36660
rect 2228 35148 2280 35154
rect 2228 35090 2280 35096
rect 2240 34202 2268 35090
rect 2412 34400 2464 34406
rect 2412 34342 2464 34348
rect 2228 34196 2280 34202
rect 2228 34138 2280 34144
rect 2226 33960 2282 33969
rect 2148 33918 2226 33946
rect 2226 33895 2282 33904
rect 2320 33924 2372 33930
rect 2320 33866 2372 33872
rect 2228 33856 2280 33862
rect 2228 33798 2280 33804
rect 2134 32600 2190 32609
rect 2134 32535 2190 32544
rect 2148 32366 2176 32535
rect 2136 32360 2188 32366
rect 2136 32302 2188 32308
rect 2240 31686 2268 33798
rect 2228 31680 2280 31686
rect 2226 31648 2228 31657
rect 2280 31648 2282 31657
rect 2226 31583 2282 31592
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 2226 30832 2282 30841
rect 2226 30767 2282 30776
rect 1952 30728 2004 30734
rect 1952 30670 2004 30676
rect 1964 29850 1992 30670
rect 2134 30424 2190 30433
rect 2134 30359 2190 30368
rect 2148 30190 2176 30359
rect 2136 30184 2188 30190
rect 2136 30126 2188 30132
rect 2136 30048 2188 30054
rect 2136 29990 2188 29996
rect 1952 29844 2004 29850
rect 1952 29786 2004 29792
rect 2148 29481 2176 29990
rect 2240 29730 2268 30767
rect 2332 29850 2360 33866
rect 2424 32366 2452 34342
rect 2516 33930 2544 37606
rect 2700 36174 2728 38218
rect 2792 37369 2820 38898
rect 2884 37913 2912 39086
rect 2870 37904 2926 37913
rect 2870 37839 2926 37848
rect 2778 37360 2834 37369
rect 2778 37295 2834 37304
rect 2780 37256 2832 37262
rect 2780 37198 2832 37204
rect 2688 36168 2740 36174
rect 2688 36110 2740 36116
rect 2688 36032 2740 36038
rect 2688 35974 2740 35980
rect 2700 35698 2728 35974
rect 2688 35692 2740 35698
rect 2688 35634 2740 35640
rect 2700 34202 2728 35634
rect 2792 35465 2820 37198
rect 2872 36780 2924 36786
rect 2872 36722 2924 36728
rect 2778 35456 2834 35465
rect 2778 35391 2834 35400
rect 2780 35080 2832 35086
rect 2780 35022 2832 35028
rect 2792 34746 2820 35022
rect 2780 34740 2832 34746
rect 2780 34682 2832 34688
rect 2884 34649 2912 36722
rect 2870 34640 2926 34649
rect 2870 34575 2926 34584
rect 2872 34536 2924 34542
rect 2872 34478 2924 34484
rect 2688 34196 2740 34202
rect 2688 34138 2740 34144
rect 2780 33992 2832 33998
rect 2780 33934 2832 33940
rect 2504 33924 2556 33930
rect 2504 33866 2556 33872
rect 2688 33856 2740 33862
rect 2688 33798 2740 33804
rect 2700 33590 2728 33798
rect 2688 33584 2740 33590
rect 2688 33526 2740 33532
rect 2504 33516 2556 33522
rect 2504 33458 2556 33464
rect 2516 32881 2544 33458
rect 2596 33448 2648 33454
rect 2648 33408 2728 33436
rect 2596 33390 2648 33396
rect 2502 32872 2558 32881
rect 2502 32807 2558 32816
rect 2596 32768 2648 32774
rect 2700 32745 2728 33408
rect 2792 33017 2820 33934
rect 2884 33318 2912 34478
rect 2872 33312 2924 33318
rect 2872 33254 2924 33260
rect 2778 33008 2834 33017
rect 2778 32943 2834 32952
rect 2778 32872 2834 32881
rect 2778 32807 2834 32816
rect 2596 32710 2648 32716
rect 2686 32736 2742 32745
rect 2608 32570 2636 32710
rect 2686 32671 2742 32680
rect 2596 32564 2648 32570
rect 2596 32506 2648 32512
rect 2412 32360 2464 32366
rect 2412 32302 2464 32308
rect 2596 32360 2648 32366
rect 2596 32302 2648 32308
rect 2424 29850 2452 32302
rect 2608 32026 2636 32302
rect 2596 32020 2648 32026
rect 2596 31962 2648 31968
rect 2792 31906 2820 32807
rect 2884 32570 2912 33254
rect 2872 32564 2924 32570
rect 2872 32506 2924 32512
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 2700 31878 2820 31906
rect 2596 31340 2648 31346
rect 2596 31282 2648 31288
rect 2504 30728 2556 30734
rect 2504 30670 2556 30676
rect 2320 29844 2372 29850
rect 2320 29786 2372 29792
rect 2412 29844 2464 29850
rect 2412 29786 2464 29792
rect 2240 29702 2360 29730
rect 2228 29640 2280 29646
rect 2228 29582 2280 29588
rect 2134 29472 2190 29481
rect 2134 29407 2190 29416
rect 1872 29158 2176 29186
rect 1860 29028 1912 29034
rect 1860 28970 1912 28976
rect 2044 29028 2096 29034
rect 2044 28970 2096 28976
rect 1768 28076 1820 28082
rect 1768 28018 1820 28024
rect 1582 27976 1638 27985
rect 1582 27911 1638 27920
rect 1596 27402 1624 27911
rect 1584 27396 1636 27402
rect 1584 27338 1636 27344
rect 1596 26790 1624 27338
rect 1674 27160 1730 27169
rect 1674 27095 1730 27104
rect 1584 26784 1636 26790
rect 1584 26726 1636 26732
rect 1228 26438 1532 26466
rect 1584 26512 1636 26518
rect 1584 26454 1636 26460
rect 1122 23080 1178 23089
rect 1122 23015 1178 23024
rect 1228 22778 1256 26438
rect 1400 26376 1452 26382
rect 1596 26353 1624 26454
rect 1688 26382 1716 27095
rect 1676 26376 1728 26382
rect 1400 26318 1452 26324
rect 1582 26344 1638 26353
rect 1412 25673 1440 26318
rect 1676 26318 1728 26324
rect 1582 26279 1638 26288
rect 1676 26240 1728 26246
rect 1676 26182 1728 26188
rect 1492 25900 1544 25906
rect 1492 25842 1544 25848
rect 1398 25664 1454 25673
rect 1398 25599 1454 25608
rect 1504 25514 1532 25842
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1320 25486 1532 25514
rect 1596 25498 1624 25638
rect 1584 25492 1636 25498
rect 1320 24857 1348 25486
rect 1584 25434 1636 25440
rect 1688 25378 1716 26182
rect 1504 25350 1716 25378
rect 1306 24848 1362 24857
rect 1306 24783 1362 24792
rect 1400 24812 1452 24818
rect 1504 24800 1532 25350
rect 1676 25288 1728 25294
rect 1676 25230 1728 25236
rect 1584 25152 1636 25158
rect 1582 25120 1584 25129
rect 1636 25120 1638 25129
rect 1582 25055 1638 25064
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1452 24772 1532 24800
rect 1400 24754 1452 24760
rect 1308 24608 1360 24614
rect 1306 24576 1308 24585
rect 1360 24576 1362 24585
rect 1306 24511 1362 24520
rect 1308 23792 1360 23798
rect 1308 23734 1360 23740
rect 1320 23497 1348 23734
rect 1412 23662 1440 24754
rect 1492 23724 1544 23730
rect 1492 23666 1544 23672
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1306 23488 1362 23497
rect 1306 23423 1362 23432
rect 1412 23186 1440 23598
rect 1400 23180 1452 23186
rect 1400 23122 1452 23128
rect 1308 23044 1360 23050
rect 1308 22986 1360 22992
rect 1320 22953 1348 22986
rect 1306 22944 1362 22953
rect 1306 22879 1362 22888
rect 1216 22772 1268 22778
rect 1216 22714 1268 22720
rect 1044 22066 1164 22094
rect 846 21856 902 21865
rect 846 21791 902 21800
rect 860 21486 888 21791
rect 1032 21616 1084 21622
rect 1030 21584 1032 21593
rect 1084 21584 1086 21593
rect 1030 21519 1086 21528
rect 848 21480 900 21486
rect 848 21422 900 21428
rect 938 21312 994 21321
rect 938 21247 994 21256
rect 952 20942 980 21247
rect 940 20936 992 20942
rect 940 20878 992 20884
rect 768 19638 1072 19666
rect 938 19544 994 19553
rect 860 19502 938 19530
rect 754 19136 810 19145
rect 754 19071 810 19080
rect 768 18766 796 19071
rect 756 18760 808 18766
rect 756 18702 808 18708
rect 754 18592 810 18601
rect 754 18527 810 18536
rect 768 18358 796 18527
rect 756 18352 808 18358
rect 756 18294 808 18300
rect 860 17218 888 19502
rect 938 19479 994 19488
rect 938 18864 994 18873
rect 938 18799 940 18808
rect 992 18799 994 18808
rect 940 18770 992 18776
rect 938 17504 994 17513
rect 938 17439 994 17448
rect 952 17338 980 17439
rect 940 17332 992 17338
rect 940 17274 992 17280
rect 676 17190 796 17218
rect 860 17190 980 17218
rect 664 17128 716 17134
rect 664 17070 716 17076
rect 768 17082 796 17190
rect 572 2984 624 2990
rect 572 2926 624 2932
rect 676 2774 704 17070
rect 768 17054 888 17082
rect 756 16856 808 16862
rect 756 16798 808 16804
rect 768 11218 796 16798
rect 756 11212 808 11218
rect 756 11154 808 11160
rect 860 2774 888 17054
rect 952 6225 980 17190
rect 1044 13410 1072 19638
rect 1136 18986 1164 22066
rect 1228 20602 1256 22714
rect 1412 22642 1440 23122
rect 1504 22681 1532 23666
rect 1596 22692 1624 24890
rect 1688 24041 1716 25230
rect 1674 24032 1730 24041
rect 1674 23967 1730 23976
rect 1674 23760 1730 23769
rect 1674 23695 1676 23704
rect 1728 23695 1730 23704
rect 1676 23666 1728 23672
rect 1780 22794 1808 28018
rect 1872 27674 1900 28970
rect 1952 28756 2004 28762
rect 1952 28698 2004 28704
rect 1964 28422 1992 28698
rect 1952 28416 2004 28422
rect 1952 28358 2004 28364
rect 1860 27668 1912 27674
rect 1860 27610 1912 27616
rect 1872 24954 1900 27610
rect 1964 26466 1992 28358
rect 2056 28218 2084 28970
rect 2148 28937 2176 29158
rect 2134 28928 2190 28937
rect 2134 28863 2190 28872
rect 2044 28212 2096 28218
rect 2044 28154 2096 28160
rect 2148 28014 2176 28863
rect 2240 28150 2268 29582
rect 2332 29170 2360 29702
rect 2320 29164 2372 29170
rect 2320 29106 2372 29112
rect 2516 28994 2544 30670
rect 2608 29594 2636 31282
rect 2700 30734 2728 31878
rect 2780 31816 2832 31822
rect 2780 31758 2832 31764
rect 2792 31385 2820 31758
rect 2778 31376 2834 31385
rect 2778 31311 2834 31320
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2688 30728 2740 30734
rect 2688 30670 2740 30676
rect 2792 30394 2820 31214
rect 2780 30388 2832 30394
rect 2780 30330 2832 30336
rect 2688 30320 2740 30326
rect 2688 30262 2740 30268
rect 2700 29782 2728 30262
rect 2780 30252 2832 30258
rect 2780 30194 2832 30200
rect 2688 29776 2740 29782
rect 2792 29753 2820 30194
rect 2688 29718 2740 29724
rect 2778 29744 2834 29753
rect 2778 29679 2834 29688
rect 2608 29566 2728 29594
rect 2700 29510 2728 29566
rect 2596 29504 2648 29510
rect 2596 29446 2648 29452
rect 2688 29504 2740 29510
rect 2688 29446 2740 29452
rect 2608 29170 2636 29446
rect 2596 29164 2648 29170
rect 2596 29106 2648 29112
rect 2424 28966 2544 28994
rect 2320 28552 2372 28558
rect 2320 28494 2372 28500
rect 2228 28144 2280 28150
rect 2228 28086 2280 28092
rect 2136 28008 2188 28014
rect 2136 27950 2188 27956
rect 2332 27878 2360 28494
rect 2424 28257 2452 28966
rect 2504 28552 2556 28558
rect 2504 28494 2556 28500
rect 2688 28552 2740 28558
rect 2688 28494 2740 28500
rect 2410 28248 2466 28257
rect 2410 28183 2466 28192
rect 2516 28082 2544 28494
rect 2596 28416 2648 28422
rect 2596 28358 2648 28364
rect 2504 28076 2556 28082
rect 2504 28018 2556 28024
rect 2412 28008 2464 28014
rect 2412 27950 2464 27956
rect 2136 27872 2188 27878
rect 2136 27814 2188 27820
rect 2320 27872 2372 27878
rect 2320 27814 2372 27820
rect 2148 27130 2176 27814
rect 2228 27464 2280 27470
rect 2228 27406 2280 27412
rect 2136 27124 2188 27130
rect 2136 27066 2188 27072
rect 2044 26988 2096 26994
rect 2044 26930 2096 26936
rect 2136 26988 2188 26994
rect 2136 26930 2188 26936
rect 2056 26761 2084 26930
rect 2042 26752 2098 26761
rect 2042 26687 2098 26696
rect 2148 26586 2176 26930
rect 2240 26625 2268 27406
rect 2226 26616 2282 26625
rect 2136 26580 2188 26586
rect 2226 26551 2282 26560
rect 2136 26522 2188 26528
rect 2134 26480 2190 26489
rect 1964 26438 2084 26466
rect 1952 25288 2004 25294
rect 1952 25230 2004 25236
rect 1860 24948 1912 24954
rect 1860 24890 1912 24896
rect 1858 24848 1914 24857
rect 1858 24783 1914 24792
rect 1872 24138 1900 24783
rect 1964 24313 1992 25230
rect 1950 24304 2006 24313
rect 1950 24239 2006 24248
rect 2056 24154 2084 26438
rect 2134 26415 2190 26424
rect 2148 26042 2176 26415
rect 2136 26036 2188 26042
rect 2136 25978 2188 25984
rect 2134 25936 2190 25945
rect 2134 25871 2190 25880
rect 2228 25900 2280 25906
rect 2148 25430 2176 25871
rect 2228 25842 2280 25848
rect 2240 25809 2268 25842
rect 2226 25800 2282 25809
rect 2226 25735 2282 25744
rect 2332 25702 2360 27814
rect 2424 27418 2452 27950
rect 2608 27946 2636 28358
rect 2596 27940 2648 27946
rect 2596 27882 2648 27888
rect 2594 27568 2650 27577
rect 2594 27503 2650 27512
rect 2424 27390 2544 27418
rect 2412 27328 2464 27334
rect 2412 27270 2464 27276
rect 2424 26926 2452 27270
rect 2516 27112 2544 27390
rect 2608 27334 2636 27503
rect 2596 27328 2648 27334
rect 2596 27270 2648 27276
rect 2516 27084 2636 27112
rect 2504 26988 2556 26994
rect 2504 26930 2556 26936
rect 2412 26920 2464 26926
rect 2516 26897 2544 26930
rect 2412 26862 2464 26868
rect 2502 26888 2558 26897
rect 2502 26823 2558 26832
rect 2502 26208 2558 26217
rect 2502 26143 2558 26152
rect 2516 25906 2544 26143
rect 2504 25900 2556 25906
rect 2504 25842 2556 25848
rect 2410 25800 2466 25809
rect 2410 25735 2412 25744
rect 2464 25735 2466 25744
rect 2412 25706 2464 25712
rect 2228 25696 2280 25702
rect 2228 25638 2280 25644
rect 2320 25696 2372 25702
rect 2320 25638 2372 25644
rect 2136 25424 2188 25430
rect 2136 25366 2188 25372
rect 2240 24954 2268 25638
rect 2332 25430 2360 25638
rect 2320 25424 2372 25430
rect 2320 25366 2372 25372
rect 2228 24948 2280 24954
rect 2608 24936 2636 27084
rect 2700 26042 2728 28494
rect 2780 28076 2832 28082
rect 2780 28018 2832 28024
rect 2792 27305 2820 28018
rect 2884 27606 2912 32399
rect 2872 27600 2924 27606
rect 2872 27542 2924 27548
rect 2976 27554 3004 39986
rect 3068 39574 3096 42570
rect 3252 42362 3280 42570
rect 3240 42356 3292 42362
rect 3240 42298 3292 42304
rect 3240 40996 3292 41002
rect 3240 40938 3292 40944
rect 3252 40594 3280 40938
rect 3240 40588 3292 40594
rect 3240 40530 3292 40536
rect 3240 40384 3292 40390
rect 3240 40326 3292 40332
rect 3148 40180 3200 40186
rect 3148 40122 3200 40128
rect 3056 39568 3108 39574
rect 3056 39510 3108 39516
rect 3160 39370 3188 40122
rect 3252 39982 3280 40326
rect 3436 40118 3464 43658
rect 3528 43450 3556 43998
rect 3608 43852 3660 43858
rect 3608 43794 3660 43800
rect 3516 43444 3568 43450
rect 3516 43386 3568 43392
rect 3620 43314 3648 43794
rect 3608 43308 3660 43314
rect 3608 43250 3660 43256
rect 3608 42220 3660 42226
rect 3608 42162 3660 42168
rect 3516 41132 3568 41138
rect 3516 41074 3568 41080
rect 3424 40112 3476 40118
rect 3424 40054 3476 40060
rect 3332 40044 3384 40050
rect 3332 39986 3384 39992
rect 3240 39976 3292 39982
rect 3240 39918 3292 39924
rect 3148 39364 3200 39370
rect 3148 39306 3200 39312
rect 3056 39296 3108 39302
rect 3056 39238 3108 39244
rect 3068 38894 3096 39238
rect 3148 39092 3200 39098
rect 3148 39034 3200 39040
rect 3056 38888 3108 38894
rect 3056 38830 3108 38836
rect 3056 38412 3108 38418
rect 3056 38354 3108 38360
rect 3068 36281 3096 38354
rect 3160 37806 3188 39034
rect 3344 38978 3372 39986
rect 3436 39098 3464 40054
rect 3528 39522 3556 41074
rect 3620 40730 3648 42162
rect 3712 41698 3740 44934
rect 3790 44840 3846 45000
rect 4066 44840 4122 45000
rect 4342 44840 4398 45000
rect 4618 44840 4674 45000
rect 4894 44840 4950 45000
rect 5170 44840 5226 45000
rect 5446 44840 5502 45000
rect 5722 44840 5778 45000
rect 5998 44840 6054 45000
rect 6274 44840 6330 45000
rect 6550 44840 6606 45000
rect 6826 44962 6882 45000
rect 6748 44934 6882 44962
rect 3804 42566 3832 44840
rect 3976 43648 4028 43654
rect 3976 43590 4028 43596
rect 3988 43450 4016 43590
rect 3976 43444 4028 43450
rect 3976 43386 4028 43392
rect 4080 43194 4108 44840
rect 4356 44010 4384 44840
rect 4632 44062 4660 44840
rect 4620 44056 4672 44062
rect 4356 43982 4568 44010
rect 4620 43998 4672 44004
rect 4540 43314 4568 43982
rect 4804 43784 4856 43790
rect 4804 43726 4856 43732
rect 4160 43308 4212 43314
rect 4528 43308 4580 43314
rect 4212 43268 4476 43296
rect 4160 43250 4212 43256
rect 4080 43166 4292 43194
rect 3917 43004 4225 43013
rect 3917 43002 3923 43004
rect 3979 43002 4003 43004
rect 4059 43002 4083 43004
rect 4139 43002 4163 43004
rect 4219 43002 4225 43004
rect 3979 42950 3981 43002
rect 4161 42950 4163 43002
rect 3917 42948 3923 42950
rect 3979 42948 4003 42950
rect 4059 42948 4083 42950
rect 4139 42948 4163 42950
rect 4219 42948 4225 42950
rect 3917 42939 4225 42948
rect 4264 42922 4292 43166
rect 4264 42906 4384 42922
rect 4264 42900 4396 42906
rect 4264 42894 4344 42900
rect 4344 42842 4396 42848
rect 3792 42560 3844 42566
rect 3792 42502 3844 42508
rect 4448 42344 4476 43268
rect 4528 43250 4580 43256
rect 4620 43308 4672 43314
rect 4620 43250 4672 43256
rect 4528 42696 4580 42702
rect 4528 42638 4580 42644
rect 4264 42316 4476 42344
rect 3792 42220 3844 42226
rect 3792 42162 3844 42168
rect 3804 41818 3832 42162
rect 3917 41916 4225 41925
rect 3917 41914 3923 41916
rect 3979 41914 4003 41916
rect 4059 41914 4083 41916
rect 4139 41914 4163 41916
rect 4219 41914 4225 41916
rect 3979 41862 3981 41914
rect 4161 41862 4163 41914
rect 3917 41860 3923 41862
rect 3979 41860 4003 41862
rect 4059 41860 4083 41862
rect 4139 41860 4163 41862
rect 4219 41860 4225 41862
rect 3917 41851 4225 41860
rect 3792 41812 3844 41818
rect 3792 41754 3844 41760
rect 3884 41812 3936 41818
rect 3884 41754 3936 41760
rect 3896 41698 3924 41754
rect 3712 41670 3924 41698
rect 3700 41608 3752 41614
rect 3700 41550 3752 41556
rect 3884 41608 3936 41614
rect 3884 41550 3936 41556
rect 3608 40724 3660 40730
rect 3608 40666 3660 40672
rect 3606 39536 3662 39545
rect 3528 39494 3606 39522
rect 3606 39471 3662 39480
rect 3424 39092 3476 39098
rect 3424 39034 3476 39040
rect 3422 38992 3478 39001
rect 3240 38956 3292 38962
rect 3344 38950 3422 38978
rect 3478 38936 3648 38944
rect 3422 38927 3424 38936
rect 3240 38898 3292 38904
rect 3476 38916 3648 38936
rect 3424 38898 3476 38904
rect 3252 38654 3280 38898
rect 3252 38626 3556 38654
rect 3528 38350 3556 38626
rect 3240 38344 3292 38350
rect 3238 38312 3240 38321
rect 3516 38344 3568 38350
rect 3292 38312 3294 38321
rect 3516 38286 3568 38292
rect 3238 38247 3294 38256
rect 3332 37868 3384 37874
rect 3252 37828 3332 37856
rect 3148 37800 3200 37806
rect 3148 37742 3200 37748
rect 3148 37664 3200 37670
rect 3148 37606 3200 37612
rect 3054 36272 3110 36281
rect 3054 36207 3110 36216
rect 3056 36168 3108 36174
rect 3056 36110 3108 36116
rect 3068 35698 3096 36110
rect 3056 35692 3108 35698
rect 3056 35634 3108 35640
rect 3068 34542 3096 35634
rect 3160 35290 3188 37606
rect 3252 36553 3280 37828
rect 3332 37810 3384 37816
rect 3424 37800 3476 37806
rect 3424 37742 3476 37748
rect 3436 36922 3464 37742
rect 3528 37330 3556 38286
rect 3516 37324 3568 37330
rect 3516 37266 3568 37272
rect 3424 36916 3476 36922
rect 3424 36858 3476 36864
rect 3332 36712 3384 36718
rect 3332 36654 3384 36660
rect 3238 36544 3294 36553
rect 3238 36479 3294 36488
rect 3344 36378 3372 36654
rect 3332 36372 3384 36378
rect 3332 36314 3384 36320
rect 3436 36258 3464 36858
rect 3252 36230 3464 36258
rect 3148 35284 3200 35290
rect 3148 35226 3200 35232
rect 3160 35057 3188 35226
rect 3146 35048 3202 35057
rect 3146 34983 3202 34992
rect 3148 34740 3200 34746
rect 3252 34728 3280 36230
rect 3528 35986 3556 37266
rect 3620 36854 3648 38916
rect 3608 36848 3660 36854
rect 3608 36790 3660 36796
rect 3528 35958 3648 35986
rect 3516 35828 3568 35834
rect 3516 35770 3568 35776
rect 3332 35624 3384 35630
rect 3332 35566 3384 35572
rect 3200 34700 3280 34728
rect 3148 34682 3200 34688
rect 3056 34536 3108 34542
rect 3056 34478 3108 34484
rect 3056 33380 3108 33386
rect 3056 33322 3108 33328
rect 3068 32978 3096 33322
rect 3056 32972 3108 32978
rect 3056 32914 3108 32920
rect 3056 32836 3108 32842
rect 3056 32778 3108 32784
rect 3068 31249 3096 32778
rect 3054 31240 3110 31249
rect 3054 31175 3110 31184
rect 3056 31136 3108 31142
rect 3056 31078 3108 31084
rect 3068 30190 3096 31078
rect 3056 30184 3108 30190
rect 3056 30126 3108 30132
rect 3056 29640 3108 29646
rect 3056 29582 3108 29588
rect 3068 28393 3096 29582
rect 3054 28384 3110 28393
rect 3054 28319 3110 28328
rect 3056 28144 3108 28150
rect 3056 28086 3108 28092
rect 3068 27713 3096 28086
rect 3054 27704 3110 27713
rect 3054 27639 3110 27648
rect 2976 27526 3096 27554
rect 2964 27464 3016 27470
rect 2962 27432 2964 27441
rect 3016 27432 3018 27441
rect 2962 27367 3018 27376
rect 2778 27296 2834 27305
rect 2778 27231 2834 27240
rect 2962 27296 3018 27305
rect 2962 27231 3018 27240
rect 2870 26752 2926 26761
rect 2870 26687 2926 26696
rect 2884 26586 2912 26687
rect 2872 26580 2924 26586
rect 2872 26522 2924 26528
rect 2780 26444 2832 26450
rect 2780 26386 2832 26392
rect 2688 26036 2740 26042
rect 2688 25978 2740 25984
rect 2688 25288 2740 25294
rect 2686 25256 2688 25265
rect 2740 25256 2742 25265
rect 2686 25191 2742 25200
rect 2228 24890 2280 24896
rect 2516 24908 2636 24936
rect 2228 24812 2280 24818
rect 2228 24754 2280 24760
rect 2240 24206 2268 24754
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2424 24274 2452 24550
rect 2412 24268 2464 24274
rect 2412 24210 2464 24216
rect 1860 24132 1912 24138
rect 1860 24074 1912 24080
rect 1964 24126 2084 24154
rect 2228 24200 2280 24206
rect 2228 24142 2280 24148
rect 2136 24132 2188 24138
rect 1964 22930 1992 24126
rect 2136 24074 2188 24080
rect 2148 23866 2176 24074
rect 2228 24064 2280 24070
rect 2228 24006 2280 24012
rect 2136 23860 2188 23866
rect 2136 23802 2188 23808
rect 1964 22902 2084 22930
rect 1780 22766 1992 22794
rect 1490 22672 1546 22681
rect 1400 22636 1452 22642
rect 1596 22664 1808 22692
rect 1490 22607 1546 22616
rect 1400 22578 1452 22584
rect 1306 22264 1362 22273
rect 1306 22199 1308 22208
rect 1360 22199 1362 22208
rect 1308 22170 1360 22176
rect 1306 22128 1362 22137
rect 1306 22063 1362 22072
rect 1320 21978 1348 22063
rect 1674 21992 1730 22001
rect 1320 21950 1440 21978
rect 1412 21554 1440 21950
rect 1674 21927 1730 21936
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1688 21146 1716 21927
rect 1676 21140 1728 21146
rect 1676 21082 1728 21088
rect 1582 21040 1638 21049
rect 1582 20975 1638 20984
rect 1492 20868 1544 20874
rect 1492 20810 1544 20816
rect 1398 20768 1454 20777
rect 1398 20703 1454 20712
rect 1216 20596 1268 20602
rect 1216 20538 1268 20544
rect 1412 20466 1440 20703
rect 1504 20641 1532 20810
rect 1490 20632 1546 20641
rect 1490 20567 1546 20576
rect 1400 20460 1452 20466
rect 1400 20402 1452 20408
rect 1216 20392 1268 20398
rect 1216 20334 1268 20340
rect 1228 20233 1256 20334
rect 1214 20224 1270 20233
rect 1214 20159 1270 20168
rect 1306 19952 1362 19961
rect 1306 19887 1362 19896
rect 1320 19786 1348 19887
rect 1596 19854 1624 20975
rect 1780 20058 1808 22664
rect 1860 21956 1912 21962
rect 1860 21898 1912 21904
rect 1768 20052 1820 20058
rect 1768 19994 1820 20000
rect 1872 20040 1900 21898
rect 1964 20924 1992 22766
rect 2056 21962 2084 22902
rect 2044 21956 2096 21962
rect 2044 21898 2096 21904
rect 2136 21616 2188 21622
rect 2136 21558 2188 21564
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 2056 21078 2084 21490
rect 2148 21457 2176 21558
rect 2134 21448 2190 21457
rect 2134 21383 2190 21392
rect 2136 21344 2188 21350
rect 2136 21286 2188 21292
rect 2044 21072 2096 21078
rect 2044 21014 2096 21020
rect 2044 20936 2096 20942
rect 1964 20896 2044 20924
rect 2148 20913 2176 21286
rect 2044 20878 2096 20884
rect 2134 20904 2190 20913
rect 1952 20052 2004 20058
rect 1872 20012 1952 20040
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1676 19848 1728 19854
rect 1728 19796 1808 19802
rect 1676 19790 1808 19796
rect 1308 19780 1360 19786
rect 1688 19774 1808 19790
rect 1308 19722 1360 19728
rect 1584 19712 1636 19718
rect 1584 19654 1636 19660
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1308 19508 1360 19514
rect 1308 19450 1360 19456
rect 1320 19417 1348 19450
rect 1596 19417 1624 19654
rect 1306 19408 1362 19417
rect 1306 19343 1362 19352
rect 1582 19408 1638 19417
rect 1582 19343 1584 19352
rect 1636 19343 1638 19352
rect 1584 19314 1636 19320
rect 1136 18958 1256 18986
rect 1228 17082 1256 18958
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 1398 18048 1454 18057
rect 1398 17983 1454 17992
rect 1306 17776 1362 17785
rect 1306 17711 1362 17720
rect 1320 17270 1348 17711
rect 1308 17264 1360 17270
rect 1308 17206 1360 17212
rect 1136 17054 1256 17082
rect 1308 17060 1360 17066
rect 1136 16289 1164 17054
rect 1308 17002 1360 17008
rect 1320 16969 1348 17002
rect 1306 16960 1362 16969
rect 1306 16895 1362 16904
rect 1308 16788 1360 16794
rect 1308 16730 1360 16736
rect 1320 16697 1348 16730
rect 1306 16688 1362 16697
rect 1306 16623 1362 16632
rect 1122 16280 1178 16289
rect 1122 16215 1178 16224
rect 1412 15910 1440 17983
rect 1504 16182 1532 18906
rect 1582 18728 1638 18737
rect 1582 18663 1638 18672
rect 1596 18630 1624 18663
rect 1584 18624 1636 18630
rect 1584 18566 1636 18572
rect 1688 18358 1716 19654
rect 1780 19378 1808 19774
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1676 18352 1728 18358
rect 1676 18294 1728 18300
rect 1780 17864 1808 19314
rect 1872 18290 1900 20012
rect 1952 19994 2004 20000
rect 1952 18896 2004 18902
rect 1950 18864 1952 18873
rect 2004 18864 2006 18873
rect 1950 18799 2006 18808
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1688 17836 1808 17864
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1596 16810 1624 17478
rect 1688 16969 1716 17836
rect 1872 17814 1900 18226
rect 1964 18193 1992 18226
rect 1950 18184 2006 18193
rect 1950 18119 2006 18128
rect 1860 17808 1912 17814
rect 1766 17776 1822 17785
rect 1912 17768 1992 17796
rect 1860 17750 1912 17756
rect 1766 17711 1822 17720
rect 1780 17678 1808 17711
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1780 16998 1808 17614
rect 1860 17332 1912 17338
rect 1860 17274 1912 17280
rect 1872 17241 1900 17274
rect 1858 17232 1914 17241
rect 1858 17167 1914 17176
rect 1768 16992 1820 16998
rect 1674 16960 1730 16969
rect 1768 16934 1820 16940
rect 1674 16895 1730 16904
rect 1596 16782 1900 16810
rect 1676 16720 1728 16726
rect 1674 16688 1676 16697
rect 1728 16688 1730 16697
rect 1674 16623 1730 16632
rect 1686 16612 1716 16623
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1596 16250 1624 16526
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1492 16176 1544 16182
rect 1492 16118 1544 16124
rect 1582 16144 1638 16153
rect 1582 16079 1638 16088
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1398 15464 1454 15473
rect 1398 15399 1454 15408
rect 1308 14544 1360 14550
rect 1306 14512 1308 14521
rect 1360 14512 1362 14521
rect 1306 14447 1362 14456
rect 1308 14340 1360 14346
rect 1308 14282 1360 14288
rect 1320 13977 1348 14282
rect 1412 14074 1440 15399
rect 1490 14784 1546 14793
rect 1490 14719 1546 14728
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1306 13968 1362 13977
rect 1306 13903 1362 13912
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1306 13832 1362 13841
rect 1412 13818 1440 13874
rect 1504 13841 1532 14719
rect 1596 14618 1624 16079
rect 1688 14958 1716 16612
rect 1766 16416 1822 16425
rect 1766 16351 1822 16360
rect 1780 15162 1808 16351
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 1766 15056 1822 15065
rect 1766 14991 1822 15000
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1688 14328 1716 14894
rect 1596 14300 1716 14328
rect 1362 13790 1440 13818
rect 1490 13832 1546 13841
rect 1306 13767 1362 13776
rect 1490 13767 1546 13776
rect 1400 13728 1452 13734
rect 1400 13670 1452 13676
rect 1306 13424 1362 13433
rect 1044 13382 1306 13410
rect 1306 13359 1362 13368
rect 1412 12442 1440 13670
rect 1596 13394 1624 14300
rect 1674 14240 1730 14249
rect 1674 14175 1730 14184
rect 1584 13388 1636 13394
rect 1504 13348 1584 13376
rect 1400 12436 1452 12442
rect 1400 12378 1452 12384
rect 1504 12306 1532 13348
rect 1584 13330 1636 13336
rect 1688 12986 1716 14175
rect 1780 13530 1808 14991
rect 1872 14006 1900 16782
rect 1964 15638 1992 17768
rect 2056 16590 2084 20878
rect 2134 20839 2190 20848
rect 2136 20800 2188 20806
rect 2136 20742 2188 20748
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2056 15706 2084 16526
rect 2148 15994 2176 20742
rect 2240 20369 2268 24006
rect 2516 23322 2544 24908
rect 2594 24848 2650 24857
rect 2594 24783 2650 24792
rect 2608 23730 2636 24783
rect 2596 23724 2648 23730
rect 2596 23666 2648 23672
rect 2504 23316 2556 23322
rect 2504 23258 2556 23264
rect 2700 23118 2728 25191
rect 2792 24177 2820 26386
rect 2872 25696 2924 25702
rect 2872 25638 2924 25644
rect 2884 24274 2912 25638
rect 2976 24290 3004 27231
rect 3068 27130 3096 27526
rect 3056 27124 3108 27130
rect 3056 27066 3108 27072
rect 3056 25288 3108 25294
rect 3056 25230 3108 25236
rect 3068 24886 3096 25230
rect 3056 24880 3108 24886
rect 3056 24822 3108 24828
rect 3054 24712 3110 24721
rect 3054 24647 3110 24656
rect 3068 24410 3096 24647
rect 3160 24596 3188 34682
rect 3238 34096 3294 34105
rect 3238 34031 3294 34040
rect 3252 32570 3280 34031
rect 3240 32564 3292 32570
rect 3240 32506 3292 32512
rect 3344 31793 3372 35566
rect 3424 35488 3476 35494
rect 3424 35430 3476 35436
rect 3436 35154 3464 35430
rect 3424 35148 3476 35154
rect 3424 35090 3476 35096
rect 3424 34944 3476 34950
rect 3424 34886 3476 34892
rect 3436 34746 3464 34886
rect 3424 34740 3476 34746
rect 3424 34682 3476 34688
rect 3528 33096 3556 35770
rect 3620 34134 3648 35958
rect 3712 35290 3740 41550
rect 3896 41177 3924 41550
rect 4160 41540 4212 41546
rect 4160 41482 4212 41488
rect 4172 41274 4200 41482
rect 4160 41268 4212 41274
rect 4160 41210 4212 41216
rect 3882 41168 3938 41177
rect 3882 41103 3938 41112
rect 3792 40928 3844 40934
rect 3792 40870 3844 40876
rect 3804 40186 3832 40870
rect 3917 40828 4225 40837
rect 3917 40826 3923 40828
rect 3979 40826 4003 40828
rect 4059 40826 4083 40828
rect 4139 40826 4163 40828
rect 4219 40826 4225 40828
rect 3979 40774 3981 40826
rect 4161 40774 4163 40826
rect 3917 40772 3923 40774
rect 3979 40772 4003 40774
rect 4059 40772 4083 40774
rect 4139 40772 4163 40774
rect 4219 40772 4225 40774
rect 3917 40763 4225 40772
rect 4264 40730 4292 42316
rect 4436 42220 4488 42226
rect 4436 42162 4488 42168
rect 4344 41608 4396 41614
rect 4344 41550 4396 41556
rect 4252 40724 4304 40730
rect 4252 40666 4304 40672
rect 3976 40520 4028 40526
rect 3882 40488 3938 40497
rect 4252 40520 4304 40526
rect 3976 40462 4028 40468
rect 4158 40488 4214 40497
rect 3882 40423 3938 40432
rect 3896 40186 3924 40423
rect 3792 40180 3844 40186
rect 3792 40122 3844 40128
rect 3884 40180 3936 40186
rect 3884 40122 3936 40128
rect 3792 40044 3844 40050
rect 3792 39986 3844 39992
rect 3804 39098 3832 39986
rect 3988 39953 4016 40462
rect 4252 40462 4304 40468
rect 4158 40423 4160 40432
rect 4212 40423 4214 40432
rect 4160 40394 4212 40400
rect 4160 40180 4212 40186
rect 4160 40122 4212 40128
rect 3974 39944 4030 39953
rect 3974 39879 4030 39888
rect 4172 39828 4200 40122
rect 4264 40089 4292 40462
rect 4250 40080 4306 40089
rect 4250 40015 4306 40024
rect 4172 39800 4292 39828
rect 3917 39740 4225 39749
rect 3917 39738 3923 39740
rect 3979 39738 4003 39740
rect 4059 39738 4083 39740
rect 4139 39738 4163 39740
rect 4219 39738 4225 39740
rect 3979 39686 3981 39738
rect 4161 39686 4163 39738
rect 3917 39684 3923 39686
rect 3979 39684 4003 39686
rect 4059 39684 4083 39686
rect 4139 39684 4163 39686
rect 4219 39684 4225 39686
rect 3917 39675 4225 39684
rect 4264 39522 4292 39800
rect 4356 39642 4384 41550
rect 4448 41070 4476 42162
rect 4540 42090 4568 42638
rect 4528 42084 4580 42090
rect 4528 42026 4580 42032
rect 4632 41818 4660 43250
rect 4712 42696 4764 42702
rect 4816 42684 4844 43726
rect 4908 42752 4936 44840
rect 5184 43450 5212 44840
rect 5264 43648 5316 43654
rect 5264 43590 5316 43596
rect 5172 43444 5224 43450
rect 5172 43386 5224 43392
rect 4988 42764 5040 42770
rect 4908 42724 4988 42752
rect 4988 42706 5040 42712
rect 4816 42656 4936 42684
rect 4712 42638 4764 42644
rect 4620 41812 4672 41818
rect 4620 41754 4672 41760
rect 4724 41721 4752 42638
rect 4804 42016 4856 42022
rect 4804 41958 4856 41964
rect 4710 41712 4766 41721
rect 4528 41676 4580 41682
rect 4710 41647 4766 41656
rect 4528 41618 4580 41624
rect 4436 41064 4488 41070
rect 4436 41006 4488 41012
rect 4540 40118 4568 41618
rect 4620 41608 4672 41614
rect 4620 41550 4672 41556
rect 4528 40112 4580 40118
rect 4528 40054 4580 40060
rect 4344 39636 4396 39642
rect 4344 39578 4396 39584
rect 4436 39568 4488 39574
rect 4264 39494 4384 39522
rect 4436 39510 4488 39516
rect 4252 39432 4304 39438
rect 4252 39374 4304 39380
rect 3792 39092 3844 39098
rect 3792 39034 3844 39040
rect 3804 38962 3832 39034
rect 3792 38956 3844 38962
rect 3792 38898 3844 38904
rect 3804 36786 3832 38898
rect 4264 38894 4292 39374
rect 4356 39030 4384 39494
rect 4344 39024 4396 39030
rect 4344 38966 4396 38972
rect 4252 38888 4304 38894
rect 4252 38830 4304 38836
rect 3917 38652 4225 38661
rect 3917 38650 3923 38652
rect 3979 38650 4003 38652
rect 4059 38650 4083 38652
rect 4139 38650 4163 38652
rect 4219 38650 4225 38652
rect 3979 38598 3981 38650
rect 4161 38598 4163 38650
rect 3917 38596 3923 38598
rect 3979 38596 4003 38598
rect 4059 38596 4083 38598
rect 4139 38596 4163 38598
rect 4219 38596 4225 38598
rect 3917 38587 4225 38596
rect 4068 38344 4120 38350
rect 4068 38286 4120 38292
rect 4080 37913 4108 38286
rect 4066 37904 4122 37913
rect 4066 37839 4068 37848
rect 4120 37839 4122 37848
rect 4068 37810 4120 37816
rect 4160 37800 4212 37806
rect 4158 37768 4160 37777
rect 4212 37768 4214 37777
rect 4158 37703 4214 37712
rect 3917 37564 4225 37573
rect 3917 37562 3923 37564
rect 3979 37562 4003 37564
rect 4059 37562 4083 37564
rect 4139 37562 4163 37564
rect 4219 37562 4225 37564
rect 3979 37510 3981 37562
rect 4161 37510 4163 37562
rect 3917 37508 3923 37510
rect 3979 37508 4003 37510
rect 4059 37508 4083 37510
rect 4139 37508 4163 37510
rect 4219 37508 4225 37510
rect 3917 37499 4225 37508
rect 4356 37398 4384 38966
rect 4448 38740 4476 39510
rect 4528 39500 4580 39506
rect 4528 39442 4580 39448
rect 4540 39030 4568 39442
rect 4528 39024 4580 39030
rect 4528 38966 4580 38972
rect 4528 38752 4580 38758
rect 4448 38712 4528 38740
rect 4528 38694 4580 38700
rect 4540 37890 4568 38694
rect 4632 38049 4660 41550
rect 4816 41546 4844 41958
rect 4804 41540 4856 41546
rect 4804 41482 4856 41488
rect 4908 41414 4936 42656
rect 5172 41608 5224 41614
rect 5170 41576 5172 41585
rect 5224 41576 5226 41585
rect 5170 41511 5226 41520
rect 4816 41386 4936 41414
rect 4816 41274 4844 41386
rect 5276 41274 5304 43590
rect 5460 43450 5488 44840
rect 5736 43450 5764 44840
rect 6012 43738 6040 44840
rect 6012 43710 6132 43738
rect 5448 43444 5500 43450
rect 5448 43386 5500 43392
rect 5724 43444 5776 43450
rect 5724 43386 5776 43392
rect 5448 43308 5500 43314
rect 5448 43250 5500 43256
rect 5460 41818 5488 43250
rect 5540 43104 5592 43110
rect 5540 43046 5592 43052
rect 5552 42702 5580 43046
rect 6104 42906 6132 43710
rect 6092 42900 6144 42906
rect 6092 42842 6144 42848
rect 5540 42696 5592 42702
rect 5540 42638 5592 42644
rect 6000 42628 6052 42634
rect 6000 42570 6052 42576
rect 5540 42560 5592 42566
rect 5540 42502 5592 42508
rect 5448 41812 5500 41818
rect 5448 41754 5500 41760
rect 5552 41274 5580 42502
rect 5632 42356 5684 42362
rect 5632 42298 5684 42304
rect 5644 41414 5672 42298
rect 5816 42288 5868 42294
rect 5816 42230 5868 42236
rect 5724 42016 5776 42022
rect 5724 41958 5776 41964
rect 5736 41818 5764 41958
rect 5828 41818 5856 42230
rect 5908 42084 5960 42090
rect 5908 42026 5960 42032
rect 5724 41812 5776 41818
rect 5724 41754 5776 41760
rect 5816 41812 5868 41818
rect 5816 41754 5868 41760
rect 5920 41546 5948 42026
rect 6012 41818 6040 42570
rect 6288 42566 6316 44840
rect 6368 43852 6420 43858
rect 6368 43794 6420 43800
rect 6380 43330 6408 43794
rect 6564 43738 6592 44840
rect 6564 43710 6684 43738
rect 6380 43302 6500 43330
rect 6368 43240 6420 43246
rect 6368 43182 6420 43188
rect 6276 42560 6328 42566
rect 6276 42502 6328 42508
rect 6092 42220 6144 42226
rect 6092 42162 6144 42168
rect 6184 42220 6236 42226
rect 6184 42162 6236 42168
rect 6000 41812 6052 41818
rect 6000 41754 6052 41760
rect 6000 41608 6052 41614
rect 6000 41550 6052 41556
rect 5908 41540 5960 41546
rect 5908 41482 5960 41488
rect 5644 41386 5856 41414
rect 5828 41274 5856 41386
rect 4804 41268 4856 41274
rect 4804 41210 4856 41216
rect 5264 41268 5316 41274
rect 5264 41210 5316 41216
rect 5540 41268 5592 41274
rect 5540 41210 5592 41216
rect 5816 41268 5868 41274
rect 5816 41210 5868 41216
rect 5080 41132 5132 41138
rect 4908 41092 5080 41120
rect 4712 41064 4764 41070
rect 4712 41006 4764 41012
rect 4618 38040 4674 38049
rect 4618 37975 4674 37984
rect 4540 37862 4660 37890
rect 4528 37800 4580 37806
rect 4528 37742 4580 37748
rect 4436 37664 4488 37670
rect 4436 37606 4488 37612
rect 4344 37392 4396 37398
rect 4344 37334 4396 37340
rect 3884 37256 3936 37262
rect 3884 37198 3936 37204
rect 3896 36825 3924 37198
rect 4356 36854 4384 37334
rect 4160 36848 4212 36854
rect 3882 36816 3938 36825
rect 3792 36780 3844 36786
rect 4344 36848 4396 36854
rect 4212 36796 4292 36802
rect 4160 36790 4292 36796
rect 4344 36790 4396 36796
rect 4172 36774 4292 36790
rect 4448 36786 4476 37606
rect 4540 37330 4568 37742
rect 4528 37324 4580 37330
rect 4528 37266 4580 37272
rect 4528 37188 4580 37194
rect 4528 37130 4580 37136
rect 3882 36751 3938 36760
rect 3792 36722 3844 36728
rect 3804 36258 3832 36722
rect 3917 36476 4225 36485
rect 3917 36474 3923 36476
rect 3979 36474 4003 36476
rect 4059 36474 4083 36476
rect 4139 36474 4163 36476
rect 4219 36474 4225 36476
rect 3979 36422 3981 36474
rect 4161 36422 4163 36474
rect 3917 36420 3923 36422
rect 3979 36420 4003 36422
rect 4059 36420 4083 36422
rect 4139 36420 4163 36422
rect 4219 36420 4225 36422
rect 3917 36411 4225 36420
rect 3804 36230 3924 36258
rect 3792 36168 3844 36174
rect 3792 36110 3844 36116
rect 3804 35873 3832 36110
rect 3896 35986 3924 36230
rect 4068 36100 4120 36106
rect 4068 36042 4120 36048
rect 3974 36000 4030 36009
rect 3896 35958 3974 35986
rect 3974 35935 4030 35944
rect 3790 35864 3846 35873
rect 3790 35799 3846 35808
rect 4080 35601 4108 36042
rect 4160 36032 4212 36038
rect 4160 35974 4212 35980
rect 4172 35630 4200 35974
rect 4160 35624 4212 35630
rect 4066 35592 4122 35601
rect 4160 35566 4212 35572
rect 4066 35527 4122 35536
rect 3917 35388 4225 35397
rect 3917 35386 3923 35388
rect 3979 35386 4003 35388
rect 4059 35386 4083 35388
rect 4139 35386 4163 35388
rect 4219 35386 4225 35388
rect 3979 35334 3981 35386
rect 4161 35334 4163 35386
rect 3917 35332 3923 35334
rect 3979 35332 4003 35334
rect 4059 35332 4083 35334
rect 4139 35332 4163 35334
rect 4219 35332 4225 35334
rect 3917 35323 4225 35332
rect 3700 35284 3752 35290
rect 3700 35226 3752 35232
rect 4264 35086 4292 36774
rect 4436 36780 4488 36786
rect 4436 36722 4488 36728
rect 4344 36644 4396 36650
rect 4344 36586 4396 36592
rect 4356 36378 4384 36586
rect 4436 36576 4488 36582
rect 4436 36518 4488 36524
rect 4344 36372 4396 36378
rect 4344 36314 4396 36320
rect 4448 36310 4476 36518
rect 4436 36304 4488 36310
rect 4342 36272 4398 36281
rect 4398 36252 4436 36258
rect 4540 36281 4568 37130
rect 4632 36310 4660 37862
rect 4620 36304 4672 36310
rect 4398 36246 4488 36252
rect 4526 36272 4582 36281
rect 4398 36230 4476 36246
rect 4342 36207 4398 36216
rect 4620 36246 4672 36252
rect 4526 36207 4582 36216
rect 4344 36168 4396 36174
rect 4344 36110 4396 36116
rect 4436 36168 4488 36174
rect 4436 36110 4488 36116
rect 4356 35737 4384 36110
rect 4342 35728 4398 35737
rect 4342 35663 4398 35672
rect 4068 35080 4120 35086
rect 3790 35048 3846 35057
rect 3712 35006 3790 35034
rect 3608 34128 3660 34134
rect 3608 34070 3660 34076
rect 3436 33068 3556 33096
rect 3330 31784 3386 31793
rect 3330 31719 3386 31728
rect 3240 31680 3292 31686
rect 3240 31622 3292 31628
rect 3252 30433 3280 31622
rect 3332 30592 3384 30598
rect 3332 30534 3384 30540
rect 3238 30424 3294 30433
rect 3344 30394 3372 30534
rect 3238 30359 3294 30368
rect 3332 30388 3384 30394
rect 3436 30376 3464 33068
rect 3606 33008 3662 33017
rect 3516 32972 3568 32978
rect 3606 32943 3662 32952
rect 3516 32914 3568 32920
rect 3528 30598 3556 32914
rect 3620 32910 3648 32943
rect 3608 32904 3660 32910
rect 3608 32846 3660 32852
rect 3712 32774 3740 35006
rect 4068 35022 4120 35028
rect 4252 35080 4304 35086
rect 4252 35022 4304 35028
rect 3790 34983 3846 34992
rect 4080 34678 4108 35022
rect 4160 35012 4212 35018
rect 4160 34954 4212 34960
rect 4172 34746 4200 34954
rect 4160 34740 4212 34746
rect 4160 34682 4212 34688
rect 4068 34672 4120 34678
rect 4068 34614 4120 34620
rect 4344 34604 4396 34610
rect 4344 34546 4396 34552
rect 3917 34300 4225 34309
rect 3917 34298 3923 34300
rect 3979 34298 4003 34300
rect 4059 34298 4083 34300
rect 4139 34298 4163 34300
rect 4219 34298 4225 34300
rect 3979 34246 3981 34298
rect 4161 34246 4163 34298
rect 3917 34244 3923 34246
rect 3979 34244 4003 34246
rect 4059 34244 4083 34246
rect 4139 34244 4163 34246
rect 4219 34244 4225 34246
rect 3917 34235 4225 34244
rect 3792 33992 3844 33998
rect 3792 33934 3844 33940
rect 3884 33992 3936 33998
rect 3884 33934 3936 33940
rect 3804 33425 3832 33934
rect 3896 33833 3924 33934
rect 4252 33924 4304 33930
rect 4252 33866 4304 33872
rect 3882 33824 3938 33833
rect 3882 33759 3938 33768
rect 3790 33416 3846 33425
rect 4264 33402 4292 33866
rect 4356 33522 4384 34546
rect 4344 33516 4396 33522
rect 4344 33458 4396 33464
rect 4264 33374 4384 33402
rect 3790 33351 3846 33360
rect 3884 33312 3936 33318
rect 3804 33272 3884 33300
rect 3804 32978 3832 33272
rect 3884 33254 3936 33260
rect 4252 33312 4304 33318
rect 4252 33254 4304 33260
rect 3917 33212 4225 33221
rect 3917 33210 3923 33212
rect 3979 33210 4003 33212
rect 4059 33210 4083 33212
rect 4139 33210 4163 33212
rect 4219 33210 4225 33212
rect 3979 33158 3981 33210
rect 4161 33158 4163 33210
rect 3917 33156 3923 33158
rect 3979 33156 4003 33158
rect 4059 33156 4083 33158
rect 4139 33156 4163 33158
rect 4219 33156 4225 33158
rect 3917 33147 4225 33156
rect 3792 32972 3844 32978
rect 3792 32914 3844 32920
rect 4264 32910 4292 33254
rect 4356 33153 4384 33374
rect 4342 33144 4398 33153
rect 4342 33079 4398 33088
rect 3884 32904 3936 32910
rect 4252 32904 4304 32910
rect 3884 32846 3936 32852
rect 3974 32872 4030 32881
rect 3608 32768 3660 32774
rect 3608 32710 3660 32716
rect 3700 32768 3752 32774
rect 3700 32710 3752 32716
rect 3620 32570 3648 32710
rect 3608 32564 3660 32570
rect 3608 32506 3660 32512
rect 3896 32212 3924 32846
rect 4252 32846 4304 32852
rect 4344 32904 4396 32910
rect 4344 32846 4396 32852
rect 3974 32807 4030 32816
rect 3988 32434 4016 32807
rect 4356 32570 4384 32846
rect 4344 32564 4396 32570
rect 4344 32506 4396 32512
rect 4252 32496 4304 32502
rect 4252 32438 4304 32444
rect 3976 32428 4028 32434
rect 3976 32370 4028 32376
rect 4264 32337 4292 32438
rect 4250 32328 4306 32337
rect 4250 32263 4306 32272
rect 3804 32184 3924 32212
rect 3608 30932 3660 30938
rect 3608 30874 3660 30880
rect 3516 30592 3568 30598
rect 3620 30569 3648 30874
rect 3516 30534 3568 30540
rect 3606 30560 3662 30569
rect 3606 30495 3662 30504
rect 3436 30348 3740 30376
rect 3332 30330 3384 30336
rect 3240 30252 3292 30258
rect 3240 30194 3292 30200
rect 3424 30252 3476 30258
rect 3424 30194 3476 30200
rect 3252 25362 3280 30194
rect 3436 29322 3464 30194
rect 3608 29844 3660 29850
rect 3608 29786 3660 29792
rect 3516 29708 3568 29714
rect 3516 29650 3568 29656
rect 3344 29294 3464 29322
rect 3344 26450 3372 29294
rect 3528 29220 3556 29650
rect 3620 29628 3648 29786
rect 3712 29696 3740 30348
rect 3804 29850 3832 32184
rect 3917 32124 4225 32133
rect 3917 32122 3923 32124
rect 3979 32122 4003 32124
rect 4059 32122 4083 32124
rect 4139 32122 4163 32124
rect 4219 32122 4225 32124
rect 3979 32070 3981 32122
rect 4161 32070 4163 32122
rect 3917 32068 3923 32070
rect 3979 32068 4003 32070
rect 4059 32068 4083 32070
rect 4139 32068 4163 32070
rect 4219 32068 4225 32070
rect 3917 32059 4225 32068
rect 3884 31476 3936 31482
rect 3884 31418 3936 31424
rect 3896 31385 3924 31418
rect 3882 31376 3938 31385
rect 3882 31311 3938 31320
rect 3917 31036 4225 31045
rect 3917 31034 3923 31036
rect 3979 31034 4003 31036
rect 4059 31034 4083 31036
rect 4139 31034 4163 31036
rect 4219 31034 4225 31036
rect 3979 30982 3981 31034
rect 4161 30982 4163 31034
rect 3917 30980 3923 30982
rect 3979 30980 4003 30982
rect 4059 30980 4083 30982
rect 4139 30980 4163 30982
rect 4219 30980 4225 30982
rect 3917 30971 4225 30980
rect 3976 30728 4028 30734
rect 3976 30670 4028 30676
rect 3988 30394 4016 30670
rect 4068 30592 4120 30598
rect 4068 30534 4120 30540
rect 3976 30388 4028 30394
rect 3976 30330 4028 30336
rect 4080 30036 4108 30534
rect 4264 30326 4292 32263
rect 4344 31748 4396 31754
rect 4344 31690 4396 31696
rect 4252 30320 4304 30326
rect 4252 30262 4304 30268
rect 4080 30008 4292 30036
rect 3917 29948 4225 29957
rect 3917 29946 3923 29948
rect 3979 29946 4003 29948
rect 4059 29946 4083 29948
rect 4139 29946 4163 29948
rect 4219 29946 4225 29948
rect 3979 29894 3981 29946
rect 4161 29894 4163 29946
rect 3917 29892 3923 29894
rect 3979 29892 4003 29894
rect 4059 29892 4083 29894
rect 4139 29892 4163 29894
rect 4219 29892 4225 29894
rect 3917 29883 4225 29892
rect 3792 29844 3844 29850
rect 3792 29786 3844 29792
rect 4068 29708 4120 29714
rect 3712 29668 3924 29696
rect 3620 29600 3832 29628
rect 3700 29504 3752 29510
rect 3700 29446 3752 29452
rect 3436 29192 3556 29220
rect 3332 26444 3384 26450
rect 3332 26386 3384 26392
rect 3240 25356 3292 25362
rect 3240 25298 3292 25304
rect 3332 25152 3384 25158
rect 3332 25094 3384 25100
rect 3344 24750 3372 25094
rect 3436 24886 3464 29192
rect 3516 28960 3568 28966
rect 3516 28902 3568 28908
rect 3608 28960 3660 28966
rect 3608 28902 3660 28908
rect 3528 28218 3556 28902
rect 3620 28762 3648 28902
rect 3608 28756 3660 28762
rect 3608 28698 3660 28704
rect 3516 28212 3568 28218
rect 3516 28154 3568 28160
rect 3606 28112 3662 28121
rect 3528 28070 3606 28098
rect 3424 24880 3476 24886
rect 3424 24822 3476 24828
rect 3332 24744 3384 24750
rect 3332 24686 3384 24692
rect 3160 24568 3372 24596
rect 3056 24404 3108 24410
rect 3056 24346 3108 24352
rect 3148 24404 3200 24410
rect 3148 24346 3200 24352
rect 2872 24268 2924 24274
rect 2976 24262 3096 24290
rect 2872 24210 2924 24216
rect 2778 24168 2834 24177
rect 2778 24103 2834 24112
rect 2792 23526 2820 24103
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2688 23112 2740 23118
rect 2688 23054 2740 23060
rect 2412 22976 2464 22982
rect 2412 22918 2464 22924
rect 2424 22522 2452 22918
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2792 22545 2820 22578
rect 2332 22494 2452 22522
rect 2778 22536 2834 22545
rect 2332 22098 2360 22494
rect 2778 22471 2834 22480
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2424 22030 2452 22374
rect 2686 22264 2742 22273
rect 2742 22234 2820 22250
rect 2742 22228 2832 22234
rect 2742 22222 2780 22228
rect 2686 22199 2742 22208
rect 2780 22170 2832 22176
rect 2412 22024 2464 22030
rect 2412 21966 2464 21972
rect 2412 21888 2464 21894
rect 2412 21830 2464 21836
rect 2778 21856 2834 21865
rect 2320 21344 2372 21350
rect 2424 21332 2452 21830
rect 2778 21791 2834 21800
rect 2596 21616 2648 21622
rect 2596 21558 2648 21564
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 2372 21304 2452 21332
rect 2320 21286 2372 21292
rect 2424 20584 2452 21304
rect 2516 20806 2544 21490
rect 2608 20874 2636 21558
rect 2596 20868 2648 20874
rect 2596 20810 2648 20816
rect 2688 20868 2740 20874
rect 2688 20810 2740 20816
rect 2504 20800 2556 20806
rect 2504 20742 2556 20748
rect 2596 20596 2648 20602
rect 2424 20556 2596 20584
rect 2596 20538 2648 20544
rect 2700 20482 2728 20810
rect 2792 20534 2820 21791
rect 2884 21010 2912 24210
rect 2964 24132 3016 24138
rect 2964 24074 3016 24080
rect 2976 22506 3004 24074
rect 2964 22500 3016 22506
rect 2964 22442 3016 22448
rect 2976 21894 3004 22442
rect 2964 21888 3016 21894
rect 2964 21830 3016 21836
rect 3068 21554 3096 24262
rect 3160 22642 3188 24346
rect 3240 24064 3292 24070
rect 3240 24006 3292 24012
rect 3148 22636 3200 22642
rect 3148 22578 3200 22584
rect 3252 21865 3280 24006
rect 3238 21856 3294 21865
rect 3238 21791 3294 21800
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 3056 20800 3108 20806
rect 3056 20742 3108 20748
rect 2608 20454 2728 20482
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 2964 20460 3016 20466
rect 2226 20360 2282 20369
rect 2226 20295 2282 20304
rect 2608 19417 2636 20454
rect 2964 20402 3016 20408
rect 2688 19984 2740 19990
rect 2688 19926 2740 19932
rect 2594 19408 2650 19417
rect 2594 19343 2650 19352
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2228 18352 2280 18358
rect 2228 18294 2280 18300
rect 2240 17542 2268 18294
rect 2332 18222 2360 19110
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2332 17660 2360 18158
rect 2424 17814 2452 19110
rect 2608 18698 2636 19343
rect 2596 18692 2648 18698
rect 2596 18634 2648 18640
rect 2700 18034 2728 19926
rect 2872 19372 2924 19378
rect 2872 19314 2924 19320
rect 2780 18624 2832 18630
rect 2884 18601 2912 19314
rect 2976 18850 3004 20402
rect 3068 20398 3096 20742
rect 3252 20466 3280 21286
rect 3344 20534 3372 24568
rect 3436 23866 3464 24822
rect 3528 23866 3556 28070
rect 3606 28047 3662 28056
rect 3712 27674 3740 29446
rect 3804 28422 3832 29600
rect 3896 29170 3924 29668
rect 4120 29668 4200 29696
rect 4068 29650 4120 29656
rect 3884 29164 3936 29170
rect 3884 29106 3936 29112
rect 4172 29102 4200 29668
rect 4264 29646 4292 30008
rect 4252 29640 4304 29646
rect 4252 29582 4304 29588
rect 4160 29096 4212 29102
rect 4160 29038 4212 29044
rect 3917 28860 4225 28869
rect 3917 28858 3923 28860
rect 3979 28858 4003 28860
rect 4059 28858 4083 28860
rect 4139 28858 4163 28860
rect 4219 28858 4225 28860
rect 3979 28806 3981 28858
rect 4161 28806 4163 28858
rect 3917 28804 3923 28806
rect 3979 28804 4003 28806
rect 4059 28804 4083 28806
rect 4139 28804 4163 28806
rect 4219 28804 4225 28806
rect 3917 28795 4225 28804
rect 4356 28608 4384 31690
rect 4264 28580 4384 28608
rect 3882 28520 3938 28529
rect 3882 28455 3884 28464
rect 3936 28455 3938 28464
rect 3884 28426 3936 28432
rect 3792 28416 3844 28422
rect 3792 28358 3844 28364
rect 4264 28098 4292 28580
rect 4344 28484 4396 28490
rect 4344 28426 4396 28432
rect 4356 28218 4384 28426
rect 4344 28212 4396 28218
rect 4344 28154 4396 28160
rect 4264 28070 4384 28098
rect 4252 27872 4304 27878
rect 3790 27840 3846 27849
rect 4252 27814 4304 27820
rect 3790 27775 3846 27784
rect 3608 27668 3660 27674
rect 3608 27610 3660 27616
rect 3700 27668 3752 27674
rect 3700 27610 3752 27616
rect 3620 27577 3648 27610
rect 3606 27568 3662 27577
rect 3606 27503 3662 27512
rect 3804 27470 3832 27775
rect 3917 27772 4225 27781
rect 3917 27770 3923 27772
rect 3979 27770 4003 27772
rect 4059 27770 4083 27772
rect 4139 27770 4163 27772
rect 4219 27770 4225 27772
rect 3979 27718 3981 27770
rect 4161 27718 4163 27770
rect 3917 27716 3923 27718
rect 3979 27716 4003 27718
rect 4059 27716 4083 27718
rect 4139 27716 4163 27718
rect 4219 27716 4225 27718
rect 3917 27707 4225 27716
rect 4160 27532 4212 27538
rect 4160 27474 4212 27480
rect 3792 27464 3844 27470
rect 3792 27406 3844 27412
rect 4172 26994 4200 27474
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 3917 26684 4225 26693
rect 3917 26682 3923 26684
rect 3979 26682 4003 26684
rect 4059 26682 4083 26684
rect 4139 26682 4163 26684
rect 4219 26682 4225 26684
rect 3979 26630 3981 26682
rect 4161 26630 4163 26682
rect 3917 26628 3923 26630
rect 3979 26628 4003 26630
rect 4059 26628 4083 26630
rect 4139 26628 4163 26630
rect 4219 26628 4225 26630
rect 3917 26619 4225 26628
rect 3606 26072 3662 26081
rect 4158 26072 4214 26081
rect 3662 26030 3740 26058
rect 3606 26007 3662 26016
rect 3608 25356 3660 25362
rect 3608 25298 3660 25304
rect 3620 24290 3648 25298
rect 3712 24818 3740 26030
rect 4158 26007 4214 26016
rect 4068 25968 4120 25974
rect 4172 25956 4200 26007
rect 4264 25974 4292 27814
rect 4356 27538 4384 28070
rect 4448 27878 4476 36110
rect 4724 35834 4752 41006
rect 4804 40452 4856 40458
rect 4804 40394 4856 40400
rect 4816 39982 4844 40394
rect 4804 39976 4856 39982
rect 4804 39918 4856 39924
rect 4804 38956 4856 38962
rect 4804 38898 4856 38904
rect 4816 38554 4844 38898
rect 4804 38548 4856 38554
rect 4804 38490 4856 38496
rect 4802 36000 4858 36009
rect 4802 35935 4858 35944
rect 4712 35828 4764 35834
rect 4712 35770 4764 35776
rect 4528 35624 4580 35630
rect 4528 35566 4580 35572
rect 4540 34950 4568 35566
rect 4620 35556 4672 35562
rect 4672 35516 4752 35544
rect 4620 35498 4672 35504
rect 4618 35048 4674 35057
rect 4618 34983 4674 34992
rect 4528 34944 4580 34950
rect 4528 34886 4580 34892
rect 4632 34746 4660 34983
rect 4620 34740 4672 34746
rect 4620 34682 4672 34688
rect 4528 34604 4580 34610
rect 4528 34546 4580 34552
rect 4540 31142 4568 34546
rect 4620 34196 4672 34202
rect 4620 34138 4672 34144
rect 4632 32065 4660 34138
rect 4618 32056 4674 32065
rect 4618 31991 4674 32000
rect 4632 31754 4660 31991
rect 4620 31748 4672 31754
rect 4620 31690 4672 31696
rect 4618 31512 4674 31521
rect 4618 31447 4620 31456
rect 4672 31447 4674 31456
rect 4620 31418 4672 31424
rect 4620 31204 4672 31210
rect 4620 31146 4672 31152
rect 4528 31136 4580 31142
rect 4632 31113 4660 31146
rect 4528 31078 4580 31084
rect 4618 31104 4674 31113
rect 4540 29594 4568 31078
rect 4618 31039 4674 31048
rect 4724 30376 4752 35516
rect 4816 35018 4844 35935
rect 4804 35012 4856 35018
rect 4804 34954 4856 34960
rect 4816 34921 4844 34954
rect 4802 34912 4858 34921
rect 4802 34847 4858 34856
rect 4804 34672 4856 34678
rect 4804 34614 4856 34620
rect 4816 33386 4844 34614
rect 4804 33380 4856 33386
rect 4804 33322 4856 33328
rect 4804 31748 4856 31754
rect 4804 31690 4856 31696
rect 4816 31346 4844 31690
rect 4804 31340 4856 31346
rect 4804 31282 4856 31288
rect 4804 31136 4856 31142
rect 4804 31078 4856 31084
rect 4816 30938 4844 31078
rect 4804 30932 4856 30938
rect 4804 30874 4856 30880
rect 4802 30832 4858 30841
rect 4802 30767 4858 30776
rect 4816 30598 4844 30767
rect 4908 30734 4936 41092
rect 5080 41074 5132 41080
rect 5448 41132 5500 41138
rect 5448 41074 5500 41080
rect 5540 41132 5592 41138
rect 5540 41074 5592 41080
rect 5264 40520 5316 40526
rect 5264 40462 5316 40468
rect 5276 40361 5304 40462
rect 5356 40384 5408 40390
rect 5262 40352 5318 40361
rect 5356 40326 5408 40332
rect 5262 40287 5318 40296
rect 5276 40186 5304 40287
rect 5264 40180 5316 40186
rect 5264 40122 5316 40128
rect 4988 40112 5040 40118
rect 4988 40054 5040 40060
rect 5000 37398 5028 40054
rect 5172 39840 5224 39846
rect 5172 39782 5224 39788
rect 5184 39438 5212 39782
rect 5368 39642 5396 40326
rect 5460 40225 5488 41074
rect 5446 40216 5502 40225
rect 5446 40151 5502 40160
rect 5356 39636 5408 39642
rect 5356 39578 5408 39584
rect 5172 39432 5224 39438
rect 5092 39392 5172 39420
rect 4988 37392 5040 37398
rect 4988 37334 5040 37340
rect 4988 36848 5040 36854
rect 4988 36790 5040 36796
rect 5000 35034 5028 36790
rect 5092 36174 5120 39392
rect 5172 39374 5224 39380
rect 5356 38956 5408 38962
rect 5356 38898 5408 38904
rect 5368 38486 5396 38898
rect 5356 38480 5408 38486
rect 5356 38422 5408 38428
rect 5172 37188 5224 37194
rect 5172 37130 5224 37136
rect 5184 36854 5212 37130
rect 5264 37120 5316 37126
rect 5264 37062 5316 37068
rect 5172 36848 5224 36854
rect 5172 36790 5224 36796
rect 5080 36168 5132 36174
rect 5080 36110 5132 36116
rect 5170 36136 5226 36145
rect 5170 36071 5172 36080
rect 5224 36071 5226 36080
rect 5172 36042 5224 36048
rect 5276 35986 5304 37062
rect 5448 36848 5500 36854
rect 5448 36790 5500 36796
rect 5184 35958 5304 35986
rect 5184 35086 5212 35958
rect 5264 35624 5316 35630
rect 5264 35566 5316 35572
rect 5356 35624 5408 35630
rect 5356 35566 5408 35572
rect 5172 35080 5224 35086
rect 5000 35006 5120 35034
rect 5172 35022 5224 35028
rect 5092 34950 5120 35006
rect 4988 34944 5040 34950
rect 4988 34886 5040 34892
rect 5080 34944 5132 34950
rect 5080 34886 5132 34892
rect 5172 34944 5224 34950
rect 5276 34932 5304 35566
rect 5224 34904 5304 34932
rect 5172 34886 5224 34892
rect 5000 33454 5028 34886
rect 4988 33448 5040 33454
rect 4988 33390 5040 33396
rect 5000 32774 5028 33390
rect 5092 33289 5120 34886
rect 5078 33280 5134 33289
rect 5078 33215 5134 33224
rect 5080 32972 5132 32978
rect 5080 32914 5132 32920
rect 4988 32768 5040 32774
rect 4988 32710 5040 32716
rect 4896 30728 4948 30734
rect 4896 30670 4948 30676
rect 4804 30592 4856 30598
rect 4804 30534 4856 30540
rect 4724 30348 4936 30376
rect 4802 30288 4858 30297
rect 4802 30223 4858 30232
rect 4816 30122 4844 30223
rect 4804 30116 4856 30122
rect 4804 30058 4856 30064
rect 4712 30048 4764 30054
rect 4908 30002 4936 30348
rect 4712 29990 4764 29996
rect 4540 29566 4660 29594
rect 4528 29096 4580 29102
rect 4528 29038 4580 29044
rect 4436 27872 4488 27878
rect 4436 27814 4488 27820
rect 4344 27532 4396 27538
rect 4344 27474 4396 27480
rect 4344 27056 4396 27062
rect 4344 26998 4396 27004
rect 4356 26314 4384 26998
rect 4344 26308 4396 26314
rect 4344 26250 4396 26256
rect 4120 25928 4200 25956
rect 4252 25968 4304 25974
rect 4068 25910 4120 25916
rect 4252 25910 4304 25916
rect 3792 25900 3844 25906
rect 3792 25842 3844 25848
rect 3804 24954 3832 25842
rect 3917 25596 4225 25605
rect 3917 25594 3923 25596
rect 3979 25594 4003 25596
rect 4059 25594 4083 25596
rect 4139 25594 4163 25596
rect 4219 25594 4225 25596
rect 3979 25542 3981 25594
rect 4161 25542 4163 25594
rect 3917 25540 3923 25542
rect 3979 25540 4003 25542
rect 4059 25540 4083 25542
rect 4139 25540 4163 25542
rect 4219 25540 4225 25542
rect 3917 25531 4225 25540
rect 3792 24948 3844 24954
rect 3792 24890 3844 24896
rect 4264 24886 4292 25910
rect 4356 25362 4384 26250
rect 4344 25356 4396 25362
rect 4344 25298 4396 25304
rect 4356 24886 4384 25298
rect 4252 24880 4304 24886
rect 4252 24822 4304 24828
rect 4344 24880 4396 24886
rect 4344 24822 4396 24828
rect 3700 24812 3752 24818
rect 3700 24754 3752 24760
rect 3792 24812 3844 24818
rect 3792 24754 3844 24760
rect 3712 24410 3740 24754
rect 3804 24410 3832 24754
rect 3917 24508 4225 24517
rect 3917 24506 3923 24508
rect 3979 24506 4003 24508
rect 4059 24506 4083 24508
rect 4139 24506 4163 24508
rect 4219 24506 4225 24508
rect 3979 24454 3981 24506
rect 4161 24454 4163 24506
rect 3917 24452 3923 24454
rect 3979 24452 4003 24454
rect 4059 24452 4083 24454
rect 4139 24452 4163 24454
rect 4219 24452 4225 24454
rect 3917 24443 4225 24452
rect 3700 24404 3752 24410
rect 3700 24346 3752 24352
rect 3792 24404 3844 24410
rect 3792 24346 3844 24352
rect 3620 24262 3832 24290
rect 3424 23860 3476 23866
rect 3424 23802 3476 23808
rect 3516 23860 3568 23866
rect 3516 23802 3568 23808
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 3436 23225 3464 23666
rect 3422 23216 3478 23225
rect 3422 23151 3478 23160
rect 3804 22953 3832 24262
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4172 23508 4200 24142
rect 4264 23730 4292 24822
rect 4252 23724 4304 23730
rect 4252 23666 4304 23672
rect 4172 23480 4292 23508
rect 3917 23420 4225 23429
rect 3917 23418 3923 23420
rect 3979 23418 4003 23420
rect 4059 23418 4083 23420
rect 4139 23418 4163 23420
rect 4219 23418 4225 23420
rect 3979 23366 3981 23418
rect 4161 23366 4163 23418
rect 3917 23364 3923 23366
rect 3979 23364 4003 23366
rect 4059 23364 4083 23366
rect 4139 23364 4163 23366
rect 4219 23364 4225 23366
rect 3917 23355 4225 23364
rect 3974 23080 4030 23089
rect 3974 23015 4030 23024
rect 3790 22944 3846 22953
rect 3790 22879 3846 22888
rect 3804 22001 3832 22879
rect 3988 22438 4016 23015
rect 4264 22710 4292 23480
rect 4344 23044 4396 23050
rect 4344 22986 4396 22992
rect 4252 22704 4304 22710
rect 4066 22672 4122 22681
rect 4252 22646 4304 22652
rect 4066 22607 4068 22616
rect 4120 22607 4122 22616
rect 4068 22578 4120 22584
rect 4252 22568 4304 22574
rect 4252 22510 4304 22516
rect 3976 22432 4028 22438
rect 3976 22374 4028 22380
rect 3917 22332 4225 22341
rect 3917 22330 3923 22332
rect 3979 22330 4003 22332
rect 4059 22330 4083 22332
rect 4139 22330 4163 22332
rect 4219 22330 4225 22332
rect 3979 22278 3981 22330
rect 4161 22278 4163 22330
rect 3917 22276 3923 22278
rect 3979 22276 4003 22278
rect 4059 22276 4083 22278
rect 4139 22276 4163 22278
rect 4219 22276 4225 22278
rect 3917 22267 4225 22276
rect 3884 22092 3936 22098
rect 4264 22094 4292 22510
rect 4356 22234 4384 22986
rect 4448 22642 4476 27814
rect 4540 27062 4568 29038
rect 4632 28218 4660 29566
rect 4724 29306 4752 29990
rect 4816 29974 4936 30002
rect 4712 29300 4764 29306
rect 4712 29242 4764 29248
rect 4620 28212 4672 28218
rect 4620 28154 4672 28160
rect 4632 27985 4660 28154
rect 4618 27976 4674 27985
rect 4618 27911 4674 27920
rect 4618 27840 4674 27849
rect 4618 27775 4674 27784
rect 4632 27606 4660 27775
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 4528 27056 4580 27062
rect 4528 26998 4580 27004
rect 4620 26988 4672 26994
rect 4620 26930 4672 26936
rect 4528 26240 4580 26246
rect 4528 26182 4580 26188
rect 4540 25974 4568 26182
rect 4528 25968 4580 25974
rect 4528 25910 4580 25916
rect 4632 25786 4660 26930
rect 4540 25758 4660 25786
rect 4540 24834 4568 25758
rect 4724 25684 4752 29242
rect 4816 28404 4844 29974
rect 4896 29640 4948 29646
rect 4896 29582 4948 29588
rect 4908 29481 4936 29582
rect 4894 29472 4950 29481
rect 4894 29407 4950 29416
rect 4894 29336 4950 29345
rect 4894 29271 4950 29280
rect 4908 29170 4936 29271
rect 4896 29164 4948 29170
rect 4896 29106 4948 29112
rect 4894 28792 4950 28801
rect 4894 28727 4950 28736
rect 4908 28529 4936 28727
rect 4894 28520 4950 28529
rect 4894 28455 4950 28464
rect 4896 28416 4948 28422
rect 4816 28376 4896 28404
rect 4896 28358 4948 28364
rect 4908 28257 4936 28358
rect 4894 28248 4950 28257
rect 4894 28183 4950 28192
rect 4804 27464 4856 27470
rect 4804 27406 4856 27412
rect 4816 27062 4844 27406
rect 4804 27056 4856 27062
rect 4804 26998 4856 27004
rect 4804 26784 4856 26790
rect 4804 26726 4856 26732
rect 4816 25838 4844 26726
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4724 25656 4844 25684
rect 4540 24806 4660 24834
rect 4528 23724 4580 23730
rect 4528 23666 4580 23672
rect 4540 22794 4568 23666
rect 4632 22982 4660 24806
rect 4710 24712 4766 24721
rect 4710 24647 4712 24656
rect 4764 24647 4766 24656
rect 4712 24618 4764 24624
rect 4816 23474 4844 25656
rect 4908 25158 4936 28183
rect 5000 26450 5028 32710
rect 5092 31890 5120 32914
rect 5080 31884 5132 31890
rect 5080 31826 5132 31832
rect 5080 31680 5132 31686
rect 5080 31622 5132 31628
rect 5092 30802 5120 31622
rect 5080 30796 5132 30802
rect 5080 30738 5132 30744
rect 5078 30696 5134 30705
rect 5078 30631 5080 30640
rect 5132 30631 5134 30640
rect 5080 30602 5132 30608
rect 5184 30410 5212 34886
rect 5368 34610 5396 35566
rect 5356 34604 5408 34610
rect 5356 34546 5408 34552
rect 5264 33992 5316 33998
rect 5264 33934 5316 33940
rect 5276 33114 5304 33934
rect 5356 33516 5408 33522
rect 5356 33458 5408 33464
rect 5264 33108 5316 33114
rect 5264 33050 5316 33056
rect 5264 32768 5316 32774
rect 5264 32710 5316 32716
rect 5276 32570 5304 32710
rect 5264 32564 5316 32570
rect 5264 32506 5316 32512
rect 5368 32348 5396 33458
rect 5460 32502 5488 36790
rect 5552 32502 5580 41074
rect 6012 41002 6040 41550
rect 6000 40996 6052 41002
rect 6000 40938 6052 40944
rect 6000 40724 6052 40730
rect 6000 40666 6052 40672
rect 5908 39840 5960 39846
rect 5908 39782 5960 39788
rect 5920 39642 5948 39782
rect 6012 39642 6040 40666
rect 6104 39658 6132 42162
rect 6196 41857 6224 42162
rect 6276 42016 6328 42022
rect 6276 41958 6328 41964
rect 6182 41848 6238 41857
rect 6182 41783 6238 41792
rect 6288 41614 6316 41958
rect 6380 41818 6408 43182
rect 6368 41812 6420 41818
rect 6368 41754 6420 41760
rect 6276 41608 6328 41614
rect 6276 41550 6328 41556
rect 6184 41540 6236 41546
rect 6184 41482 6236 41488
rect 6196 41414 6224 41482
rect 6472 41414 6500 43302
rect 6552 43308 6604 43314
rect 6552 43250 6604 43256
rect 6564 42362 6592 43250
rect 6656 42906 6684 43710
rect 6748 43432 6776 44934
rect 6826 44840 6882 44934
rect 7102 44962 7158 45000
rect 7102 44934 7328 44962
rect 7102 44840 7158 44934
rect 6884 43548 7192 43557
rect 6884 43546 6890 43548
rect 6946 43546 6970 43548
rect 7026 43546 7050 43548
rect 7106 43546 7130 43548
rect 7186 43546 7192 43548
rect 6946 43494 6948 43546
rect 7128 43494 7130 43546
rect 6884 43492 6890 43494
rect 6946 43492 6970 43494
rect 7026 43492 7050 43494
rect 7106 43492 7130 43494
rect 7186 43492 7192 43494
rect 6884 43483 7192 43492
rect 6828 43444 6880 43450
rect 6748 43404 6828 43432
rect 7300 43432 7328 44934
rect 7378 44840 7434 45000
rect 7654 44840 7710 45000
rect 7930 44840 7986 45000
rect 8206 44840 8262 45000
rect 8482 44962 8538 45000
rect 8312 44934 8538 44962
rect 6828 43386 6880 43392
rect 7208 43404 7328 43432
rect 7208 42906 7236 43404
rect 6644 42900 6696 42906
rect 6644 42842 6696 42848
rect 7196 42900 7248 42906
rect 7196 42842 7248 42848
rect 6736 42628 6788 42634
rect 6736 42570 6788 42576
rect 7288 42628 7340 42634
rect 7288 42570 7340 42576
rect 6552 42356 6604 42362
rect 6552 42298 6604 42304
rect 6644 42220 6696 42226
rect 6644 42162 6696 42168
rect 6656 41857 6684 42162
rect 6748 42106 6776 42570
rect 6884 42460 7192 42469
rect 6884 42458 6890 42460
rect 6946 42458 6970 42460
rect 7026 42458 7050 42460
rect 7106 42458 7130 42460
rect 7186 42458 7192 42460
rect 6946 42406 6948 42458
rect 7128 42406 7130 42458
rect 6884 42404 6890 42406
rect 6946 42404 6970 42406
rect 7026 42404 7050 42406
rect 7106 42404 7130 42406
rect 7186 42404 7192 42406
rect 6884 42395 7192 42404
rect 7196 42220 7248 42226
rect 7196 42162 7248 42168
rect 6748 42078 6868 42106
rect 6736 42016 6788 42022
rect 6736 41958 6788 41964
rect 6642 41848 6698 41857
rect 6748 41818 6776 41958
rect 6840 41818 6868 42078
rect 7208 42022 7236 42162
rect 7196 42016 7248 42022
rect 7196 41958 7248 41964
rect 7300 41818 7328 42570
rect 7392 42362 7420 44840
rect 7472 43308 7524 43314
rect 7472 43250 7524 43256
rect 7380 42356 7432 42362
rect 7380 42298 7432 42304
rect 7380 42016 7432 42022
rect 7380 41958 7432 41964
rect 7392 41857 7420 41958
rect 7378 41848 7434 41857
rect 6642 41783 6698 41792
rect 6736 41812 6788 41818
rect 6736 41754 6788 41760
rect 6828 41812 6880 41818
rect 6828 41754 6880 41760
rect 7288 41812 7340 41818
rect 7378 41783 7434 41792
rect 7288 41754 7340 41760
rect 6736 41608 6788 41614
rect 6734 41576 6736 41585
rect 6788 41576 6790 41585
rect 6734 41511 6790 41520
rect 7484 41478 7512 43250
rect 7564 42696 7616 42702
rect 7564 42638 7616 42644
rect 7576 41818 7604 42638
rect 7668 42634 7696 44840
rect 7944 43450 7972 44840
rect 8220 43602 8248 44840
rect 8128 43574 8248 43602
rect 7932 43444 7984 43450
rect 7932 43386 7984 43392
rect 8128 43330 8156 43574
rect 8208 43444 8260 43450
rect 8312 43432 8340 44934
rect 8482 44840 8538 44934
rect 8758 44840 8814 45000
rect 9034 44840 9090 45000
rect 9310 44962 9366 45000
rect 9310 44934 9536 44962
rect 9310 44840 9366 44934
rect 8260 43404 8340 43432
rect 8208 43386 8260 43392
rect 8128 43302 8248 43330
rect 8116 42696 8168 42702
rect 8116 42638 8168 42644
rect 7656 42628 7708 42634
rect 7656 42570 7708 42576
rect 7840 42628 7892 42634
rect 7840 42570 7892 42576
rect 7852 42344 7880 42570
rect 7932 42560 7984 42566
rect 7932 42502 7984 42508
rect 7668 42316 7880 42344
rect 7564 41812 7616 41818
rect 7564 41754 7616 41760
rect 7472 41472 7524 41478
rect 7472 41414 7524 41420
rect 6196 41386 6316 41414
rect 6472 41386 6592 41414
rect 6288 41070 6316 41386
rect 6564 41274 6592 41386
rect 6884 41372 7192 41381
rect 6884 41370 6890 41372
rect 6946 41370 6970 41372
rect 7026 41370 7050 41372
rect 7106 41370 7130 41372
rect 7186 41370 7192 41372
rect 6946 41318 6948 41370
rect 7128 41318 7130 41370
rect 6884 41316 6890 41318
rect 6946 41316 6970 41318
rect 7026 41316 7050 41318
rect 7106 41316 7130 41318
rect 7186 41316 7192 41318
rect 6884 41307 7192 41316
rect 6552 41268 6604 41274
rect 6552 41210 6604 41216
rect 6552 41132 6604 41138
rect 6552 41074 6604 41080
rect 7380 41132 7432 41138
rect 7380 41074 7432 41080
rect 6276 41064 6328 41070
rect 6276 41006 6328 41012
rect 6368 41064 6420 41070
rect 6368 41006 6420 41012
rect 5908 39636 5960 39642
rect 5908 39578 5960 39584
rect 6000 39636 6052 39642
rect 6104 39630 6224 39658
rect 6000 39578 6052 39584
rect 6092 39296 6144 39302
rect 6092 39238 6144 39244
rect 6104 39098 6132 39238
rect 6092 39092 6144 39098
rect 6092 39034 6144 39040
rect 6000 38208 6052 38214
rect 6000 38150 6052 38156
rect 5816 37732 5868 37738
rect 5816 37674 5868 37680
rect 5632 37664 5684 37670
rect 5632 37606 5684 37612
rect 5644 36310 5672 37606
rect 5724 36916 5776 36922
rect 5724 36858 5776 36864
rect 5736 36718 5764 36858
rect 5724 36712 5776 36718
rect 5724 36654 5776 36660
rect 5632 36304 5684 36310
rect 5632 36246 5684 36252
rect 5644 35494 5672 36246
rect 5724 36236 5776 36242
rect 5724 36178 5776 36184
rect 5632 35488 5684 35494
rect 5632 35430 5684 35436
rect 5736 35306 5764 36178
rect 5644 35278 5764 35306
rect 5828 35290 5856 37674
rect 5908 36168 5960 36174
rect 5908 36110 5960 36116
rect 5816 35284 5868 35290
rect 5644 33386 5672 35278
rect 5816 35226 5868 35232
rect 5724 34944 5776 34950
rect 5724 34886 5776 34892
rect 5736 34746 5764 34886
rect 5724 34740 5776 34746
rect 5920 34728 5948 36110
rect 5724 34682 5776 34688
rect 5828 34700 5948 34728
rect 5724 33992 5776 33998
rect 5724 33934 5776 33940
rect 5736 33658 5764 33934
rect 5724 33652 5776 33658
rect 5724 33594 5776 33600
rect 5632 33380 5684 33386
rect 5632 33322 5684 33328
rect 5448 32496 5500 32502
rect 5448 32438 5500 32444
rect 5540 32496 5592 32502
rect 5540 32438 5592 32444
rect 5368 32320 5488 32348
rect 5356 31884 5408 31890
rect 5356 31826 5408 31832
rect 5264 31340 5316 31346
rect 5264 31282 5316 31288
rect 5276 31249 5304 31282
rect 5262 31240 5318 31249
rect 5262 31175 5318 31184
rect 5184 30382 5304 30410
rect 5172 30252 5224 30258
rect 5172 30194 5224 30200
rect 5184 30025 5212 30194
rect 5170 30016 5226 30025
rect 5170 29951 5226 29960
rect 5080 29776 5132 29782
rect 5080 29718 5132 29724
rect 5092 28014 5120 29718
rect 5276 28490 5304 30382
rect 5368 30054 5396 31826
rect 5460 31249 5488 32320
rect 5538 31512 5594 31521
rect 5538 31447 5540 31456
rect 5592 31447 5594 31456
rect 5540 31418 5592 31424
rect 5540 31340 5592 31346
rect 5540 31282 5592 31288
rect 5446 31240 5502 31249
rect 5446 31175 5502 31184
rect 5356 30048 5408 30054
rect 5356 29990 5408 29996
rect 5356 29572 5408 29578
rect 5356 29514 5408 29520
rect 5368 28529 5396 29514
rect 5354 28520 5410 28529
rect 5172 28484 5224 28490
rect 5172 28426 5224 28432
rect 5264 28484 5316 28490
rect 5354 28455 5410 28464
rect 5264 28426 5316 28432
rect 5184 28150 5212 28426
rect 5172 28144 5224 28150
rect 5172 28086 5224 28092
rect 5276 28064 5304 28426
rect 5460 28064 5488 31175
rect 5552 30258 5580 31282
rect 5540 30252 5592 30258
rect 5540 30194 5592 30200
rect 5540 28960 5592 28966
rect 5540 28902 5592 28908
rect 5552 28558 5580 28902
rect 5540 28552 5592 28558
rect 5540 28494 5592 28500
rect 5276 28036 5396 28064
rect 5460 28036 5580 28064
rect 5080 28008 5132 28014
rect 5080 27950 5132 27956
rect 5170 27976 5226 27985
rect 5368 27928 5396 28036
rect 5170 27911 5226 27920
rect 5184 27441 5212 27911
rect 5276 27900 5396 27928
rect 5170 27432 5226 27441
rect 5170 27367 5226 27376
rect 4988 26444 5040 26450
rect 4988 26386 5040 26392
rect 4896 25152 4948 25158
rect 4896 25094 4948 25100
rect 5000 23866 5028 26386
rect 5080 25900 5132 25906
rect 5080 25842 5132 25848
rect 5092 23866 5120 25842
rect 5172 25220 5224 25226
rect 5172 25162 5224 25168
rect 4988 23860 5040 23866
rect 4988 23802 5040 23808
rect 5080 23860 5132 23866
rect 5080 23802 5132 23808
rect 4988 23588 5040 23594
rect 4988 23530 5040 23536
rect 4724 23446 4844 23474
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4540 22766 4660 22794
rect 4436 22636 4488 22642
rect 4436 22578 4488 22584
rect 4344 22228 4396 22234
rect 4344 22170 4396 22176
rect 4264 22066 4384 22094
rect 3884 22034 3936 22040
rect 3790 21992 3846 22001
rect 3608 21956 3660 21962
rect 3790 21927 3846 21936
rect 3608 21898 3660 21904
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3528 21010 3556 21422
rect 3516 21004 3568 21010
rect 3516 20946 3568 20952
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3332 20528 3384 20534
rect 3332 20470 3384 20476
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 3160 19446 3188 20402
rect 3422 20360 3478 20369
rect 3422 20295 3478 20304
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 3344 19689 3372 19790
rect 3330 19680 3386 19689
rect 3330 19615 3386 19624
rect 3148 19440 3200 19446
rect 3054 19408 3110 19417
rect 3148 19382 3200 19388
rect 3054 19343 3110 19352
rect 3068 19242 3096 19343
rect 3436 19334 3464 20295
rect 3528 20058 3556 20742
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 3528 19689 3556 19790
rect 3620 19718 3648 21898
rect 3896 21690 3924 22034
rect 3884 21684 3936 21690
rect 3884 21626 3936 21632
rect 4252 21616 4304 21622
rect 4252 21558 4304 21564
rect 3792 21548 3844 21554
rect 3792 21490 3844 21496
rect 3700 21004 3752 21010
rect 3700 20946 3752 20952
rect 3608 19712 3660 19718
rect 3514 19680 3570 19689
rect 3608 19654 3660 19660
rect 3514 19615 3570 19624
rect 3528 19378 3556 19615
rect 3606 19408 3662 19417
rect 3160 19306 3464 19334
rect 3516 19372 3568 19378
rect 3606 19343 3662 19352
rect 3516 19314 3568 19320
rect 3056 19236 3108 19242
rect 3056 19178 3108 19184
rect 2976 18822 3096 18850
rect 2780 18566 2832 18572
rect 2870 18592 2926 18601
rect 2792 18154 2820 18566
rect 2870 18527 2926 18536
rect 3068 18170 3096 18822
rect 2780 18148 2832 18154
rect 2780 18090 2832 18096
rect 2976 18142 3096 18170
rect 2700 18006 2912 18034
rect 2412 17808 2464 17814
rect 2412 17750 2464 17756
rect 2884 17746 2912 18006
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2780 17672 2832 17678
rect 2332 17632 2728 17660
rect 2228 17536 2280 17542
rect 2228 17478 2280 17484
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2226 17232 2282 17241
rect 2226 17167 2228 17176
rect 2280 17167 2282 17176
rect 2228 17138 2280 17144
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2148 15966 2268 15994
rect 2136 15904 2188 15910
rect 2136 15846 2188 15852
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 1952 15632 2004 15638
rect 1952 15574 2004 15580
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 1860 14000 1912 14006
rect 1860 13942 1912 13948
rect 1858 13832 1914 13841
rect 1858 13767 1914 13776
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1582 12880 1638 12889
rect 1582 12815 1638 12824
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1308 12164 1360 12170
rect 1308 12106 1360 12112
rect 1320 12073 1348 12106
rect 1306 12064 1362 12073
rect 1306 11999 1362 12008
rect 1504 11898 1532 12242
rect 1492 11892 1544 11898
rect 1320 11852 1492 11880
rect 1320 9178 1348 11852
rect 1492 11834 1544 11840
rect 1400 11008 1452 11014
rect 1400 10950 1452 10956
rect 1412 10062 1440 10950
rect 1596 10470 1624 12815
rect 1674 12608 1730 12617
rect 1674 12543 1730 12552
rect 1584 10464 1636 10470
rect 1490 10432 1546 10441
rect 1584 10406 1636 10412
rect 1490 10367 1546 10376
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1398 9888 1454 9897
rect 1398 9823 1454 9832
rect 1308 9172 1360 9178
rect 1228 9132 1308 9160
rect 1228 7954 1256 9132
rect 1308 9114 1360 9120
rect 1306 9072 1362 9081
rect 1306 9007 1362 9016
rect 1320 8906 1348 9007
rect 1308 8900 1360 8906
rect 1308 8842 1360 8848
rect 1412 8566 1440 9823
rect 1400 8560 1452 8566
rect 1400 8502 1452 8508
rect 1504 8090 1532 10367
rect 1688 10198 1716 12543
rect 1780 11354 1808 13126
rect 1872 11694 1900 13767
rect 1964 12782 1992 15438
rect 2056 14906 2084 15506
rect 2148 15094 2176 15846
rect 2240 15162 2268 15966
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 2136 15088 2188 15094
rect 2136 15030 2188 15036
rect 2056 14878 2176 14906
rect 2148 14822 2176 14878
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 2056 13326 2084 14214
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1766 11248 1822 11257
rect 1766 11183 1822 11192
rect 1676 10192 1728 10198
rect 1676 10134 1728 10140
rect 1780 9722 1808 11183
rect 1872 11150 1900 11290
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1858 8936 1914 8945
rect 1688 8634 1716 8910
rect 1858 8871 1914 8880
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1582 8528 1638 8537
rect 1582 8463 1638 8472
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1216 7948 1268 7954
rect 1216 7890 1268 7896
rect 1228 6984 1256 7890
rect 1492 7812 1544 7818
rect 1492 7754 1544 7760
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 1320 7546 1348 7647
rect 1308 7540 1360 7546
rect 1308 7482 1360 7488
rect 1398 7304 1454 7313
rect 1308 7268 1360 7274
rect 1398 7239 1454 7248
rect 1308 7210 1360 7216
rect 1320 7177 1348 7210
rect 1306 7168 1362 7177
rect 1306 7103 1362 7112
rect 1228 6956 1348 6984
rect 1216 6860 1268 6866
rect 1216 6802 1268 6808
rect 1228 6361 1256 6802
rect 1214 6352 1270 6361
rect 1320 6322 1348 6956
rect 1214 6287 1270 6296
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 938 6216 994 6225
rect 938 6151 994 6160
rect 1122 5536 1178 5545
rect 1122 5471 1178 5480
rect 1136 4486 1164 5471
rect 1412 5370 1440 7239
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 1124 4480 1176 4486
rect 1124 4422 1176 4428
rect 1504 3738 1532 7754
rect 1596 6458 1624 8463
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1688 6712 1716 8366
rect 1766 8120 1822 8129
rect 1766 8055 1822 8064
rect 1780 7002 1808 8055
rect 1872 7478 1900 8871
rect 1964 8090 1992 12582
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1860 7472 1912 7478
rect 1860 7414 1912 7420
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1964 7002 1992 7346
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2056 6882 2084 12922
rect 2148 12782 2176 14758
rect 2226 14512 2282 14521
rect 2226 14447 2282 14456
rect 2240 14414 2268 14447
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2332 13977 2360 16050
rect 2318 13968 2374 13977
rect 2318 13903 2374 13912
rect 2424 13818 2452 17478
rect 2700 16980 2728 17632
rect 2832 17620 2912 17626
rect 2780 17614 2912 17620
rect 2792 17598 2912 17614
rect 2700 16952 2820 16980
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2516 15638 2544 16390
rect 2686 16144 2742 16153
rect 2686 16079 2688 16088
rect 2740 16079 2742 16088
rect 2688 16050 2740 16056
rect 2504 15632 2556 15638
rect 2504 15574 2556 15580
rect 2594 15600 2650 15609
rect 2594 15535 2650 15544
rect 2608 15366 2636 15535
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2608 14770 2636 15302
rect 2700 15178 2728 16050
rect 2792 15910 2820 16952
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2884 15570 2912 17598
rect 2976 17542 3004 18142
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 3068 17270 3096 18022
rect 3056 17264 3108 17270
rect 3056 17206 3108 17212
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2700 15150 2912 15178
rect 2976 15162 3004 15438
rect 2884 14770 2912 15150
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2608 14742 2820 14770
rect 2884 14742 3096 14770
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2792 14362 2820 14742
rect 2240 13790 2452 13818
rect 2240 13530 2268 13790
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 13569 2360 13670
rect 2318 13560 2374 13569
rect 2228 13524 2280 13530
rect 2318 13495 2374 13504
rect 2228 13466 2280 13472
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 2136 11824 2188 11830
rect 2136 11766 2188 11772
rect 2148 9489 2176 11766
rect 2240 11354 2268 13466
rect 2412 12708 2464 12714
rect 2412 12650 2464 12656
rect 2318 12336 2374 12345
rect 2424 12306 2452 12650
rect 2318 12271 2374 12280
rect 2412 12300 2464 12306
rect 2332 12238 2360 12271
rect 2412 12242 2464 12248
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2424 10606 2452 11494
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2318 10160 2374 10169
rect 2318 10095 2374 10104
rect 2332 9722 2360 10095
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2424 9602 2452 10542
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2332 9574 2452 9602
rect 2134 9480 2190 9489
rect 2134 9415 2190 9424
rect 2240 9178 2268 9522
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2332 9058 2360 9574
rect 2240 9030 2360 9058
rect 2136 7880 2188 7886
rect 2134 7848 2136 7857
rect 2188 7848 2190 7857
rect 2134 7783 2190 7792
rect 2240 7698 2268 9030
rect 2318 8936 2374 8945
rect 2318 8871 2374 8880
rect 2332 8430 2360 8871
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 1872 6854 2084 6882
rect 2148 7670 2268 7698
rect 1688 6684 1808 6712
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1582 6080 1638 6089
rect 1582 6015 1638 6024
rect 1596 4826 1624 6015
rect 1780 5778 1808 6684
rect 1872 6322 1900 6854
rect 2148 6798 2176 7670
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1860 6180 1912 6186
rect 1860 6122 1912 6128
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1676 5704 1728 5710
rect 1674 5672 1676 5681
rect 1728 5672 1730 5681
rect 1674 5607 1730 5616
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1582 4312 1638 4321
rect 1582 4247 1584 4256
rect 1636 4247 1638 4256
rect 1584 4218 1636 4224
rect 1492 3732 1544 3738
rect 1492 3674 1544 3680
rect 1780 3641 1808 5714
rect 1872 4146 1900 6122
rect 1964 4690 1992 6666
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2134 6624 2190 6633
rect 2056 5302 2084 6598
rect 2134 6559 2190 6568
rect 2148 5370 2176 6559
rect 2240 5914 2268 6666
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2332 5778 2360 8366
rect 2516 8090 2544 14350
rect 2792 14334 2912 14362
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2594 13424 2650 13433
rect 2594 13359 2650 13368
rect 2608 10674 2636 13359
rect 2700 12986 2728 14010
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2792 12782 2820 14214
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2884 12764 2912 14334
rect 2964 14340 3016 14346
rect 2964 14282 3016 14288
rect 2976 13734 3004 14282
rect 3068 13938 3096 14742
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3068 13841 3096 13874
rect 3054 13832 3110 13841
rect 3054 13767 3110 13776
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 3068 13326 3096 13670
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3068 12850 3096 12922
rect 3056 12844 3108 12850
rect 3160 12832 3188 19306
rect 3528 19281 3556 19314
rect 3514 19272 3570 19281
rect 3514 19207 3570 19216
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3252 18290 3280 19110
rect 3620 18698 3648 19343
rect 3712 18834 3740 20946
rect 3804 20942 3832 21490
rect 3917 21244 4225 21253
rect 3917 21242 3923 21244
rect 3979 21242 4003 21244
rect 4059 21242 4083 21244
rect 4139 21242 4163 21244
rect 4219 21242 4225 21244
rect 3979 21190 3981 21242
rect 4161 21190 4163 21242
rect 3917 21188 3923 21190
rect 3979 21188 4003 21190
rect 4059 21188 4083 21190
rect 4139 21188 4163 21190
rect 4219 21188 4225 21190
rect 3917 21179 4225 21188
rect 3792 20936 3844 20942
rect 3792 20878 3844 20884
rect 3804 20505 3832 20878
rect 4264 20534 4292 21558
rect 4252 20528 4304 20534
rect 3790 20496 3846 20505
rect 4252 20470 4304 20476
rect 3790 20431 3846 20440
rect 4264 20369 4292 20470
rect 4250 20360 4306 20369
rect 4250 20295 4306 20304
rect 4160 20256 4212 20262
rect 4212 20216 4292 20244
rect 4160 20198 4212 20204
rect 3917 20156 4225 20165
rect 3917 20154 3923 20156
rect 3979 20154 4003 20156
rect 4059 20154 4083 20156
rect 4139 20154 4163 20156
rect 4219 20154 4225 20156
rect 3979 20102 3981 20154
rect 4161 20102 4163 20154
rect 3917 20100 3923 20102
rect 3979 20100 4003 20102
rect 4059 20100 4083 20102
rect 4139 20100 4163 20102
rect 4219 20100 4225 20102
rect 3917 20091 4225 20100
rect 3792 19848 3844 19854
rect 3792 19790 3844 19796
rect 3804 19514 3832 19790
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3896 19514 3924 19654
rect 4264 19553 4292 20216
rect 4250 19544 4306 19553
rect 3792 19508 3844 19514
rect 3792 19450 3844 19456
rect 3884 19508 3936 19514
rect 4250 19479 4306 19488
rect 3884 19450 3936 19456
rect 3917 19068 4225 19077
rect 3917 19066 3923 19068
rect 3979 19066 4003 19068
rect 4059 19066 4083 19068
rect 4139 19066 4163 19068
rect 4219 19066 4225 19068
rect 3979 19014 3981 19066
rect 4161 19014 4163 19066
rect 3917 19012 3923 19014
rect 3979 19012 4003 19014
rect 4059 19012 4083 19014
rect 4139 19012 4163 19014
rect 4219 19012 4225 19014
rect 3917 19003 4225 19012
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 3608 18692 3660 18698
rect 3608 18634 3660 18640
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3528 18329 3556 18362
rect 3514 18320 3570 18329
rect 3240 18284 3292 18290
rect 3514 18255 3570 18264
rect 3240 18226 3292 18232
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3344 17882 3372 18022
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3516 17536 3568 17542
rect 3568 17496 3648 17524
rect 3516 17478 3568 17484
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3252 13394 3280 15846
rect 3424 15632 3476 15638
rect 3424 15574 3476 15580
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3252 13025 3280 13126
rect 3238 13016 3294 13025
rect 3344 12986 3372 15506
rect 3436 14482 3464 15574
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 3528 14278 3556 16730
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3514 13696 3570 13705
rect 3514 13631 3570 13640
rect 3528 13530 3556 13631
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3514 13152 3570 13161
rect 3514 13087 3570 13096
rect 3528 12986 3556 13087
rect 3238 12951 3294 12960
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3160 12804 3280 12832
rect 3056 12786 3108 12792
rect 2964 12776 3016 12782
rect 2884 12736 2964 12764
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 2700 12442 2728 12650
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2884 12322 2912 12736
rect 2964 12718 3016 12724
rect 2700 12294 2912 12322
rect 2700 11257 2728 12294
rect 2778 12200 2834 12209
rect 2778 12135 2834 12144
rect 3148 12164 3200 12170
rect 2686 11248 2742 11257
rect 2686 11183 2742 11192
rect 2700 11150 2728 11183
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2792 10130 2820 12135
rect 3148 12106 3200 12112
rect 3160 11898 3188 12106
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2884 11665 2912 11698
rect 2870 11656 2926 11665
rect 3252 11608 3280 12804
rect 3344 12209 3372 12922
rect 3422 12608 3478 12617
rect 3422 12543 3478 12552
rect 3330 12200 3386 12209
rect 3330 12135 3386 12144
rect 2870 11591 2926 11600
rect 3160 11580 3280 11608
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 3068 11354 3096 11494
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 3160 11234 3188 11580
rect 3238 11520 3294 11529
rect 3238 11455 3294 11464
rect 3068 11206 3188 11234
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2976 10810 3004 11086
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2884 10010 2912 10406
rect 2884 9994 3004 10010
rect 2688 9988 2740 9994
rect 2884 9988 3016 9994
rect 2884 9982 2964 9988
rect 2688 9930 2740 9936
rect 2964 9930 3016 9936
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2608 9110 2636 9522
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2608 8430 2636 8910
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2504 7404 2556 7410
rect 2424 7364 2504 7392
rect 2424 6118 2452 7364
rect 2504 7346 2556 7352
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2516 6202 2544 6666
rect 2516 6174 2636 6202
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2044 5296 2096 5302
rect 2044 5238 2096 5244
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 2332 4622 2360 5510
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1766 3632 1822 3641
rect 1766 3567 1822 3576
rect 1872 3534 1900 4082
rect 2424 3738 2452 5714
rect 2502 5536 2558 5545
rect 2502 5471 2558 5480
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1596 3194 1624 3470
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 584 2746 704 2774
rect 768 2746 888 2774
rect 386 1456 442 1465
rect 386 1391 442 1400
rect 584 814 612 2746
rect 768 2378 796 2746
rect 1964 2650 1992 3062
rect 2516 2774 2544 5471
rect 2608 5370 2636 6174
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2608 4826 2636 5170
rect 2700 4826 2728 9930
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2884 9625 2912 9862
rect 2870 9616 2926 9625
rect 2870 9551 2926 9560
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2976 9178 3004 9522
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2870 8800 2926 8809
rect 2792 8430 2820 8774
rect 2870 8735 2926 8744
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2884 7478 2912 8735
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2976 7290 3004 8366
rect 3068 8072 3096 11206
rect 3146 10704 3202 10713
rect 3146 10639 3202 10648
rect 3160 9654 3188 10639
rect 3252 10266 3280 11455
rect 3344 11218 3372 12135
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3330 10976 3386 10985
rect 3330 10911 3386 10920
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3344 9926 3372 10911
rect 3436 10656 3464 12543
rect 3620 12374 3648 17496
rect 3712 16658 3740 18770
rect 4356 18630 4384 22066
rect 4434 21992 4490 22001
rect 4434 21927 4436 21936
rect 4488 21927 4490 21936
rect 4436 21898 4488 21904
rect 4436 21412 4488 21418
rect 4436 21354 4488 21360
rect 4448 21146 4476 21354
rect 4528 21344 4580 21350
rect 4528 21286 4580 21292
rect 4436 21140 4488 21146
rect 4436 21082 4488 21088
rect 4434 19952 4490 19961
rect 4434 19887 4490 19896
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 4356 18290 4384 18566
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 4160 18216 4212 18222
rect 4212 18176 4292 18204
rect 4160 18158 4212 18164
rect 3700 16652 3752 16658
rect 3700 16594 3752 16600
rect 3712 16114 3740 16594
rect 3804 16114 3832 18158
rect 3917 17980 4225 17989
rect 3917 17978 3923 17980
rect 3979 17978 4003 17980
rect 4059 17978 4083 17980
rect 4139 17978 4163 17980
rect 4219 17978 4225 17980
rect 3979 17926 3981 17978
rect 4161 17926 4163 17978
rect 3917 17924 3923 17926
rect 3979 17924 4003 17926
rect 4059 17924 4083 17926
rect 4139 17924 4163 17926
rect 4219 17924 4225 17926
rect 3917 17915 4225 17924
rect 4264 17785 4292 18176
rect 4448 18170 4476 19887
rect 4540 18222 4568 21286
rect 4632 20534 4660 22766
rect 4724 22137 4752 23446
rect 5000 22574 5028 23530
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 4988 22568 5040 22574
rect 4988 22510 5040 22516
rect 4804 22500 4856 22506
rect 4804 22442 4856 22448
rect 4710 22128 4766 22137
rect 4710 22063 4766 22072
rect 4620 20528 4672 20534
rect 4620 20470 4672 20476
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4724 19990 4752 20402
rect 4712 19984 4764 19990
rect 4712 19926 4764 19932
rect 4618 19000 4674 19009
rect 4618 18935 4674 18944
rect 4632 18766 4660 18935
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4356 18142 4476 18170
rect 4528 18216 4580 18222
rect 4528 18158 4580 18164
rect 4250 17776 4306 17785
rect 4250 17711 4306 17720
rect 3917 16892 4225 16901
rect 3917 16890 3923 16892
rect 3979 16890 4003 16892
rect 4059 16890 4083 16892
rect 4139 16890 4163 16892
rect 4219 16890 4225 16892
rect 3979 16838 3981 16890
rect 4161 16838 4163 16890
rect 3917 16836 3923 16838
rect 3979 16836 4003 16838
rect 4059 16836 4083 16838
rect 4139 16836 4163 16838
rect 4219 16836 4225 16838
rect 3917 16827 4225 16836
rect 4250 16688 4306 16697
rect 4250 16623 4306 16632
rect 4264 16590 4292 16623
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 3698 15872 3754 15881
rect 3698 15807 3754 15816
rect 3712 15162 3740 15807
rect 3917 15804 4225 15813
rect 3917 15802 3923 15804
rect 3979 15802 4003 15804
rect 4059 15802 4083 15804
rect 4139 15802 4163 15804
rect 4219 15802 4225 15804
rect 3979 15750 3981 15802
rect 4161 15750 4163 15802
rect 3917 15748 3923 15750
rect 3979 15748 4003 15750
rect 4059 15748 4083 15750
rect 4139 15748 4163 15750
rect 4219 15748 4225 15750
rect 3917 15739 4225 15748
rect 4264 15688 4292 16526
rect 3988 15660 4292 15688
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3700 14884 3752 14890
rect 3700 14826 3752 14832
rect 3712 14074 3740 14826
rect 3804 14414 3832 14962
rect 3988 14890 4016 15660
rect 4066 15328 4122 15337
rect 4122 15286 4292 15314
rect 4066 15263 4122 15272
rect 3976 14884 4028 14890
rect 3976 14826 4028 14832
rect 3917 14716 4225 14725
rect 3917 14714 3923 14716
rect 3979 14714 4003 14716
rect 4059 14714 4083 14716
rect 4139 14714 4163 14716
rect 4219 14714 4225 14716
rect 3979 14662 3981 14714
rect 4161 14662 4163 14714
rect 3917 14660 3923 14662
rect 3979 14660 4003 14662
rect 4059 14660 4083 14662
rect 4139 14660 4163 14662
rect 4219 14660 4225 14662
rect 3917 14651 4225 14660
rect 4160 14544 4212 14550
rect 4264 14498 4292 15286
rect 4212 14492 4292 14498
rect 4160 14486 4292 14492
rect 4172 14470 4292 14486
rect 3792 14408 3844 14414
rect 4356 14396 4384 18142
rect 4816 16114 4844 22442
rect 4908 22098 4936 22510
rect 5000 22234 5028 22510
rect 4988 22228 5040 22234
rect 4988 22170 5040 22176
rect 4896 22092 4948 22098
rect 4896 22034 4948 22040
rect 4908 20466 4936 22034
rect 4988 21140 5040 21146
rect 4988 21082 5040 21088
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 5000 20097 5028 21082
rect 4986 20088 5042 20097
rect 4986 20023 5042 20032
rect 5000 19922 5028 20023
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 5000 18290 5028 18566
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4712 16040 4764 16046
rect 4618 16008 4674 16017
rect 4712 15982 4764 15988
rect 4618 15943 4674 15952
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4540 15706 4568 15846
rect 4632 15706 4660 15943
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4540 15026 4568 15642
rect 4724 15434 4752 15982
rect 4620 15428 4672 15434
rect 4620 15370 4672 15376
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4632 15337 4660 15370
rect 4618 15328 4674 15337
rect 4618 15263 4674 15272
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4632 14906 4660 15263
rect 3792 14350 3844 14356
rect 4264 14368 4384 14396
rect 4448 14878 4660 14906
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3700 13728 3752 13734
rect 3700 13670 3752 13676
rect 3712 13462 3740 13670
rect 3804 13512 3832 13806
rect 3917 13628 4225 13637
rect 3917 13626 3923 13628
rect 3979 13626 4003 13628
rect 4059 13626 4083 13628
rect 4139 13626 4163 13628
rect 4219 13626 4225 13628
rect 3979 13574 3981 13626
rect 4161 13574 4163 13626
rect 3917 13572 3923 13574
rect 3979 13572 4003 13574
rect 4059 13572 4083 13574
rect 4139 13572 4163 13574
rect 4219 13572 4225 13574
rect 3917 13563 4225 13572
rect 3804 13484 3924 13512
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 3700 13320 3752 13326
rect 3752 13280 3832 13308
rect 3700 13262 3752 13268
rect 3700 12640 3752 12646
rect 3804 12617 3832 13280
rect 3896 12918 3924 13484
rect 3974 13016 4030 13025
rect 3974 12951 4030 12960
rect 3884 12912 3936 12918
rect 3884 12854 3936 12860
rect 3988 12850 4016 12951
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3700 12582 3752 12588
rect 3790 12608 3846 12617
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 3712 11234 3740 12582
rect 3790 12543 3846 12552
rect 3917 12540 4225 12549
rect 3917 12538 3923 12540
rect 3979 12538 4003 12540
rect 4059 12538 4083 12540
rect 4139 12538 4163 12540
rect 4219 12538 4225 12540
rect 3979 12486 3981 12538
rect 4161 12486 4163 12538
rect 3917 12484 3923 12486
rect 3979 12484 4003 12486
rect 4059 12484 4083 12486
rect 4139 12484 4163 12486
rect 4219 12484 4225 12486
rect 3917 12475 4225 12484
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11801 4016 12038
rect 3974 11792 4030 11801
rect 4264 11778 4292 14368
rect 4264 11762 4384 11778
rect 3974 11727 4030 11736
rect 4068 11756 4120 11762
rect 4264 11756 4396 11762
rect 4264 11750 4344 11756
rect 4068 11698 4120 11704
rect 4344 11698 4396 11704
rect 4080 11665 4108 11698
rect 4066 11656 4122 11665
rect 4066 11591 4122 11600
rect 4160 11552 4212 11558
rect 4212 11512 4292 11540
rect 4160 11494 4212 11500
rect 3917 11452 4225 11461
rect 3917 11450 3923 11452
rect 3979 11450 4003 11452
rect 4059 11450 4083 11452
rect 4139 11450 4163 11452
rect 4219 11450 4225 11452
rect 3979 11398 3981 11450
rect 4161 11398 4163 11450
rect 3917 11396 3923 11398
rect 3979 11396 4003 11398
rect 4059 11396 4083 11398
rect 4139 11396 4163 11398
rect 4219 11396 4225 11398
rect 3917 11387 4225 11396
rect 4264 11336 4292 11512
rect 4172 11308 4384 11336
rect 3712 11206 4108 11234
rect 3884 11144 3936 11150
rect 3804 11104 3884 11132
rect 3804 10962 3832 11104
rect 3884 11086 3936 11092
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3620 10934 3832 10962
rect 3436 10628 3556 10656
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3436 9586 3464 10474
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 3436 9110 3464 9386
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3422 8936 3478 8945
rect 3528 8922 3556 10628
rect 3620 8974 3648 10934
rect 3988 10826 4016 11086
rect 3804 10798 4016 10826
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3478 8894 3556 8922
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3422 8871 3478 8880
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3330 8528 3386 8537
rect 3240 8492 3292 8498
rect 3330 8463 3386 8472
rect 3240 8434 3292 8440
rect 3252 8090 3280 8434
rect 3240 8084 3292 8090
rect 3068 8044 3188 8072
rect 3054 7984 3110 7993
rect 3054 7919 3110 7928
rect 2884 7274 3004 7290
rect 2884 7268 3016 7274
rect 2884 7262 2964 7268
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 2792 6458 2820 6666
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2884 6338 2912 7262
rect 2964 7210 3016 7216
rect 2964 6928 3016 6934
rect 2964 6870 3016 6876
rect 2792 6310 2912 6338
rect 2792 5914 2820 6310
rect 2976 6304 3004 6870
rect 3068 6866 3096 7919
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2976 6276 3096 6304
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2778 5808 2834 5817
rect 2884 5778 2912 5850
rect 2976 5778 3004 6054
rect 2778 5743 2834 5752
rect 2872 5772 2924 5778
rect 2792 5370 2820 5743
rect 2872 5714 2924 5720
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 3068 5114 3096 6276
rect 2884 5086 3096 5114
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2884 4622 2912 5086
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 3068 4826 3096 4966
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 2962 4720 3018 4729
rect 2962 4655 3018 4664
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2608 4049 2636 4082
rect 2594 4040 2650 4049
rect 2594 3975 2650 3984
rect 2976 3534 3004 4655
rect 2964 3528 3016 3534
rect 2870 3496 2926 3505
rect 2964 3470 3016 3476
rect 2870 3431 2926 3440
rect 2516 2746 2636 2774
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 756 2372 808 2378
rect 756 2314 808 2320
rect 848 1896 900 1902
rect 676 1856 848 1884
rect 572 808 624 814
rect 572 750 624 756
rect 202 0 258 160
rect 478 82 534 160
rect 676 82 704 1856
rect 848 1838 900 1844
rect 478 54 704 82
rect 754 82 810 160
rect 952 82 980 2382
rect 1032 1828 1084 1834
rect 1032 1770 1084 1776
rect 1044 160 1072 1770
rect 1504 1442 1532 2382
rect 1320 1414 1532 1442
rect 1320 160 1348 1414
rect 1676 1352 1728 1358
rect 1674 1320 1676 1329
rect 2044 1352 2096 1358
rect 1728 1320 1730 1329
rect 1584 1284 1636 1290
rect 2042 1320 2044 1329
rect 2228 1352 2280 1358
rect 2096 1320 2098 1329
rect 1674 1255 1730 1264
rect 1952 1284 2004 1290
rect 1584 1226 1636 1232
rect 2516 1306 2544 2382
rect 2608 1358 2636 2746
rect 2884 2038 2912 3431
rect 3160 2774 3188 8044
rect 3240 8026 3292 8032
rect 3344 7886 3372 8463
rect 3436 8430 3464 8774
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3330 6896 3386 6905
rect 3330 6831 3332 6840
rect 3384 6831 3386 6840
rect 3332 6802 3384 6808
rect 3332 6656 3384 6662
rect 3252 6616 3332 6644
rect 3252 4146 3280 6616
rect 3332 6598 3384 6604
rect 3330 6488 3386 6497
rect 3330 6423 3386 6432
rect 3344 5030 3372 6423
rect 3436 5914 3464 8366
rect 3712 7410 3740 10542
rect 3804 8956 3832 10798
rect 3974 10704 4030 10713
rect 3974 10639 3976 10648
rect 4028 10639 4030 10648
rect 3976 10610 4028 10616
rect 4080 10606 4108 11206
rect 4172 10674 4200 11308
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3917 10364 4225 10373
rect 3917 10362 3923 10364
rect 3979 10362 4003 10364
rect 4059 10362 4083 10364
rect 4139 10362 4163 10364
rect 4219 10362 4225 10364
rect 3979 10310 3981 10362
rect 4161 10310 4163 10362
rect 3917 10308 3923 10310
rect 3979 10308 4003 10310
rect 4059 10308 4083 10310
rect 4139 10308 4163 10310
rect 4219 10308 4225 10310
rect 3917 10299 4225 10308
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 3896 9722 3924 9930
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3917 9276 4225 9285
rect 3917 9274 3923 9276
rect 3979 9274 4003 9276
rect 4059 9274 4083 9276
rect 4139 9274 4163 9276
rect 4219 9274 4225 9276
rect 3979 9222 3981 9274
rect 4161 9222 4163 9274
rect 3917 9220 3923 9222
rect 3979 9220 4003 9222
rect 4059 9220 4083 9222
rect 4139 9220 4163 9222
rect 4219 9220 4225 9222
rect 3917 9211 4225 9220
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 3976 8968 4028 8974
rect 3804 8928 3976 8956
rect 3976 8910 4028 8916
rect 3988 8537 4016 8910
rect 3790 8528 3846 8537
rect 3974 8528 4030 8537
rect 3846 8486 3924 8514
rect 3790 8463 3846 8472
rect 3896 8412 3924 8486
rect 3974 8463 4030 8472
rect 3976 8424 4028 8430
rect 3790 8392 3846 8401
rect 3896 8384 3976 8412
rect 3976 8366 4028 8372
rect 3790 8327 3846 8336
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3700 7268 3752 7274
rect 3700 7210 3752 7216
rect 3712 6798 3740 7210
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3700 6656 3752 6662
rect 3698 6624 3700 6633
rect 3752 6624 3754 6633
rect 3698 6559 3754 6568
rect 3712 6322 3740 6559
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3528 5642 3556 6190
rect 3620 5914 3648 6258
rect 3698 6216 3754 6225
rect 3698 6151 3754 6160
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3712 5710 3740 6151
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3424 4616 3476 4622
rect 3422 4584 3424 4593
rect 3476 4584 3478 4593
rect 3422 4519 3478 4528
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3344 4282 3372 4422
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3528 4146 3556 5578
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3712 2774 3740 4218
rect 3068 2746 3188 2774
rect 3620 2746 3740 2774
rect 3068 2106 3096 2746
rect 3620 2106 3648 2746
rect 3056 2100 3108 2106
rect 3056 2042 3108 2048
rect 3608 2100 3660 2106
rect 3608 2042 3660 2048
rect 2872 2032 2924 2038
rect 2872 1974 2924 1980
rect 2780 1964 2832 1970
rect 2700 1924 2780 1952
rect 2228 1294 2280 1300
rect 2042 1255 2098 1264
rect 1952 1226 2004 1232
rect 1596 160 1624 1226
rect 754 54 980 82
rect 478 0 534 54
rect 754 0 810 54
rect 1030 0 1086 160
rect 1306 0 1362 160
rect 1582 0 1638 160
rect 1858 82 1914 160
rect 1964 82 1992 1226
rect 1858 54 1992 82
rect 2134 82 2190 160
rect 2240 82 2268 1294
rect 2424 1278 2544 1306
rect 2596 1352 2648 1358
rect 2596 1294 2648 1300
rect 2424 160 2452 1278
rect 2700 160 2728 1924
rect 2780 1906 2832 1912
rect 3056 1964 3108 1970
rect 3516 1964 3568 1970
rect 3108 1924 3280 1952
rect 3056 1906 3108 1912
rect 2964 1284 3016 1290
rect 2964 1226 3016 1232
rect 2976 160 3004 1226
rect 3252 160 3280 1924
rect 3516 1906 3568 1912
rect 3700 1964 3752 1970
rect 3700 1906 3752 1912
rect 3332 1760 3384 1766
rect 3332 1702 3384 1708
rect 3344 1562 3372 1702
rect 3332 1556 3384 1562
rect 3332 1498 3384 1504
rect 3528 160 3556 1906
rect 2134 54 2268 82
rect 1858 0 1914 54
rect 2134 0 2190 54
rect 2410 0 2466 160
rect 2686 0 2742 160
rect 2962 0 3018 160
rect 3238 0 3294 160
rect 3514 0 3570 160
rect 3712 82 3740 1906
rect 3804 1358 3832 8327
rect 4172 8294 4200 9046
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 3917 8188 4225 8197
rect 3917 8186 3923 8188
rect 3979 8186 4003 8188
rect 4059 8186 4083 8188
rect 4139 8186 4163 8188
rect 4219 8186 4225 8188
rect 3979 8134 3981 8186
rect 4161 8134 4163 8186
rect 3917 8132 3923 8134
rect 3979 8132 4003 8134
rect 4059 8132 4083 8134
rect 4139 8132 4163 8134
rect 4219 8132 4225 8134
rect 3917 8123 4225 8132
rect 4264 7546 4292 11154
rect 4356 10130 4384 11308
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4356 9178 4384 9522
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4356 8090 4384 9114
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4448 7392 4476 14878
rect 4724 14482 4752 14894
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4712 14340 4764 14346
rect 4712 14282 4764 14288
rect 4724 13394 4752 14282
rect 4816 13394 4844 16050
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4540 12986 4568 13330
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4618 12880 4674 12889
rect 4618 12815 4620 12824
rect 4672 12815 4674 12824
rect 4620 12786 4672 12792
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4540 9586 4568 12378
rect 4632 12345 4660 12786
rect 4618 12336 4674 12345
rect 4618 12271 4674 12280
rect 4724 12288 4752 13330
rect 4724 12260 4844 12288
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4632 11694 4660 12174
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4632 11354 4660 11494
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4540 9178 4568 9318
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4632 9058 4660 9318
rect 4724 9178 4752 12106
rect 4816 11626 4844 12260
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 4802 11248 4858 11257
rect 4802 11183 4804 11192
rect 4856 11183 4858 11192
rect 4804 11154 4856 11160
rect 4802 10160 4858 10169
rect 4802 10095 4858 10104
rect 4816 10062 4844 10095
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4540 9042 4660 9058
rect 4528 9036 4660 9042
rect 4580 9030 4660 9036
rect 4528 8978 4580 8984
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4724 8838 4752 8910
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4264 7364 4476 7392
rect 3917 7100 4225 7109
rect 3917 7098 3923 7100
rect 3979 7098 4003 7100
rect 4059 7098 4083 7100
rect 4139 7098 4163 7100
rect 4219 7098 4225 7100
rect 3979 7046 3981 7098
rect 4161 7046 4163 7098
rect 3917 7044 3923 7046
rect 3979 7044 4003 7046
rect 4059 7044 4083 7046
rect 4139 7044 4163 7046
rect 4219 7044 4225 7046
rect 3917 7035 4225 7044
rect 3917 6012 4225 6021
rect 3917 6010 3923 6012
rect 3979 6010 4003 6012
rect 4059 6010 4083 6012
rect 4139 6010 4163 6012
rect 4219 6010 4225 6012
rect 3979 5958 3981 6010
rect 4161 5958 4163 6010
rect 3917 5956 3923 5958
rect 3979 5956 4003 5958
rect 4059 5956 4083 5958
rect 4139 5956 4163 5958
rect 4219 5956 4225 5958
rect 3917 5947 4225 5956
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4080 5370 4108 5646
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4080 5166 4108 5306
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3917 4924 4225 4933
rect 3917 4922 3923 4924
rect 3979 4922 4003 4924
rect 4059 4922 4083 4924
rect 4139 4922 4163 4924
rect 4219 4922 4225 4924
rect 3979 4870 3981 4922
rect 4161 4870 4163 4922
rect 3917 4868 3923 4870
rect 3979 4868 4003 4870
rect 4059 4868 4083 4870
rect 4139 4868 4163 4870
rect 4219 4868 4225 4870
rect 3917 4859 4225 4868
rect 4066 4720 4122 4729
rect 4066 4655 4122 4664
rect 4080 4486 4108 4655
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3917 3836 4225 3845
rect 3917 3834 3923 3836
rect 3979 3834 4003 3836
rect 4059 3834 4083 3836
rect 4139 3834 4163 3836
rect 4219 3834 4225 3836
rect 3979 3782 3981 3834
rect 4161 3782 4163 3834
rect 3917 3780 3923 3782
rect 3979 3780 4003 3782
rect 4059 3780 4083 3782
rect 4139 3780 4163 3782
rect 4219 3780 4225 3782
rect 3917 3771 4225 3780
rect 3917 2748 4225 2757
rect 3917 2746 3923 2748
rect 3979 2746 4003 2748
rect 4059 2746 4083 2748
rect 4139 2746 4163 2748
rect 4219 2746 4225 2748
rect 3979 2694 3981 2746
rect 4161 2694 4163 2746
rect 3917 2692 3923 2694
rect 3979 2692 4003 2694
rect 4059 2692 4083 2694
rect 4139 2692 4163 2694
rect 4219 2692 4225 2694
rect 3917 2683 4225 2692
rect 4068 2304 4120 2310
rect 3974 2272 4030 2281
rect 4068 2246 4120 2252
rect 3974 2207 4030 2216
rect 3988 2106 4016 2207
rect 4080 2106 4108 2246
rect 4264 2106 4292 7364
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4356 6458 4384 6598
rect 4632 6497 4660 6598
rect 4618 6488 4674 6497
rect 4344 6452 4396 6458
rect 4618 6423 4674 6432
rect 4344 6394 4396 6400
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4436 6248 4488 6254
rect 4632 6225 4660 6258
rect 4436 6190 4488 6196
rect 4618 6216 4674 6225
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4356 5370 4384 6122
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4448 4146 4476 6190
rect 4618 6151 4674 6160
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4540 5234 4568 5510
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4724 4826 4752 6938
rect 4816 5234 4844 9998
rect 4908 9042 4936 18022
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 5000 16114 5028 16390
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 5000 13394 5028 13670
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5092 13240 5120 23802
rect 5184 22234 5212 25162
rect 5276 23730 5304 27900
rect 5552 27860 5580 28036
rect 5368 27832 5580 27860
rect 5368 26246 5396 27832
rect 5540 27668 5592 27674
rect 5540 27610 5592 27616
rect 5448 27464 5500 27470
rect 5446 27432 5448 27441
rect 5500 27432 5502 27441
rect 5446 27367 5502 27376
rect 5448 27328 5500 27334
rect 5448 27270 5500 27276
rect 5460 26586 5488 27270
rect 5448 26580 5500 26586
rect 5448 26522 5500 26528
rect 5448 26444 5500 26450
rect 5448 26386 5500 26392
rect 5356 26240 5408 26246
rect 5356 26182 5408 26188
rect 5368 24682 5396 26182
rect 5460 25906 5488 26386
rect 5448 25900 5500 25906
rect 5448 25842 5500 25848
rect 5446 25800 5502 25809
rect 5446 25735 5502 25744
rect 5460 24818 5488 25735
rect 5448 24812 5500 24818
rect 5448 24754 5500 24760
rect 5356 24676 5408 24682
rect 5356 24618 5408 24624
rect 5356 23860 5408 23866
rect 5356 23802 5408 23808
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5172 22228 5224 22234
rect 5172 22170 5224 22176
rect 5172 20460 5224 20466
rect 5172 20402 5224 20408
rect 5184 20058 5212 20402
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 5184 18290 5212 18566
rect 5172 18284 5224 18290
rect 5172 18226 5224 18232
rect 5276 18086 5304 23666
rect 5368 22642 5396 23802
rect 5552 23746 5580 27610
rect 5644 26081 5672 33322
rect 5828 33318 5856 34700
rect 6012 34660 6040 38150
rect 6090 37904 6146 37913
rect 6196 37890 6224 39630
rect 6276 39092 6328 39098
rect 6276 39034 6328 39040
rect 6146 37862 6224 37890
rect 6090 37839 6146 37848
rect 6184 37120 6236 37126
rect 6184 37062 6236 37068
rect 6196 36242 6224 37062
rect 6184 36236 6236 36242
rect 6184 36178 6236 36184
rect 6196 35698 6224 36178
rect 6184 35692 6236 35698
rect 6184 35634 6236 35640
rect 6184 35284 6236 35290
rect 6184 35226 6236 35232
rect 5920 34632 6040 34660
rect 5920 33998 5948 34632
rect 6196 34610 6224 35226
rect 6184 34604 6236 34610
rect 6184 34546 6236 34552
rect 6288 34490 6316 39034
rect 6012 34462 6316 34490
rect 5908 33992 5960 33998
rect 5908 33934 5960 33940
rect 5816 33312 5868 33318
rect 5816 33254 5868 33260
rect 5722 32872 5778 32881
rect 5722 32807 5724 32816
rect 5776 32807 5778 32816
rect 5724 32778 5776 32784
rect 5722 32328 5778 32337
rect 5722 32263 5778 32272
rect 5736 31657 5764 32263
rect 5908 31680 5960 31686
rect 5722 31648 5778 31657
rect 5908 31622 5960 31628
rect 5722 31583 5778 31592
rect 5736 31346 5764 31583
rect 5724 31340 5776 31346
rect 5724 31282 5776 31288
rect 5920 31226 5948 31622
rect 5828 31198 5948 31226
rect 5724 30660 5776 30666
rect 5724 30602 5776 30608
rect 5630 26072 5686 26081
rect 5630 26007 5686 26016
rect 5644 25838 5672 26007
rect 5632 25832 5684 25838
rect 5632 25774 5684 25780
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5644 25129 5672 25230
rect 5630 25120 5686 25129
rect 5630 25055 5686 25064
rect 5552 23718 5672 23746
rect 5540 23656 5592 23662
rect 5540 23598 5592 23604
rect 5446 23352 5502 23361
rect 5552 23322 5580 23598
rect 5446 23287 5502 23296
rect 5540 23316 5592 23322
rect 5460 23118 5488 23287
rect 5540 23258 5592 23264
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5356 22636 5408 22642
rect 5356 22578 5408 22584
rect 5460 22094 5488 22918
rect 5552 22574 5580 23258
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 5540 22432 5592 22438
rect 5540 22374 5592 22380
rect 5552 22098 5580 22374
rect 5368 22066 5488 22094
rect 5540 22092 5592 22098
rect 5368 20890 5396 22066
rect 5644 22094 5672 23718
rect 5736 22817 5764 30602
rect 5722 22808 5778 22817
rect 5722 22743 5778 22752
rect 5828 22094 5856 31198
rect 5908 31136 5960 31142
rect 5908 31078 5960 31084
rect 5920 30802 5948 31078
rect 5908 30796 5960 30802
rect 5908 30738 5960 30744
rect 5908 30592 5960 30598
rect 5906 30560 5908 30569
rect 5960 30560 5962 30569
rect 5906 30495 5962 30504
rect 5908 30048 5960 30054
rect 5908 29990 5960 29996
rect 5920 29714 5948 29990
rect 5908 29708 5960 29714
rect 5908 29650 5960 29656
rect 5908 29504 5960 29510
rect 5908 29446 5960 29452
rect 5920 29209 5948 29446
rect 5906 29200 5962 29209
rect 5906 29135 5962 29144
rect 5906 28792 5962 28801
rect 5906 28727 5908 28736
rect 5960 28727 5962 28736
rect 5908 28698 5960 28704
rect 5908 28552 5960 28558
rect 5908 28494 5960 28500
rect 5920 28082 5948 28494
rect 5908 28076 5960 28082
rect 5908 28018 5960 28024
rect 5906 27976 5962 27985
rect 5906 27911 5908 27920
rect 5960 27911 5962 27920
rect 5908 27882 5960 27888
rect 5908 27532 5960 27538
rect 5908 27474 5960 27480
rect 5920 27441 5948 27474
rect 5906 27432 5962 27441
rect 5906 27367 5962 27376
rect 5906 27160 5962 27169
rect 5906 27095 5962 27104
rect 5920 24857 5948 27095
rect 5906 24848 5962 24857
rect 5906 24783 5908 24792
rect 5960 24783 5962 24792
rect 5908 24754 5960 24760
rect 6012 22098 6040 34462
rect 6092 34400 6144 34406
rect 6092 34342 6144 34348
rect 6184 34400 6236 34406
rect 6184 34342 6236 34348
rect 6104 33930 6132 34342
rect 6092 33924 6144 33930
rect 6092 33866 6144 33872
rect 6196 33454 6224 34342
rect 6184 33448 6236 33454
rect 6184 33390 6236 33396
rect 6276 33448 6328 33454
rect 6276 33390 6328 33396
rect 6092 33312 6144 33318
rect 6092 33254 6144 33260
rect 6104 30977 6132 33254
rect 6182 31784 6238 31793
rect 6182 31719 6184 31728
rect 6236 31719 6238 31728
rect 6184 31690 6236 31696
rect 6182 31104 6238 31113
rect 6288 31090 6316 33390
rect 6380 31210 6408 41006
rect 6460 40384 6512 40390
rect 6460 40326 6512 40332
rect 6472 39982 6500 40326
rect 6460 39976 6512 39982
rect 6460 39918 6512 39924
rect 6472 39098 6500 39918
rect 6460 39092 6512 39098
rect 6460 39034 6512 39040
rect 6460 37732 6512 37738
rect 6460 37674 6512 37680
rect 6472 37330 6500 37674
rect 6460 37324 6512 37330
rect 6460 37266 6512 37272
rect 6460 35760 6512 35766
rect 6460 35702 6512 35708
rect 6472 32842 6500 35702
rect 6564 34105 6592 41074
rect 6826 40624 6882 40633
rect 6826 40559 6882 40568
rect 6840 40526 6868 40559
rect 6828 40520 6880 40526
rect 6920 40520 6972 40526
rect 6828 40462 6880 40468
rect 6918 40488 6920 40497
rect 6972 40488 6974 40497
rect 6918 40423 6974 40432
rect 6736 40384 6788 40390
rect 6736 40326 6788 40332
rect 6748 39574 6776 40326
rect 6884 40284 7192 40293
rect 6884 40282 6890 40284
rect 6946 40282 6970 40284
rect 7026 40282 7050 40284
rect 7106 40282 7130 40284
rect 7186 40282 7192 40284
rect 6946 40230 6948 40282
rect 7128 40230 7130 40282
rect 6884 40228 6890 40230
rect 6946 40228 6970 40230
rect 7026 40228 7050 40230
rect 7106 40228 7130 40230
rect 7186 40228 7192 40230
rect 6884 40219 7192 40228
rect 6828 40044 6880 40050
rect 6828 39986 6880 39992
rect 6736 39568 6788 39574
rect 6840 39545 6868 39986
rect 6736 39510 6788 39516
rect 6826 39536 6882 39545
rect 6644 39500 6696 39506
rect 6826 39471 6882 39480
rect 7010 39536 7066 39545
rect 7010 39471 7066 39480
rect 6644 39442 6696 39448
rect 6656 39098 6684 39442
rect 6840 39420 6868 39471
rect 7024 39438 7052 39471
rect 6748 39392 6868 39420
rect 7012 39432 7064 39438
rect 6644 39092 6696 39098
rect 6644 39034 6696 39040
rect 6656 39001 6684 39034
rect 6642 38992 6698 39001
rect 6642 38927 6698 38936
rect 6748 38554 6776 39392
rect 7012 39374 7064 39380
rect 7196 39432 7248 39438
rect 7196 39374 7248 39380
rect 7208 39302 7236 39374
rect 7196 39296 7248 39302
rect 7196 39238 7248 39244
rect 6884 39196 7192 39205
rect 6884 39194 6890 39196
rect 6946 39194 6970 39196
rect 7026 39194 7050 39196
rect 7106 39194 7130 39196
rect 7186 39194 7192 39196
rect 6946 39142 6948 39194
rect 7128 39142 7130 39194
rect 6884 39140 6890 39142
rect 6946 39140 6970 39142
rect 7026 39140 7050 39142
rect 7106 39140 7130 39142
rect 7186 39140 7192 39142
rect 6884 39131 7192 39140
rect 7286 38992 7342 39001
rect 7196 38956 7248 38962
rect 7248 38936 7286 38944
rect 7248 38927 7342 38936
rect 7248 38916 7328 38927
rect 7196 38898 7248 38904
rect 7392 38593 7420 41074
rect 7472 40520 7524 40526
rect 7524 40480 7604 40508
rect 7472 40462 7524 40468
rect 7472 39840 7524 39846
rect 7472 39782 7524 39788
rect 7484 39506 7512 39782
rect 7472 39500 7524 39506
rect 7472 39442 7524 39448
rect 7576 39386 7604 40480
rect 7484 39358 7604 39386
rect 7378 38584 7434 38593
rect 6736 38548 6788 38554
rect 7378 38519 7434 38528
rect 6736 38490 6788 38496
rect 7288 38344 7340 38350
rect 7484 38332 7512 39358
rect 7340 38304 7512 38332
rect 7288 38286 7340 38292
rect 6884 38108 7192 38117
rect 6884 38106 6890 38108
rect 6946 38106 6970 38108
rect 7026 38106 7050 38108
rect 7106 38106 7130 38108
rect 7186 38106 7192 38108
rect 6946 38054 6948 38106
rect 7128 38054 7130 38106
rect 6884 38052 6890 38054
rect 6946 38052 6970 38054
rect 7026 38052 7050 38054
rect 7106 38052 7130 38054
rect 7186 38052 7192 38054
rect 6884 38043 7192 38052
rect 6736 38004 6788 38010
rect 6736 37946 6788 37952
rect 6644 37732 6696 37738
rect 6644 37674 6696 37680
rect 6656 37194 6684 37674
rect 6644 37188 6696 37194
rect 6644 37130 6696 37136
rect 6748 37126 6776 37946
rect 7300 37126 7328 38286
rect 7668 38026 7696 42316
rect 7748 42220 7800 42226
rect 7748 42162 7800 42168
rect 7392 37998 7696 38026
rect 6736 37120 6788 37126
rect 6736 37062 6788 37068
rect 7288 37120 7340 37126
rect 7288 37062 7340 37068
rect 6642 35592 6698 35601
rect 6642 35527 6698 35536
rect 6656 34678 6684 35527
rect 6644 34672 6696 34678
rect 6642 34640 6644 34649
rect 6696 34640 6698 34649
rect 6642 34575 6698 34584
rect 6642 34504 6698 34513
rect 6642 34439 6698 34448
rect 6550 34096 6606 34105
rect 6550 34031 6606 34040
rect 6552 33856 6604 33862
rect 6552 33798 6604 33804
rect 6564 32978 6592 33798
rect 6552 32972 6604 32978
rect 6552 32914 6604 32920
rect 6460 32836 6512 32842
rect 6460 32778 6512 32784
rect 6552 32836 6604 32842
rect 6552 32778 6604 32784
rect 6564 32026 6592 32778
rect 6460 32020 6512 32026
rect 6460 31962 6512 31968
rect 6552 32020 6604 32026
rect 6552 31962 6604 31968
rect 6472 31822 6500 31962
rect 6460 31816 6512 31822
rect 6460 31758 6512 31764
rect 6368 31204 6420 31210
rect 6368 31146 6420 31152
rect 6288 31062 6408 31090
rect 6182 31039 6238 31048
rect 6090 30968 6146 30977
rect 6090 30903 6092 30912
rect 6144 30903 6146 30912
rect 6092 30874 6144 30880
rect 6196 30394 6224 31039
rect 6184 30388 6236 30394
rect 6184 30330 6236 30336
rect 6276 30252 6328 30258
rect 6276 30194 6328 30200
rect 6184 30184 6236 30190
rect 6288 30161 6316 30194
rect 6184 30126 6236 30132
rect 6274 30152 6330 30161
rect 6092 29164 6144 29170
rect 6092 29106 6144 29112
rect 6104 27674 6132 29106
rect 6092 27668 6144 27674
rect 6092 27610 6144 27616
rect 6092 25696 6144 25702
rect 6092 25638 6144 25644
rect 6104 25226 6132 25638
rect 6196 25378 6224 30126
rect 6274 30087 6330 30096
rect 6274 28792 6330 28801
rect 6274 28727 6330 28736
rect 6288 28558 6316 28727
rect 6276 28552 6328 28558
rect 6276 28494 6328 28500
rect 6288 27062 6316 28494
rect 6276 27056 6328 27062
rect 6276 26998 6328 27004
rect 6276 26240 6328 26246
rect 6276 26182 6328 26188
rect 6288 25498 6316 26182
rect 6276 25492 6328 25498
rect 6276 25434 6328 25440
rect 6274 25392 6330 25401
rect 6196 25350 6274 25378
rect 6274 25327 6330 25336
rect 6092 25220 6144 25226
rect 6092 25162 6144 25168
rect 6276 25152 6328 25158
rect 6276 25094 6328 25100
rect 6092 24676 6144 24682
rect 6092 24618 6144 24624
rect 5644 22066 5764 22094
rect 5828 22066 5948 22094
rect 5540 22034 5592 22040
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 5368 20862 5580 20890
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5356 20460 5408 20466
rect 5356 20402 5408 20408
rect 5368 19786 5396 20402
rect 5460 20398 5488 20742
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5552 20244 5580 20862
rect 5460 20216 5580 20244
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 5354 19408 5410 19417
rect 5354 19343 5410 19352
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5172 17672 5224 17678
rect 5368 17660 5396 19343
rect 5224 17632 5396 17660
rect 5172 17614 5224 17620
rect 5025 13212 5120 13240
rect 5025 13138 5053 13212
rect 5000 13110 5053 13138
rect 5000 11218 5028 13110
rect 5184 12442 5212 17614
rect 5460 17218 5488 20216
rect 5644 19553 5672 21966
rect 5630 19544 5686 19553
rect 5630 19479 5686 19488
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5552 18766 5580 19246
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5368 17190 5488 17218
rect 5368 16590 5396 17190
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5264 15496 5316 15502
rect 5262 15464 5264 15473
rect 5316 15464 5318 15473
rect 5262 15399 5318 15408
rect 5368 15042 5396 16526
rect 5460 16522 5488 17070
rect 5448 16516 5500 16522
rect 5448 16458 5500 16464
rect 5552 16182 5580 18022
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 5644 15978 5672 19479
rect 5736 16114 5764 22066
rect 5920 21185 5948 22066
rect 6000 22092 6052 22098
rect 6000 22034 6052 22040
rect 6000 21956 6052 21962
rect 6000 21898 6052 21904
rect 5906 21176 5962 21185
rect 5906 21111 5962 21120
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5920 19334 5948 20334
rect 5828 19306 5948 19334
rect 5828 17678 5856 19306
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5920 18086 5948 18362
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 6012 17898 6040 21898
rect 6104 20380 6132 24618
rect 6184 23520 6236 23526
rect 6184 23462 6236 23468
rect 6196 23118 6224 23462
rect 6288 23338 6316 25094
rect 6380 23497 6408 31062
rect 6460 30932 6512 30938
rect 6512 30892 6592 30920
rect 6460 30874 6512 30880
rect 6564 28994 6592 30892
rect 6656 29646 6684 34439
rect 6748 33590 6776 37062
rect 6884 37020 7192 37029
rect 6884 37018 6890 37020
rect 6946 37018 6970 37020
rect 7026 37018 7050 37020
rect 7106 37018 7130 37020
rect 7186 37018 7192 37020
rect 6946 36966 6948 37018
rect 7128 36966 7130 37018
rect 6884 36964 6890 36966
rect 6946 36964 6970 36966
rect 7026 36964 7050 36966
rect 7106 36964 7130 36966
rect 7186 36964 7192 36966
rect 6884 36955 7192 36964
rect 7196 36916 7248 36922
rect 7300 36904 7328 37062
rect 7248 36876 7328 36904
rect 7196 36858 7248 36864
rect 7196 36780 7248 36786
rect 7196 36722 7248 36728
rect 7208 36378 7236 36722
rect 7196 36372 7248 36378
rect 7196 36314 7248 36320
rect 7288 36168 7340 36174
rect 7288 36110 7340 36116
rect 6884 35932 7192 35941
rect 6884 35930 6890 35932
rect 6946 35930 6970 35932
rect 7026 35930 7050 35932
rect 7106 35930 7130 35932
rect 7186 35930 7192 35932
rect 6946 35878 6948 35930
rect 7128 35878 7130 35930
rect 6884 35876 6890 35878
rect 6946 35876 6970 35878
rect 7026 35876 7050 35878
rect 7106 35876 7130 35878
rect 7186 35876 7192 35878
rect 6884 35867 7192 35876
rect 7300 35834 7328 36110
rect 7288 35828 7340 35834
rect 7288 35770 7340 35776
rect 7392 35766 7420 37998
rect 7564 37868 7616 37874
rect 7564 37810 7616 37816
rect 7472 37392 7524 37398
rect 7472 37334 7524 37340
rect 7380 35760 7432 35766
rect 7380 35702 7432 35708
rect 6884 34844 7192 34853
rect 6884 34842 6890 34844
rect 6946 34842 6970 34844
rect 7026 34842 7050 34844
rect 7106 34842 7130 34844
rect 7186 34842 7192 34844
rect 6946 34790 6948 34842
rect 7128 34790 7130 34842
rect 6884 34788 6890 34790
rect 6946 34788 6970 34790
rect 7026 34788 7050 34790
rect 7106 34788 7130 34790
rect 7186 34788 7192 34790
rect 6884 34779 7192 34788
rect 6828 34400 6880 34406
rect 6828 34342 6880 34348
rect 6840 34066 6868 34342
rect 6828 34060 6880 34066
rect 6828 34002 6880 34008
rect 6840 33844 6868 34002
rect 6822 33816 6868 33844
rect 7380 33856 7432 33862
rect 6822 33640 6850 33816
rect 7380 33798 7432 33804
rect 6884 33756 7192 33765
rect 6884 33754 6890 33756
rect 6946 33754 6970 33756
rect 7026 33754 7050 33756
rect 7106 33754 7130 33756
rect 7186 33754 7192 33756
rect 6946 33702 6948 33754
rect 7128 33702 7130 33754
rect 6884 33700 6890 33702
rect 6946 33700 6970 33702
rect 7026 33700 7050 33702
rect 7106 33700 7130 33702
rect 7186 33700 7192 33702
rect 6884 33691 7192 33700
rect 6822 33612 6868 33640
rect 6736 33584 6788 33590
rect 6736 33526 6788 33532
rect 6840 33522 6868 33612
rect 6828 33516 6880 33522
rect 6828 33458 6880 33464
rect 6840 32756 6868 33458
rect 7102 33008 7158 33017
rect 7102 32943 7158 32952
rect 7288 32972 7340 32978
rect 6918 32872 6974 32881
rect 7116 32842 7144 32943
rect 7288 32914 7340 32920
rect 6918 32807 6920 32816
rect 6972 32807 6974 32816
rect 7104 32836 7156 32842
rect 6920 32778 6972 32784
rect 7104 32778 7156 32784
rect 6822 32728 6868 32756
rect 6734 32600 6790 32609
rect 6734 32535 6790 32544
rect 6822 32552 6850 32728
rect 6884 32668 7192 32677
rect 6884 32666 6890 32668
rect 6946 32666 6970 32668
rect 7026 32666 7050 32668
rect 7106 32666 7130 32668
rect 7186 32666 7192 32668
rect 6946 32614 6948 32666
rect 7128 32614 7130 32666
rect 6884 32612 6890 32614
rect 6946 32612 6970 32614
rect 7026 32612 7050 32614
rect 7106 32612 7130 32614
rect 7186 32612 7192 32614
rect 6884 32603 7192 32612
rect 7300 32552 7328 32914
rect 6748 32502 6776 32535
rect 6822 32524 6960 32552
rect 6736 32496 6788 32502
rect 6736 32438 6788 32444
rect 6932 31890 6960 32524
rect 7208 32524 7328 32552
rect 6920 31884 6972 31890
rect 6920 31826 6972 31832
rect 6828 31816 6880 31822
rect 6748 31776 6828 31804
rect 6644 29640 6696 29646
rect 6644 29582 6696 29588
rect 6644 29096 6696 29102
rect 6644 29038 6696 29044
rect 6472 28966 6592 28994
rect 6472 27470 6500 28966
rect 6656 28558 6684 29038
rect 6552 28552 6604 28558
rect 6552 28494 6604 28500
rect 6644 28552 6696 28558
rect 6644 28494 6696 28500
rect 6564 28393 6592 28494
rect 6550 28384 6606 28393
rect 6550 28319 6606 28328
rect 6550 28248 6606 28257
rect 6550 28183 6552 28192
rect 6604 28183 6606 28192
rect 6552 28154 6604 28160
rect 6644 28008 6696 28014
rect 6644 27950 6696 27956
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 6472 26625 6500 27406
rect 6458 26616 6514 26625
rect 6458 26551 6514 26560
rect 6460 26512 6512 26518
rect 6460 26454 6512 26460
rect 6472 25158 6500 26454
rect 6656 26450 6684 27950
rect 6748 26489 6776 31776
rect 6828 31758 6880 31764
rect 7208 31668 7236 32524
rect 7208 31640 7328 31668
rect 6884 31580 7192 31589
rect 6884 31578 6890 31580
rect 6946 31578 6970 31580
rect 7026 31578 7050 31580
rect 7106 31578 7130 31580
rect 7186 31578 7192 31580
rect 6946 31526 6948 31578
rect 7128 31526 7130 31578
rect 6884 31524 6890 31526
rect 6946 31524 6970 31526
rect 7026 31524 7050 31526
rect 7106 31524 7130 31526
rect 7186 31524 7192 31526
rect 6884 31515 7192 31524
rect 7300 30734 7328 31640
rect 7392 30938 7420 33798
rect 7484 33114 7512 37334
rect 7576 36922 7604 37810
rect 7656 37800 7708 37806
rect 7656 37742 7708 37748
rect 7668 37466 7696 37742
rect 7656 37460 7708 37466
rect 7656 37402 7708 37408
rect 7668 37262 7696 37402
rect 7760 37369 7788 42162
rect 7840 42152 7892 42158
rect 7840 42094 7892 42100
rect 7852 41414 7880 42094
rect 7944 41818 7972 42502
rect 8024 42220 8076 42226
rect 8024 42162 8076 42168
rect 7932 41812 7984 41818
rect 7932 41754 7984 41760
rect 7852 41386 7972 41414
rect 7840 41268 7892 41274
rect 7840 41210 7892 41216
rect 7746 37360 7802 37369
rect 7746 37295 7802 37304
rect 7656 37256 7708 37262
rect 7656 37198 7708 37204
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 7564 36916 7616 36922
rect 7564 36858 7616 36864
rect 7656 36780 7708 36786
rect 7656 36722 7708 36728
rect 7564 36712 7616 36718
rect 7564 36654 7616 36660
rect 7576 35086 7604 36654
rect 7668 36378 7696 36722
rect 7656 36372 7708 36378
rect 7656 36314 7708 36320
rect 7760 35290 7788 37062
rect 7748 35284 7800 35290
rect 7748 35226 7800 35232
rect 7564 35080 7616 35086
rect 7564 35022 7616 35028
rect 7564 34944 7616 34950
rect 7564 34886 7616 34892
rect 7472 33108 7524 33114
rect 7472 33050 7524 33056
rect 7472 32768 7524 32774
rect 7472 32710 7524 32716
rect 7484 32502 7512 32710
rect 7472 32496 7524 32502
rect 7576 32473 7604 34886
rect 7760 34610 7788 35226
rect 7748 34604 7800 34610
rect 7748 34546 7800 34552
rect 7656 33652 7708 33658
rect 7656 33594 7708 33600
rect 7668 33046 7696 33594
rect 7656 33040 7708 33046
rect 7656 32982 7708 32988
rect 7748 32496 7800 32502
rect 7472 32438 7524 32444
rect 7562 32464 7618 32473
rect 7748 32438 7800 32444
rect 7562 32399 7618 32408
rect 7562 31920 7618 31929
rect 7472 31884 7524 31890
rect 7562 31855 7618 31864
rect 7472 31826 7524 31832
rect 7484 31346 7512 31826
rect 7576 31754 7604 31855
rect 7656 31816 7708 31822
rect 7656 31758 7708 31764
rect 7564 31748 7616 31754
rect 7564 31690 7616 31696
rect 7564 31408 7616 31414
rect 7564 31350 7616 31356
rect 7472 31340 7524 31346
rect 7472 31282 7524 31288
rect 7380 30932 7432 30938
rect 7380 30874 7432 30880
rect 7484 30802 7512 31282
rect 7472 30796 7524 30802
rect 7472 30738 7524 30744
rect 7288 30728 7340 30734
rect 7288 30670 7340 30676
rect 6884 30492 7192 30501
rect 6884 30490 6890 30492
rect 6946 30490 6970 30492
rect 7026 30490 7050 30492
rect 7106 30490 7130 30492
rect 7186 30490 7192 30492
rect 6946 30438 6948 30490
rect 7128 30438 7130 30490
rect 6884 30436 6890 30438
rect 6946 30436 6970 30438
rect 7026 30436 7050 30438
rect 7106 30436 7130 30438
rect 7186 30436 7192 30438
rect 6884 30427 7192 30436
rect 7194 29880 7250 29889
rect 7194 29815 7250 29824
rect 7208 29578 7236 29815
rect 7196 29572 7248 29578
rect 7196 29514 7248 29520
rect 6884 29404 7192 29413
rect 6884 29402 6890 29404
rect 6946 29402 6970 29404
rect 7026 29402 7050 29404
rect 7106 29402 7130 29404
rect 7186 29402 7192 29404
rect 6946 29350 6948 29402
rect 7128 29350 7130 29402
rect 6884 29348 6890 29350
rect 6946 29348 6970 29350
rect 7026 29348 7050 29350
rect 7106 29348 7130 29350
rect 7186 29348 7192 29350
rect 6884 29339 7192 29348
rect 7300 29034 7328 30670
rect 7380 30048 7432 30054
rect 7380 29990 7432 29996
rect 7392 29646 7420 29990
rect 7380 29640 7432 29646
rect 7380 29582 7432 29588
rect 7380 29096 7432 29102
rect 7380 29038 7432 29044
rect 7288 29028 7340 29034
rect 7288 28970 7340 28976
rect 7288 28416 7340 28422
rect 7288 28358 7340 28364
rect 6884 28316 7192 28325
rect 6884 28314 6890 28316
rect 6946 28314 6970 28316
rect 7026 28314 7050 28316
rect 7106 28314 7130 28316
rect 7186 28314 7192 28316
rect 6946 28262 6948 28314
rect 7128 28262 7130 28314
rect 6884 28260 6890 28262
rect 6946 28260 6970 28262
rect 7026 28260 7050 28262
rect 7106 28260 7130 28262
rect 7186 28260 7192 28262
rect 6884 28251 7192 28260
rect 6918 28112 6974 28121
rect 6918 28047 6974 28056
rect 6932 27402 6960 28047
rect 7300 27470 7328 28358
rect 7392 28150 7420 29038
rect 7484 28801 7512 30738
rect 7576 30598 7604 31350
rect 7564 30592 7616 30598
rect 7564 30534 7616 30540
rect 7668 30410 7696 31758
rect 7760 31521 7788 32438
rect 7746 31512 7802 31521
rect 7746 31447 7802 31456
rect 7852 30705 7880 41210
rect 7944 40730 7972 41386
rect 7932 40724 7984 40730
rect 7932 40666 7984 40672
rect 7932 39364 7984 39370
rect 7932 39306 7984 39312
rect 7944 38962 7972 39306
rect 7932 38956 7984 38962
rect 7932 38898 7984 38904
rect 7944 37738 7972 38898
rect 8036 37777 8064 42162
rect 8128 42129 8156 42638
rect 8220 42362 8248 43302
rect 8300 43308 8352 43314
rect 8300 43250 8352 43256
rect 8312 42906 8340 43250
rect 8300 42900 8352 42906
rect 8300 42842 8352 42848
rect 8772 42770 8800 44840
rect 8944 44804 8996 44810
rect 8944 44746 8996 44752
rect 8956 43450 8984 44746
rect 9048 43450 9076 44840
rect 9508 44554 9536 44934
rect 9586 44840 9642 45000
rect 9862 44840 9918 45000
rect 10138 44962 10194 45000
rect 10414 44962 10470 45000
rect 9968 44934 10194 44962
rect 9600 44810 9628 44840
rect 9588 44804 9640 44810
rect 9588 44746 9640 44752
rect 9508 44526 9628 44554
rect 9128 43648 9180 43654
rect 9128 43590 9180 43596
rect 8944 43444 8996 43450
rect 8944 43386 8996 43392
rect 9036 43444 9088 43450
rect 9036 43386 9088 43392
rect 9140 42786 9168 43590
rect 8760 42764 8812 42770
rect 8760 42706 8812 42712
rect 8956 42758 9168 42786
rect 9600 42786 9628 44526
rect 9876 43450 9904 44840
rect 9864 43444 9916 43450
rect 9864 43386 9916 43392
rect 9968 43314 9996 44934
rect 10138 44840 10194 44934
rect 10336 44934 10470 44962
rect 10336 43314 10364 44934
rect 10414 44840 10470 44934
rect 10690 44840 10746 45000
rect 10966 44840 11022 45000
rect 11242 44840 11298 45000
rect 11518 44962 11574 45000
rect 11794 44962 11850 45000
rect 11518 44934 11652 44962
rect 11518 44840 11574 44934
rect 10508 43716 10560 43722
rect 10508 43658 10560 43664
rect 10520 43450 10548 43658
rect 10508 43444 10560 43450
rect 10508 43386 10560 43392
rect 10704 43314 10732 44840
rect 10980 44146 11008 44840
rect 10980 44118 11100 44146
rect 11072 43314 11100 44118
rect 11256 43382 11284 44840
rect 11244 43376 11296 43382
rect 11244 43318 11296 43324
rect 9956 43308 10008 43314
rect 9956 43250 10008 43256
rect 10324 43308 10376 43314
rect 10324 43250 10376 43256
rect 10692 43308 10744 43314
rect 10692 43250 10744 43256
rect 11060 43308 11112 43314
rect 11060 43250 11112 43256
rect 10324 43172 10376 43178
rect 10324 43114 10376 43120
rect 9772 43104 9824 43110
rect 9772 43046 9824 43052
rect 9784 42838 9812 43046
rect 9851 43004 10159 43013
rect 9851 43002 9857 43004
rect 9913 43002 9937 43004
rect 9993 43002 10017 43004
rect 10073 43002 10097 43004
rect 10153 43002 10159 43004
rect 9913 42950 9915 43002
rect 10095 42950 10097 43002
rect 9851 42948 9857 42950
rect 9913 42948 9937 42950
rect 9993 42948 10017 42950
rect 10073 42948 10097 42950
rect 10153 42948 10159 42950
rect 9851 42939 10159 42948
rect 9772 42832 9824 42838
rect 9312 42764 9364 42770
rect 8300 42560 8352 42566
rect 8300 42502 8352 42508
rect 8208 42356 8260 42362
rect 8208 42298 8260 42304
rect 8312 42294 8340 42502
rect 8852 42356 8904 42362
rect 8852 42298 8904 42304
rect 8300 42288 8352 42294
rect 8300 42230 8352 42236
rect 8392 42220 8444 42226
rect 8392 42162 8444 42168
rect 8668 42220 8720 42226
rect 8668 42162 8720 42168
rect 8114 42120 8170 42129
rect 8114 42055 8170 42064
rect 8208 42084 8260 42090
rect 8208 42026 8260 42032
rect 8220 41818 8248 42026
rect 8300 42016 8352 42022
rect 8300 41958 8352 41964
rect 8312 41818 8340 41958
rect 8404 41818 8432 42162
rect 8208 41812 8260 41818
rect 8208 41754 8260 41760
rect 8300 41812 8352 41818
rect 8300 41754 8352 41760
rect 8392 41812 8444 41818
rect 8392 41754 8444 41760
rect 8576 41744 8628 41750
rect 8220 41692 8576 41698
rect 8220 41686 8628 41692
rect 8220 41670 8616 41686
rect 8220 41274 8248 41670
rect 8208 41268 8260 41274
rect 8208 41210 8260 41216
rect 8116 41132 8168 41138
rect 8116 41074 8168 41080
rect 8208 41132 8260 41138
rect 8208 41074 8260 41080
rect 8022 37768 8078 37777
rect 7932 37732 7984 37738
rect 8022 37703 8078 37712
rect 7932 37674 7984 37680
rect 7944 36009 7972 37674
rect 8128 37262 8156 41074
rect 8220 40089 8248 41074
rect 8576 40724 8628 40730
rect 8680 40712 8708 42162
rect 8628 40684 8708 40712
rect 8576 40666 8628 40672
rect 8300 40520 8352 40526
rect 8298 40488 8300 40497
rect 8352 40488 8354 40497
rect 8354 40446 8432 40474
rect 8298 40423 8354 40432
rect 8404 40186 8432 40446
rect 8484 40384 8536 40390
rect 8484 40326 8536 40332
rect 8392 40180 8444 40186
rect 8392 40122 8444 40128
rect 8300 40112 8352 40118
rect 8206 40080 8262 40089
rect 8300 40054 8352 40060
rect 8206 40015 8262 40024
rect 8208 39500 8260 39506
rect 8208 39442 8260 39448
rect 8220 39001 8248 39442
rect 8312 39030 8340 40054
rect 8496 39982 8524 40326
rect 8588 40050 8616 40666
rect 8576 40044 8628 40050
rect 8576 39986 8628 39992
rect 8760 40044 8812 40050
rect 8760 39986 8812 39992
rect 8484 39976 8536 39982
rect 8772 39930 8800 39986
rect 8484 39918 8536 39924
rect 8680 39902 8800 39930
rect 8392 39636 8444 39642
rect 8392 39578 8444 39584
rect 8404 39098 8432 39578
rect 8392 39092 8444 39098
rect 8392 39034 8444 39040
rect 8300 39024 8352 39030
rect 8206 38992 8262 39001
rect 8300 38966 8352 38972
rect 8206 38927 8262 38936
rect 8206 38312 8262 38321
rect 8206 38247 8208 38256
rect 8260 38247 8262 38256
rect 8208 38218 8260 38224
rect 8312 37942 8340 38966
rect 8680 38962 8708 39902
rect 8668 38956 8720 38962
rect 8668 38898 8720 38904
rect 8392 38752 8444 38758
rect 8392 38694 8444 38700
rect 8404 38554 8432 38694
rect 8392 38548 8444 38554
rect 8392 38490 8444 38496
rect 8484 38208 8536 38214
rect 8484 38150 8536 38156
rect 8300 37936 8352 37942
rect 8300 37878 8352 37884
rect 8208 37664 8260 37670
rect 8208 37606 8260 37612
rect 8220 37330 8248 37606
rect 8208 37324 8260 37330
rect 8208 37266 8260 37272
rect 8024 37256 8076 37262
rect 8024 37198 8076 37204
rect 8116 37256 8168 37262
rect 8116 37198 8168 37204
rect 8036 36922 8064 37198
rect 8024 36916 8076 36922
rect 8024 36858 8076 36864
rect 8116 36372 8168 36378
rect 8116 36314 8168 36320
rect 8022 36136 8078 36145
rect 8022 36071 8078 36080
rect 7930 36000 7986 36009
rect 7930 35935 7986 35944
rect 8036 35086 8064 36071
rect 7932 35080 7984 35086
rect 7932 35022 7984 35028
rect 8024 35080 8076 35086
rect 8024 35022 8076 35028
rect 7944 33454 7972 35022
rect 8024 34672 8076 34678
rect 8128 34660 8156 36314
rect 8208 35760 8260 35766
rect 8312 35714 8340 37878
rect 8496 37806 8524 38150
rect 8680 37942 8708 38898
rect 8668 37936 8720 37942
rect 8668 37878 8720 37884
rect 8484 37800 8536 37806
rect 8484 37742 8536 37748
rect 8392 37120 8444 37126
rect 8392 37062 8444 37068
rect 8404 36038 8432 37062
rect 8392 36032 8444 36038
rect 8392 35974 8444 35980
rect 8680 35816 8708 37878
rect 8260 35708 8340 35714
rect 8208 35702 8340 35708
rect 8220 35686 8340 35702
rect 8496 35788 8708 35816
rect 8496 35698 8524 35788
rect 8208 35624 8260 35630
rect 8208 35566 8260 35572
rect 8220 35290 8248 35566
rect 8208 35284 8260 35290
rect 8208 35226 8260 35232
rect 8312 35086 8340 35686
rect 8392 35692 8444 35698
rect 8392 35634 8444 35640
rect 8484 35692 8536 35698
rect 8484 35634 8536 35640
rect 8668 35692 8720 35698
rect 8668 35634 8720 35640
rect 8760 35692 8812 35698
rect 8760 35634 8812 35640
rect 8300 35080 8352 35086
rect 8300 35022 8352 35028
rect 8404 34746 8432 35634
rect 8680 35476 8708 35634
rect 8772 35601 8800 35634
rect 8758 35592 8814 35601
rect 8758 35527 8814 35536
rect 8680 35448 8800 35476
rect 8668 35284 8720 35290
rect 8668 35226 8720 35232
rect 8484 35080 8536 35086
rect 8484 35022 8536 35028
rect 8300 34740 8352 34746
rect 8300 34682 8352 34688
rect 8392 34740 8444 34746
rect 8392 34682 8444 34688
rect 8076 34632 8156 34660
rect 8024 34614 8076 34620
rect 8312 34626 8340 34682
rect 7932 33448 7984 33454
rect 7930 33416 7932 33425
rect 7984 33416 7986 33425
rect 7930 33351 7986 33360
rect 8036 33300 8064 34614
rect 8312 34598 8432 34626
rect 8116 33856 8168 33862
rect 8116 33798 8168 33804
rect 8128 33454 8156 33798
rect 8116 33448 8168 33454
rect 8116 33390 8168 33396
rect 8298 33416 8354 33425
rect 7944 33272 8064 33300
rect 7944 32337 7972 33272
rect 8024 33108 8076 33114
rect 8024 33050 8076 33056
rect 7930 32328 7986 32337
rect 7930 32263 7986 32272
rect 7838 30696 7894 30705
rect 7838 30631 7894 30640
rect 7748 30592 7800 30598
rect 7748 30534 7800 30540
rect 7932 30592 7984 30598
rect 7932 30534 7984 30540
rect 7576 30382 7696 30410
rect 7470 28792 7526 28801
rect 7470 28727 7526 28736
rect 7484 28626 7512 28727
rect 7472 28620 7524 28626
rect 7472 28562 7524 28568
rect 7380 28144 7432 28150
rect 7380 28086 7432 28092
rect 7378 27568 7434 27577
rect 7378 27503 7434 27512
rect 7288 27464 7340 27470
rect 7288 27406 7340 27412
rect 6920 27396 6972 27402
rect 6972 27356 7144 27384
rect 6920 27338 6972 27344
rect 7116 27316 7144 27356
rect 7392 27334 7420 27503
rect 7576 27470 7604 30382
rect 7656 30252 7708 30258
rect 7656 30194 7708 30200
rect 7564 27464 7616 27470
rect 7564 27406 7616 27412
rect 7380 27328 7432 27334
rect 7116 27288 7328 27316
rect 6884 27228 7192 27237
rect 6884 27226 6890 27228
rect 6946 27226 6970 27228
rect 7026 27226 7050 27228
rect 7106 27226 7130 27228
rect 7186 27226 7192 27228
rect 6946 27174 6948 27226
rect 7128 27174 7130 27226
rect 6884 27172 6890 27174
rect 6946 27172 6970 27174
rect 7026 27172 7050 27174
rect 7106 27172 7130 27174
rect 7186 27172 7192 27174
rect 6884 27163 7192 27172
rect 6918 26752 6974 26761
rect 6918 26687 6974 26696
rect 6734 26480 6790 26489
rect 6644 26444 6696 26450
rect 6734 26415 6790 26424
rect 6644 26386 6696 26392
rect 6552 26036 6604 26042
rect 6552 25978 6604 25984
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6460 24200 6512 24206
rect 6460 24142 6512 24148
rect 6366 23488 6422 23497
rect 6366 23423 6422 23432
rect 6288 23310 6408 23338
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 6184 22976 6236 22982
rect 6184 22918 6236 22924
rect 6196 22574 6224 22918
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 6184 22432 6236 22438
rect 6184 22374 6236 22380
rect 6196 21962 6224 22374
rect 6184 21956 6236 21962
rect 6184 21898 6236 21904
rect 6184 21480 6236 21486
rect 6184 21422 6236 21428
rect 6196 20534 6224 21422
rect 6276 20936 6328 20942
rect 6276 20878 6328 20884
rect 6184 20528 6236 20534
rect 6184 20470 6236 20476
rect 6104 20352 6224 20380
rect 6196 20262 6224 20352
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6104 19825 6132 20198
rect 6090 19816 6146 19825
rect 6090 19751 6146 19760
rect 6090 19680 6146 19689
rect 6090 19615 6146 19624
rect 5920 17870 6040 17898
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5920 17270 5948 17870
rect 5998 17776 6054 17785
rect 5998 17711 6054 17720
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5460 15178 5488 15574
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 5460 15150 5764 15178
rect 5828 15162 5856 15506
rect 6012 15502 6040 17711
rect 6104 17678 6132 19615
rect 6288 19334 6316 20878
rect 6196 19306 6316 19334
rect 6196 18630 6224 19306
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 6196 17218 6224 18566
rect 6380 18086 6408 23310
rect 6472 21593 6500 24142
rect 6458 21584 6514 21593
rect 6458 21519 6514 21528
rect 6472 18306 6500 21519
rect 6564 18426 6592 25978
rect 6656 22438 6684 26386
rect 6932 26228 6960 26687
rect 7196 26512 7248 26518
rect 7196 26454 7248 26460
rect 7208 26314 7236 26454
rect 7196 26308 7248 26314
rect 7196 26250 7248 26256
rect 6748 26200 6960 26228
rect 6748 25922 6776 26200
rect 6884 26140 7192 26149
rect 6884 26138 6890 26140
rect 6946 26138 6970 26140
rect 7026 26138 7050 26140
rect 7106 26138 7130 26140
rect 7186 26138 7192 26140
rect 6946 26086 6948 26138
rect 7128 26086 7130 26138
rect 6884 26084 6890 26086
rect 6946 26084 6970 26086
rect 7026 26084 7050 26086
rect 7106 26084 7130 26086
rect 7186 26084 7192 26086
rect 6884 26075 7192 26084
rect 6748 25894 6960 25922
rect 6932 25140 6960 25894
rect 7300 25242 7328 27288
rect 7380 27270 7432 27276
rect 7472 27328 7524 27334
rect 7472 27270 7524 27276
rect 7208 25226 7328 25242
rect 7392 25226 7420 27270
rect 7484 27033 7512 27270
rect 7564 27056 7616 27062
rect 7470 27024 7526 27033
rect 7564 26998 7616 27004
rect 7470 26959 7526 26968
rect 7576 26897 7604 26998
rect 7562 26888 7618 26897
rect 7562 26823 7618 26832
rect 7576 25922 7604 26823
rect 7668 26042 7696 30194
rect 7760 29628 7788 30534
rect 7944 30054 7972 30534
rect 8036 30394 8064 33050
rect 8128 32298 8156 33390
rect 8298 33351 8354 33360
rect 8208 33312 8260 33318
rect 8312 33300 8340 33351
rect 8260 33272 8340 33300
rect 8208 33254 8260 33260
rect 8208 32768 8260 32774
rect 8208 32710 8260 32716
rect 8116 32292 8168 32298
rect 8116 32234 8168 32240
rect 8116 30592 8168 30598
rect 8116 30534 8168 30540
rect 8024 30388 8076 30394
rect 8024 30330 8076 30336
rect 8128 30190 8156 30534
rect 8220 30326 8248 32710
rect 8208 30320 8260 30326
rect 8208 30262 8260 30268
rect 8116 30184 8168 30190
rect 8116 30126 8168 30132
rect 7932 30048 7984 30054
rect 7932 29990 7984 29996
rect 7838 29880 7894 29889
rect 8114 29880 8170 29889
rect 7894 29838 7972 29866
rect 7838 29815 7894 29824
rect 7760 29600 7880 29628
rect 7748 29504 7800 29510
rect 7748 29446 7800 29452
rect 7760 29306 7788 29446
rect 7748 29300 7800 29306
rect 7748 29242 7800 29248
rect 7748 29028 7800 29034
rect 7748 28970 7800 28976
rect 7760 26761 7788 28970
rect 7852 27538 7880 29600
rect 7840 27532 7892 27538
rect 7840 27474 7892 27480
rect 7840 27328 7892 27334
rect 7840 27270 7892 27276
rect 7852 27062 7880 27270
rect 7840 27056 7892 27062
rect 7840 26998 7892 27004
rect 7746 26752 7802 26761
rect 7746 26687 7802 26696
rect 7852 26432 7880 26998
rect 7760 26404 7880 26432
rect 7760 26314 7788 26404
rect 7748 26308 7800 26314
rect 7748 26250 7800 26256
rect 7840 26308 7892 26314
rect 7840 26250 7892 26256
rect 7656 26036 7708 26042
rect 7656 25978 7708 25984
rect 7576 25894 7788 25922
rect 7470 25664 7526 25673
rect 7470 25599 7526 25608
rect 7484 25498 7512 25599
rect 7472 25492 7524 25498
rect 7472 25434 7524 25440
rect 7562 25256 7618 25265
rect 7196 25220 7328 25226
rect 7248 25214 7328 25220
rect 7380 25220 7432 25226
rect 7196 25162 7248 25168
rect 7562 25191 7618 25200
rect 7380 25162 7432 25168
rect 7576 25158 7604 25191
rect 6748 25112 6960 25140
rect 7288 25152 7340 25158
rect 6748 24834 6776 25112
rect 7288 25094 7340 25100
rect 7564 25152 7616 25158
rect 7564 25094 7616 25100
rect 6884 25052 7192 25061
rect 6884 25050 6890 25052
rect 6946 25050 6970 25052
rect 7026 25050 7050 25052
rect 7106 25050 7130 25052
rect 7186 25050 7192 25052
rect 6946 24998 6948 25050
rect 7128 24998 7130 25050
rect 6884 24996 6890 24998
rect 6946 24996 6970 24998
rect 7026 24996 7050 24998
rect 7106 24996 7130 24998
rect 7186 24996 7192 24998
rect 6884 24987 7192 24996
rect 7300 24954 7328 25094
rect 7288 24948 7340 24954
rect 7288 24890 7340 24896
rect 6748 24806 6960 24834
rect 6736 24608 6788 24614
rect 6736 24550 6788 24556
rect 6748 23186 6776 24550
rect 6932 24138 6960 24806
rect 6920 24132 6972 24138
rect 6920 24074 6972 24080
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 6884 23964 7192 23973
rect 6884 23962 6890 23964
rect 6946 23962 6970 23964
rect 7026 23962 7050 23964
rect 7106 23962 7130 23964
rect 7186 23962 7192 23964
rect 6946 23910 6948 23962
rect 7128 23910 7130 23962
rect 6884 23908 6890 23910
rect 6946 23908 6970 23910
rect 7026 23908 7050 23910
rect 7106 23908 7130 23910
rect 7186 23908 7192 23910
rect 6884 23899 7192 23908
rect 7562 23896 7618 23905
rect 7562 23831 7618 23840
rect 7116 23446 7420 23474
rect 6736 23180 6788 23186
rect 6736 23122 6788 23128
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 6748 21690 6776 23122
rect 7116 23118 7144 23446
rect 7196 23316 7248 23322
rect 7248 23276 7328 23304
rect 7196 23258 7248 23264
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 6884 22876 7192 22885
rect 6884 22874 6890 22876
rect 6946 22874 6970 22876
rect 7026 22874 7050 22876
rect 7106 22874 7130 22876
rect 7186 22874 7192 22876
rect 6946 22822 6948 22874
rect 7128 22822 7130 22874
rect 6884 22820 6890 22822
rect 6946 22820 6970 22822
rect 7026 22820 7050 22822
rect 7106 22820 7130 22822
rect 7186 22820 7192 22822
rect 6884 22811 7192 22820
rect 7196 22432 7248 22438
rect 7196 22374 7248 22380
rect 7208 22098 7236 22374
rect 7196 22092 7248 22098
rect 7196 22034 7248 22040
rect 7300 22030 7328 23276
rect 7392 22438 7420 23446
rect 7576 23118 7604 23831
rect 7564 23112 7616 23118
rect 7564 23054 7616 23060
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7380 22432 7432 22438
rect 7380 22374 7432 22380
rect 7380 22160 7432 22166
rect 7378 22128 7380 22137
rect 7432 22128 7434 22137
rect 7378 22063 7434 22072
rect 7484 22030 7512 22918
rect 7576 22234 7604 22918
rect 7564 22228 7616 22234
rect 7564 22170 7616 22176
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7472 22024 7524 22030
rect 7472 21966 7524 21972
rect 6884 21788 7192 21797
rect 6884 21786 6890 21788
rect 6946 21786 6970 21788
rect 7026 21786 7050 21788
rect 7106 21786 7130 21788
rect 7186 21786 7192 21788
rect 6946 21734 6948 21786
rect 7128 21734 7130 21786
rect 6884 21732 6890 21734
rect 6946 21732 6970 21734
rect 7026 21732 7050 21734
rect 7106 21732 7130 21734
rect 7186 21732 7192 21734
rect 6884 21723 7192 21732
rect 6736 21684 6788 21690
rect 6736 21626 6788 21632
rect 6644 21480 6696 21486
rect 6748 21468 6776 21626
rect 7668 21622 7696 24074
rect 7656 21616 7708 21622
rect 7656 21558 7708 21564
rect 7760 21554 7788 25894
rect 7852 25702 7880 26250
rect 7840 25696 7892 25702
rect 7840 25638 7892 25644
rect 7852 23769 7880 25638
rect 7838 23760 7894 23769
rect 7838 23695 7894 23704
rect 7852 23662 7880 23695
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7838 23352 7894 23361
rect 7838 23287 7894 23296
rect 7852 22642 7880 23287
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7748 21548 7800 21554
rect 7748 21490 7800 21496
rect 6696 21440 6776 21468
rect 6644 21422 6696 21428
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6656 19514 6684 20402
rect 6748 20398 6776 21440
rect 7194 21448 7250 21457
rect 7378 21448 7434 21457
rect 7194 21383 7250 21392
rect 7300 21406 7378 21434
rect 7208 20788 7236 21383
rect 7300 21078 7328 21406
rect 7378 21383 7434 21392
rect 7576 21321 7604 21490
rect 7656 21344 7708 21350
rect 7562 21312 7618 21321
rect 7656 21286 7708 21292
rect 7562 21247 7618 21256
rect 7380 21140 7432 21146
rect 7432 21100 7512 21128
rect 7380 21082 7432 21088
rect 7288 21072 7340 21078
rect 7288 21014 7340 21020
rect 7484 20942 7512 21100
rect 7576 20942 7604 21247
rect 7668 21010 7696 21286
rect 7656 21004 7708 21010
rect 7656 20946 7708 20952
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7300 20788 7328 20878
rect 7748 20868 7800 20874
rect 7748 20810 7800 20816
rect 7208 20760 7328 20788
rect 6884 20700 7192 20709
rect 6884 20698 6890 20700
rect 6946 20698 6970 20700
rect 7026 20698 7050 20700
rect 7106 20698 7130 20700
rect 7186 20698 7192 20700
rect 6946 20646 6948 20698
rect 7128 20646 7130 20698
rect 6884 20644 6890 20646
rect 6946 20644 6970 20646
rect 7026 20644 7050 20646
rect 7106 20644 7130 20646
rect 7186 20644 7192 20646
rect 6884 20635 7192 20644
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6884 19612 7192 19621
rect 6884 19610 6890 19612
rect 6946 19610 6970 19612
rect 7026 19610 7050 19612
rect 7106 19610 7130 19612
rect 7186 19610 7192 19612
rect 6946 19558 6948 19610
rect 7128 19558 7130 19610
rect 6884 19556 6890 19558
rect 6946 19556 6970 19558
rect 7026 19556 7050 19558
rect 7106 19556 7130 19558
rect 7186 19556 7192 19558
rect 6884 19547 7192 19556
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 7194 19408 7250 19417
rect 7194 19343 7250 19352
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6656 18358 6684 18906
rect 7208 18873 7236 19343
rect 7194 18864 7250 18873
rect 7194 18799 7250 18808
rect 7300 18766 7328 20760
rect 7760 20602 7788 20810
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7288 18760 7340 18766
rect 6734 18728 6790 18737
rect 7288 18702 7340 18708
rect 6734 18663 6790 18672
rect 6748 18426 6776 18663
rect 6884 18524 7192 18533
rect 6884 18522 6890 18524
rect 6946 18522 6970 18524
rect 7026 18522 7050 18524
rect 7106 18522 7130 18524
rect 7186 18522 7192 18524
rect 6946 18470 6948 18522
rect 7128 18470 7130 18522
rect 6884 18468 6890 18470
rect 6946 18468 6970 18470
rect 7026 18468 7050 18470
rect 7106 18468 7130 18470
rect 7186 18468 7192 18470
rect 6884 18459 7192 18468
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6644 18352 6696 18358
rect 6472 18278 6592 18306
rect 6644 18294 6696 18300
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6104 17190 6224 17218
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 5368 15014 5672 15042
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5552 14278 5580 14418
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5446 13968 5502 13977
rect 5446 13903 5502 13912
rect 5172 12436 5224 12442
rect 5460 12434 5488 13903
rect 5538 12744 5594 12753
rect 5538 12679 5594 12688
rect 5552 12442 5580 12679
rect 5172 12378 5224 12384
rect 5276 12406 5488 12434
rect 5540 12436 5592 12442
rect 5170 12336 5226 12345
rect 5170 12271 5172 12280
rect 5224 12271 5226 12280
rect 5172 12242 5224 12248
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5092 11778 5120 12174
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5184 11898 5212 12038
rect 5276 11898 5304 12406
rect 5540 12378 5592 12384
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5092 11750 5304 11778
rect 5080 11620 5132 11626
rect 5132 11580 5212 11608
rect 5080 11562 5132 11568
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 5000 10810 5028 10950
rect 5092 10810 5120 11086
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5184 10690 5212 11580
rect 5092 10662 5212 10690
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5000 8634 5028 8910
rect 5092 8838 5120 10662
rect 5170 9616 5226 9625
rect 5170 9551 5172 9560
rect 5224 9551 5226 9560
rect 5172 9522 5224 9528
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5276 8634 5304 11750
rect 5368 9586 5396 12310
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5460 9926 5488 11698
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5552 10810 5580 11630
rect 5644 11218 5672 15014
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5552 10266 5580 10474
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5460 8378 5488 9862
rect 5644 9636 5672 11018
rect 5736 10146 5764 15150
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5828 14618 5856 14758
rect 5920 14618 5948 15438
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5920 12442 5948 12582
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 5908 12232 5960 12238
rect 5906 12200 5908 12209
rect 5960 12200 5962 12209
rect 5906 12135 5962 12144
rect 6012 11898 6040 12378
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5828 10674 5856 11290
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5920 10266 5948 10746
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5736 10118 5948 10146
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5552 9625 5672 9636
rect 5538 9616 5672 9625
rect 5594 9608 5672 9616
rect 5736 9568 5764 9658
rect 5538 9551 5594 9560
rect 5644 9540 5764 9568
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5552 8634 5580 8842
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5276 8350 5488 8378
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4908 5914 4936 6258
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4618 4040 4674 4049
rect 4540 3738 4568 4014
rect 4618 3975 4674 3984
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4356 2961 4384 3062
rect 4342 2952 4398 2961
rect 4342 2887 4398 2896
rect 4448 2774 4476 3062
rect 4632 2990 4660 3975
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4802 2816 4858 2825
rect 4448 2760 4802 2774
rect 4448 2751 4858 2760
rect 4448 2746 4844 2751
rect 4448 2650 4476 2746
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4908 2530 4936 2926
rect 5000 2650 5028 6802
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 4908 2502 5028 2530
rect 4620 2440 4672 2446
rect 4434 2408 4490 2417
rect 4620 2382 4672 2388
rect 4712 2440 4764 2446
rect 4764 2400 4936 2428
rect 4712 2382 4764 2388
rect 4434 2343 4490 2352
rect 4528 2372 4580 2378
rect 4448 2106 4476 2343
rect 4528 2314 4580 2320
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 4252 2100 4304 2106
rect 4252 2042 4304 2048
rect 4436 2100 4488 2106
rect 4436 2042 4488 2048
rect 4068 1896 4120 1902
rect 4120 1856 4292 1884
rect 4068 1838 4120 1844
rect 3917 1660 4225 1669
rect 3917 1658 3923 1660
rect 3979 1658 4003 1660
rect 4059 1658 4083 1660
rect 4139 1658 4163 1660
rect 4219 1658 4225 1660
rect 3979 1606 3981 1658
rect 4161 1606 4163 1658
rect 3917 1604 3923 1606
rect 3979 1604 4003 1606
rect 4059 1604 4083 1606
rect 4139 1604 4163 1606
rect 4219 1604 4225 1606
rect 3917 1595 4225 1604
rect 3792 1352 3844 1358
rect 3792 1294 3844 1300
rect 3884 1216 3936 1222
rect 3884 1158 3936 1164
rect 4068 1216 4120 1222
rect 4068 1158 4120 1164
rect 3896 950 3924 1158
rect 3884 944 3936 950
rect 3884 886 3936 892
rect 4080 160 4108 1158
rect 3790 82 3846 160
rect 3712 54 3846 82
rect 3790 0 3846 54
rect 4066 0 4122 160
rect 4264 82 4292 1856
rect 4434 1728 4490 1737
rect 4434 1663 4490 1672
rect 4448 1562 4476 1663
rect 4540 1562 4568 2314
rect 4436 1556 4488 1562
rect 4436 1498 4488 1504
rect 4528 1556 4580 1562
rect 4528 1498 4580 1504
rect 4436 1352 4488 1358
rect 4434 1320 4436 1329
rect 4488 1320 4490 1329
rect 4434 1255 4490 1264
rect 4632 160 4660 2382
rect 4804 1760 4856 1766
rect 4804 1702 4856 1708
rect 4816 1601 4844 1702
rect 4802 1592 4858 1601
rect 4802 1527 4858 1536
rect 4908 160 4936 2400
rect 5000 1952 5028 2502
rect 5092 2106 5120 7142
rect 5184 5574 5212 8298
rect 5276 6225 5304 8350
rect 5552 7886 5580 8570
rect 5644 7886 5672 9540
rect 5828 9450 5856 9930
rect 5920 9586 5948 10118
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5736 8634 5764 9318
rect 5906 9208 5962 9217
rect 5906 9143 5962 9152
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5262 6216 5318 6225
rect 5262 6151 5318 6160
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5184 4282 5212 4558
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5276 3942 5304 6151
rect 5368 5710 5396 6394
rect 5446 6352 5502 6361
rect 5446 6287 5502 6296
rect 5460 6254 5488 6287
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5552 5710 5580 7822
rect 5644 5846 5672 7822
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5184 2650 5212 3674
rect 5552 3369 5580 3946
rect 5920 3738 5948 9143
rect 6012 7954 6040 11154
rect 6104 9654 6132 17190
rect 6288 15994 6316 17274
rect 6196 15966 6316 15994
rect 6196 9976 6224 15966
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6288 10826 6316 15370
rect 6380 11150 6408 18022
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6288 10798 6408 10826
rect 6276 9988 6328 9994
rect 6196 9948 6276 9976
rect 6276 9930 6328 9936
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 6104 8362 6132 9590
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6196 7954 6224 8842
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6012 7410 6040 7890
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6104 6934 6132 7278
rect 6196 7274 6224 7890
rect 6184 7268 6236 7274
rect 6184 7210 6236 7216
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6196 6118 6224 7210
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6104 5914 6132 6054
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6196 5370 6224 5714
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6288 5234 6316 9930
rect 6380 6866 6408 10798
rect 6472 8922 6500 17614
rect 6564 17338 6592 18278
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 7288 18284 7340 18290
rect 7392 18272 7420 20538
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7484 18358 7512 20402
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 7576 19514 7604 19994
rect 7656 19780 7708 19786
rect 7656 19722 7708 19728
rect 7668 19514 7696 19722
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7760 18766 7788 19450
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7656 18760 7708 18766
rect 7656 18702 7708 18708
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7472 18352 7524 18358
rect 7472 18294 7524 18300
rect 7340 18244 7420 18272
rect 7288 18226 7340 18232
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6748 17882 6776 18158
rect 6932 17882 6960 18226
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6884 17436 7192 17445
rect 6884 17434 6890 17436
rect 6946 17434 6970 17436
rect 7026 17434 7050 17436
rect 7106 17434 7130 17436
rect 7186 17434 7192 17436
rect 6946 17382 6948 17434
rect 7128 17382 7130 17434
rect 6884 17380 6890 17382
rect 6946 17380 6970 17382
rect 7026 17380 7050 17382
rect 7106 17380 7130 17382
rect 7186 17380 7192 17382
rect 6884 17371 7192 17380
rect 6552 17332 6604 17338
rect 7576 17320 7604 18702
rect 7668 17746 7696 18702
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 7760 17338 7788 18158
rect 7748 17332 7800 17338
rect 7576 17292 7696 17320
rect 6552 17274 6604 17280
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 6748 16250 6776 17138
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7208 16658 7236 17070
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 6884 16348 7192 16357
rect 6884 16346 6890 16348
rect 6946 16346 6970 16348
rect 7026 16346 7050 16348
rect 7106 16346 7130 16348
rect 7186 16346 7192 16348
rect 6946 16294 6948 16346
rect 7128 16294 7130 16346
rect 6884 16292 6890 16294
rect 6946 16292 6970 16294
rect 7026 16292 7050 16294
rect 7106 16292 7130 16294
rect 7186 16292 7192 16294
rect 6884 16283 7192 16292
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6564 13734 6592 16050
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6826 15600 6882 15609
rect 6932 15570 6960 15914
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 6826 15535 6828 15544
rect 6880 15535 6882 15544
rect 6920 15564 6972 15570
rect 6828 15506 6880 15512
rect 6920 15506 6972 15512
rect 6644 15360 6696 15366
rect 6642 15328 6644 15337
rect 6932 15348 6960 15506
rect 7208 15502 7236 15846
rect 7196 15496 7248 15502
rect 7380 15496 7432 15502
rect 7196 15438 7248 15444
rect 7300 15444 7380 15450
rect 7300 15438 7432 15444
rect 6696 15328 6698 15337
rect 6642 15263 6698 15272
rect 6748 15320 6960 15348
rect 7300 15422 7420 15438
rect 6748 15042 6776 15320
rect 6884 15260 7192 15269
rect 6884 15258 6890 15260
rect 6946 15258 6970 15260
rect 7026 15258 7050 15260
rect 7106 15258 7130 15260
rect 7186 15258 7192 15260
rect 6946 15206 6948 15258
rect 7128 15206 7130 15258
rect 6884 15204 6890 15206
rect 6946 15204 6970 15206
rect 7026 15204 7050 15206
rect 7106 15204 7130 15206
rect 7186 15204 7192 15206
rect 6884 15195 7192 15204
rect 6748 15014 6868 15042
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6656 13938 6684 14418
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6564 12918 6592 13670
rect 6656 13394 6684 13874
rect 6748 13734 6776 14894
rect 6840 14482 6868 15014
rect 7300 14958 7328 15422
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7392 14958 7420 15302
rect 7484 14958 7512 15982
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7576 14804 7604 17138
rect 7668 16232 7696 17292
rect 7748 17274 7800 17280
rect 7760 17134 7788 17274
rect 7852 17202 7880 20198
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7944 16454 7972 29838
rect 8114 29815 8170 29824
rect 8024 28756 8076 28762
rect 8024 28698 8076 28704
rect 8036 28422 8064 28698
rect 8024 28416 8076 28422
rect 8024 28358 8076 28364
rect 8024 27464 8076 27470
rect 8024 27406 8076 27412
rect 8036 26382 8064 27406
rect 8024 26376 8076 26382
rect 8024 26318 8076 26324
rect 8128 26217 8156 29815
rect 8208 29776 8260 29782
rect 8208 29718 8260 29724
rect 8220 28642 8248 29718
rect 8312 28966 8340 33272
rect 8404 29034 8432 34598
rect 8392 29028 8444 29034
rect 8392 28970 8444 28976
rect 8300 28960 8352 28966
rect 8300 28902 8352 28908
rect 8220 28614 8432 28642
rect 8208 28552 8260 28558
rect 8208 28494 8260 28500
rect 8220 28082 8248 28494
rect 8208 28076 8260 28082
rect 8208 28018 8260 28024
rect 8220 27713 8248 28018
rect 8300 27872 8352 27878
rect 8300 27814 8352 27820
rect 8206 27704 8262 27713
rect 8206 27639 8262 27648
rect 8208 27532 8260 27538
rect 8208 27474 8260 27480
rect 8114 26208 8170 26217
rect 8114 26143 8170 26152
rect 8116 26036 8168 26042
rect 8116 25978 8168 25984
rect 8024 25696 8076 25702
rect 8024 25638 8076 25644
rect 8036 24750 8064 25638
rect 8024 24744 8076 24750
rect 8024 24686 8076 24692
rect 8024 23656 8076 23662
rect 8024 23598 8076 23604
rect 8036 20058 8064 23598
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 8024 19780 8076 19786
rect 8024 19722 8076 19728
rect 7932 16448 7984 16454
rect 7932 16390 7984 16396
rect 7668 16204 7880 16232
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7668 15162 7696 15846
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7300 14776 7604 14804
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6884 14172 7192 14181
rect 6884 14170 6890 14172
rect 6946 14170 6970 14172
rect 7026 14170 7050 14172
rect 7106 14170 7130 14172
rect 7186 14170 7192 14172
rect 6946 14118 6948 14170
rect 7128 14118 7130 14170
rect 6884 14116 6890 14118
rect 6946 14116 6970 14118
rect 7026 14116 7050 14118
rect 7106 14116 7130 14118
rect 7186 14116 7192 14118
rect 6884 14107 7192 14116
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6564 11898 6592 12854
rect 6656 12646 6684 13330
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6644 12368 6696 12374
rect 6642 12336 6644 12345
rect 6696 12336 6698 12345
rect 6642 12271 6698 12280
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6656 11218 6684 12271
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6564 10606 6592 11018
rect 6748 10674 6776 13670
rect 6884 13084 7192 13093
rect 6884 13082 6890 13084
rect 6946 13082 6970 13084
rect 7026 13082 7050 13084
rect 7106 13082 7130 13084
rect 7186 13082 7192 13084
rect 6946 13030 6948 13082
rect 7128 13030 7130 13082
rect 6884 13028 6890 13030
rect 6946 13028 6970 13030
rect 7026 13028 7050 13030
rect 7106 13028 7130 13030
rect 7186 13028 7192 13030
rect 6884 13019 7192 13028
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7116 12434 7144 12582
rect 7024 12406 7144 12434
rect 7024 12306 7052 12406
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6884 11996 7192 12005
rect 6884 11994 6890 11996
rect 6946 11994 6970 11996
rect 7026 11994 7050 11996
rect 7106 11994 7130 11996
rect 7186 11994 7192 11996
rect 6946 11942 6948 11994
rect 7128 11942 7130 11994
rect 6884 11940 6890 11942
rect 6946 11940 6970 11942
rect 7026 11940 7050 11942
rect 7106 11940 7130 11942
rect 7186 11940 7192 11942
rect 6884 11931 7192 11940
rect 6884 10908 7192 10917
rect 6884 10906 6890 10908
rect 6946 10906 6970 10908
rect 7026 10906 7050 10908
rect 7106 10906 7130 10908
rect 7186 10906 7192 10908
rect 6946 10854 6948 10906
rect 7128 10854 7130 10906
rect 6884 10852 6890 10854
rect 6946 10852 6970 10854
rect 7026 10852 7050 10854
rect 7106 10852 7130 10854
rect 7186 10852 7192 10854
rect 6884 10843 7192 10852
rect 7300 10792 7328 14776
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 7392 13326 7420 13942
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7378 12880 7434 12889
rect 7378 12815 7434 12824
rect 7392 11830 7420 12815
rect 7470 12744 7526 12753
rect 7470 12679 7526 12688
rect 7484 12306 7512 12679
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7576 11898 7604 12310
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7380 11280 7432 11286
rect 7668 11234 7696 15098
rect 7760 15026 7788 16050
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7852 14346 7880 16204
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7944 15434 7972 15846
rect 7932 15428 7984 15434
rect 7932 15370 7984 15376
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7944 14618 7972 14894
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7746 13696 7802 13705
rect 7746 13631 7802 13640
rect 7380 11222 7432 11228
rect 7116 10764 7328 10792
rect 6826 10704 6882 10713
rect 6736 10668 6788 10674
rect 6826 10639 6882 10648
rect 6736 10610 6788 10616
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6564 9722 6592 10542
rect 6840 10266 6868 10639
rect 7116 10452 7144 10764
rect 7288 10600 7340 10606
rect 7208 10577 7288 10588
rect 7194 10568 7288 10577
rect 7250 10560 7288 10568
rect 7288 10542 7340 10548
rect 7194 10503 7250 10512
rect 7116 10424 7328 10452
rect 6918 10296 6974 10305
rect 6828 10260 6880 10266
rect 6918 10231 6920 10240
rect 6828 10202 6880 10208
rect 6972 10231 6974 10240
rect 6920 10202 6972 10208
rect 6884 9820 7192 9829
rect 6884 9818 6890 9820
rect 6946 9818 6970 9820
rect 7026 9818 7050 9820
rect 7106 9818 7130 9820
rect 7186 9818 7192 9820
rect 6946 9766 6948 9818
rect 7128 9766 7130 9818
rect 6884 9764 6890 9766
rect 6946 9764 6970 9766
rect 7026 9764 7050 9766
rect 7106 9764 7130 9766
rect 7186 9764 7192 9766
rect 6884 9755 7192 9764
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6472 8894 6592 8922
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6472 7954 6500 8774
rect 6564 8498 6592 8894
rect 6748 8634 6776 9386
rect 7208 9178 7236 9454
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 6918 9072 6974 9081
rect 6918 9007 6920 9016
rect 6972 9007 6974 9016
rect 6920 8978 6972 8984
rect 6884 8732 7192 8741
rect 6884 8730 6890 8732
rect 6946 8730 6970 8732
rect 7026 8730 7050 8732
rect 7106 8730 7130 8732
rect 7186 8730 7192 8732
rect 6946 8678 6948 8730
rect 7128 8678 7130 8730
rect 6884 8676 6890 8678
rect 6946 8676 6970 8678
rect 7026 8676 7050 8678
rect 7106 8676 7130 8678
rect 7186 8676 7192 8678
rect 6884 8667 7192 8676
rect 7300 8634 7328 10424
rect 7392 9217 7420 11222
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7576 11206 7696 11234
rect 7378 9208 7434 9217
rect 7378 9143 7434 9152
rect 7362 9104 7414 9110
rect 7414 9052 7420 9092
rect 7484 9081 7512 11154
rect 7576 11082 7604 11206
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 10305 7604 10610
rect 7668 10577 7696 11086
rect 7654 10568 7710 10577
rect 7654 10503 7710 10512
rect 7562 10296 7618 10305
rect 7562 10231 7618 10240
rect 7362 9046 7420 9052
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6564 8401 6592 8434
rect 6644 8424 6696 8430
rect 6550 8392 6606 8401
rect 6644 8366 6696 8372
rect 6550 8327 6606 8336
rect 6460 7948 6512 7954
rect 6512 7908 6592 7936
rect 6460 7890 6512 7896
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5658 6408 6054
rect 6564 5778 6592 7908
rect 6656 6934 6684 8366
rect 6748 7392 6776 8570
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6840 8090 6868 8230
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 7208 7818 7236 8570
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 6884 7644 7192 7653
rect 6884 7642 6890 7644
rect 6946 7642 6970 7644
rect 7026 7642 7050 7644
rect 7106 7642 7130 7644
rect 7186 7642 7192 7644
rect 6946 7590 6948 7642
rect 7128 7590 7130 7642
rect 6884 7588 6890 7590
rect 6946 7588 6970 7590
rect 7026 7588 7050 7590
rect 7106 7588 7130 7590
rect 7186 7588 7192 7590
rect 6884 7579 7192 7588
rect 7300 7546 7328 7958
rect 7392 7546 7420 9046
rect 7470 9072 7526 9081
rect 7668 9042 7696 10503
rect 7470 9007 7526 9016
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 7857 7512 8774
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7576 7886 7604 8570
rect 7656 8560 7708 8566
rect 7654 8528 7656 8537
rect 7708 8528 7710 8537
rect 7654 8463 7710 8472
rect 7564 7880 7616 7886
rect 7470 7848 7526 7857
rect 7564 7822 7616 7828
rect 7470 7783 7526 7792
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 6828 7404 6880 7410
rect 6748 7364 6828 7392
rect 6828 7346 6880 7352
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6734 6896 6790 6905
rect 6734 6831 6790 6840
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6656 6118 6684 6734
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6460 5704 6512 5710
rect 6380 5652 6460 5658
rect 6380 5646 6512 5652
rect 6380 5630 6500 5646
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5538 3360 5594 3369
rect 5538 3295 5594 3304
rect 6656 3176 6684 3878
rect 6748 3534 6776 6831
rect 6884 6556 7192 6565
rect 6884 6554 6890 6556
rect 6946 6554 6970 6556
rect 7026 6554 7050 6556
rect 7106 6554 7130 6556
rect 7186 6554 7192 6556
rect 6946 6502 6948 6554
rect 7128 6502 7130 6554
rect 6884 6500 6890 6502
rect 6946 6500 6970 6502
rect 7026 6500 7050 6502
rect 7106 6500 7130 6502
rect 7186 6500 7192 6502
rect 6884 6491 7192 6500
rect 6884 5468 7192 5477
rect 6884 5466 6890 5468
rect 6946 5466 6970 5468
rect 7026 5466 7050 5468
rect 7106 5466 7130 5468
rect 7186 5466 7192 5468
rect 6946 5414 6948 5466
rect 7128 5414 7130 5466
rect 6884 5412 6890 5414
rect 6946 5412 6970 5414
rect 7026 5412 7050 5414
rect 7106 5412 7130 5414
rect 7186 5412 7192 5414
rect 6884 5403 7192 5412
rect 7300 5234 7328 7346
rect 7380 6792 7432 6798
rect 7564 6792 7616 6798
rect 7432 6740 7512 6746
rect 7380 6734 7512 6740
rect 7564 6734 7616 6740
rect 7392 6718 7512 6734
rect 7484 6662 7512 6718
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7392 5914 7420 6598
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7392 5370 7420 5714
rect 7576 5642 7604 6734
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7300 4622 7328 5170
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 4690 7420 4966
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 6884 4380 7192 4389
rect 6884 4378 6890 4380
rect 6946 4378 6970 4380
rect 7026 4378 7050 4380
rect 7106 4378 7130 4380
rect 7186 4378 7192 4380
rect 6946 4326 6948 4378
rect 7128 4326 7130 4378
rect 6884 4324 6890 4326
rect 6946 4324 6970 4326
rect 7026 4324 7050 4326
rect 7106 4324 7130 4326
rect 7186 4324 7192 4326
rect 6884 4315 7192 4324
rect 7300 3602 7328 4558
rect 7484 4486 7512 5306
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6884 3292 7192 3301
rect 6884 3290 6890 3292
rect 6946 3290 6970 3292
rect 7026 3290 7050 3292
rect 7106 3290 7130 3292
rect 7186 3290 7192 3292
rect 6946 3238 6948 3290
rect 7128 3238 7130 3290
rect 6884 3236 6890 3238
rect 6946 3236 6970 3238
rect 7026 3236 7050 3238
rect 7106 3236 7130 3238
rect 7186 3236 7192 3238
rect 6884 3227 7192 3236
rect 7300 3176 7328 3538
rect 6656 3148 6868 3176
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5906 2816 5962 2825
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5368 2514 5396 2790
rect 5906 2751 5962 2760
rect 5722 2544 5778 2553
rect 5356 2508 5408 2514
rect 5722 2479 5778 2488
rect 5356 2450 5408 2456
rect 5736 2446 5764 2479
rect 5920 2446 5948 2751
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 5080 2100 5132 2106
rect 5080 2042 5132 2048
rect 5172 2100 5224 2106
rect 5172 2042 5224 2048
rect 5080 1964 5132 1970
rect 5000 1924 5080 1952
rect 5184 1952 5212 2042
rect 5132 1924 5212 1952
rect 5080 1906 5132 1912
rect 5080 1216 5132 1222
rect 5080 1158 5132 1164
rect 5092 1018 5120 1158
rect 5080 1012 5132 1018
rect 5080 954 5132 960
rect 4342 82 4398 160
rect 4264 54 4398 82
rect 4342 0 4398 54
rect 4618 0 4674 160
rect 4894 0 4950 160
rect 5170 82 5226 160
rect 5276 82 5304 2314
rect 5540 2304 5592 2310
rect 5592 2264 5764 2292
rect 5540 2246 5592 2252
rect 5632 2032 5684 2038
rect 5538 2000 5594 2009
rect 5632 1974 5684 1980
rect 5538 1935 5594 1944
rect 5356 1760 5408 1766
rect 5408 1720 5488 1748
rect 5356 1702 5408 1708
rect 5460 160 5488 1720
rect 5552 1222 5580 1935
rect 5540 1216 5592 1222
rect 5540 1158 5592 1164
rect 5644 1034 5672 1974
rect 5736 1902 5764 2264
rect 5828 2106 5856 2314
rect 5816 2100 5868 2106
rect 5816 2042 5868 2048
rect 6000 2100 6052 2106
rect 6000 2042 6052 2048
rect 6012 2009 6040 2042
rect 5998 2000 6054 2009
rect 5998 1935 6054 1944
rect 5724 1896 5776 1902
rect 5724 1838 5776 1844
rect 5816 1352 5868 1358
rect 5816 1294 5868 1300
rect 5644 1006 5764 1034
rect 5736 160 5764 1006
rect 5828 542 5856 1294
rect 6000 1284 6052 1290
rect 6000 1226 6052 1232
rect 5816 536 5868 542
rect 5816 478 5868 484
rect 6012 160 6040 1226
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 6104 785 6132 1158
rect 6090 776 6146 785
rect 6196 746 6224 3062
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 6380 1970 6408 2246
rect 6368 1964 6420 1970
rect 6368 1906 6420 1912
rect 6472 1426 6500 2790
rect 6564 2038 6592 2858
rect 6552 2032 6604 2038
rect 6552 1974 6604 1980
rect 6460 1420 6512 1426
rect 6460 1362 6512 1368
rect 6276 1352 6328 1358
rect 6276 1294 6328 1300
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 6090 711 6146 720
rect 6184 740 6236 746
rect 6184 682 6236 688
rect 6288 160 6316 1294
rect 6380 610 6408 1294
rect 6460 1216 6512 1222
rect 6460 1158 6512 1164
rect 6552 1216 6604 1222
rect 6552 1158 6604 1164
rect 6472 882 6500 1158
rect 6460 876 6512 882
rect 6460 818 6512 824
rect 6368 604 6420 610
rect 6368 546 6420 552
rect 6564 160 6592 1158
rect 5170 54 5304 82
rect 5170 0 5226 54
rect 5446 0 5502 160
rect 5722 0 5778 160
rect 5998 0 6054 160
rect 6274 0 6330 160
rect 6550 0 6606 160
rect 6656 82 6684 2994
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6748 1358 6776 2790
rect 6840 2650 6868 3148
rect 7116 3148 7328 3176
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 7116 2446 7144 3148
rect 7196 3052 7248 3058
rect 7248 3012 7420 3040
rect 7196 2994 7248 3000
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 6884 2204 7192 2213
rect 6884 2202 6890 2204
rect 6946 2202 6970 2204
rect 7026 2202 7050 2204
rect 7106 2202 7130 2204
rect 7186 2202 7192 2204
rect 6946 2150 6948 2202
rect 7128 2150 7130 2202
rect 6884 2148 6890 2150
rect 6946 2148 6970 2150
rect 7026 2148 7050 2150
rect 7106 2148 7130 2150
rect 7186 2148 7192 2150
rect 6884 2139 7192 2148
rect 7012 2100 7064 2106
rect 7012 2042 7064 2048
rect 7024 2009 7052 2042
rect 7300 2038 7328 2790
rect 7288 2032 7340 2038
rect 7010 2000 7066 2009
rect 7288 1974 7340 1980
rect 7010 1935 7066 1944
rect 6918 1592 6974 1601
rect 6918 1527 6974 1536
rect 6932 1426 6960 1527
rect 6920 1420 6972 1426
rect 6920 1362 6972 1368
rect 6736 1352 6788 1358
rect 6736 1294 6788 1300
rect 6918 1320 6974 1329
rect 6918 1255 6974 1264
rect 6932 1222 6960 1255
rect 6736 1216 6788 1222
rect 6736 1158 6788 1164
rect 6920 1216 6972 1222
rect 6920 1158 6972 1164
rect 6748 406 6776 1158
rect 6884 1116 7192 1125
rect 6884 1114 6890 1116
rect 6946 1114 6970 1116
rect 7026 1114 7050 1116
rect 7106 1114 7130 1116
rect 7186 1114 7192 1116
rect 6946 1062 6948 1114
rect 7128 1062 7130 1114
rect 6884 1060 6890 1062
rect 6946 1060 6970 1062
rect 7026 1060 7050 1062
rect 7106 1060 7130 1062
rect 7186 1060 7192 1062
rect 6884 1051 7192 1060
rect 7104 740 7156 746
rect 7104 682 7156 688
rect 6736 400 6788 406
rect 6736 342 6788 348
rect 7116 160 7144 682
rect 7392 160 7420 3012
rect 7576 2446 7604 5578
rect 7668 4049 7696 7482
rect 7654 4040 7710 4049
rect 7654 3975 7710 3984
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7472 1964 7524 1970
rect 7472 1906 7524 1912
rect 7484 950 7512 1906
rect 7564 1216 7616 1222
rect 7564 1158 7616 1164
rect 7472 944 7524 950
rect 7472 886 7524 892
rect 7576 746 7604 1158
rect 7564 740 7616 746
rect 7564 682 7616 688
rect 7668 160 7696 2926
rect 7760 2774 7788 13631
rect 7852 12238 7880 14282
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7944 9194 7972 13194
rect 8036 11778 8064 19722
rect 8128 17354 8156 25978
rect 8220 24818 8248 27474
rect 8312 27062 8340 27814
rect 8404 27334 8432 28614
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8300 27056 8352 27062
rect 8300 26998 8352 27004
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 8312 26586 8340 26862
rect 8300 26580 8352 26586
rect 8300 26522 8352 26528
rect 8298 25392 8354 25401
rect 8298 25327 8354 25336
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 8312 23050 8340 25327
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8404 23866 8432 24754
rect 8392 23860 8444 23866
rect 8392 23802 8444 23808
rect 8300 23044 8352 23050
rect 8300 22986 8352 22992
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 8300 22636 8352 22642
rect 8300 22578 8352 22584
rect 8312 22094 8340 22578
rect 8404 22574 8432 22918
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 8312 22066 8432 22094
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 8220 21690 8248 21898
rect 8404 21690 8432 22066
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8390 21584 8446 21593
rect 8390 21519 8392 21528
rect 8444 21519 8446 21528
rect 8392 21490 8444 21496
rect 8206 20904 8262 20913
rect 8390 20904 8446 20913
rect 8206 20839 8262 20848
rect 8300 20868 8352 20874
rect 8220 18766 8248 20839
rect 8390 20839 8446 20848
rect 8300 20810 8352 20816
rect 8312 19009 8340 20810
rect 8298 19000 8354 19009
rect 8298 18935 8354 18944
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8128 17326 8248 17354
rect 8220 16046 8248 17326
rect 8404 16794 8432 20839
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8312 16046 8340 16662
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8128 15706 8156 15846
rect 8116 15700 8168 15706
rect 8116 15642 8168 15648
rect 8404 14634 8432 16390
rect 8312 14606 8432 14634
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8128 11898 8156 12174
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8036 11750 8156 11778
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 7852 9166 7972 9194
rect 7852 7460 7880 9166
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7944 8634 7972 8910
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7944 8401 7972 8434
rect 7930 8392 7986 8401
rect 7930 8327 7986 8336
rect 7932 7472 7984 7478
rect 7852 7432 7932 7460
rect 7932 7414 7984 7420
rect 8036 6866 8064 11086
rect 8128 10606 8156 11750
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8220 9058 8248 12038
rect 8312 11286 8340 14606
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8404 13938 8432 14486
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8128 9042 8248 9058
rect 8116 9036 8248 9042
rect 8168 9030 8248 9036
rect 8116 8978 8168 8984
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 8036 6662 8064 6802
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8220 6322 8248 6598
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7852 5914 7880 6190
rect 8312 6186 8340 9998
rect 8392 9104 8444 9110
rect 8390 9072 8392 9081
rect 8444 9072 8446 9081
rect 8496 9042 8524 35022
rect 8680 33522 8708 35226
rect 8772 34388 8800 35448
rect 8864 34513 8892 42298
rect 8956 40050 8984 42758
rect 9232 42724 9312 42752
rect 9128 42696 9180 42702
rect 9128 42638 9180 42644
rect 9036 42016 9088 42022
rect 9036 41958 9088 41964
rect 9048 40118 9076 41958
rect 9140 41818 9168 42638
rect 9128 41812 9180 41818
rect 9128 41754 9180 41760
rect 9232 41274 9260 42724
rect 9600 42758 9720 42786
rect 9772 42774 9824 42780
rect 9312 42706 9364 42712
rect 9692 42634 9720 42758
rect 10336 42702 10364 43114
rect 10416 43104 10468 43110
rect 10416 43046 10468 43052
rect 10876 43104 10928 43110
rect 10876 43046 10928 43052
rect 11244 43104 11296 43110
rect 11244 43046 11296 43052
rect 10428 42945 10456 43046
rect 10414 42936 10470 42945
rect 10414 42871 10470 42880
rect 10888 42786 10916 43046
rect 10704 42758 10916 42786
rect 10324 42696 10376 42702
rect 10324 42638 10376 42644
rect 10508 42696 10560 42702
rect 10508 42638 10560 42644
rect 9496 42628 9548 42634
rect 9496 42570 9548 42576
rect 9680 42628 9732 42634
rect 9680 42570 9732 42576
rect 9404 42288 9456 42294
rect 9324 42248 9404 42276
rect 9220 41268 9272 41274
rect 9220 41210 9272 41216
rect 9126 41168 9182 41177
rect 9324 41154 9352 42248
rect 9404 42230 9456 42236
rect 9508 41970 9536 42570
rect 9588 42560 9640 42566
rect 9588 42502 9640 42508
rect 9600 42294 9628 42502
rect 9588 42288 9640 42294
rect 9588 42230 9640 42236
rect 9772 42152 9824 42158
rect 9772 42094 9824 42100
rect 9508 41942 9628 41970
rect 9404 41472 9456 41478
rect 9402 41440 9404 41449
rect 9456 41440 9458 41449
rect 9402 41375 9458 41384
rect 9182 41126 9352 41154
rect 9600 41138 9628 41942
rect 9784 41614 9812 42094
rect 9851 41916 10159 41925
rect 9851 41914 9857 41916
rect 9913 41914 9937 41916
rect 9993 41914 10017 41916
rect 10073 41914 10097 41916
rect 10153 41914 10159 41916
rect 9913 41862 9915 41914
rect 10095 41862 10097 41914
rect 9851 41860 9857 41862
rect 9913 41860 9937 41862
rect 9993 41860 10017 41862
rect 10073 41860 10097 41862
rect 10153 41860 10159 41862
rect 9851 41851 10159 41860
rect 9772 41608 9824 41614
rect 9772 41550 9824 41556
rect 9784 41414 9812 41550
rect 10048 41540 10100 41546
rect 10048 41482 10100 41488
rect 10060 41414 10088 41482
rect 9784 41386 9904 41414
rect 10060 41386 10272 41414
rect 9772 41268 9824 41274
rect 9772 41210 9824 41216
rect 9588 41132 9640 41138
rect 9126 41103 9182 41112
rect 9588 41074 9640 41080
rect 9680 41132 9732 41138
rect 9680 41074 9732 41080
rect 9128 40928 9180 40934
rect 9128 40870 9180 40876
rect 9036 40112 9088 40118
rect 9036 40054 9088 40060
rect 8944 40044 8996 40050
rect 8944 39986 8996 39992
rect 9140 39574 9168 40870
rect 9312 40112 9364 40118
rect 9692 40089 9720 41074
rect 9784 40662 9812 41210
rect 9876 41138 9904 41386
rect 10244 41177 10272 41386
rect 10230 41168 10286 41177
rect 9864 41132 9916 41138
rect 10230 41103 10286 41112
rect 10324 41132 10376 41138
rect 9864 41074 9916 41080
rect 9851 40828 10159 40837
rect 9851 40826 9857 40828
rect 9913 40826 9937 40828
rect 9993 40826 10017 40828
rect 10073 40826 10097 40828
rect 10153 40826 10159 40828
rect 9913 40774 9915 40826
rect 10095 40774 10097 40826
rect 9851 40772 9857 40774
rect 9913 40772 9937 40774
rect 9993 40772 10017 40774
rect 10073 40772 10097 40774
rect 10153 40772 10159 40774
rect 9851 40763 10159 40772
rect 9772 40656 9824 40662
rect 9772 40598 9824 40604
rect 9772 40520 9824 40526
rect 10244 40497 10272 41103
rect 10324 41074 10376 41080
rect 10336 40730 10364 41074
rect 10324 40724 10376 40730
rect 10324 40666 10376 40672
rect 9772 40462 9824 40468
rect 10230 40488 10286 40497
rect 9312 40054 9364 40060
rect 9678 40080 9734 40089
rect 9220 40044 9272 40050
rect 9220 39986 9272 39992
rect 9128 39568 9180 39574
rect 9128 39510 9180 39516
rect 9232 38962 9260 39986
rect 9220 38956 9272 38962
rect 9220 38898 9272 38904
rect 9232 38554 9260 38898
rect 9220 38548 9272 38554
rect 9220 38490 9272 38496
rect 8944 38480 8996 38486
rect 8944 38422 8996 38428
rect 8956 35170 8984 38422
rect 9232 37874 9260 38490
rect 9324 38486 9352 40054
rect 9784 40050 9812 40462
rect 10230 40423 10286 40432
rect 10244 40089 10272 40423
rect 10336 40361 10364 40666
rect 10322 40352 10378 40361
rect 10322 40287 10378 40296
rect 10230 40080 10286 40089
rect 9678 40015 9734 40024
rect 9772 40044 9824 40050
rect 10230 40015 10286 40024
rect 9772 39986 9824 39992
rect 9402 39536 9458 39545
rect 9402 39471 9458 39480
rect 9416 39030 9444 39471
rect 9496 39432 9548 39438
rect 9496 39374 9548 39380
rect 9404 39024 9456 39030
rect 9404 38966 9456 38972
rect 9312 38480 9364 38486
rect 9312 38422 9364 38428
rect 9508 38010 9536 39374
rect 9680 38956 9732 38962
rect 9784 38944 9812 39986
rect 10232 39840 10284 39846
rect 10232 39782 10284 39788
rect 9851 39740 10159 39749
rect 9851 39738 9857 39740
rect 9913 39738 9937 39740
rect 9993 39738 10017 39740
rect 10073 39738 10097 39740
rect 10153 39738 10159 39740
rect 9913 39686 9915 39738
rect 10095 39686 10097 39738
rect 9851 39684 9857 39686
rect 9913 39684 9937 39686
rect 9993 39684 10017 39686
rect 10073 39684 10097 39686
rect 10153 39684 10159 39686
rect 9851 39675 10159 39684
rect 10244 39522 10272 39782
rect 10152 39494 10272 39522
rect 10152 39302 10180 39494
rect 10140 39296 10192 39302
rect 10140 39238 10192 39244
rect 10232 39296 10284 39302
rect 10232 39238 10284 39244
rect 10244 39098 10272 39238
rect 10232 39092 10284 39098
rect 10232 39034 10284 39040
rect 9732 38916 9812 38944
rect 10232 38956 10284 38962
rect 9680 38898 9732 38904
rect 10232 38898 10284 38904
rect 9692 38026 9720 38898
rect 9851 38652 10159 38661
rect 9851 38650 9857 38652
rect 9913 38650 9937 38652
rect 9993 38650 10017 38652
rect 10073 38650 10097 38652
rect 10153 38650 10159 38652
rect 9913 38598 9915 38650
rect 10095 38598 10097 38650
rect 9851 38596 9857 38598
rect 9913 38596 9937 38598
rect 9993 38596 10017 38598
rect 10073 38596 10097 38598
rect 10153 38596 10159 38598
rect 9851 38587 10159 38596
rect 10244 38536 10272 38898
rect 10152 38508 10272 38536
rect 10152 38350 10180 38508
rect 10140 38344 10192 38350
rect 10336 38298 10364 40287
rect 10416 39840 10468 39846
rect 10416 39782 10468 39788
rect 10140 38286 10192 38292
rect 10244 38270 10364 38298
rect 9772 38208 9824 38214
rect 9772 38150 9824 38156
rect 9496 38004 9548 38010
rect 9496 37946 9548 37952
rect 9600 37998 9720 38026
rect 9600 37942 9628 37998
rect 9784 37942 9812 38150
rect 9588 37936 9640 37942
rect 9588 37878 9640 37884
rect 9772 37936 9824 37942
rect 9772 37878 9824 37884
rect 9220 37868 9272 37874
rect 9220 37810 9272 37816
rect 9128 37256 9180 37262
rect 9128 37198 9180 37204
rect 9140 36922 9168 37198
rect 9128 36916 9180 36922
rect 9128 36858 9180 36864
rect 9232 35698 9260 37810
rect 9312 37256 9364 37262
rect 9312 37198 9364 37204
rect 9324 37126 9352 37198
rect 9404 37188 9456 37194
rect 9404 37130 9456 37136
rect 9312 37120 9364 37126
rect 9312 37062 9364 37068
rect 9416 36922 9444 37130
rect 9404 36916 9456 36922
rect 9404 36858 9456 36864
rect 9404 35828 9456 35834
rect 9404 35770 9456 35776
rect 9220 35692 9272 35698
rect 9220 35634 9272 35640
rect 9312 35488 9364 35494
rect 9312 35430 9364 35436
rect 8956 35142 9076 35170
rect 8944 34536 8996 34542
rect 8850 34504 8906 34513
rect 8944 34478 8996 34484
rect 8850 34439 8906 34448
rect 8772 34360 8892 34388
rect 8668 33516 8720 33522
rect 8668 33458 8720 33464
rect 8760 33516 8812 33522
rect 8760 33458 8812 33464
rect 8680 33114 8708 33458
rect 8668 33108 8720 33114
rect 8668 33050 8720 33056
rect 8666 32872 8722 32881
rect 8666 32807 8722 32816
rect 8680 31906 8708 32807
rect 8772 32434 8800 33458
rect 8760 32428 8812 32434
rect 8760 32370 8812 32376
rect 8772 32026 8800 32370
rect 8760 32020 8812 32026
rect 8760 31962 8812 31968
rect 8680 31878 8800 31906
rect 8666 31240 8722 31249
rect 8666 31175 8722 31184
rect 8576 31136 8628 31142
rect 8576 31078 8628 31084
rect 8588 30326 8616 31078
rect 8680 30734 8708 31175
rect 8668 30728 8720 30734
rect 8668 30670 8720 30676
rect 8576 30320 8628 30326
rect 8576 30262 8628 30268
rect 8668 30252 8720 30258
rect 8668 30194 8720 30200
rect 8576 29640 8628 29646
rect 8576 29582 8628 29588
rect 8588 27849 8616 29582
rect 8680 28937 8708 30194
rect 8666 28928 8722 28937
rect 8666 28863 8722 28872
rect 8668 28688 8720 28694
rect 8668 28630 8720 28636
rect 8680 28150 8708 28630
rect 8668 28144 8720 28150
rect 8668 28086 8720 28092
rect 8574 27840 8630 27849
rect 8574 27775 8630 27784
rect 8668 26512 8720 26518
rect 8668 26454 8720 26460
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 8588 24410 8616 26318
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8576 24268 8628 24274
rect 8576 24210 8628 24216
rect 8588 22098 8616 24210
rect 8680 23361 8708 26454
rect 8666 23352 8722 23361
rect 8666 23287 8722 23296
rect 8668 23248 8720 23254
rect 8668 23190 8720 23196
rect 8680 22642 8708 23190
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8668 22024 8720 22030
rect 8574 21992 8630 22001
rect 8668 21966 8720 21972
rect 8574 21927 8630 21936
rect 8588 21622 8616 21927
rect 8576 21616 8628 21622
rect 8576 21558 8628 21564
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8588 19174 8616 19654
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8588 18630 8616 19110
rect 8680 18850 8708 21966
rect 8772 19281 8800 31878
rect 8864 31686 8892 34360
rect 8852 31680 8904 31686
rect 8852 31622 8904 31628
rect 8850 31512 8906 31521
rect 8956 31498 8984 34478
rect 9048 31754 9076 35142
rect 9128 34468 9180 34474
rect 9128 34410 9180 34416
rect 9140 34134 9168 34410
rect 9220 34196 9272 34202
rect 9220 34138 9272 34144
rect 9128 34128 9180 34134
rect 9128 34070 9180 34076
rect 9128 33992 9180 33998
rect 9126 33960 9128 33969
rect 9180 33960 9182 33969
rect 9126 33895 9182 33904
rect 9232 33561 9260 34138
rect 9218 33552 9274 33561
rect 9218 33487 9274 33496
rect 9232 31754 9260 33487
rect 9324 32230 9352 35430
rect 9416 35222 9444 35770
rect 9600 35766 9628 37878
rect 9680 37868 9732 37874
rect 9680 37810 9732 37816
rect 9692 37466 9720 37810
rect 9851 37564 10159 37573
rect 9851 37562 9857 37564
rect 9913 37562 9937 37564
rect 9993 37562 10017 37564
rect 10073 37562 10097 37564
rect 10153 37562 10159 37564
rect 9913 37510 9915 37562
rect 10095 37510 10097 37562
rect 9851 37508 9857 37510
rect 9913 37508 9937 37510
rect 9993 37508 10017 37510
rect 10073 37508 10097 37510
rect 10153 37508 10159 37510
rect 9851 37499 10159 37508
rect 9680 37460 9732 37466
rect 9680 37402 9732 37408
rect 10140 36916 10192 36922
rect 10140 36858 10192 36864
rect 10152 36786 10180 36858
rect 10140 36780 10192 36786
rect 10140 36722 10192 36728
rect 9851 36476 10159 36485
rect 9851 36474 9857 36476
rect 9913 36474 9937 36476
rect 9993 36474 10017 36476
rect 10073 36474 10097 36476
rect 10153 36474 10159 36476
rect 9913 36422 9915 36474
rect 10095 36422 10097 36474
rect 9851 36420 9857 36422
rect 9913 36420 9937 36422
rect 9993 36420 10017 36422
rect 10073 36420 10097 36422
rect 10153 36420 10159 36422
rect 9851 36411 10159 36420
rect 10244 36258 10272 38270
rect 10324 38208 10376 38214
rect 10324 38150 10376 38156
rect 10152 36230 10272 36258
rect 10048 36168 10100 36174
rect 10048 36110 10100 36116
rect 9956 36032 10008 36038
rect 10060 36009 10088 36110
rect 9956 35974 10008 35980
rect 10046 36000 10102 36009
rect 9588 35760 9640 35766
rect 9588 35702 9640 35708
rect 9968 35562 9996 35974
rect 10046 35935 10102 35944
rect 9956 35556 10008 35562
rect 9956 35498 10008 35504
rect 9496 35488 9548 35494
rect 10152 35476 10180 36230
rect 10336 36106 10364 38150
rect 10324 36100 10376 36106
rect 10324 36042 10376 36048
rect 10232 35828 10284 35834
rect 10232 35770 10284 35776
rect 10244 35630 10272 35770
rect 10428 35698 10456 39782
rect 10520 35748 10548 42638
rect 10704 40474 10732 42758
rect 10876 42696 10928 42702
rect 10876 42638 10928 42644
rect 10784 42628 10836 42634
rect 10784 42570 10836 42576
rect 10796 42362 10824 42570
rect 10784 42356 10836 42362
rect 10784 42298 10836 42304
rect 10784 41472 10836 41478
rect 10784 41414 10836 41420
rect 10888 41414 10916 42638
rect 11152 42560 11204 42566
rect 11152 42502 11204 42508
rect 11164 42362 11192 42502
rect 11152 42356 11204 42362
rect 11152 42298 11204 42304
rect 11256 41414 11284 43046
rect 11624 42702 11652 44934
rect 11794 44934 11928 44962
rect 11794 44840 11850 44934
rect 11796 43172 11848 43178
rect 11796 43114 11848 43120
rect 11612 42696 11664 42702
rect 11612 42638 11664 42644
rect 11336 42560 11388 42566
rect 11336 42502 11388 42508
rect 11348 41818 11376 42502
rect 11336 41812 11388 41818
rect 11336 41754 11388 41760
rect 10796 40730 10824 41414
rect 10888 41386 11008 41414
rect 11256 41386 11468 41414
rect 10876 40996 10928 41002
rect 10876 40938 10928 40944
rect 10784 40724 10836 40730
rect 10784 40666 10836 40672
rect 10888 40610 10916 40938
rect 10796 40594 10916 40610
rect 10784 40588 10916 40594
rect 10836 40582 10916 40588
rect 10784 40530 10836 40536
rect 10876 40520 10928 40526
rect 10704 40468 10876 40474
rect 10704 40462 10928 40468
rect 10704 40446 10916 40462
rect 10888 40186 10916 40446
rect 10876 40180 10928 40186
rect 10876 40122 10928 40128
rect 10690 40080 10746 40089
rect 10690 40015 10746 40024
rect 10600 38276 10652 38282
rect 10600 38218 10652 38224
rect 10612 38010 10640 38218
rect 10600 38004 10652 38010
rect 10600 37946 10652 37952
rect 10518 35720 10548 35748
rect 10416 35692 10468 35698
rect 10416 35634 10468 35640
rect 10232 35624 10284 35630
rect 10284 35584 10364 35612
rect 10232 35566 10284 35572
rect 10152 35448 10272 35476
rect 9496 35430 9548 35436
rect 9404 35216 9456 35222
rect 9404 35158 9456 35164
rect 9508 34950 9536 35430
rect 9851 35388 10159 35397
rect 9851 35386 9857 35388
rect 9913 35386 9937 35388
rect 9993 35386 10017 35388
rect 10073 35386 10097 35388
rect 10153 35386 10159 35388
rect 9913 35334 9915 35386
rect 10095 35334 10097 35386
rect 9851 35332 9857 35334
rect 9913 35332 9937 35334
rect 9993 35332 10017 35334
rect 10073 35332 10097 35334
rect 10153 35332 10159 35334
rect 9851 35323 10159 35332
rect 10048 35080 10100 35086
rect 10048 35022 10100 35028
rect 9864 35012 9916 35018
rect 9864 34954 9916 34960
rect 9496 34944 9548 34950
rect 9496 34886 9548 34892
rect 9876 34746 9904 34954
rect 10060 34950 10088 35022
rect 10048 34944 10100 34950
rect 10048 34886 10100 34892
rect 9864 34740 9916 34746
rect 9864 34682 9916 34688
rect 9494 34504 9550 34513
rect 9494 34439 9550 34448
rect 9588 34468 9640 34474
rect 9404 33856 9456 33862
rect 9402 33824 9404 33833
rect 9456 33824 9458 33833
rect 9402 33759 9458 33768
rect 9404 33516 9456 33522
rect 9404 33458 9456 33464
rect 9416 33114 9444 33458
rect 9508 33454 9536 34439
rect 9588 34410 9640 34416
rect 9600 34202 9628 34410
rect 9851 34300 10159 34309
rect 9851 34298 9857 34300
rect 9913 34298 9937 34300
rect 9993 34298 10017 34300
rect 10073 34298 10097 34300
rect 10153 34298 10159 34300
rect 9913 34246 9915 34298
rect 10095 34246 10097 34298
rect 9851 34244 9857 34246
rect 9913 34244 9937 34246
rect 9993 34244 10017 34246
rect 10073 34244 10097 34246
rect 10153 34244 10159 34246
rect 9851 34235 10159 34244
rect 9588 34196 9640 34202
rect 9588 34138 9640 34144
rect 10140 33992 10192 33998
rect 10140 33934 10192 33940
rect 10048 33924 10100 33930
rect 9784 33884 10048 33912
rect 9680 33856 9732 33862
rect 9600 33804 9680 33810
rect 9784 33833 9812 33884
rect 10048 33866 10100 33872
rect 9600 33798 9732 33804
rect 9770 33824 9826 33833
rect 9600 33782 9720 33798
rect 9600 33658 9628 33782
rect 9954 33824 10010 33833
rect 9770 33759 9826 33768
rect 9876 33782 9954 33810
rect 9770 33688 9826 33697
rect 9588 33652 9640 33658
rect 9588 33594 9640 33600
rect 9692 33646 9770 33674
rect 9496 33448 9548 33454
rect 9496 33390 9548 33396
rect 9586 33280 9642 33289
rect 9586 33215 9642 33224
rect 9404 33108 9456 33114
rect 9404 33050 9456 33056
rect 9496 32904 9548 32910
rect 9496 32846 9548 32852
rect 9508 32570 9536 32846
rect 9496 32564 9548 32570
rect 9496 32506 9548 32512
rect 9494 32464 9550 32473
rect 9494 32399 9550 32408
rect 9508 32366 9536 32399
rect 9496 32360 9548 32366
rect 9496 32302 9548 32308
rect 9600 32314 9628 33215
rect 9692 32978 9720 33646
rect 9770 33623 9826 33632
rect 9876 33318 9904 33782
rect 9954 33759 10010 33768
rect 10152 33658 10180 33934
rect 10140 33652 10192 33658
rect 10140 33594 10192 33600
rect 9954 33416 10010 33425
rect 9954 33351 10010 33360
rect 9968 33318 9996 33351
rect 9864 33312 9916 33318
rect 9784 33272 9864 33300
rect 9680 32972 9732 32978
rect 9680 32914 9732 32920
rect 9692 32434 9720 32914
rect 9680 32428 9732 32434
rect 9680 32370 9732 32376
rect 9312 32224 9364 32230
rect 9312 32166 9364 32172
rect 9048 31726 9168 31754
rect 9232 31726 9352 31754
rect 8906 31470 8984 31498
rect 8850 31447 8906 31456
rect 8864 30258 8892 31447
rect 9034 31376 9090 31385
rect 8944 31340 8996 31346
rect 9034 31311 9090 31320
rect 8944 31282 8996 31288
rect 8956 30666 8984 31282
rect 9048 31278 9076 31311
rect 9036 31272 9088 31278
rect 9036 31214 9088 31220
rect 9140 31124 9168 31726
rect 9220 31136 9272 31142
rect 9140 31096 9220 31124
rect 9034 30832 9090 30841
rect 9034 30767 9090 30776
rect 9048 30666 9076 30767
rect 8944 30660 8996 30666
rect 8944 30602 8996 30608
rect 9036 30660 9088 30666
rect 9036 30602 9088 30608
rect 9140 30410 9168 31096
rect 9220 31078 9272 31084
rect 8956 30382 9168 30410
rect 8852 30252 8904 30258
rect 8852 30194 8904 30200
rect 8864 29617 8892 30194
rect 8850 29608 8906 29617
rect 8850 29543 8906 29552
rect 8852 29504 8904 29510
rect 8852 29446 8904 29452
rect 8864 29170 8892 29446
rect 8852 29164 8904 29170
rect 8852 29106 8904 29112
rect 8852 28960 8904 28966
rect 8852 28902 8904 28908
rect 8864 26994 8892 28902
rect 8852 26988 8904 26994
rect 8852 26930 8904 26936
rect 8864 19417 8892 26930
rect 8956 24993 8984 30382
rect 9036 30320 9088 30326
rect 9034 30288 9036 30297
rect 9088 30288 9090 30297
rect 9034 30223 9090 30232
rect 9036 30184 9088 30190
rect 9036 30126 9088 30132
rect 9048 29102 9076 30126
rect 9220 30048 9272 30054
rect 9220 29990 9272 29996
rect 9232 29617 9260 29990
rect 9218 29608 9274 29617
rect 9218 29543 9274 29552
rect 9036 29096 9088 29102
rect 9036 29038 9088 29044
rect 9128 27872 9180 27878
rect 9128 27814 9180 27820
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 8942 24984 8998 24993
rect 8942 24919 8998 24928
rect 8944 24812 8996 24818
rect 8944 24754 8996 24760
rect 8956 23798 8984 24754
rect 8944 23792 8996 23798
rect 8944 23734 8996 23740
rect 9048 23610 9076 26930
rect 9140 26926 9168 27814
rect 9220 26988 9272 26994
rect 9324 26976 9352 31726
rect 9404 31680 9456 31686
rect 9404 31622 9456 31628
rect 9416 29578 9444 31622
rect 9508 30598 9536 32302
rect 9600 32286 9720 32314
rect 9586 32056 9642 32065
rect 9586 31991 9642 32000
rect 9600 31686 9628 31991
rect 9588 31680 9640 31686
rect 9588 31622 9640 31628
rect 9496 30592 9548 30598
rect 9496 30534 9548 30540
rect 9494 30288 9550 30297
rect 9494 30223 9550 30232
rect 9508 29782 9536 30223
rect 9496 29776 9548 29782
rect 9496 29718 9548 29724
rect 9496 29640 9548 29646
rect 9496 29582 9548 29588
rect 9404 29572 9456 29578
rect 9404 29514 9456 29520
rect 9272 26948 9352 26976
rect 9220 26930 9272 26936
rect 9128 26920 9180 26926
rect 9128 26862 9180 26868
rect 9140 26314 9168 26862
rect 9232 26518 9260 26930
rect 9220 26512 9272 26518
rect 9220 26454 9272 26460
rect 9128 26308 9180 26314
rect 9128 26250 9180 26256
rect 9508 26042 9536 29582
rect 9600 29306 9628 31622
rect 9692 31142 9720 32286
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 9680 30932 9732 30938
rect 9680 30874 9732 30880
rect 9692 30394 9720 30874
rect 9680 30388 9732 30394
rect 9680 30330 9732 30336
rect 9680 30184 9732 30190
rect 9680 30126 9732 30132
rect 9588 29300 9640 29306
rect 9588 29242 9640 29248
rect 9692 29238 9720 30126
rect 9784 29782 9812 33272
rect 9864 33254 9916 33260
rect 9956 33312 10008 33318
rect 9956 33254 10008 33260
rect 9851 33212 10159 33221
rect 9851 33210 9857 33212
rect 9913 33210 9937 33212
rect 9993 33210 10017 33212
rect 10073 33210 10097 33212
rect 10153 33210 10159 33212
rect 9913 33158 9915 33210
rect 10095 33158 10097 33210
rect 9851 33156 9857 33158
rect 9913 33156 9937 33158
rect 9993 33156 10017 33158
rect 10073 33156 10097 33158
rect 10153 33156 10159 33158
rect 9851 33147 10159 33156
rect 10046 33008 10102 33017
rect 10046 32943 10102 32952
rect 10060 32910 10088 32943
rect 10048 32904 10100 32910
rect 10048 32846 10100 32852
rect 9864 32836 9916 32842
rect 9864 32778 9916 32784
rect 9876 32502 9904 32778
rect 9864 32496 9916 32502
rect 9864 32438 9916 32444
rect 10244 32434 10272 35448
rect 10336 35290 10364 35584
rect 10324 35284 10376 35290
rect 10324 35226 10376 35232
rect 10322 35184 10378 35193
rect 10322 35119 10378 35128
rect 10336 33590 10364 35119
rect 10428 34542 10456 35634
rect 10518 35612 10546 35720
rect 10518 35584 10548 35612
rect 10416 34536 10468 34542
rect 10416 34478 10468 34484
rect 10520 34202 10548 35584
rect 10600 34604 10652 34610
rect 10600 34546 10652 34552
rect 10508 34196 10560 34202
rect 10508 34138 10560 34144
rect 10506 33960 10562 33969
rect 10506 33895 10562 33904
rect 10520 33862 10548 33895
rect 10508 33856 10560 33862
rect 10612 33833 10640 34546
rect 10508 33798 10560 33804
rect 10598 33824 10654 33833
rect 10520 33658 10548 33798
rect 10598 33759 10654 33768
rect 10508 33652 10560 33658
rect 10508 33594 10560 33600
rect 10324 33584 10376 33590
rect 10324 33526 10376 33532
rect 10324 33448 10376 33454
rect 10324 33390 10376 33396
rect 10232 32428 10284 32434
rect 10232 32370 10284 32376
rect 9851 32124 10159 32133
rect 9851 32122 9857 32124
rect 9913 32122 9937 32124
rect 9993 32122 10017 32124
rect 10073 32122 10097 32124
rect 10153 32122 10159 32124
rect 9913 32070 9915 32122
rect 10095 32070 10097 32122
rect 9851 32068 9857 32070
rect 9913 32068 9937 32070
rect 9993 32068 10017 32070
rect 10073 32068 10097 32070
rect 10153 32068 10159 32070
rect 9851 32059 10159 32068
rect 10232 32020 10284 32026
rect 10336 32008 10364 33390
rect 10416 33312 10468 33318
rect 10416 33254 10468 33260
rect 10284 31980 10364 32008
rect 10232 31962 10284 31968
rect 10428 31890 10456 33254
rect 10506 33008 10562 33017
rect 10704 32994 10732 40015
rect 10784 36712 10836 36718
rect 10784 36654 10836 36660
rect 10796 36378 10824 36654
rect 10876 36576 10928 36582
rect 10876 36518 10928 36524
rect 10784 36372 10836 36378
rect 10784 36314 10836 36320
rect 10796 33697 10824 36314
rect 10888 35222 10916 36518
rect 10876 35216 10928 35222
rect 10876 35158 10928 35164
rect 10980 34490 11008 41386
rect 11060 40928 11112 40934
rect 11060 40870 11112 40876
rect 11072 40594 11100 40870
rect 11060 40588 11112 40594
rect 11060 40530 11112 40536
rect 11152 40384 11204 40390
rect 11152 40326 11204 40332
rect 11336 40384 11388 40390
rect 11336 40326 11388 40332
rect 11164 38350 11192 40326
rect 11348 40118 11376 40326
rect 11336 40112 11388 40118
rect 11336 40054 11388 40060
rect 11336 39364 11388 39370
rect 11336 39306 11388 39312
rect 11348 38962 11376 39306
rect 11336 38956 11388 38962
rect 11336 38898 11388 38904
rect 11348 38729 11376 38898
rect 11334 38720 11390 38729
rect 11334 38655 11390 38664
rect 11152 38344 11204 38350
rect 11152 38286 11204 38292
rect 11060 37664 11112 37670
rect 11060 37606 11112 37612
rect 11072 35086 11100 37606
rect 11164 35086 11192 38286
rect 11244 38208 11296 38214
rect 11244 38150 11296 38156
rect 11256 35630 11284 38150
rect 11336 36032 11388 36038
rect 11336 35974 11388 35980
rect 11244 35624 11296 35630
rect 11244 35566 11296 35572
rect 11348 35086 11376 35974
rect 11060 35080 11112 35086
rect 11060 35022 11112 35028
rect 11152 35080 11204 35086
rect 11152 35022 11204 35028
rect 11336 35080 11388 35086
rect 11336 35022 11388 35028
rect 11072 34610 11100 35022
rect 11164 34678 11192 35022
rect 11152 34672 11204 34678
rect 11152 34614 11204 34620
rect 11334 34640 11390 34649
rect 11060 34604 11112 34610
rect 11334 34575 11390 34584
rect 11060 34546 11112 34552
rect 10980 34462 11192 34490
rect 10782 33688 10838 33697
rect 10782 33623 10838 33632
rect 10968 33584 11020 33590
rect 10968 33526 11020 33532
rect 10562 32966 10732 32994
rect 10506 32943 10562 32952
rect 10784 32768 10836 32774
rect 10784 32710 10836 32716
rect 10692 32428 10744 32434
rect 10692 32370 10744 32376
rect 10508 32224 10560 32230
rect 10508 32166 10560 32172
rect 10416 31884 10468 31890
rect 10416 31826 10468 31832
rect 10520 31804 10548 32166
rect 10704 31890 10732 32370
rect 10796 32026 10824 32710
rect 10784 32020 10836 32026
rect 10784 31962 10836 31968
rect 10692 31884 10744 31890
rect 10744 31844 10916 31872
rect 10692 31826 10744 31832
rect 10600 31816 10652 31822
rect 10520 31776 10600 31804
rect 10600 31758 10652 31764
rect 10612 31226 10640 31758
rect 10612 31198 10824 31226
rect 10692 31136 10744 31142
rect 10692 31078 10744 31084
rect 9851 31036 10159 31045
rect 9851 31034 9857 31036
rect 9913 31034 9937 31036
rect 9993 31034 10017 31036
rect 10073 31034 10097 31036
rect 10153 31034 10159 31036
rect 9913 30982 9915 31034
rect 10095 30982 10097 31034
rect 9851 30980 9857 30982
rect 9913 30980 9937 30982
rect 9993 30980 10017 30982
rect 10073 30980 10097 30982
rect 10153 30980 10159 30982
rect 9851 30971 10159 30980
rect 10508 30932 10560 30938
rect 10560 30892 10640 30920
rect 10508 30874 10560 30880
rect 9956 30796 10008 30802
rect 9956 30738 10008 30744
rect 9968 30433 9996 30738
rect 10508 30592 10560 30598
rect 10508 30534 10560 30540
rect 9954 30424 10010 30433
rect 9876 30382 9954 30410
rect 9876 30258 9904 30382
rect 9954 30359 10010 30368
rect 10046 30288 10102 30297
rect 9864 30252 9916 30258
rect 10046 30223 10102 30232
rect 9864 30194 9916 30200
rect 10060 30190 10088 30223
rect 10520 30190 10548 30534
rect 10048 30184 10100 30190
rect 10508 30184 10560 30190
rect 10048 30126 10100 30132
rect 10428 30132 10508 30138
rect 10428 30126 10560 30132
rect 10232 30116 10284 30122
rect 10232 30058 10284 30064
rect 10428 30110 10548 30126
rect 9851 29948 10159 29957
rect 9851 29946 9857 29948
rect 9913 29946 9937 29948
rect 9993 29946 10017 29948
rect 10073 29946 10097 29948
rect 10153 29946 10159 29948
rect 9913 29894 9915 29946
rect 10095 29894 10097 29946
rect 9851 29892 9857 29894
rect 9913 29892 9937 29894
rect 9993 29892 10017 29894
rect 10073 29892 10097 29894
rect 10153 29892 10159 29894
rect 9851 29883 10159 29892
rect 9772 29776 9824 29782
rect 9772 29718 9824 29724
rect 10140 29708 10192 29714
rect 10244 29696 10272 30058
rect 10428 30025 10456 30110
rect 10612 30036 10640 30892
rect 10414 30016 10470 30025
rect 10414 29951 10470 29960
rect 10520 30008 10640 30036
rect 10192 29668 10272 29696
rect 10140 29650 10192 29656
rect 9864 29640 9916 29646
rect 9864 29582 9916 29588
rect 9680 29232 9732 29238
rect 9586 29200 9642 29209
rect 9680 29174 9732 29180
rect 9586 29135 9588 29144
rect 9640 29135 9642 29144
rect 9588 29116 9640 29122
rect 9876 28966 9904 29582
rect 10152 29306 10180 29650
rect 10140 29300 10192 29306
rect 10140 29242 10192 29248
rect 10232 29028 10284 29034
rect 10232 28970 10284 28976
rect 9864 28960 9916 28966
rect 9864 28902 9916 28908
rect 9851 28860 10159 28869
rect 9851 28858 9857 28860
rect 9913 28858 9937 28860
rect 9993 28858 10017 28860
rect 10073 28858 10097 28860
rect 10153 28858 10159 28860
rect 9913 28806 9915 28858
rect 10095 28806 10097 28858
rect 9851 28804 9857 28806
rect 9913 28804 9937 28806
rect 9993 28804 10017 28806
rect 10073 28804 10097 28806
rect 10153 28804 10159 28806
rect 9678 28792 9734 28801
rect 9851 28795 10159 28804
rect 9734 28750 9812 28778
rect 9678 28727 9734 28736
rect 9680 27872 9732 27878
rect 9680 27814 9732 27820
rect 9692 27538 9720 27814
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 9588 27396 9640 27402
rect 9588 27338 9640 27344
rect 9680 27396 9732 27402
rect 9680 27338 9732 27344
rect 9496 26036 9548 26042
rect 9496 25978 9548 25984
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 9128 24744 9180 24750
rect 9128 24686 9180 24692
rect 8956 23582 9076 23610
rect 8956 20874 8984 23582
rect 9140 23474 9168 24686
rect 9232 24274 9260 25774
rect 9402 24984 9458 24993
rect 9402 24919 9458 24928
rect 9220 24268 9272 24274
rect 9220 24210 9272 24216
rect 9048 23446 9168 23474
rect 9310 23488 9366 23497
rect 9048 21350 9076 23446
rect 9416 23474 9444 24919
rect 9496 24744 9548 24750
rect 9496 24686 9548 24692
rect 9508 24410 9536 24686
rect 9496 24404 9548 24410
rect 9496 24346 9548 24352
rect 9416 23446 9536 23474
rect 9310 23423 9366 23432
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 9128 23112 9180 23118
rect 9128 23054 9180 23060
rect 9140 22778 9168 23054
rect 9232 22778 9260 23258
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 9220 22772 9272 22778
rect 9220 22714 9272 22720
rect 9128 22636 9180 22642
rect 9128 22578 9180 22584
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 9048 21146 9076 21286
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 8944 20868 8996 20874
rect 8944 20810 8996 20816
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 8942 20496 8998 20505
rect 9048 20466 9076 20742
rect 8942 20431 8998 20440
rect 9036 20460 9088 20466
rect 8956 19718 8984 20431
rect 9036 20402 9088 20408
rect 9034 20088 9090 20097
rect 9034 20023 9090 20032
rect 9048 19922 9076 20023
rect 9036 19916 9088 19922
rect 9036 19858 9088 19864
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 9048 19530 9076 19858
rect 8956 19502 9076 19530
rect 8850 19408 8906 19417
rect 8956 19378 8984 19502
rect 9140 19428 9168 22578
rect 9220 22092 9272 22098
rect 9220 22034 9272 22040
rect 9232 21010 9260 22034
rect 9324 22030 9352 23423
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9416 22098 9444 22374
rect 9404 22092 9456 22098
rect 9404 22034 9456 22040
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 9324 21457 9352 21490
rect 9310 21448 9366 21457
rect 9310 21383 9366 21392
rect 9310 21176 9366 21185
rect 9310 21111 9366 21120
rect 9220 21004 9272 21010
rect 9220 20946 9272 20952
rect 9232 19922 9260 20946
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 9232 19514 9260 19654
rect 9218 19508 9270 19514
rect 9218 19450 9270 19456
rect 9048 19400 9168 19428
rect 8850 19343 8906 19352
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 9048 19334 9076 19400
rect 9048 19306 9168 19334
rect 8758 19272 8814 19281
rect 8758 19207 8814 19216
rect 8852 19236 8904 19242
rect 8852 19178 8904 19184
rect 8864 18970 8892 19178
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 8680 18822 8800 18850
rect 8666 18728 8722 18737
rect 8666 18663 8722 18672
rect 8680 18630 8708 18663
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8772 16130 8800 18822
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 9048 18290 9076 18770
rect 9036 18284 9088 18290
rect 8956 18244 9036 18272
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8588 16102 8800 16130
rect 8864 16114 8892 16934
rect 8852 16108 8904 16114
rect 8588 13705 8616 16102
rect 8852 16050 8904 16056
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8574 13696 8630 13705
rect 8574 13631 8630 13640
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8390 9007 8446 9016
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7852 4078 7880 5850
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8312 4978 8340 5034
rect 8220 4950 8340 4978
rect 8220 4128 8248 4950
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8128 4100 8248 4128
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7852 2990 7880 4014
rect 8128 4010 8156 4100
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8128 2990 8156 3946
rect 8220 3738 8248 3946
rect 8312 3738 8340 4762
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8404 3466 8432 7890
rect 8588 6882 8616 13330
rect 8680 8022 8708 13874
rect 8772 12102 8800 15982
rect 8956 13530 8984 18244
rect 9036 18226 9088 18232
rect 9036 17672 9088 17678
rect 9140 17660 9168 19306
rect 9088 17632 9168 17660
rect 9036 17614 9088 17620
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 9048 12730 9076 17614
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 8956 12702 9076 12730
rect 8956 12434 8984 12702
rect 9140 12434 9168 17478
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9232 15706 9260 17274
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9232 15162 9260 15642
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9232 13870 9260 14010
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 8864 12406 8984 12434
rect 9048 12406 9168 12434
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8760 11824 8812 11830
rect 8760 11766 8812 11772
rect 8772 11218 8800 11766
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8588 6854 8708 6882
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8588 6225 8616 6666
rect 8574 6216 8630 6225
rect 8574 6151 8630 6160
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8496 4690 8524 5170
rect 8680 5098 8708 6854
rect 8772 5896 8800 9998
rect 8864 9636 8892 12406
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8956 11150 8984 11562
rect 8944 11144 8996 11150
rect 9048 11132 9076 12406
rect 9232 11558 9260 12582
rect 9324 12434 9352 21111
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 9416 19514 9444 19858
rect 9508 19786 9536 23446
rect 9600 22094 9628 27338
rect 9692 27130 9720 27338
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9784 26217 9812 28750
rect 9851 27772 10159 27781
rect 9851 27770 9857 27772
rect 9913 27770 9937 27772
rect 9993 27770 10017 27772
rect 10073 27770 10097 27772
rect 10153 27770 10159 27772
rect 9913 27718 9915 27770
rect 10095 27718 10097 27770
rect 9851 27716 9857 27718
rect 9913 27716 9937 27718
rect 9993 27716 10017 27718
rect 10073 27716 10097 27718
rect 10153 27716 10159 27718
rect 9851 27707 10159 27716
rect 10244 27520 10272 28970
rect 10324 27872 10376 27878
rect 10324 27814 10376 27820
rect 10152 27492 10272 27520
rect 10048 27396 10100 27402
rect 10152 27384 10180 27492
rect 10336 27418 10364 27814
rect 10520 27690 10548 30008
rect 10600 28756 10652 28762
rect 10600 28698 10652 28704
rect 10612 28529 10640 28698
rect 10598 28520 10654 28529
rect 10598 28455 10654 28464
rect 10612 28150 10640 28455
rect 10600 28144 10652 28150
rect 10600 28086 10652 28092
rect 10612 27849 10640 28086
rect 10598 27840 10654 27849
rect 10598 27775 10654 27784
rect 10520 27662 10640 27690
rect 10506 27568 10562 27577
rect 10506 27503 10562 27512
rect 10100 27356 10180 27384
rect 10048 27338 10100 27344
rect 10152 26994 10180 27356
rect 10244 27390 10364 27418
rect 10140 26988 10192 26994
rect 10140 26930 10192 26936
rect 9851 26684 10159 26693
rect 9851 26682 9857 26684
rect 9913 26682 9937 26684
rect 9993 26682 10017 26684
rect 10073 26682 10097 26684
rect 10153 26682 10159 26684
rect 9913 26630 9915 26682
rect 10095 26630 10097 26682
rect 9851 26628 9857 26630
rect 9913 26628 9937 26630
rect 9993 26628 10017 26630
rect 10073 26628 10097 26630
rect 10153 26628 10159 26630
rect 9851 26619 10159 26628
rect 9770 26208 9826 26217
rect 9770 26143 9826 26152
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 9680 24744 9732 24750
rect 9680 24686 9732 24692
rect 9692 24070 9720 24686
rect 9784 24138 9812 25978
rect 10140 25900 10192 25906
rect 10244 25888 10272 27390
rect 10324 27328 10376 27334
rect 10324 27270 10376 27276
rect 10416 27328 10468 27334
rect 10416 27270 10468 27276
rect 10192 25860 10272 25888
rect 10140 25842 10192 25848
rect 9851 25596 10159 25605
rect 9851 25594 9857 25596
rect 9913 25594 9937 25596
rect 9993 25594 10017 25596
rect 10073 25594 10097 25596
rect 10153 25594 10159 25596
rect 9913 25542 9915 25594
rect 10095 25542 10097 25594
rect 9851 25540 9857 25542
rect 9913 25540 9937 25542
rect 9993 25540 10017 25542
rect 10073 25540 10097 25542
rect 10153 25540 10159 25542
rect 9851 25531 10159 25540
rect 10048 25356 10100 25362
rect 10048 25298 10100 25304
rect 10060 24750 10088 25298
rect 10336 24834 10364 27270
rect 10428 26926 10456 27270
rect 10416 26920 10468 26926
rect 10416 26862 10468 26868
rect 10428 25362 10456 26862
rect 10416 25356 10468 25362
rect 10416 25298 10468 25304
rect 10520 24954 10548 27503
rect 10612 25378 10640 27662
rect 10704 26042 10732 31078
rect 10796 29306 10824 31198
rect 10888 29714 10916 31844
rect 10980 31142 11008 33526
rect 11060 32224 11112 32230
rect 11060 32166 11112 32172
rect 11072 31890 11100 32166
rect 11060 31884 11112 31890
rect 11060 31826 11112 31832
rect 10968 31136 11020 31142
rect 10968 31078 11020 31084
rect 11060 30592 11112 30598
rect 11060 30534 11112 30540
rect 11072 30190 11100 30534
rect 11060 30184 11112 30190
rect 11060 30126 11112 30132
rect 10876 29708 10928 29714
rect 10876 29650 10928 29656
rect 10888 29510 10916 29650
rect 10968 29640 11020 29646
rect 11072 29628 11100 30126
rect 11020 29600 11100 29628
rect 10968 29582 11020 29588
rect 10876 29504 10928 29510
rect 10876 29446 10928 29452
rect 10784 29300 10836 29306
rect 10784 29242 10836 29248
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10612 25362 10732 25378
rect 10612 25356 10744 25362
rect 10612 25350 10692 25356
rect 10692 25298 10744 25304
rect 10600 25288 10652 25294
rect 10600 25230 10652 25236
rect 10612 24954 10640 25230
rect 10508 24948 10560 24954
rect 10508 24890 10560 24896
rect 10600 24948 10652 24954
rect 10600 24890 10652 24896
rect 10336 24818 10548 24834
rect 10336 24812 10560 24818
rect 10336 24806 10508 24812
rect 10048 24744 10100 24750
rect 10100 24692 10272 24698
rect 10048 24686 10272 24692
rect 10060 24670 10272 24686
rect 9851 24508 10159 24517
rect 9851 24506 9857 24508
rect 9913 24506 9937 24508
rect 9993 24506 10017 24508
rect 10073 24506 10097 24508
rect 10153 24506 10159 24508
rect 9913 24454 9915 24506
rect 10095 24454 10097 24506
rect 9851 24452 9857 24454
rect 9913 24452 9937 24454
rect 9993 24452 10017 24454
rect 10073 24452 10097 24454
rect 10153 24452 10159 24454
rect 9851 24443 10159 24452
rect 10244 24410 10272 24670
rect 10232 24404 10284 24410
rect 10232 24346 10284 24352
rect 9772 24132 9824 24138
rect 9772 24074 9824 24080
rect 9680 24064 9732 24070
rect 9680 24006 9732 24012
rect 10230 23488 10286 23497
rect 9851 23420 10159 23429
rect 10230 23423 10286 23432
rect 9851 23418 9857 23420
rect 9913 23418 9937 23420
rect 9993 23418 10017 23420
rect 10073 23418 10097 23420
rect 10153 23418 10159 23420
rect 9913 23366 9915 23418
rect 10095 23366 10097 23418
rect 9851 23364 9857 23366
rect 9913 23364 9937 23366
rect 9993 23364 10017 23366
rect 10073 23364 10097 23366
rect 10153 23364 10159 23366
rect 9851 23355 10159 23364
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 9784 22982 9812 23054
rect 9772 22976 9824 22982
rect 9772 22918 9824 22924
rect 9784 22438 9812 22918
rect 10152 22817 10180 23054
rect 10138 22808 10194 22817
rect 10138 22743 10194 22752
rect 10244 22710 10272 23423
rect 10232 22704 10284 22710
rect 10232 22646 10284 22652
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9600 22066 9720 22094
rect 9692 20466 9720 22066
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9494 19680 9550 19689
rect 9494 19615 9550 19624
rect 9508 19514 9536 19615
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9600 18766 9628 20402
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9692 18630 9720 20402
rect 9784 20312 9812 22374
rect 9851 22332 10159 22341
rect 9851 22330 9857 22332
rect 9913 22330 9937 22332
rect 9993 22330 10017 22332
rect 10073 22330 10097 22332
rect 10153 22330 10159 22332
rect 9913 22278 9915 22330
rect 10095 22278 10097 22330
rect 9851 22276 9857 22278
rect 9913 22276 9937 22278
rect 9993 22276 10017 22278
rect 10073 22276 10097 22278
rect 10153 22276 10159 22278
rect 9851 22267 10159 22276
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 9851 21244 10159 21253
rect 9851 21242 9857 21244
rect 9913 21242 9937 21244
rect 9993 21242 10017 21244
rect 10073 21242 10097 21244
rect 10153 21242 10159 21244
rect 9913 21190 9915 21242
rect 10095 21190 10097 21242
rect 9851 21188 9857 21190
rect 9913 21188 9937 21190
rect 9993 21188 10017 21190
rect 10073 21188 10097 21190
rect 10153 21188 10159 21190
rect 9851 21179 10159 21188
rect 10244 20380 10272 21966
rect 10336 20602 10364 24806
rect 10508 24754 10560 24760
rect 10416 24744 10468 24750
rect 10416 24686 10468 24692
rect 10428 24426 10456 24686
rect 10520 24585 10548 24754
rect 10506 24576 10562 24585
rect 10506 24511 10562 24520
rect 10506 24440 10562 24449
rect 10428 24398 10506 24426
rect 10506 24375 10562 24384
rect 10612 24256 10640 24890
rect 10704 24614 10732 25298
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10520 24228 10640 24256
rect 10520 24018 10548 24228
rect 10428 23990 10548 24018
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10428 22642 10456 23990
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 10508 22568 10560 22574
rect 10508 22510 10560 22516
rect 10414 22400 10470 22409
rect 10414 22335 10470 22344
rect 10428 22030 10456 22335
rect 10520 22234 10548 22510
rect 10508 22228 10560 22234
rect 10508 22170 10560 22176
rect 10416 22024 10468 22030
rect 10416 21966 10468 21972
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10428 20534 10456 20742
rect 10416 20528 10468 20534
rect 10416 20470 10468 20476
rect 10508 20528 10560 20534
rect 10508 20470 10560 20476
rect 10244 20352 10364 20380
rect 9782 20284 9812 20312
rect 9782 19938 9810 20284
rect 9851 20156 10159 20165
rect 9851 20154 9857 20156
rect 9913 20154 9937 20156
rect 9993 20154 10017 20156
rect 10073 20154 10097 20156
rect 10153 20154 10159 20156
rect 9913 20102 9915 20154
rect 10095 20102 10097 20154
rect 9851 20100 9857 20102
rect 9913 20100 9937 20102
rect 9993 20100 10017 20102
rect 10073 20100 10097 20102
rect 10153 20100 10159 20102
rect 9851 20091 10159 20100
rect 9954 19952 10010 19961
rect 9782 19910 9812 19938
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9692 17814 9720 18226
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9678 17640 9734 17649
rect 9678 17575 9734 17584
rect 9692 17338 9720 17575
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9588 17264 9640 17270
rect 9508 17224 9588 17252
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9416 16182 9444 16390
rect 9404 16176 9456 16182
rect 9404 16118 9456 16124
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 9416 12646 9444 14962
rect 9508 13938 9536 17224
rect 9588 17206 9640 17212
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9692 17105 9720 17138
rect 9678 17096 9734 17105
rect 9678 17031 9734 17040
rect 9588 16992 9640 16998
rect 9640 16952 9720 16980
rect 9588 16934 9640 16940
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9600 16250 9628 16458
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9600 15706 9628 15982
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9600 13410 9628 15438
rect 9692 14822 9720 16952
rect 9784 16658 9812 19910
rect 10336 19938 10364 20352
rect 10414 20360 10470 20369
rect 10414 20295 10470 20304
rect 9954 19887 10010 19896
rect 10244 19910 10364 19938
rect 9968 19786 9996 19887
rect 9956 19780 10008 19786
rect 9956 19722 10008 19728
rect 9851 19068 10159 19077
rect 9851 19066 9857 19068
rect 9913 19066 9937 19068
rect 9993 19066 10017 19068
rect 10073 19066 10097 19068
rect 10153 19066 10159 19068
rect 9913 19014 9915 19066
rect 10095 19014 10097 19066
rect 9851 19012 9857 19014
rect 9913 19012 9937 19014
rect 9993 19012 10017 19014
rect 10073 19012 10097 19014
rect 10153 19012 10159 19014
rect 9851 19003 10159 19012
rect 10244 18834 10272 19910
rect 10322 19816 10378 19825
rect 10322 19751 10378 19760
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 9851 17980 10159 17989
rect 9851 17978 9857 17980
rect 9913 17978 9937 17980
rect 9993 17978 10017 17980
rect 10073 17978 10097 17980
rect 10153 17978 10159 17980
rect 9913 17926 9915 17978
rect 10095 17926 10097 17978
rect 9851 17924 9857 17926
rect 9913 17924 9937 17926
rect 9993 17924 10017 17926
rect 10073 17924 10097 17926
rect 10153 17924 10159 17926
rect 9851 17915 10159 17924
rect 10244 17864 10272 18362
rect 10152 17836 10272 17864
rect 10152 17678 10180 17836
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10232 17672 10284 17678
rect 10336 17649 10364 19751
rect 10232 17614 10284 17620
rect 10322 17640 10378 17649
rect 10152 17218 10180 17614
rect 10244 17338 10272 17614
rect 10322 17575 10378 17584
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10336 17270 10364 17575
rect 10324 17264 10376 17270
rect 10152 17190 10272 17218
rect 10324 17206 10376 17212
rect 9851 16892 10159 16901
rect 9851 16890 9857 16892
rect 9913 16890 9937 16892
rect 9993 16890 10017 16892
rect 10073 16890 10097 16892
rect 10153 16890 10159 16892
rect 9913 16838 9915 16890
rect 10095 16838 10097 16890
rect 9851 16836 9857 16838
rect 9913 16836 9937 16838
rect 9993 16836 10017 16838
rect 10073 16836 10097 16838
rect 10153 16836 10159 16838
rect 9851 16827 10159 16836
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 10244 16522 10272 17190
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 9784 15502 9812 16458
rect 10336 15858 10364 16594
rect 10244 15830 10364 15858
rect 9851 15804 10159 15813
rect 9851 15802 9857 15804
rect 9913 15802 9937 15804
rect 9993 15802 10017 15804
rect 10073 15802 10097 15804
rect 10153 15802 10159 15804
rect 9913 15750 9915 15802
rect 10095 15750 10097 15802
rect 9851 15748 9857 15750
rect 9913 15748 9937 15750
rect 9993 15748 10017 15750
rect 10073 15748 10097 15750
rect 10153 15748 10159 15750
rect 9851 15739 10159 15748
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9692 13530 9720 14010
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9508 13394 9628 13410
rect 9496 13388 9628 13394
rect 9548 13382 9628 13388
rect 9496 13330 9548 13336
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9508 12782 9536 13126
rect 9600 12850 9628 13382
rect 9680 13388 9732 13394
rect 9784 13376 9812 15438
rect 9851 14716 10159 14725
rect 9851 14714 9857 14716
rect 9913 14714 9937 14716
rect 9993 14714 10017 14716
rect 10073 14714 10097 14716
rect 10153 14714 10159 14716
rect 9913 14662 9915 14714
rect 10095 14662 10097 14714
rect 9851 14660 9857 14662
rect 9913 14660 9937 14662
rect 9993 14660 10017 14662
rect 10073 14660 10097 14662
rect 10153 14660 10159 14662
rect 9851 14651 10159 14660
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 10152 13716 10180 14486
rect 10244 14278 10272 15830
rect 10428 15722 10456 20295
rect 10520 18970 10548 20470
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10612 18426 10640 24006
rect 10692 22636 10744 22642
rect 10692 22578 10744 22584
rect 10704 20369 10732 22578
rect 10796 22012 10824 29242
rect 11164 28642 11192 34462
rect 11348 33930 11376 34575
rect 11336 33924 11388 33930
rect 11336 33866 11388 33872
rect 11244 33380 11296 33386
rect 11244 33322 11296 33328
rect 11256 32473 11284 33322
rect 11242 32464 11298 32473
rect 11242 32399 11298 32408
rect 11244 31884 11296 31890
rect 11244 31826 11296 31832
rect 11256 31793 11284 31826
rect 11242 31784 11298 31793
rect 11242 31719 11298 31728
rect 11336 30048 11388 30054
rect 11336 29990 11388 29996
rect 11348 29306 11376 29990
rect 11336 29300 11388 29306
rect 11336 29242 11388 29248
rect 11164 28614 11284 28642
rect 11256 28218 11284 28614
rect 10968 28212 11020 28218
rect 10968 28154 11020 28160
rect 11244 28212 11296 28218
rect 11244 28154 11296 28160
rect 10980 27538 11008 28154
rect 11058 28112 11114 28121
rect 11058 28047 11114 28056
rect 10968 27532 11020 27538
rect 10968 27474 11020 27480
rect 11072 27062 11100 28047
rect 11244 27872 11296 27878
rect 11244 27814 11296 27820
rect 11256 27674 11284 27814
rect 11244 27668 11296 27674
rect 11244 27610 11296 27616
rect 11152 27464 11204 27470
rect 11152 27406 11204 27412
rect 11164 27130 11192 27406
rect 11152 27124 11204 27130
rect 11152 27066 11204 27072
rect 11060 27056 11112 27062
rect 11060 26998 11112 27004
rect 11060 26784 11112 26790
rect 11060 26726 11112 26732
rect 10876 25696 10928 25702
rect 10876 25638 10928 25644
rect 10888 25362 10916 25638
rect 11072 25401 11100 26726
rect 11058 25392 11114 25401
rect 10876 25356 10928 25362
rect 11058 25327 11114 25336
rect 10876 25298 10928 25304
rect 10888 24750 10916 25298
rect 11334 24848 11390 24857
rect 11334 24783 11390 24792
rect 10876 24744 10928 24750
rect 10876 24686 10928 24692
rect 10876 24608 10928 24614
rect 10876 24550 10928 24556
rect 10888 22080 10916 24550
rect 11244 23724 11296 23730
rect 11244 23666 11296 23672
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 10968 22976 11020 22982
rect 10968 22918 11020 22924
rect 10980 22710 11008 22918
rect 10968 22704 11020 22710
rect 10968 22646 11020 22652
rect 11072 22166 11100 23598
rect 11152 22704 11204 22710
rect 11150 22672 11152 22681
rect 11204 22672 11206 22681
rect 11150 22607 11206 22616
rect 11256 22556 11284 23666
rect 11348 23050 11376 24783
rect 11336 23044 11388 23050
rect 11336 22986 11388 22992
rect 11164 22528 11284 22556
rect 11060 22160 11112 22166
rect 11060 22102 11112 22108
rect 10888 22052 11008 22080
rect 10796 21984 10916 22012
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 10690 20360 10746 20369
rect 10690 20295 10746 20304
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10612 17898 10640 18226
rect 10704 18193 10732 20198
rect 10690 18184 10746 18193
rect 10690 18119 10746 18128
rect 10612 17882 10732 17898
rect 10612 17876 10744 17882
rect 10612 17870 10692 17876
rect 10692 17818 10744 17824
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10704 16658 10732 17070
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10690 16552 10746 16561
rect 10690 16487 10746 16496
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10336 15694 10456 15722
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10152 13688 10272 13716
rect 9851 13628 10159 13637
rect 9851 13626 9857 13628
rect 9913 13626 9937 13628
rect 9993 13626 10017 13628
rect 10073 13626 10097 13628
rect 10153 13626 10159 13628
rect 9913 13574 9915 13626
rect 10095 13574 10097 13626
rect 9851 13572 9857 13574
rect 9913 13572 9937 13574
rect 9993 13572 10017 13574
rect 10073 13572 10097 13574
rect 10153 13572 10159 13574
rect 9851 13563 10159 13572
rect 10244 13530 10272 13688
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10152 13394 10180 13466
rect 10336 13433 10364 15694
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10322 13424 10378 13433
rect 9732 13348 9812 13376
rect 10140 13388 10192 13394
rect 9680 13330 9732 13336
rect 10322 13359 10378 13368
rect 10140 13330 10192 13336
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9324 12406 9444 12434
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9324 11370 9352 12242
rect 9232 11342 9352 11370
rect 9048 11104 9168 11132
rect 8944 11086 8996 11092
rect 9140 10577 9168 11104
rect 9126 10568 9182 10577
rect 9126 10503 9182 10512
rect 9140 10130 9168 10503
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9036 9648 9088 9654
rect 8864 9608 9036 9636
rect 8864 6322 8892 9608
rect 9036 9590 9088 9596
rect 9232 9466 9260 11342
rect 9416 9674 9444 12406
rect 9508 12306 9536 12718
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9692 12170 9720 13330
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9876 13190 9904 13262
rect 9864 13184 9916 13190
rect 9784 13144 9864 13172
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9588 11688 9640 11694
rect 9640 11636 9720 11642
rect 9588 11630 9720 11636
rect 9600 11614 9720 11630
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9048 9438 9260 9466
rect 9324 9646 9444 9674
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8956 6458 8984 9318
rect 9048 6769 9076 9438
rect 9128 8968 9180 8974
rect 9324 8956 9352 9646
rect 9508 9602 9536 11018
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9600 9722 9628 10066
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9508 9574 9628 9602
rect 9402 9480 9458 9489
rect 9402 9415 9458 9424
rect 9180 8928 9352 8956
rect 9128 8910 9180 8916
rect 9034 6760 9090 6769
rect 9034 6695 9090 6704
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 9048 6322 9076 6598
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9140 6202 9168 8910
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 7886 9260 8230
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9324 7818 9352 8366
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9416 7546 9444 9415
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9048 6174 9168 6202
rect 8852 5908 8904 5914
rect 8772 5868 8852 5896
rect 8852 5850 8904 5856
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8772 4978 8800 5646
rect 8864 5137 8892 5850
rect 8850 5128 8906 5137
rect 8850 5063 8906 5072
rect 8772 4950 8892 4978
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8864 4486 8892 4950
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8772 4146 8800 4422
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8588 3466 8616 3878
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8390 3088 8446 3097
rect 8390 3023 8446 3032
rect 8484 3052 8536 3058
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 7760 2746 8064 2774
rect 7932 2304 7984 2310
rect 7746 2272 7802 2281
rect 7932 2246 7984 2252
rect 7746 2207 7802 2216
rect 7760 2106 7788 2207
rect 7944 2106 7972 2246
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 7932 2100 7984 2106
rect 7932 2042 7984 2048
rect 8036 1902 8064 2746
rect 8220 2650 8248 2858
rect 8404 2650 8432 3023
rect 8588 3040 8616 3402
rect 8680 3058 8708 4014
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8772 3058 8800 3334
rect 8536 3012 8616 3040
rect 8668 3052 8720 3058
rect 8484 2994 8536 3000
rect 8668 2994 8720 3000
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8484 2440 8536 2446
rect 8404 2400 8484 2428
rect 8114 2272 8170 2281
rect 8114 2207 8170 2216
rect 8128 2106 8156 2207
rect 8116 2100 8168 2106
rect 8116 2042 8168 2048
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 8024 1896 8076 1902
rect 8024 1838 8076 1844
rect 7748 1488 7800 1494
rect 7748 1430 7800 1436
rect 6826 82 6882 160
rect 6656 54 6882 82
rect 6826 0 6882 54
rect 7102 0 7158 160
rect 7378 0 7434 160
rect 7654 0 7710 160
rect 7760 82 7788 1430
rect 8208 1352 8260 1358
rect 8208 1294 8260 1300
rect 7932 1216 7984 1222
rect 7932 1158 7984 1164
rect 7944 921 7972 1158
rect 7930 912 7986 921
rect 7930 847 7986 856
rect 8220 160 8248 1294
rect 8312 1018 8340 1906
rect 8404 1306 8432 2400
rect 8484 2382 8536 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 8576 2304 8628 2310
rect 8482 2272 8538 2281
rect 8576 2246 8628 2252
rect 8482 2207 8538 2216
rect 8496 2106 8524 2207
rect 8588 2106 8616 2246
rect 8484 2100 8536 2106
rect 8484 2042 8536 2048
rect 8576 2100 8628 2106
rect 8576 2042 8628 2048
rect 8404 1278 8524 1306
rect 8300 1012 8352 1018
rect 8300 954 8352 960
rect 8496 160 8524 1278
rect 8680 1018 8708 2314
rect 8668 1012 8720 1018
rect 8668 954 8720 960
rect 8772 160 8800 2382
rect 8850 2272 8906 2281
rect 8850 2207 8906 2216
rect 8864 2106 8892 2207
rect 8852 2100 8904 2106
rect 8852 2042 8904 2048
rect 8956 2038 8984 3334
rect 8944 2032 8996 2038
rect 8944 1974 8996 1980
rect 9048 1562 9076 6174
rect 9232 6100 9260 7210
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9140 6072 9260 6100
rect 9140 5710 9168 6072
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9140 5234 9168 5646
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9140 4758 9168 5170
rect 9128 4752 9180 4758
rect 9128 4694 9180 4700
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9140 2774 9168 3470
rect 9324 2922 9352 5646
rect 9416 4672 9444 6666
rect 9508 5234 9536 8230
rect 9600 6905 9628 9574
rect 9692 7970 9720 11614
rect 9784 10248 9812 13144
rect 9864 13126 9916 13132
rect 10428 12782 10456 15438
rect 10416 12776 10468 12782
rect 10414 12744 10416 12753
rect 10468 12744 10470 12753
rect 10048 12708 10100 12714
rect 10100 12668 10272 12696
rect 10414 12679 10470 12688
rect 10048 12650 10100 12656
rect 9851 12540 10159 12549
rect 9851 12538 9857 12540
rect 9913 12538 9937 12540
rect 9993 12538 10017 12540
rect 10073 12538 10097 12540
rect 10153 12538 10159 12540
rect 9913 12486 9915 12538
rect 10095 12486 10097 12538
rect 9851 12484 9857 12486
rect 9913 12484 9937 12486
rect 9993 12484 10017 12486
rect 10073 12484 10097 12486
rect 10153 12484 10159 12486
rect 9851 12475 10159 12484
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10060 11898 10088 12174
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9851 11452 10159 11461
rect 9851 11450 9857 11452
rect 9913 11450 9937 11452
rect 9993 11450 10017 11452
rect 10073 11450 10097 11452
rect 10153 11450 10159 11452
rect 9913 11398 9915 11450
rect 10095 11398 10097 11450
rect 9851 11396 9857 11398
rect 9913 11396 9937 11398
rect 9993 11396 10017 11398
rect 10073 11396 10097 11398
rect 10153 11396 10159 11398
rect 9851 11387 10159 11396
rect 10244 11354 10272 12668
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10152 10742 10180 11154
rect 10336 10962 10364 11834
rect 10520 11082 10548 16050
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10612 15706 10640 15846
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10612 15162 10640 15438
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10612 11898 10640 12718
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10244 10934 10364 10962
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 9851 10364 10159 10373
rect 9851 10362 9857 10364
rect 9913 10362 9937 10364
rect 9993 10362 10017 10364
rect 10073 10362 10097 10364
rect 10153 10362 10159 10364
rect 9913 10310 9915 10362
rect 10095 10310 10097 10362
rect 9851 10308 9857 10310
rect 9913 10308 9937 10310
rect 9993 10308 10017 10310
rect 10073 10308 10097 10310
rect 10153 10308 10159 10310
rect 9851 10299 10159 10308
rect 9784 10220 9904 10248
rect 9876 10130 9904 10220
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10152 9722 10180 9998
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 9851 9276 10159 9285
rect 9851 9274 9857 9276
rect 9913 9274 9937 9276
rect 9993 9274 10017 9276
rect 10073 9274 10097 9276
rect 10153 9274 10159 9276
rect 9913 9222 9915 9274
rect 10095 9222 10097 9274
rect 9851 9220 9857 9222
rect 9913 9220 9937 9222
rect 9993 9220 10017 9222
rect 10073 9220 10097 9222
rect 10153 9220 10159 9222
rect 9851 9211 10159 9220
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9784 8090 9812 9046
rect 10244 8838 10272 10934
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10428 9674 10456 9862
rect 10336 9646 10456 9674
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 9851 8188 10159 8197
rect 9851 8186 9857 8188
rect 9913 8186 9937 8188
rect 9993 8186 10017 8188
rect 10073 8186 10097 8188
rect 10153 8186 10159 8188
rect 9913 8134 9915 8186
rect 10095 8134 10097 8186
rect 9851 8132 9857 8134
rect 9913 8132 9937 8134
rect 9993 8132 10017 8134
rect 10073 8132 10097 8134
rect 10153 8132 10159 8134
rect 9851 8123 10159 8132
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9692 7942 9812 7970
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9586 6896 9642 6905
rect 9586 6831 9642 6840
rect 9692 6458 9720 7346
rect 9784 6769 9812 7942
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9876 7478 9904 7754
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9851 7100 10159 7109
rect 9851 7098 9857 7100
rect 9913 7098 9937 7100
rect 9993 7098 10017 7100
rect 10073 7098 10097 7100
rect 10153 7098 10159 7100
rect 9913 7046 9915 7098
rect 10095 7046 10097 7098
rect 9851 7044 9857 7046
rect 9913 7044 9937 7046
rect 9993 7044 10017 7046
rect 10073 7044 10097 7046
rect 10153 7044 10159 7046
rect 9851 7035 10159 7044
rect 9770 6760 9826 6769
rect 9770 6695 9826 6704
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9586 5400 9642 5409
rect 9586 5335 9588 5344
rect 9640 5335 9642 5344
rect 9588 5306 9640 5312
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9692 4826 9720 5102
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9416 4644 9536 4672
rect 9402 4584 9458 4593
rect 9402 4519 9458 4528
rect 9416 4282 9444 4519
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9508 3942 9536 4644
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9508 3534 9536 3878
rect 9496 3528 9548 3534
rect 9692 3505 9720 4762
rect 9784 4622 9812 6695
rect 9851 6012 10159 6021
rect 9851 6010 9857 6012
rect 9913 6010 9937 6012
rect 9993 6010 10017 6012
rect 10073 6010 10097 6012
rect 10153 6010 10159 6012
rect 9913 5958 9915 6010
rect 10095 5958 10097 6010
rect 9851 5956 9857 5958
rect 9913 5956 9937 5958
rect 9993 5956 10017 5958
rect 10073 5956 10097 5958
rect 10153 5956 10159 5958
rect 9851 5947 10159 5956
rect 10244 5710 10272 8774
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10152 5166 10180 5510
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 9851 4924 10159 4933
rect 9851 4922 9857 4924
rect 9913 4922 9937 4924
rect 9993 4922 10017 4924
rect 10073 4922 10097 4924
rect 10153 4922 10159 4924
rect 9913 4870 9915 4922
rect 10095 4870 10097 4922
rect 9851 4868 9857 4870
rect 9913 4868 9937 4870
rect 9993 4868 10017 4870
rect 10073 4868 10097 4870
rect 10153 4868 10159 4870
rect 9851 4859 10159 4868
rect 10048 4752 10100 4758
rect 10046 4720 10048 4729
rect 10100 4720 10102 4729
rect 10046 4655 10102 4664
rect 10140 4684 10192 4690
rect 10244 4672 10272 5510
rect 10192 4644 10272 4672
rect 10140 4626 10192 4632
rect 10336 4622 10364 9646
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10428 6866 10456 8910
rect 10520 8634 10548 8910
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10428 6322 10456 6802
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10520 6458 10548 6734
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10414 6080 10470 6089
rect 10414 6015 10470 6024
rect 10428 5166 10456 6015
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10520 4622 10548 5578
rect 10612 5234 10640 8570
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9784 3602 9812 3946
rect 9851 3836 10159 3845
rect 9851 3834 9857 3836
rect 9913 3834 9937 3836
rect 9993 3834 10017 3836
rect 10073 3834 10097 3836
rect 10153 3834 10159 3836
rect 9913 3782 9915 3834
rect 10095 3782 10097 3834
rect 9851 3780 9857 3782
rect 9913 3780 9937 3782
rect 9993 3780 10017 3782
rect 10073 3780 10097 3782
rect 10153 3780 10159 3782
rect 9851 3771 10159 3780
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9496 3470 9548 3476
rect 9678 3496 9734 3505
rect 9678 3431 9734 3440
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9416 2961 9444 2994
rect 9402 2952 9458 2961
rect 9312 2916 9364 2922
rect 9402 2887 9458 2896
rect 9312 2858 9364 2864
rect 9140 2746 9352 2774
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9036 1556 9088 1562
rect 9036 1498 9088 1504
rect 9140 1465 9168 2382
rect 9126 1456 9182 1465
rect 9126 1391 9182 1400
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 8944 1216 8996 1222
rect 8944 1158 8996 1164
rect 8956 950 8984 1158
rect 8944 944 8996 950
rect 8944 886 8996 892
rect 9048 746 9076 1294
rect 9036 740 9088 746
rect 9036 682 9088 688
rect 9036 536 9088 542
rect 9036 478 9088 484
rect 9048 160 9076 478
rect 9324 160 9352 2746
rect 9402 2680 9458 2689
rect 9402 2615 9404 2624
rect 9456 2615 9458 2624
rect 9784 2632 9812 3538
rect 10138 3496 10194 3505
rect 10138 3431 10194 3440
rect 10152 3126 10180 3431
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10244 3126 10272 3334
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 9851 2748 10159 2757
rect 9851 2746 9857 2748
rect 9913 2746 9937 2748
rect 9993 2746 10017 2748
rect 10073 2746 10097 2748
rect 10153 2746 10159 2748
rect 9913 2694 9915 2746
rect 10095 2694 10097 2746
rect 9851 2692 9857 2694
rect 9913 2692 9937 2694
rect 9993 2692 10017 2694
rect 10073 2692 10097 2694
rect 10153 2692 10159 2694
rect 9851 2683 10159 2692
rect 9784 2604 9904 2632
rect 9404 2586 9456 2592
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9770 2544 9826 2553
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9404 1964 9456 1970
rect 9404 1906 9456 1912
rect 9416 1737 9444 1906
rect 9402 1728 9458 1737
rect 9402 1663 9458 1672
rect 9600 1358 9628 2246
rect 9692 1358 9720 2518
rect 9770 2479 9826 2488
rect 9784 2446 9812 2479
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9876 2106 9904 2604
rect 10138 2408 10194 2417
rect 10138 2343 10194 2352
rect 9864 2100 9916 2106
rect 9864 2042 9916 2048
rect 10152 1748 10180 2343
rect 10244 2106 10272 2926
rect 10232 2100 10284 2106
rect 10232 2042 10284 2048
rect 10336 2038 10364 4558
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10324 2032 10376 2038
rect 10324 1974 10376 1980
rect 10428 1970 10456 3062
rect 10704 2632 10732 16487
rect 10796 14074 10824 20538
rect 10888 16522 10916 21984
rect 10980 20466 11008 22052
rect 11072 21486 11100 22102
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 11164 21010 11192 22528
rect 11336 22500 11388 22506
rect 11336 22442 11388 22448
rect 11348 22094 11376 22442
rect 11256 22066 11376 22094
rect 11256 21457 11284 22066
rect 11242 21448 11298 21457
rect 11242 21383 11298 21392
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10980 20330 11008 20402
rect 11058 20360 11114 20369
rect 10968 20324 11020 20330
rect 11058 20295 11114 20304
rect 10968 20266 11020 20272
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 10980 18834 11008 19994
rect 11072 19786 11100 20295
rect 11164 19922 11192 20946
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11060 19780 11112 19786
rect 11060 19722 11112 19728
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 11164 19281 11192 19722
rect 11150 19272 11206 19281
rect 11150 19207 11206 19216
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 11072 18290 11100 18634
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 10980 18193 11008 18226
rect 10966 18184 11022 18193
rect 10966 18119 11022 18128
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10980 17202 11008 18022
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10980 17105 11008 17138
rect 10966 17096 11022 17105
rect 10966 17031 11022 17040
rect 10876 16516 10928 16522
rect 10876 16458 10928 16464
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11164 15706 11192 16050
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11256 15570 11284 21383
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11348 19922 11376 21082
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 11440 16250 11468 41386
rect 11612 39432 11664 39438
rect 11612 39374 11664 39380
rect 11520 38888 11572 38894
rect 11520 38830 11572 38836
rect 11532 32366 11560 38830
rect 11624 37126 11652 39374
rect 11704 38888 11756 38894
rect 11808 38865 11836 43114
rect 11900 42702 11928 44934
rect 12070 44840 12126 45000
rect 12346 44840 12402 45000
rect 12622 44840 12678 45000
rect 12898 44962 12954 45000
rect 12728 44934 12954 44962
rect 12084 43314 12112 44840
rect 12360 44146 12388 44840
rect 12360 44118 12480 44146
rect 12452 43382 12480 44118
rect 12636 43382 12664 44840
rect 12440 43376 12492 43382
rect 12440 43318 12492 43324
rect 12624 43376 12676 43382
rect 12624 43318 12676 43324
rect 12072 43308 12124 43314
rect 12072 43250 12124 43256
rect 12164 43308 12216 43314
rect 12164 43250 12216 43256
rect 11888 42696 11940 42702
rect 11888 42638 11940 42644
rect 12176 39642 12204 43250
rect 12256 43104 12308 43110
rect 12256 43046 12308 43052
rect 12268 42945 12296 43046
rect 12254 42936 12310 42945
rect 12254 42871 12310 42880
rect 12728 42702 12756 44934
rect 12898 44840 12954 44934
rect 13174 44840 13230 45000
rect 13450 44840 13506 45000
rect 13726 44840 13782 45000
rect 14002 44962 14058 45000
rect 14278 44962 14334 45000
rect 14554 44962 14610 45000
rect 14002 44934 14136 44962
rect 14002 44840 14058 44934
rect 12818 43548 13126 43557
rect 12818 43546 12824 43548
rect 12880 43546 12904 43548
rect 12960 43546 12984 43548
rect 13040 43546 13064 43548
rect 13120 43546 13126 43548
rect 12880 43494 12882 43546
rect 13062 43494 13064 43546
rect 12818 43492 12824 43494
rect 12880 43492 12904 43494
rect 12960 43492 12984 43494
rect 13040 43492 13064 43494
rect 13120 43492 13126 43494
rect 12818 43483 13126 43492
rect 13188 43450 13216 44840
rect 13176 43444 13228 43450
rect 13176 43386 13228 43392
rect 13464 43382 13492 44840
rect 13452 43376 13504 43382
rect 13452 43318 13504 43324
rect 13636 43240 13688 43246
rect 13636 43182 13688 43188
rect 13084 43172 13136 43178
rect 13084 43114 13136 43120
rect 12900 43104 12952 43110
rect 12898 43072 12900 43081
rect 13096 43081 13124 43114
rect 12952 43072 12954 43081
rect 12898 43007 12954 43016
rect 13082 43072 13138 43081
rect 13082 43007 13138 43016
rect 13648 42906 13676 43182
rect 13636 42900 13688 42906
rect 13636 42842 13688 42848
rect 13544 42764 13596 42770
rect 13740 42752 13768 44840
rect 13820 43104 13872 43110
rect 13820 43046 13872 43052
rect 13832 42945 13860 43046
rect 13818 42936 13874 42945
rect 13818 42871 13874 42880
rect 13820 42764 13872 42770
rect 13740 42724 13820 42752
rect 13544 42706 13596 42712
rect 13820 42706 13872 42712
rect 12348 42696 12400 42702
rect 12348 42638 12400 42644
rect 12716 42696 12768 42702
rect 12716 42638 12768 42644
rect 12360 41414 12388 42638
rect 13360 42628 13412 42634
rect 13360 42570 13412 42576
rect 12532 42560 12584 42566
rect 12532 42502 12584 42508
rect 13268 42560 13320 42566
rect 13268 42502 13320 42508
rect 12544 42362 12572 42502
rect 12818 42460 13126 42469
rect 12818 42458 12824 42460
rect 12880 42458 12904 42460
rect 12960 42458 12984 42460
rect 13040 42458 13064 42460
rect 13120 42458 13126 42460
rect 12880 42406 12882 42458
rect 13062 42406 13064 42458
rect 12818 42404 12824 42406
rect 12880 42404 12904 42406
rect 12960 42404 12984 42406
rect 13040 42404 13064 42406
rect 13120 42404 13126 42406
rect 12818 42395 13126 42404
rect 12532 42356 12584 42362
rect 12532 42298 12584 42304
rect 12530 41712 12586 41721
rect 12530 41647 12586 41656
rect 12268 41386 12388 41414
rect 12164 39636 12216 39642
rect 12164 39578 12216 39584
rect 12268 39098 12296 41386
rect 12440 40384 12492 40390
rect 12440 40326 12492 40332
rect 12256 39092 12308 39098
rect 12256 39034 12308 39040
rect 12452 38962 12480 40326
rect 12544 39846 12572 41647
rect 13280 41414 13308 42502
rect 13188 41386 13308 41414
rect 12818 41372 13126 41381
rect 12818 41370 12824 41372
rect 12880 41370 12904 41372
rect 12960 41370 12984 41372
rect 13040 41370 13064 41372
rect 13120 41370 13126 41372
rect 12880 41318 12882 41370
rect 13062 41318 13064 41370
rect 12818 41316 12824 41318
rect 12880 41316 12904 41318
rect 12960 41316 12984 41318
rect 13040 41316 13064 41318
rect 13120 41316 13126 41318
rect 12818 41307 13126 41316
rect 12818 40284 13126 40293
rect 12818 40282 12824 40284
rect 12880 40282 12904 40284
rect 12960 40282 12984 40284
rect 13040 40282 13064 40284
rect 13120 40282 13126 40284
rect 12880 40230 12882 40282
rect 13062 40230 13064 40282
rect 12818 40228 12824 40230
rect 12880 40228 12904 40230
rect 12960 40228 12984 40230
rect 13040 40228 13064 40230
rect 13120 40228 13126 40230
rect 12818 40219 13126 40228
rect 12532 39840 12584 39846
rect 12532 39782 12584 39788
rect 12532 39636 12584 39642
rect 12584 39596 12664 39624
rect 12532 39578 12584 39584
rect 12440 38956 12492 38962
rect 12492 38916 12572 38944
rect 12440 38898 12492 38904
rect 11704 38830 11756 38836
rect 11794 38856 11850 38865
rect 11716 38418 11744 38830
rect 11794 38791 11850 38800
rect 11796 38752 11848 38758
rect 11796 38694 11848 38700
rect 11704 38412 11756 38418
rect 11704 38354 11756 38360
rect 11612 37120 11664 37126
rect 11612 37062 11664 37068
rect 11808 35834 11836 38694
rect 12348 38412 12400 38418
rect 12348 38354 12400 38360
rect 12072 36576 12124 36582
rect 12072 36518 12124 36524
rect 11888 36100 11940 36106
rect 11888 36042 11940 36048
rect 11796 35828 11848 35834
rect 11796 35770 11848 35776
rect 11808 33386 11836 35770
rect 11900 34066 11928 36042
rect 12084 35698 12112 36518
rect 12256 36168 12308 36174
rect 12256 36110 12308 36116
rect 12164 36032 12216 36038
rect 12164 35974 12216 35980
rect 12176 35698 12204 35974
rect 12268 35698 12296 36110
rect 11980 35692 12032 35698
rect 11980 35634 12032 35640
rect 12072 35692 12124 35698
rect 12072 35634 12124 35640
rect 12164 35692 12216 35698
rect 12164 35634 12216 35640
rect 12256 35692 12308 35698
rect 12256 35634 12308 35640
rect 11992 35601 12020 35634
rect 11978 35592 12034 35601
rect 11978 35527 12034 35536
rect 12268 35170 12296 35634
rect 12072 35148 12124 35154
rect 12176 35142 12296 35170
rect 12360 35170 12388 38354
rect 12544 38214 12572 38916
rect 12636 38842 12664 39596
rect 12716 39296 12768 39302
rect 12716 39238 12768 39244
rect 12728 38962 12756 39238
rect 12818 39196 13126 39205
rect 12818 39194 12824 39196
rect 12880 39194 12904 39196
rect 12960 39194 12984 39196
rect 13040 39194 13064 39196
rect 13120 39194 13126 39196
rect 12880 39142 12882 39194
rect 13062 39142 13064 39194
rect 12818 39140 12824 39142
rect 12880 39140 12904 39142
rect 12960 39140 12984 39142
rect 13040 39140 13064 39142
rect 13120 39140 13126 39142
rect 12818 39131 13126 39140
rect 12716 38956 12768 38962
rect 12716 38898 12768 38904
rect 12636 38814 12756 38842
rect 12624 38752 12676 38758
rect 12624 38694 12676 38700
rect 12636 38554 12664 38694
rect 12624 38548 12676 38554
rect 12624 38490 12676 38496
rect 12440 38208 12492 38214
rect 12440 38150 12492 38156
rect 12532 38208 12584 38214
rect 12532 38150 12584 38156
rect 12452 37874 12480 38150
rect 12440 37868 12492 37874
rect 12440 37810 12492 37816
rect 12544 36582 12572 38150
rect 12728 37806 12756 38814
rect 13084 38344 13136 38350
rect 13084 38286 13136 38292
rect 13096 38214 13124 38286
rect 13084 38208 13136 38214
rect 13084 38150 13136 38156
rect 12818 38108 13126 38117
rect 12818 38106 12824 38108
rect 12880 38106 12904 38108
rect 12960 38106 12984 38108
rect 13040 38106 13064 38108
rect 13120 38106 13126 38108
rect 12880 38054 12882 38106
rect 13062 38054 13064 38106
rect 12818 38052 12824 38054
rect 12880 38052 12904 38054
rect 12960 38052 12984 38054
rect 13040 38052 13064 38054
rect 13120 38052 13126 38054
rect 12818 38043 13126 38052
rect 12716 37800 12768 37806
rect 12636 37748 12716 37754
rect 12636 37742 12768 37748
rect 12636 37726 12756 37742
rect 12636 37262 12664 37726
rect 12716 37664 12768 37670
rect 12716 37606 12768 37612
rect 12624 37256 12676 37262
rect 12624 37198 12676 37204
rect 12532 36576 12584 36582
rect 12532 36518 12584 36524
rect 12438 36272 12494 36281
rect 12438 36207 12494 36216
rect 12452 36174 12480 36207
rect 12440 36168 12492 36174
rect 12440 36110 12492 36116
rect 12360 35142 12572 35170
rect 12176 35136 12204 35142
rect 12124 35108 12204 35136
rect 12072 35090 12124 35096
rect 12084 34513 12112 35090
rect 12256 35080 12308 35086
rect 12176 35040 12256 35068
rect 12070 34504 12126 34513
rect 12070 34439 12126 34448
rect 11888 34060 11940 34066
rect 11940 34020 12020 34048
rect 11888 34002 11940 34008
rect 11796 33380 11848 33386
rect 11796 33322 11848 33328
rect 11992 33114 12020 34020
rect 11980 33108 12032 33114
rect 12032 33068 12112 33096
rect 11980 33050 12032 33056
rect 11702 33008 11758 33017
rect 11702 32943 11758 32952
rect 11520 32360 11572 32366
rect 11520 32302 11572 32308
rect 11716 30734 11744 32943
rect 11980 32836 12032 32842
rect 11980 32778 12032 32784
rect 11794 32464 11850 32473
rect 11794 32399 11850 32408
rect 11808 31686 11836 32399
rect 11886 32328 11942 32337
rect 11886 32263 11888 32272
rect 11940 32263 11942 32272
rect 11888 32234 11940 32240
rect 11886 31784 11942 31793
rect 11886 31719 11942 31728
rect 11796 31680 11848 31686
rect 11796 31622 11848 31628
rect 11900 31414 11928 31719
rect 11888 31408 11940 31414
rect 11888 31350 11940 31356
rect 11886 31240 11942 31249
rect 11886 31175 11942 31184
rect 11704 30728 11756 30734
rect 11704 30670 11756 30676
rect 11612 30592 11664 30598
rect 11612 30534 11664 30540
rect 11624 30433 11652 30534
rect 11610 30424 11666 30433
rect 11610 30359 11666 30368
rect 11520 30320 11572 30326
rect 11520 30262 11572 30268
rect 11610 30288 11666 30297
rect 11532 29850 11560 30262
rect 11610 30223 11666 30232
rect 11520 29844 11572 29850
rect 11520 29786 11572 29792
rect 11624 29646 11652 30223
rect 11900 29753 11928 31175
rect 11886 29744 11942 29753
rect 11886 29679 11942 29688
rect 11612 29640 11664 29646
rect 11612 29582 11664 29588
rect 11900 28994 11928 29679
rect 11992 29646 12020 32778
rect 12084 31940 12112 33068
rect 12176 32042 12204 35040
rect 12256 35022 12308 35028
rect 12360 33658 12388 35142
rect 12544 35034 12572 35142
rect 12544 35018 12664 35034
rect 12544 35012 12676 35018
rect 12544 35006 12624 35012
rect 12624 34954 12676 34960
rect 12728 33658 12756 37606
rect 12818 37020 13126 37029
rect 12818 37018 12824 37020
rect 12880 37018 12904 37020
rect 12960 37018 12984 37020
rect 13040 37018 13064 37020
rect 13120 37018 13126 37020
rect 12880 36966 12882 37018
rect 13062 36966 13064 37018
rect 12818 36964 12824 36966
rect 12880 36964 12904 36966
rect 12960 36964 12984 36966
rect 13040 36964 13064 36966
rect 13120 36964 13126 36966
rect 12818 36955 13126 36964
rect 12818 35932 13126 35941
rect 12818 35930 12824 35932
rect 12880 35930 12904 35932
rect 12960 35930 12984 35932
rect 13040 35930 13064 35932
rect 13120 35930 13126 35932
rect 12880 35878 12882 35930
rect 13062 35878 13064 35930
rect 12818 35876 12824 35878
rect 12880 35876 12904 35878
rect 12960 35876 12984 35878
rect 13040 35876 13064 35878
rect 13120 35876 13126 35878
rect 12818 35867 13126 35876
rect 12900 35760 12952 35766
rect 12900 35702 12952 35708
rect 12912 35018 12940 35702
rect 13084 35624 13136 35630
rect 13084 35566 13136 35572
rect 13096 35290 13124 35566
rect 13084 35284 13136 35290
rect 13084 35226 13136 35232
rect 12900 35012 12952 35018
rect 12900 34954 12952 34960
rect 12818 34844 13126 34853
rect 12818 34842 12824 34844
rect 12880 34842 12904 34844
rect 12960 34842 12984 34844
rect 13040 34842 13064 34844
rect 13120 34842 13126 34844
rect 12880 34790 12882 34842
rect 13062 34790 13064 34842
rect 12818 34788 12824 34790
rect 12880 34788 12904 34790
rect 12960 34788 12984 34790
rect 13040 34788 13064 34790
rect 13120 34788 13126 34790
rect 12818 34779 13126 34788
rect 13188 33946 13216 41386
rect 13268 39296 13320 39302
rect 13268 39238 13320 39244
rect 13280 38554 13308 39238
rect 13268 38548 13320 38554
rect 13268 38490 13320 38496
rect 13268 38344 13320 38350
rect 13268 38286 13320 38292
rect 13280 38010 13308 38286
rect 13268 38004 13320 38010
rect 13268 37946 13320 37952
rect 13188 33918 13308 33946
rect 13176 33856 13228 33862
rect 13176 33798 13228 33804
rect 12818 33756 13126 33765
rect 12818 33754 12824 33756
rect 12880 33754 12904 33756
rect 12960 33754 12984 33756
rect 13040 33754 13064 33756
rect 13120 33754 13126 33756
rect 12880 33702 12882 33754
rect 13062 33702 13064 33754
rect 12818 33700 12824 33702
rect 12880 33700 12904 33702
rect 12960 33700 12984 33702
rect 13040 33700 13064 33702
rect 13120 33700 13126 33702
rect 12818 33691 13126 33700
rect 12348 33652 12400 33658
rect 12348 33594 12400 33600
rect 12716 33652 12768 33658
rect 12716 33594 12768 33600
rect 13188 33454 13216 33798
rect 12624 33448 12676 33454
rect 12624 33390 12676 33396
rect 13176 33448 13228 33454
rect 13176 33390 13228 33396
rect 12256 33380 12308 33386
rect 12256 33322 12308 33328
rect 12268 33114 12296 33322
rect 12636 33318 12664 33390
rect 12624 33312 12676 33318
rect 12624 33254 12676 33260
rect 12256 33108 12308 33114
rect 12256 33050 12308 33056
rect 12532 32972 12584 32978
rect 12532 32914 12584 32920
rect 12176 32014 12388 32042
rect 12084 31912 12204 31940
rect 12072 31816 12124 31822
rect 12072 31758 12124 31764
rect 12084 31686 12112 31758
rect 12072 31680 12124 31686
rect 12072 31622 12124 31628
rect 12072 30252 12124 30258
rect 12072 30194 12124 30200
rect 12084 29850 12112 30194
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 11980 29640 12032 29646
rect 11980 29582 12032 29588
rect 12176 29073 12204 31912
rect 12256 31204 12308 31210
rect 12256 31146 12308 31152
rect 12268 30938 12296 31146
rect 12256 30932 12308 30938
rect 12256 30874 12308 30880
rect 12162 29064 12218 29073
rect 12162 28999 12218 29008
rect 12256 29028 12308 29034
rect 11716 28966 11928 28994
rect 11612 28620 11664 28626
rect 11612 28562 11664 28568
rect 11624 28082 11652 28562
rect 11520 28076 11572 28082
rect 11520 28018 11572 28024
rect 11612 28076 11664 28082
rect 11612 28018 11664 28024
rect 11532 27470 11560 28018
rect 11520 27464 11572 27470
rect 11520 27406 11572 27412
rect 11612 27464 11664 27470
rect 11612 27406 11664 27412
rect 11624 27130 11652 27406
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11612 26988 11664 26994
rect 11612 26930 11664 26936
rect 11520 26512 11572 26518
rect 11520 26454 11572 26460
rect 11532 26042 11560 26454
rect 11520 26036 11572 26042
rect 11520 25978 11572 25984
rect 11624 25514 11652 26930
rect 11532 25486 11652 25514
rect 11532 24818 11560 25486
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11624 24274 11652 25298
rect 11716 25242 11744 28966
rect 12176 28626 12204 28999
rect 12256 28970 12308 28976
rect 11888 28620 11940 28626
rect 11888 28562 11940 28568
rect 12164 28620 12216 28626
rect 12164 28562 12216 28568
rect 11796 28008 11848 28014
rect 11796 27950 11848 27956
rect 11808 27674 11836 27950
rect 11796 27668 11848 27674
rect 11796 27610 11848 27616
rect 11900 27538 11928 28562
rect 12268 27614 12296 28970
rect 12176 27586 12296 27614
rect 11888 27532 11940 27538
rect 11888 27474 11940 27480
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 11900 26382 11928 27270
rect 12072 26988 12124 26994
rect 12072 26930 12124 26936
rect 11978 26480 12034 26489
rect 11978 26415 12034 26424
rect 11888 26376 11940 26382
rect 11888 26318 11940 26324
rect 11900 25702 11928 26318
rect 11992 25906 12020 26415
rect 11980 25900 12032 25906
rect 11980 25842 12032 25848
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11900 25378 11928 25638
rect 12084 25498 12112 26930
rect 12176 26926 12204 27586
rect 12360 27334 12388 32014
rect 12544 31822 12572 32914
rect 13082 32872 13138 32881
rect 13082 32807 13084 32816
rect 13136 32807 13138 32816
rect 13084 32778 13136 32784
rect 12818 32668 13126 32677
rect 12818 32666 12824 32668
rect 12880 32666 12904 32668
rect 12960 32666 12984 32668
rect 13040 32666 13064 32668
rect 13120 32666 13126 32668
rect 12880 32614 12882 32666
rect 13062 32614 13064 32666
rect 12818 32612 12824 32614
rect 12880 32612 12904 32614
rect 12960 32612 12984 32614
rect 13040 32612 13064 32614
rect 13120 32612 13126 32614
rect 12818 32603 13126 32612
rect 13280 32502 13308 33918
rect 13268 32496 13320 32502
rect 13268 32438 13320 32444
rect 13176 31884 13228 31890
rect 13176 31826 13228 31832
rect 12532 31816 12584 31822
rect 12532 31758 12584 31764
rect 12440 31272 12492 31278
rect 12440 31214 12492 31220
rect 12452 30938 12480 31214
rect 12440 30932 12492 30938
rect 12440 30874 12492 30880
rect 12544 30802 12572 31758
rect 12716 31748 12768 31754
rect 12716 31690 12768 31696
rect 12728 31482 12756 31690
rect 12818 31580 13126 31589
rect 12818 31578 12824 31580
rect 12880 31578 12904 31580
rect 12960 31578 12984 31580
rect 13040 31578 13064 31580
rect 13120 31578 13126 31580
rect 12880 31526 12882 31578
rect 13062 31526 13064 31578
rect 12818 31524 12824 31526
rect 12880 31524 12904 31526
rect 12960 31524 12984 31526
rect 13040 31524 13064 31526
rect 13120 31524 13126 31526
rect 12818 31515 13126 31524
rect 12716 31476 12768 31482
rect 12716 31418 12768 31424
rect 12900 31476 12952 31482
rect 12900 31418 12952 31424
rect 12912 31346 12940 31418
rect 12900 31340 12952 31346
rect 12900 31282 12952 31288
rect 13084 31340 13136 31346
rect 13188 31328 13216 31826
rect 13268 31680 13320 31686
rect 13268 31622 13320 31628
rect 13136 31300 13216 31328
rect 13084 31282 13136 31288
rect 13096 31249 13124 31282
rect 13280 31278 13308 31622
rect 13268 31272 13320 31278
rect 13082 31240 13138 31249
rect 13268 31214 13320 31220
rect 13082 31175 13138 31184
rect 12624 31136 12676 31142
rect 12624 31078 12676 31084
rect 12532 30796 12584 30802
rect 12532 30738 12584 30744
rect 12532 29776 12584 29782
rect 12532 29718 12584 29724
rect 12544 29170 12572 29718
rect 12532 29164 12584 29170
rect 12532 29106 12584 29112
rect 12636 28994 12664 31078
rect 12818 30492 13126 30501
rect 12818 30490 12824 30492
rect 12880 30490 12904 30492
rect 12960 30490 12984 30492
rect 13040 30490 13064 30492
rect 13120 30490 13126 30492
rect 12880 30438 12882 30490
rect 13062 30438 13064 30490
rect 12818 30436 12824 30438
rect 12880 30436 12904 30438
rect 12960 30436 12984 30438
rect 13040 30436 13064 30438
rect 13120 30436 13126 30438
rect 12818 30427 13126 30436
rect 12716 30048 12768 30054
rect 12716 29990 12768 29996
rect 12728 29646 12756 29990
rect 12716 29640 12768 29646
rect 12716 29582 12768 29588
rect 13174 29608 13230 29617
rect 13174 29543 13230 29552
rect 12818 29404 13126 29413
rect 12818 29402 12824 29404
rect 12880 29402 12904 29404
rect 12960 29402 12984 29404
rect 13040 29402 13064 29404
rect 13120 29402 13126 29404
rect 12880 29350 12882 29402
rect 13062 29350 13064 29402
rect 12818 29348 12824 29350
rect 12880 29348 12904 29350
rect 12960 29348 12984 29350
rect 13040 29348 13064 29350
rect 13120 29348 13126 29350
rect 12818 29339 13126 29348
rect 13188 29238 13216 29543
rect 13176 29232 13228 29238
rect 12990 29200 13046 29209
rect 13176 29174 13228 29180
rect 12990 29135 12992 29144
rect 13044 29135 13046 29144
rect 12992 29106 13044 29112
rect 12636 28966 12756 28994
rect 12530 28520 12586 28529
rect 12440 28484 12492 28490
rect 12530 28455 12586 28464
rect 12440 28426 12492 28432
rect 12452 28218 12480 28426
rect 12440 28212 12492 28218
rect 12440 28154 12492 28160
rect 12544 27470 12572 28455
rect 12728 28422 12756 28966
rect 12624 28416 12676 28422
rect 12624 28358 12676 28364
rect 12716 28416 12768 28422
rect 12716 28358 12768 28364
rect 13268 28416 13320 28422
rect 13268 28358 13320 28364
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 12348 27328 12400 27334
rect 12348 27270 12400 27276
rect 12440 27124 12492 27130
rect 12440 27066 12492 27072
rect 12346 27024 12402 27033
rect 12346 26959 12348 26968
rect 12400 26959 12402 26968
rect 12348 26930 12400 26936
rect 12164 26920 12216 26926
rect 12452 26874 12480 27066
rect 12164 26862 12216 26868
rect 12176 26382 12204 26862
rect 12360 26846 12480 26874
rect 12256 26784 12308 26790
rect 12256 26726 12308 26732
rect 12268 26450 12296 26726
rect 12256 26444 12308 26450
rect 12256 26386 12308 26392
rect 12164 26376 12216 26382
rect 12164 26318 12216 26324
rect 12072 25492 12124 25498
rect 12072 25434 12124 25440
rect 11900 25350 12112 25378
rect 11716 25214 11928 25242
rect 11612 24268 11664 24274
rect 11612 24210 11664 24216
rect 11704 24132 11756 24138
rect 11704 24074 11756 24080
rect 11716 23730 11744 24074
rect 11704 23724 11756 23730
rect 11624 23684 11704 23712
rect 11520 21956 11572 21962
rect 11520 21898 11572 21904
rect 11532 20602 11560 21898
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 11532 19378 11560 20198
rect 11624 20058 11652 23684
rect 11704 23666 11756 23672
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11610 19816 11666 19825
rect 11610 19751 11666 19760
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11518 17640 11574 17649
rect 11518 17575 11520 17584
rect 11572 17575 11574 17584
rect 11520 17546 11572 17552
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11440 15473 11468 15506
rect 11426 15464 11482 15473
rect 11426 15399 11482 15408
rect 11532 15162 11560 17546
rect 11520 15156 11572 15162
rect 11256 15116 11520 15144
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 10888 14346 10916 15030
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10796 13530 10824 13874
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10888 13394 10916 14282
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10796 11694 10824 13330
rect 10888 12442 10916 13330
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10612 2604 10732 2632
rect 10416 1964 10468 1970
rect 10416 1906 10468 1912
rect 10152 1720 10272 1748
rect 9851 1660 10159 1669
rect 9851 1658 9857 1660
rect 9913 1658 9937 1660
rect 9993 1658 10017 1660
rect 10073 1658 10097 1660
rect 10153 1658 10159 1660
rect 9913 1606 9915 1658
rect 10095 1606 10097 1658
rect 9851 1604 9857 1606
rect 9913 1604 9937 1606
rect 9993 1604 10017 1606
rect 10073 1604 10097 1606
rect 10153 1604 10159 1606
rect 9851 1595 10159 1604
rect 10244 1426 10272 1720
rect 10416 1556 10468 1562
rect 10416 1498 10468 1504
rect 10232 1420 10284 1426
rect 10232 1362 10284 1368
rect 9588 1352 9640 1358
rect 9588 1294 9640 1300
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 9772 1216 9824 1222
rect 9772 1158 9824 1164
rect 9680 740 9732 746
rect 9680 682 9732 688
rect 9588 604 9640 610
rect 9588 546 9640 552
rect 9600 160 9628 546
rect 9692 354 9720 682
rect 9784 490 9812 1158
rect 9784 462 9996 490
rect 9692 326 9904 354
rect 9876 160 9904 326
rect 7930 82 7986 160
rect 7760 54 7986 82
rect 7930 0 7986 54
rect 8206 0 8262 160
rect 8482 0 8538 160
rect 8758 0 8814 160
rect 9034 0 9090 160
rect 9310 0 9366 160
rect 9586 0 9642 160
rect 9862 0 9918 160
rect 9968 82 9996 462
rect 10428 160 10456 1498
rect 10612 1222 10640 2604
rect 10796 2417 10824 11494
rect 10888 10062 10916 12378
rect 10980 11762 11008 14758
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 11072 11642 11100 14350
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 10980 11614 11100 11642
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10888 8634 10916 9998
rect 10980 9586 11008 11614
rect 11164 11218 11192 14214
rect 11256 12084 11284 15116
rect 11520 15098 11572 15104
rect 11624 15042 11652 19751
rect 11716 19334 11744 23122
rect 11900 22642 11928 25214
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 11992 24274 12020 25094
rect 11980 24268 12032 24274
rect 11980 24210 12032 24216
rect 12084 23254 12112 25350
rect 12176 24750 12204 26318
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 12268 24954 12296 25230
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12164 24744 12216 24750
rect 12164 24686 12216 24692
rect 12072 23248 12124 23254
rect 12072 23190 12124 23196
rect 11888 22636 11940 22642
rect 11888 22578 11940 22584
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11900 22273 11928 22374
rect 11886 22264 11942 22273
rect 11992 22234 12020 22578
rect 11886 22199 11942 22208
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 12176 22114 12204 24686
rect 12256 24268 12308 24274
rect 12256 24210 12308 24216
rect 12268 23866 12296 24210
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12360 23730 12388 26846
rect 12440 26784 12492 26790
rect 12440 26726 12492 26732
rect 12452 26246 12480 26726
rect 12544 26489 12572 27406
rect 12530 26480 12586 26489
rect 12530 26415 12586 26424
rect 12440 26240 12492 26246
rect 12440 26182 12492 26188
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12544 25430 12572 26182
rect 12532 25424 12584 25430
rect 12532 25366 12584 25372
rect 12636 25158 12664 28358
rect 12818 28316 13126 28325
rect 12818 28314 12824 28316
rect 12880 28314 12904 28316
rect 12960 28314 12984 28316
rect 13040 28314 13064 28316
rect 13120 28314 13126 28316
rect 12880 28262 12882 28314
rect 13062 28262 13064 28314
rect 12818 28260 12824 28262
rect 12880 28260 12904 28262
rect 12960 28260 12984 28262
rect 13040 28260 13064 28262
rect 13120 28260 13126 28262
rect 12818 28251 13126 28260
rect 13176 27532 13228 27538
rect 13176 27474 13228 27480
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12452 24154 12480 25094
rect 12728 24392 12756 27270
rect 12818 27228 13126 27237
rect 12818 27226 12824 27228
rect 12880 27226 12904 27228
rect 12960 27226 12984 27228
rect 13040 27226 13064 27228
rect 13120 27226 13126 27228
rect 12880 27174 12882 27226
rect 13062 27174 13064 27226
rect 12818 27172 12824 27174
rect 12880 27172 12904 27174
rect 12960 27172 12984 27174
rect 13040 27172 13064 27174
rect 13120 27172 13126 27174
rect 12818 27163 13126 27172
rect 13188 26874 13216 27474
rect 13096 26846 13216 26874
rect 13096 26586 13124 26846
rect 13176 26784 13228 26790
rect 13176 26726 13228 26732
rect 13188 26586 13216 26726
rect 13084 26580 13136 26586
rect 13084 26522 13136 26528
rect 13176 26580 13228 26586
rect 13176 26522 13228 26528
rect 12818 26140 13126 26149
rect 12818 26138 12824 26140
rect 12880 26138 12904 26140
rect 12960 26138 12984 26140
rect 13040 26138 13064 26140
rect 13120 26138 13126 26140
rect 12880 26086 12882 26138
rect 13062 26086 13064 26138
rect 12818 26084 12824 26086
rect 12880 26084 12904 26086
rect 12960 26084 12984 26086
rect 13040 26084 13064 26086
rect 13120 26084 13126 26086
rect 12818 26075 13126 26084
rect 13280 25702 13308 28358
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 12900 25288 12952 25294
rect 12900 25230 12952 25236
rect 13084 25288 13136 25294
rect 13136 25236 13216 25242
rect 13084 25230 13216 25236
rect 12912 25158 12940 25230
rect 13096 25214 13216 25230
rect 12900 25152 12952 25158
rect 12900 25094 12952 25100
rect 12818 25052 13126 25061
rect 12818 25050 12824 25052
rect 12880 25050 12904 25052
rect 12960 25050 12984 25052
rect 13040 25050 13064 25052
rect 13120 25050 13126 25052
rect 12880 24998 12882 25050
rect 13062 24998 13064 25050
rect 12818 24996 12824 24998
rect 12880 24996 12904 24998
rect 12960 24996 12984 24998
rect 13040 24996 13064 24998
rect 13120 24996 13126 24998
rect 12818 24987 13126 24996
rect 13188 24954 13216 25214
rect 13176 24948 13228 24954
rect 13176 24890 13228 24896
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12728 24364 12940 24392
rect 12808 24200 12860 24206
rect 12452 24126 12664 24154
rect 12912 24188 12940 24364
rect 13004 24274 13032 24550
rect 12992 24268 13044 24274
rect 12992 24210 13044 24216
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 12860 24160 12940 24188
rect 12808 24142 12860 24148
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 12532 23248 12584 23254
rect 12532 23190 12584 23196
rect 12440 23044 12492 23050
rect 12440 22986 12492 22992
rect 11900 22086 12204 22114
rect 11900 20380 11928 22086
rect 12452 22030 12480 22986
rect 12440 22024 12492 22030
rect 12346 21992 12402 22001
rect 12440 21966 12492 21972
rect 12346 21927 12402 21936
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12176 21690 12204 21830
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12268 21010 12296 21830
rect 12360 21554 12388 21927
rect 12544 21876 12572 23190
rect 12452 21848 12572 21876
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 12452 21026 12480 21848
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12544 21146 12572 21286
rect 12532 21140 12584 21146
rect 12532 21082 12584 21088
rect 12530 21040 12586 21049
rect 12256 21004 12308 21010
rect 12452 20998 12530 21026
rect 12530 20975 12586 20984
rect 12256 20946 12308 20952
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12452 20602 12480 20878
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 11808 20352 11928 20380
rect 11808 19836 11836 20352
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 11992 20058 12020 20266
rect 12084 20058 12112 20538
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 11980 19848 12032 19854
rect 11808 19808 11928 19836
rect 11716 19306 11836 19334
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 16794 11744 17682
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11808 16454 11836 19306
rect 11900 18086 11928 19808
rect 11980 19790 12032 19796
rect 11992 19689 12020 19790
rect 12084 19718 12112 19994
rect 12072 19712 12124 19718
rect 11978 19680 12034 19689
rect 12072 19654 12124 19660
rect 11978 19615 12034 19624
rect 11992 19394 12020 19615
rect 12176 19514 12204 20334
rect 12544 20330 12572 20878
rect 12532 20324 12584 20330
rect 12532 20266 12584 20272
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12268 19514 12296 19790
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 11992 19366 12204 19394
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11992 18358 12020 18566
rect 11980 18352 12032 18358
rect 12084 18329 12112 18634
rect 11980 18294 12032 18300
rect 12070 18320 12126 18329
rect 12070 18255 12126 18264
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11992 17678 12020 18022
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11888 17604 11940 17610
rect 11888 17546 11940 17552
rect 11900 17338 11928 17546
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 12176 17218 12204 19366
rect 12532 19372 12584 19378
rect 12452 19320 12532 19334
rect 12452 19314 12584 19320
rect 12452 19306 12572 19314
rect 12452 18834 12480 19306
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12268 17678 12296 18226
rect 12452 18154 12480 18566
rect 12440 18148 12492 18154
rect 12440 18090 12492 18096
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 11980 17196 12032 17202
rect 12176 17190 12296 17218
rect 12032 17156 12112 17184
rect 11980 17138 12032 17144
rect 11980 16992 12032 16998
rect 11900 16952 11980 16980
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11440 15014 11652 15042
rect 11336 12096 11388 12102
rect 11256 12056 11336 12084
rect 11336 12038 11388 12044
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11164 9674 11192 11154
rect 11348 10742 11376 12038
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11336 9988 11388 9994
rect 11336 9930 11388 9936
rect 11060 9648 11112 9654
rect 11164 9646 11284 9674
rect 11060 9590 11112 9596
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10980 7410 11008 9522
rect 11072 8294 11100 9590
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 6934 11100 7142
rect 11164 7002 11192 8774
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 11256 6662 11284 9646
rect 11348 9518 11376 9930
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11072 6186 11100 6326
rect 11060 6180 11112 6186
rect 10980 6140 11060 6168
rect 10874 5944 10930 5953
rect 10874 5879 10930 5888
rect 10888 5778 10916 5879
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10980 4078 11008 6140
rect 11060 6122 11112 6128
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10980 3074 11008 4014
rect 11072 3534 11100 5578
rect 11164 4826 11192 6122
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11256 5817 11284 5850
rect 11242 5808 11298 5817
rect 11242 5743 11298 5752
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11164 3194 11192 3470
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 10980 3046 11100 3074
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10782 2408 10838 2417
rect 10782 2343 10838 2352
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10796 2122 10824 2246
rect 10704 2094 10824 2122
rect 10600 1216 10652 1222
rect 10600 1158 10652 1164
rect 10704 160 10732 2094
rect 10980 1986 11008 2926
rect 11072 2922 11100 3046
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 11256 2650 11284 5102
rect 11334 4720 11390 4729
rect 11334 4655 11390 4664
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 10796 1958 11008 1986
rect 10796 1290 10824 1958
rect 10968 1556 11020 1562
rect 11072 1544 11100 2586
rect 11348 2514 11376 4655
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11152 1828 11204 1834
rect 11152 1770 11204 1776
rect 11020 1516 11100 1544
rect 10968 1498 11020 1504
rect 11164 1442 11192 1770
rect 10980 1414 11192 1442
rect 11336 1420 11388 1426
rect 10784 1284 10836 1290
rect 10784 1226 10836 1232
rect 10980 160 11008 1414
rect 11336 1362 11388 1368
rect 11152 1284 11204 1290
rect 11152 1226 11204 1232
rect 10138 82 10194 160
rect 9968 54 10194 82
rect 10138 0 10194 54
rect 10414 0 10470 160
rect 10690 0 10746 160
rect 10966 0 11022 160
rect 11164 82 11192 1226
rect 11244 1216 11296 1222
rect 11244 1158 11296 1164
rect 11256 1018 11284 1158
rect 11244 1012 11296 1018
rect 11244 954 11296 960
rect 11348 950 11376 1362
rect 11336 944 11388 950
rect 11336 886 11388 892
rect 11440 406 11468 15014
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11716 14618 11744 14894
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11808 14414 11836 16390
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11520 13320 11572 13326
rect 11900 13274 11928 16952
rect 11980 16934 12032 16940
rect 12084 16794 12112 17156
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 11980 15496 12032 15502
rect 11978 15464 11980 15473
rect 12084 15484 12112 16730
rect 12164 15496 12216 15502
rect 12032 15464 12034 15473
rect 12084 15456 12164 15484
rect 12164 15438 12216 15444
rect 11978 15399 12034 15408
rect 11992 15162 12020 15399
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 12084 15094 12112 15302
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11520 13262 11572 13268
rect 11532 12714 11560 13262
rect 11808 13246 11928 13274
rect 11808 13190 11836 13246
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11532 6798 11560 12650
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11624 10826 11652 12582
rect 11704 12232 11756 12238
rect 11900 12220 11928 13126
rect 11992 12238 12020 14962
rect 11756 12192 11928 12220
rect 11980 12232 12032 12238
rect 11704 12174 11756 12180
rect 11980 12174 12032 12180
rect 11624 10798 11744 10826
rect 11716 10792 11744 10798
rect 11796 10804 11848 10810
rect 11716 10764 11796 10792
rect 11796 10746 11848 10752
rect 11992 10742 12020 12174
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 10742 12112 10950
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 11624 9654 11652 10678
rect 11702 10160 11758 10169
rect 11702 10095 11758 10104
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11716 7886 11744 10095
rect 11794 10024 11850 10033
rect 11794 9959 11850 9968
rect 11808 9586 11836 9959
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11900 9518 11928 9862
rect 11992 9654 12020 10678
rect 12070 10160 12126 10169
rect 12176 10146 12204 15438
rect 12268 13258 12296 17190
rect 12360 13705 12388 18022
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12452 15162 12480 17478
rect 12544 16998 12572 18634
rect 12636 18290 12664 24126
rect 12818 23964 13126 23973
rect 12818 23962 12824 23964
rect 12880 23962 12904 23964
rect 12960 23962 12984 23964
rect 13040 23962 13064 23964
rect 13120 23962 13126 23964
rect 12880 23910 12882 23962
rect 13062 23910 13064 23962
rect 12818 23908 12824 23910
rect 12880 23908 12904 23910
rect 12960 23908 12984 23910
rect 13040 23908 13064 23910
rect 13120 23908 13126 23910
rect 12818 23899 13126 23908
rect 12818 22876 13126 22885
rect 12818 22874 12824 22876
rect 12880 22874 12904 22876
rect 12960 22874 12984 22876
rect 13040 22874 13064 22876
rect 13120 22874 13126 22876
rect 12880 22822 12882 22874
rect 13062 22822 13064 22874
rect 12818 22820 12824 22822
rect 12880 22820 12904 22822
rect 12960 22820 12984 22822
rect 13040 22820 13064 22822
rect 13120 22820 13126 22822
rect 12818 22811 13126 22820
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12728 22234 12756 22510
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12728 20262 12756 22170
rect 12818 21788 13126 21797
rect 12818 21786 12824 21788
rect 12880 21786 12904 21788
rect 12960 21786 12984 21788
rect 13040 21786 13064 21788
rect 13120 21786 13126 21788
rect 12880 21734 12882 21786
rect 13062 21734 13064 21786
rect 12818 21732 12824 21734
rect 12880 21732 12904 21734
rect 12960 21732 12984 21734
rect 13040 21732 13064 21734
rect 13120 21732 13126 21734
rect 12818 21723 13126 21732
rect 13188 21434 13216 24210
rect 13280 23526 13308 24754
rect 13268 23520 13320 23526
rect 13268 23462 13320 23468
rect 13372 23066 13400 42570
rect 13452 36576 13504 36582
rect 13452 36518 13504 36524
rect 13464 35834 13492 36518
rect 13452 35828 13504 35834
rect 13452 35770 13504 35776
rect 13452 35012 13504 35018
rect 13452 34954 13504 34960
rect 13464 34921 13492 34954
rect 13450 34912 13506 34921
rect 13450 34847 13506 34856
rect 13452 31340 13504 31346
rect 13452 31282 13504 31288
rect 13464 30938 13492 31282
rect 13452 30932 13504 30938
rect 13452 30874 13504 30880
rect 13452 30796 13504 30802
rect 13452 30738 13504 30744
rect 13464 29209 13492 30738
rect 13450 29200 13506 29209
rect 13450 29135 13506 29144
rect 13464 23866 13492 29135
rect 13556 27606 13584 42706
rect 14108 42702 14136 44934
rect 14278 44934 14412 44962
rect 14278 44840 14334 44934
rect 14280 43104 14332 43110
rect 14280 43046 14332 43052
rect 14292 42945 14320 43046
rect 14278 42936 14334 42945
rect 14278 42871 14334 42880
rect 14384 42702 14412 44934
rect 14554 44934 14780 44962
rect 14554 44840 14610 44934
rect 14752 43382 14780 44934
rect 14830 44840 14886 45000
rect 15106 44840 15162 45000
rect 15382 44840 15438 45000
rect 15658 44840 15714 45000
rect 15934 44840 15990 45000
rect 16210 44840 16266 45000
rect 16486 44840 16542 45000
rect 16762 44840 16818 45000
rect 17038 44840 17094 45000
rect 17224 44940 17276 44946
rect 17224 44882 17276 44888
rect 14844 43382 14872 44840
rect 14740 43376 14792 43382
rect 14740 43318 14792 43324
rect 14832 43376 14884 43382
rect 14832 43318 14884 43324
rect 14924 43172 14976 43178
rect 14924 43114 14976 43120
rect 14936 42945 14964 43114
rect 14922 42936 14978 42945
rect 14922 42871 14978 42880
rect 15120 42786 15148 44840
rect 15396 44146 15424 44840
rect 15396 44118 15608 44146
rect 15580 43382 15608 44118
rect 15672 43382 15700 44840
rect 15568 43376 15620 43382
rect 15568 43318 15620 43324
rect 15660 43376 15712 43382
rect 15660 43318 15712 43324
rect 15948 43330 15976 44840
rect 16224 44146 16252 44840
rect 16224 44118 16436 44146
rect 16408 43382 16436 44118
rect 16120 43376 16172 43382
rect 15948 43324 16120 43330
rect 15948 43318 16172 43324
rect 16396 43376 16448 43382
rect 16396 43318 16448 43324
rect 15948 43302 16160 43318
rect 15292 43172 15344 43178
rect 15292 43114 15344 43120
rect 16120 43172 16172 43178
rect 16120 43114 16172 43120
rect 15304 42945 15332 43114
rect 15660 43104 15712 43110
rect 15660 43046 15712 43052
rect 15290 42936 15346 42945
rect 15290 42871 15346 42880
rect 15120 42758 15240 42786
rect 14096 42696 14148 42702
rect 14096 42638 14148 42644
rect 14372 42696 14424 42702
rect 15108 42696 15160 42702
rect 14372 42638 14424 42644
rect 14936 42656 15108 42684
rect 14832 42560 14884 42566
rect 14752 42520 14832 42548
rect 13636 38752 13688 38758
rect 14280 38752 14332 38758
rect 13636 38694 13688 38700
rect 14094 38720 14150 38729
rect 13648 38418 13676 38694
rect 14280 38694 14332 38700
rect 14094 38655 14150 38664
rect 13636 38412 13688 38418
rect 13636 38354 13688 38360
rect 13820 37324 13872 37330
rect 13820 37266 13872 37272
rect 13636 37120 13688 37126
rect 13636 37062 13688 37068
rect 13648 35272 13676 37062
rect 13728 36576 13780 36582
rect 13728 36518 13780 36524
rect 13740 36174 13768 36518
rect 13728 36168 13780 36174
rect 13728 36110 13780 36116
rect 13728 35284 13780 35290
rect 13648 35244 13728 35272
rect 13728 35226 13780 35232
rect 13740 33998 13768 35226
rect 13728 33992 13780 33998
rect 13728 33934 13780 33940
rect 13728 33652 13780 33658
rect 13728 33594 13780 33600
rect 13636 32768 13688 32774
rect 13636 32710 13688 32716
rect 13648 32366 13676 32710
rect 13636 32360 13688 32366
rect 13636 32302 13688 32308
rect 13636 29572 13688 29578
rect 13636 29514 13688 29520
rect 13648 29306 13676 29514
rect 13636 29300 13688 29306
rect 13636 29242 13688 29248
rect 13740 29170 13768 33594
rect 13832 30802 13860 37266
rect 13912 35488 13964 35494
rect 13912 35430 13964 35436
rect 13924 31657 13952 35430
rect 14002 35048 14058 35057
rect 14002 34983 14058 34992
rect 14016 32910 14044 34983
rect 14108 34542 14136 38655
rect 14188 35488 14240 35494
rect 14188 35430 14240 35436
rect 14200 35018 14228 35430
rect 14188 35012 14240 35018
rect 14188 34954 14240 34960
rect 14096 34536 14148 34542
rect 14096 34478 14148 34484
rect 14108 34202 14136 34478
rect 14096 34196 14148 34202
rect 14096 34138 14148 34144
rect 14200 33504 14228 34954
rect 14108 33476 14228 33504
rect 14108 33114 14136 33476
rect 14188 33380 14240 33386
rect 14188 33322 14240 33328
rect 14096 33108 14148 33114
rect 14096 33050 14148 33056
rect 14004 32904 14056 32910
rect 14004 32846 14056 32852
rect 14004 32768 14056 32774
rect 14004 32710 14056 32716
rect 14016 32026 14044 32710
rect 14096 32496 14148 32502
rect 14096 32438 14148 32444
rect 14108 32026 14136 32438
rect 14004 32020 14056 32026
rect 14004 31962 14056 31968
rect 14096 32020 14148 32026
rect 14096 31962 14148 31968
rect 14200 31793 14228 33322
rect 14186 31784 14242 31793
rect 14186 31719 14242 31728
rect 14200 31686 14228 31719
rect 14188 31680 14240 31686
rect 13910 31648 13966 31657
rect 14188 31622 14240 31628
rect 13910 31583 13966 31592
rect 13912 31408 13964 31414
rect 13912 31350 13964 31356
rect 13820 30796 13872 30802
rect 13820 30738 13872 30744
rect 13924 30569 13952 31350
rect 14188 31272 14240 31278
rect 14188 31214 14240 31220
rect 13910 30560 13966 30569
rect 13910 30495 13966 30504
rect 14094 30424 14150 30433
rect 14094 30359 14150 30368
rect 14004 29640 14056 29646
rect 14004 29582 14056 29588
rect 14016 29209 14044 29582
rect 14002 29200 14058 29209
rect 13728 29164 13780 29170
rect 13728 29106 13780 29112
rect 13924 29158 14002 29186
rect 13924 29102 13952 29158
rect 14002 29135 14058 29144
rect 13912 29096 13964 29102
rect 13912 29038 13964 29044
rect 14004 29028 14056 29034
rect 14004 28970 14056 28976
rect 13912 28416 13964 28422
rect 13912 28358 13964 28364
rect 13818 27704 13874 27713
rect 13818 27639 13874 27648
rect 13544 27600 13596 27606
rect 13544 27542 13596 27548
rect 13636 26988 13688 26994
rect 13636 26930 13688 26936
rect 13728 26988 13780 26994
rect 13728 26930 13780 26936
rect 13544 26920 13596 26926
rect 13544 26862 13596 26868
rect 13556 26450 13584 26862
rect 13544 26444 13596 26450
rect 13544 26386 13596 26392
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13280 23038 13400 23066
rect 13280 22778 13308 23038
rect 13360 22976 13412 22982
rect 13360 22918 13412 22924
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13266 21720 13322 21729
rect 13266 21655 13322 21664
rect 13280 21554 13308 21655
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13188 21406 13308 21434
rect 12818 20700 13126 20709
rect 12818 20698 12824 20700
rect 12880 20698 12904 20700
rect 12960 20698 12984 20700
rect 13040 20698 13064 20700
rect 13120 20698 13126 20700
rect 12880 20646 12882 20698
rect 13062 20646 13064 20698
rect 12818 20644 12824 20646
rect 12880 20644 12904 20646
rect 12960 20644 12984 20646
rect 13040 20644 13064 20646
rect 13120 20644 13126 20646
rect 12818 20635 13126 20644
rect 12898 20496 12954 20505
rect 12820 20454 12898 20482
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12820 19802 12848 20454
rect 12898 20431 12954 20440
rect 12728 19774 12848 19802
rect 12728 19378 12756 19774
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 12818 19612 13126 19621
rect 12818 19610 12824 19612
rect 12880 19610 12904 19612
rect 12960 19610 12984 19612
rect 13040 19610 13064 19612
rect 13120 19610 13126 19612
rect 12880 19558 12882 19610
rect 13062 19558 13064 19610
rect 12818 19556 12824 19558
rect 12880 19556 12904 19558
rect 12960 19556 12984 19558
rect 13040 19556 13064 19558
rect 13120 19556 13126 19558
rect 12818 19547 13126 19556
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12346 13696 12402 13705
rect 12346 13631 12402 13640
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12346 12336 12402 12345
rect 12346 12271 12402 12280
rect 12360 11830 12388 12271
rect 12452 12102 12480 15098
rect 12544 13326 12572 16526
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12452 11830 12480 12038
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12440 11280 12492 11286
rect 12360 11240 12440 11268
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12268 10266 12296 10746
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12126 10118 12204 10146
rect 12070 10095 12126 10104
rect 12360 10062 12388 11240
rect 12440 11222 12492 11228
rect 12544 10418 12572 13262
rect 12636 13190 12664 17070
rect 12728 15473 12756 19314
rect 12912 18698 12940 19450
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 13004 18698 13032 19382
rect 12900 18692 12952 18698
rect 12900 18634 12952 18640
rect 12992 18692 13044 18698
rect 12992 18634 13044 18640
rect 12818 18524 13126 18533
rect 12818 18522 12824 18524
rect 12880 18522 12904 18524
rect 12960 18522 12984 18524
rect 13040 18522 13064 18524
rect 13120 18522 13126 18524
rect 12880 18470 12882 18522
rect 13062 18470 13064 18522
rect 12818 18468 12824 18470
rect 12880 18468 12904 18470
rect 12960 18468 12984 18470
rect 13040 18468 13064 18470
rect 13120 18468 13126 18470
rect 12818 18459 13126 18468
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 12912 17882 12940 18294
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12818 17436 13126 17445
rect 12818 17434 12824 17436
rect 12880 17434 12904 17436
rect 12960 17434 12984 17436
rect 13040 17434 13064 17436
rect 13120 17434 13126 17436
rect 12880 17382 12882 17434
rect 13062 17382 13064 17434
rect 12818 17380 12824 17382
rect 12880 17380 12904 17382
rect 12960 17380 12984 17382
rect 13040 17380 13064 17382
rect 13120 17380 13126 17382
rect 12818 17371 13126 17380
rect 12818 16348 13126 16357
rect 12818 16346 12824 16348
rect 12880 16346 12904 16348
rect 12960 16346 12984 16348
rect 13040 16346 13064 16348
rect 13120 16346 13126 16348
rect 12880 16294 12882 16346
rect 13062 16294 13064 16346
rect 12818 16292 12824 16294
rect 12880 16292 12904 16294
rect 12960 16292 12984 16294
rect 13040 16292 13064 16294
rect 13120 16292 13126 16294
rect 12818 16283 13126 16292
rect 12714 15464 12770 15473
rect 12714 15399 12770 15408
rect 12818 15260 13126 15269
rect 12818 15258 12824 15260
rect 12880 15258 12904 15260
rect 12960 15258 12984 15260
rect 13040 15258 13064 15260
rect 13120 15258 13126 15260
rect 12880 15206 12882 15258
rect 13062 15206 13064 15258
rect 12818 15204 12824 15206
rect 12880 15204 12904 15206
rect 12960 15204 12984 15206
rect 13040 15204 13064 15206
rect 13120 15204 13126 15206
rect 12818 15195 13126 15204
rect 13188 15178 13216 19654
rect 13280 15450 13308 21406
rect 13372 18068 13400 22918
rect 13464 19334 13492 23802
rect 13648 23730 13676 26930
rect 13740 25362 13768 26930
rect 13728 25356 13780 25362
rect 13728 25298 13780 25304
rect 13740 24206 13768 25298
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13636 23724 13688 23730
rect 13556 23684 13636 23712
rect 13556 23186 13584 23684
rect 13636 23666 13688 23672
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13556 21622 13584 21830
rect 13544 21616 13596 21622
rect 13544 21558 13596 21564
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 13556 19446 13584 20334
rect 13648 19786 13676 23462
rect 13832 22778 13860 27639
rect 13924 26926 13952 28358
rect 13912 26920 13964 26926
rect 13912 26862 13964 26868
rect 14016 26586 14044 28970
rect 14004 26580 14056 26586
rect 14004 26522 14056 26528
rect 13910 24168 13966 24177
rect 13910 24103 13966 24112
rect 13924 23186 13952 24103
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 13820 22772 13872 22778
rect 13872 22732 13952 22760
rect 13820 22714 13872 22720
rect 13728 22432 13780 22438
rect 13728 22374 13780 22380
rect 13740 21486 13768 22374
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13832 21554 13860 21830
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13464 19306 13584 19334
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13464 18222 13492 18566
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 13372 18040 13492 18068
rect 13358 17776 13414 17785
rect 13358 17711 13414 17720
rect 13372 16658 13400 17711
rect 13464 17610 13492 18040
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13556 17338 13584 19306
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 13452 16788 13504 16794
rect 13556 16776 13584 17274
rect 13648 17134 13676 19722
rect 13726 19544 13782 19553
rect 13726 19479 13782 19488
rect 13740 19446 13768 19479
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13740 18426 13768 18634
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13728 18284 13780 18290
rect 13832 18272 13860 19790
rect 13780 18244 13860 18272
rect 13728 18226 13780 18232
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13504 16748 13584 16776
rect 13452 16730 13504 16736
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13452 16584 13504 16590
rect 13358 16552 13414 16561
rect 13452 16526 13504 16532
rect 13358 16487 13414 16496
rect 13372 16182 13400 16487
rect 13464 16454 13492 16526
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 13372 15638 13400 16118
rect 13556 16114 13584 16390
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13648 16046 13676 16390
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 13280 15422 13584 15450
rect 13360 15360 13412 15366
rect 13412 15320 13492 15348
rect 13360 15302 13412 15308
rect 13188 15150 13400 15178
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12728 13870 12756 14418
rect 12818 14172 13126 14181
rect 12818 14170 12824 14172
rect 12880 14170 12904 14172
rect 12960 14170 12984 14172
rect 13040 14170 13064 14172
rect 13120 14170 13126 14172
rect 12880 14118 12882 14170
rect 13062 14118 13064 14170
rect 12818 14116 12824 14118
rect 12880 14116 12904 14118
rect 12960 14116 12984 14118
rect 13040 14116 13064 14118
rect 13120 14116 13126 14118
rect 12818 14107 13126 14116
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12728 13530 12756 13806
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12636 12442 12664 13126
rect 12818 13084 13126 13093
rect 12818 13082 12824 13084
rect 12880 13082 12904 13084
rect 12960 13082 12984 13084
rect 13040 13082 13064 13084
rect 13120 13082 13126 13084
rect 12880 13030 12882 13082
rect 13062 13030 13064 13082
rect 12818 13028 12824 13030
rect 12880 13028 12904 13030
rect 12960 13028 12984 13030
rect 13040 13028 13064 13030
rect 13120 13028 13126 13030
rect 12818 13019 13126 13028
rect 13084 12708 13136 12714
rect 13084 12650 13136 12656
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 13096 12306 13124 12650
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13188 12238 13216 14962
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13280 12782 13308 13126
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 12728 10742 12756 12174
rect 12818 11996 13126 12005
rect 12818 11994 12824 11996
rect 12880 11994 12904 11996
rect 12960 11994 12984 11996
rect 13040 11994 13064 11996
rect 13120 11994 13126 11996
rect 12880 11942 12882 11994
rect 13062 11942 13064 11994
rect 12818 11940 12824 11942
rect 12880 11940 12904 11942
rect 12960 11940 12984 11942
rect 13040 11940 13064 11942
rect 13120 11940 13126 11942
rect 12818 11931 13126 11940
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 13096 11218 13124 11562
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12818 10908 13126 10917
rect 12818 10906 12824 10908
rect 12880 10906 12904 10908
rect 12960 10906 12984 10908
rect 13040 10906 13064 10908
rect 13120 10906 13126 10908
rect 12880 10854 12882 10906
rect 13062 10854 13064 10906
rect 12818 10852 12824 10854
rect 12880 10852 12904 10854
rect 12960 10852 12984 10854
rect 13040 10852 13064 10854
rect 13120 10852 13126 10854
rect 12818 10843 13126 10852
rect 13188 10742 13216 11766
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 12452 10390 12572 10418
rect 12452 10266 12480 10390
rect 12728 10282 12756 10678
rect 12806 10432 12862 10441
rect 12806 10367 12862 10376
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12544 10254 12756 10282
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 12084 8974 12112 9862
rect 12544 9586 12572 10254
rect 12820 10180 12848 10367
rect 12636 10152 12848 10180
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12268 9178 12296 9522
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12176 9081 12204 9114
rect 12162 9072 12218 9081
rect 12162 9007 12218 9016
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 12072 8968 12124 8974
rect 12360 8922 12388 9522
rect 12072 8910 12124 8916
rect 11900 8634 11928 8910
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11716 6798 11744 7686
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11532 6304 11560 6734
rect 11612 6316 11664 6322
rect 11532 6276 11612 6304
rect 11612 6258 11664 6264
rect 11808 6254 11836 7890
rect 11900 7410 11928 8570
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11886 6896 11942 6905
rect 11886 6831 11942 6840
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11900 5710 11928 6831
rect 12084 5846 12112 8910
rect 12268 8894 12388 8922
rect 12268 8566 12296 8894
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8566 12480 8774
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12360 8242 12388 8434
rect 12360 8214 12480 8242
rect 12348 6792 12400 6798
rect 12254 6760 12310 6769
rect 12310 6740 12348 6746
rect 12310 6734 12400 6740
rect 12310 6718 12388 6734
rect 12254 6695 12310 6704
rect 12452 6662 12480 8214
rect 12544 7478 12572 9522
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12544 6730 12572 6870
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 12268 5778 12296 6598
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11888 5704 11940 5710
rect 12360 5681 12388 6598
rect 12440 6316 12492 6322
rect 12544 6304 12572 6666
rect 12492 6276 12572 6304
rect 12440 6258 12492 6264
rect 11888 5646 11940 5652
rect 12346 5672 12402 5681
rect 11624 4690 11652 5646
rect 12346 5607 12402 5616
rect 12636 5522 12664 10152
rect 12818 9820 13126 9829
rect 12818 9818 12824 9820
rect 12880 9818 12904 9820
rect 12960 9818 12984 9820
rect 13040 9818 13064 9820
rect 13120 9818 13126 9820
rect 12880 9766 12882 9818
rect 13062 9766 13064 9818
rect 12818 9764 12824 9766
rect 12880 9764 12904 9766
rect 12960 9764 12984 9766
rect 13040 9764 13064 9766
rect 13120 9764 13126 9766
rect 12818 9755 13126 9764
rect 13188 9674 13216 10678
rect 12820 9654 13216 9674
rect 12808 9648 13216 9654
rect 12728 9608 12808 9636
rect 12728 6440 12756 9608
rect 12860 9646 13216 9648
rect 12808 9590 12860 9596
rect 12818 8732 13126 8741
rect 12818 8730 12824 8732
rect 12880 8730 12904 8732
rect 12960 8730 12984 8732
rect 13040 8730 13064 8732
rect 13120 8730 13126 8732
rect 12880 8678 12882 8730
rect 13062 8678 13064 8730
rect 12818 8676 12824 8678
rect 12880 8676 12904 8678
rect 12960 8676 12984 8678
rect 13040 8676 13064 8678
rect 13120 8676 13126 8678
rect 12818 8667 13126 8676
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 13004 7818 13032 8366
rect 12992 7812 13044 7818
rect 12992 7754 13044 7760
rect 12818 7644 13126 7653
rect 12818 7642 12824 7644
rect 12880 7642 12904 7644
rect 12960 7642 12984 7644
rect 13040 7642 13064 7644
rect 13120 7642 13126 7644
rect 12880 7590 12882 7642
rect 13062 7590 13064 7642
rect 12818 7588 12824 7590
rect 12880 7588 12904 7590
rect 12960 7588 12984 7590
rect 13040 7588 13064 7590
rect 13120 7588 13126 7590
rect 12818 7579 13126 7588
rect 12818 6556 13126 6565
rect 12818 6554 12824 6556
rect 12880 6554 12904 6556
rect 12960 6554 12984 6556
rect 13040 6554 13064 6556
rect 13120 6554 13126 6556
rect 12880 6502 12882 6554
rect 13062 6502 13064 6554
rect 12818 6500 12824 6502
rect 12880 6500 12904 6502
rect 12960 6500 12984 6502
rect 13040 6500 13064 6502
rect 13120 6500 13126 6502
rect 12818 6491 13126 6500
rect 12728 6412 12848 6440
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12728 5914 12756 6190
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12820 5794 12848 6412
rect 12452 5494 12664 5522
rect 12728 5766 12848 5794
rect 12256 5160 12308 5166
rect 12308 5120 12388 5148
rect 12256 5102 12308 5108
rect 12360 4758 12388 5120
rect 12348 4752 12400 4758
rect 12346 4720 12348 4729
rect 12400 4720 12402 4729
rect 11612 4684 11664 4690
rect 12346 4655 12402 4664
rect 11612 4626 11664 4632
rect 11624 4010 11652 4626
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12164 4276 12216 4282
rect 11992 4236 12164 4264
rect 11612 4004 11664 4010
rect 11612 3946 11664 3952
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11532 3194 11560 3334
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11624 3126 11652 3946
rect 11992 3534 12020 4236
rect 12164 4218 12216 4224
rect 12360 4078 12388 4422
rect 12348 4072 12400 4078
rect 12162 4040 12218 4049
rect 12348 4014 12400 4020
rect 12162 3975 12218 3984
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 11612 3120 11664 3126
rect 11808 3097 11836 3402
rect 12084 3126 12112 3878
rect 12072 3120 12124 3126
rect 11612 3062 11664 3068
rect 11794 3088 11850 3097
rect 12072 3062 12124 3068
rect 12176 3058 12204 3975
rect 11794 3023 11850 3032
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 11796 2848 11848 2854
rect 11532 2796 11796 2802
rect 11532 2790 11848 2796
rect 11532 2774 11836 2790
rect 11532 2378 11560 2774
rect 11978 2680 12034 2689
rect 11978 2615 12034 2624
rect 11992 2446 12020 2615
rect 12452 2446 12480 5494
rect 12622 5400 12678 5409
rect 12622 5335 12678 5344
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12544 4622 12572 5238
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12636 4468 12664 5335
rect 12728 4826 12756 5766
rect 12818 5468 13126 5477
rect 12818 5466 12824 5468
rect 12880 5466 12904 5468
rect 12960 5466 12984 5468
rect 13040 5466 13064 5468
rect 13120 5466 13126 5468
rect 12880 5414 12882 5466
rect 13062 5414 13064 5466
rect 12818 5412 12824 5414
rect 12880 5412 12904 5414
rect 12960 5412 12984 5414
rect 13040 5412 13064 5414
rect 13120 5412 13126 5414
rect 12818 5403 13126 5412
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12716 4480 12768 4486
rect 12636 4440 12716 4468
rect 12716 4422 12768 4428
rect 12818 4380 13126 4389
rect 12818 4378 12824 4380
rect 12880 4378 12904 4380
rect 12960 4378 12984 4380
rect 13040 4378 13064 4380
rect 13120 4378 13126 4380
rect 12880 4326 12882 4378
rect 13062 4326 13064 4378
rect 12818 4324 12824 4326
rect 12880 4324 12904 4326
rect 12960 4324 12984 4326
rect 13040 4324 13064 4326
rect 13120 4324 13126 4326
rect 12818 4315 13126 4324
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12622 4176 12678 4185
rect 12544 3194 12572 4150
rect 12622 4111 12624 4120
rect 12676 4111 12678 4120
rect 12624 4082 12676 4088
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12728 3040 12756 3538
rect 12818 3292 13126 3301
rect 12818 3290 12824 3292
rect 12880 3290 12904 3292
rect 12960 3290 12984 3292
rect 13040 3290 13064 3292
rect 13120 3290 13126 3292
rect 12880 3238 12882 3290
rect 13062 3238 13064 3290
rect 12818 3236 12824 3238
rect 12880 3236 12904 3238
rect 12960 3236 12984 3238
rect 13040 3236 13064 3238
rect 13120 3236 13126 3238
rect 12818 3227 13126 3236
rect 12900 3052 12952 3058
rect 12728 3012 12900 3040
rect 12900 2994 12952 3000
rect 12912 2446 12940 2994
rect 13188 2774 13216 8502
rect 13280 7478 13308 12378
rect 13268 7472 13320 7478
rect 13268 7414 13320 7420
rect 13266 6216 13322 6225
rect 13266 6151 13322 6160
rect 13280 5710 13308 6151
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13266 5400 13322 5409
rect 13266 5335 13322 5344
rect 13280 3670 13308 5335
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13372 2774 13400 15150
rect 13464 11558 13492 15320
rect 13556 15162 13584 15422
rect 13544 15156 13596 15162
rect 13596 15116 13676 15144
rect 13544 15098 13596 15104
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13556 12850 13584 14010
rect 13648 12850 13676 15116
rect 13832 14278 13860 16934
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13740 12866 13768 13670
rect 13740 12850 13860 12866
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13636 12844 13688 12850
rect 13740 12844 13872 12850
rect 13740 12838 13820 12844
rect 13636 12786 13688 12792
rect 13820 12786 13872 12792
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13556 10810 13584 12786
rect 13648 12753 13676 12786
rect 13634 12744 13690 12753
rect 13634 12679 13690 12688
rect 13924 12434 13952 22732
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 14016 20466 14044 21490
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14016 18290 14044 19110
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14108 17082 14136 30359
rect 14200 30190 14228 31214
rect 14188 30184 14240 30190
rect 14188 30126 14240 30132
rect 14200 29073 14228 30126
rect 14186 29064 14242 29073
rect 14186 28999 14242 29008
rect 14200 27470 14228 28999
rect 14188 27464 14240 27470
rect 14188 27406 14240 27412
rect 14188 26784 14240 26790
rect 14188 26726 14240 26732
rect 14200 24614 14228 26726
rect 14188 24608 14240 24614
rect 14186 24576 14188 24585
rect 14240 24576 14242 24585
rect 14186 24511 14242 24520
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14200 21690 14228 24142
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 14016 17054 14136 17082
rect 14016 13705 14044 17054
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 14002 13696 14058 13705
rect 14002 13631 14058 13640
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 13740 12406 13952 12434
rect 13636 11756 13688 11762
rect 13740 11744 13768 12406
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13688 11716 13768 11744
rect 13636 11698 13688 11704
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13648 10690 13676 11698
rect 13556 10662 13676 10690
rect 13728 10736 13780 10742
rect 13832 10724 13860 12038
rect 13924 10742 13952 12106
rect 14016 11762 14044 12718
rect 14108 12102 14136 16186
rect 14200 16182 14228 16934
rect 14188 16176 14240 16182
rect 14188 16118 14240 16124
rect 14292 15094 14320 38694
rect 14556 36372 14608 36378
rect 14556 36314 14608 36320
rect 14464 35488 14516 35494
rect 14464 35430 14516 35436
rect 14372 33380 14424 33386
rect 14372 33322 14424 33328
rect 14384 33046 14412 33322
rect 14372 33040 14424 33046
rect 14372 32982 14424 32988
rect 14372 32836 14424 32842
rect 14372 32778 14424 32784
rect 14384 32434 14412 32778
rect 14476 32502 14504 35430
rect 14464 32496 14516 32502
rect 14464 32438 14516 32444
rect 14372 32428 14424 32434
rect 14372 32370 14424 32376
rect 14384 31482 14412 32370
rect 14372 31476 14424 31482
rect 14372 31418 14424 31424
rect 14464 30796 14516 30802
rect 14464 30738 14516 30744
rect 14476 30122 14504 30738
rect 14464 30116 14516 30122
rect 14464 30058 14516 30064
rect 14370 30016 14426 30025
rect 14370 29951 14426 29960
rect 14384 29510 14412 29951
rect 14568 29578 14596 36314
rect 14648 33856 14700 33862
rect 14648 33798 14700 33804
rect 14660 33454 14688 33798
rect 14648 33448 14700 33454
rect 14648 33390 14700 33396
rect 14752 30734 14780 42520
rect 14832 42502 14884 42508
rect 14936 41414 14964 42656
rect 15212 42684 15240 42758
rect 15384 42696 15436 42702
rect 15212 42656 15384 42684
rect 15108 42638 15160 42644
rect 15384 42638 15436 42644
rect 15108 42560 15160 42566
rect 14844 41386 14964 41414
rect 15028 42520 15108 42548
rect 14844 33658 14872 41386
rect 14924 33924 14976 33930
rect 14924 33866 14976 33872
rect 14832 33652 14884 33658
rect 14832 33594 14884 33600
rect 14936 33561 14964 33866
rect 14922 33552 14978 33561
rect 14922 33487 14978 33496
rect 14832 33448 14884 33454
rect 14832 33390 14884 33396
rect 14924 33448 14976 33454
rect 14924 33390 14976 33396
rect 14844 33114 14872 33390
rect 14832 33108 14884 33114
rect 14832 33050 14884 33056
rect 14832 32904 14884 32910
rect 14832 32846 14884 32852
rect 14844 32502 14872 32846
rect 14832 32496 14884 32502
rect 14832 32438 14884 32444
rect 14844 31754 14872 32438
rect 14936 32026 14964 33390
rect 14924 32020 14976 32026
rect 14924 31962 14976 31968
rect 14832 31748 14884 31754
rect 14832 31690 14884 31696
rect 14844 30938 14872 31690
rect 14832 30932 14884 30938
rect 14832 30874 14884 30880
rect 15028 30802 15056 42520
rect 15108 42502 15160 42508
rect 15292 42560 15344 42566
rect 15292 42502 15344 42508
rect 15304 42265 15332 42502
rect 15290 42256 15346 42265
rect 15290 42191 15346 42200
rect 15108 41540 15160 41546
rect 15108 41482 15160 41488
rect 15120 36310 15148 41482
rect 15200 41472 15252 41478
rect 15200 41414 15252 41420
rect 15212 40118 15240 41414
rect 15200 40112 15252 40118
rect 15200 40054 15252 40060
rect 15200 37936 15252 37942
rect 15200 37878 15252 37884
rect 15108 36304 15160 36310
rect 15108 36246 15160 36252
rect 15108 34400 15160 34406
rect 15108 34342 15160 34348
rect 15120 33522 15148 34342
rect 15108 33516 15160 33522
rect 15108 33458 15160 33464
rect 15108 31680 15160 31686
rect 15108 31622 15160 31628
rect 15016 30796 15068 30802
rect 15016 30738 15068 30744
rect 14740 30728 14792 30734
rect 14740 30670 14792 30676
rect 14832 30592 14884 30598
rect 14832 30534 14884 30540
rect 14844 29730 14872 30534
rect 14752 29702 14872 29730
rect 14556 29572 14608 29578
rect 14556 29514 14608 29520
rect 14372 29504 14424 29510
rect 14372 29446 14424 29452
rect 14648 29504 14700 29510
rect 14648 29446 14700 29452
rect 14384 29306 14412 29446
rect 14372 29300 14424 29306
rect 14372 29242 14424 29248
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14384 26772 14412 27406
rect 14556 27396 14608 27402
rect 14556 27338 14608 27344
rect 14568 26994 14596 27338
rect 14556 26988 14608 26994
rect 14556 26930 14608 26936
rect 14464 26784 14516 26790
rect 14384 26744 14464 26772
rect 14464 26726 14516 26732
rect 14372 26444 14424 26450
rect 14372 26386 14424 26392
rect 14384 24274 14412 26386
rect 14464 26376 14516 26382
rect 14568 26364 14596 26930
rect 14516 26336 14596 26364
rect 14464 26318 14516 26324
rect 14476 25362 14504 26318
rect 14554 26208 14610 26217
rect 14554 26143 14610 26152
rect 14464 25356 14516 25362
rect 14464 25298 14516 25304
rect 14568 25242 14596 26143
rect 14660 25362 14688 29446
rect 14752 28082 14780 29702
rect 14832 29640 14884 29646
rect 14832 29582 14884 29588
rect 14844 28966 14872 29582
rect 14922 29200 14978 29209
rect 15120 29186 15148 31622
rect 15212 29850 15240 37878
rect 15672 37806 15700 43046
rect 15785 43004 16093 43013
rect 15785 43002 15791 43004
rect 15847 43002 15871 43004
rect 15927 43002 15951 43004
rect 16007 43002 16031 43004
rect 16087 43002 16093 43004
rect 15847 42950 15849 43002
rect 16029 42950 16031 43002
rect 15785 42948 15791 42950
rect 15847 42948 15871 42950
rect 15927 42948 15951 42950
rect 16007 42948 16031 42950
rect 16087 42948 16093 42950
rect 15785 42939 16093 42948
rect 15785 41916 16093 41925
rect 15785 41914 15791 41916
rect 15847 41914 15871 41916
rect 15927 41914 15951 41916
rect 16007 41914 16031 41916
rect 16087 41914 16093 41916
rect 15847 41862 15849 41914
rect 16029 41862 16031 41914
rect 15785 41860 15791 41862
rect 15847 41860 15871 41862
rect 15927 41860 15951 41862
rect 16007 41860 16031 41862
rect 16087 41860 16093 41862
rect 15785 41851 16093 41860
rect 15785 40828 16093 40837
rect 15785 40826 15791 40828
rect 15847 40826 15871 40828
rect 15927 40826 15951 40828
rect 16007 40826 16031 40828
rect 16087 40826 16093 40828
rect 15847 40774 15849 40826
rect 16029 40774 16031 40826
rect 15785 40772 15791 40774
rect 15847 40772 15871 40774
rect 15927 40772 15951 40774
rect 16007 40772 16031 40774
rect 16087 40772 16093 40774
rect 15785 40763 16093 40772
rect 15785 39740 16093 39749
rect 15785 39738 15791 39740
rect 15847 39738 15871 39740
rect 15927 39738 15951 39740
rect 16007 39738 16031 39740
rect 16087 39738 16093 39740
rect 15847 39686 15849 39738
rect 16029 39686 16031 39738
rect 15785 39684 15791 39686
rect 15847 39684 15871 39686
rect 15927 39684 15951 39686
rect 16007 39684 16031 39686
rect 16087 39684 16093 39686
rect 15785 39675 16093 39684
rect 16132 38758 16160 43114
rect 16500 42702 16528 44840
rect 16776 43246 16804 44840
rect 17052 43790 17080 44840
rect 17040 43784 17092 43790
rect 17040 43726 17092 43732
rect 16856 43648 16908 43654
rect 16856 43590 16908 43596
rect 16868 43450 16896 43590
rect 16856 43444 16908 43450
rect 16856 43386 16908 43392
rect 17236 43314 17264 44882
rect 17314 44840 17370 45000
rect 17590 44840 17646 45000
rect 17866 44840 17922 45000
rect 18142 44962 18198 45000
rect 18418 44962 18474 45000
rect 18694 44962 18750 45000
rect 18064 44934 18198 44962
rect 17328 43654 17356 44840
rect 17604 43722 17632 44840
rect 17880 44792 17908 44840
rect 17880 44764 18000 44792
rect 17592 43716 17644 43722
rect 17592 43658 17644 43664
rect 17316 43648 17368 43654
rect 17316 43590 17368 43596
rect 17684 43444 17736 43450
rect 17684 43386 17736 43392
rect 17868 43444 17920 43450
rect 17868 43386 17920 43392
rect 17224 43308 17276 43314
rect 17224 43250 17276 43256
rect 17316 43308 17368 43314
rect 17316 43250 17368 43256
rect 16764 43240 16816 43246
rect 16764 43182 16816 43188
rect 17328 42906 17356 43250
rect 17408 43172 17460 43178
rect 17408 43114 17460 43120
rect 17500 43172 17552 43178
rect 17500 43114 17552 43120
rect 17420 42906 17448 43114
rect 17316 42900 17368 42906
rect 17316 42842 17368 42848
rect 17408 42900 17460 42906
rect 17408 42842 17460 42848
rect 17512 42702 17540 43114
rect 17592 43104 17644 43110
rect 17592 43046 17644 43052
rect 16488 42696 16540 42702
rect 16488 42638 16540 42644
rect 17500 42696 17552 42702
rect 17500 42638 17552 42644
rect 16396 42628 16448 42634
rect 16396 42570 16448 42576
rect 16302 42256 16358 42265
rect 16224 42226 16302 42242
rect 16212 42220 16302 42226
rect 16264 42214 16302 42220
rect 16302 42191 16358 42200
rect 16408 42208 16436 42570
rect 16764 42560 16816 42566
rect 16764 42502 16816 42508
rect 17224 42560 17276 42566
rect 17224 42502 17276 42508
rect 17316 42560 17368 42566
rect 17316 42502 17368 42508
rect 16408 42180 16528 42208
rect 16212 42162 16264 42168
rect 16396 42084 16448 42090
rect 16396 42026 16448 42032
rect 16304 42016 16356 42022
rect 16304 41958 16356 41964
rect 16316 41818 16344 41958
rect 16408 41818 16436 42026
rect 16304 41812 16356 41818
rect 16304 41754 16356 41760
rect 16396 41812 16448 41818
rect 16396 41754 16448 41760
rect 16500 41698 16528 42180
rect 16672 41812 16724 41818
rect 16672 41754 16724 41760
rect 16408 41670 16528 41698
rect 16212 41472 16264 41478
rect 16210 41440 16212 41449
rect 16264 41440 16266 41449
rect 16210 41375 16266 41384
rect 16120 38752 16172 38758
rect 16120 38694 16172 38700
rect 15785 38652 16093 38661
rect 15785 38650 15791 38652
rect 15847 38650 15871 38652
rect 15927 38650 15951 38652
rect 16007 38650 16031 38652
rect 16087 38650 16093 38652
rect 15847 38598 15849 38650
rect 16029 38598 16031 38650
rect 15785 38596 15791 38598
rect 15847 38596 15871 38598
rect 15927 38596 15951 38598
rect 16007 38596 16031 38598
rect 16087 38596 16093 38598
rect 15785 38587 16093 38596
rect 15660 37800 15712 37806
rect 15660 37742 15712 37748
rect 15785 37564 16093 37573
rect 15785 37562 15791 37564
rect 15847 37562 15871 37564
rect 15927 37562 15951 37564
rect 16007 37562 16031 37564
rect 16087 37562 16093 37564
rect 15847 37510 15849 37562
rect 16029 37510 16031 37562
rect 15785 37508 15791 37510
rect 15847 37508 15871 37510
rect 15927 37508 15951 37510
rect 16007 37508 16031 37510
rect 16087 37508 16093 37510
rect 15785 37499 16093 37508
rect 15785 36476 16093 36485
rect 15785 36474 15791 36476
rect 15847 36474 15871 36476
rect 15927 36474 15951 36476
rect 16007 36474 16031 36476
rect 16087 36474 16093 36476
rect 15847 36422 15849 36474
rect 16029 36422 16031 36474
rect 15785 36420 15791 36422
rect 15847 36420 15871 36422
rect 15927 36420 15951 36422
rect 16007 36420 16031 36422
rect 16087 36420 16093 36422
rect 15785 36411 16093 36420
rect 15290 35592 15346 35601
rect 15290 35527 15292 35536
rect 15344 35527 15346 35536
rect 15292 35498 15344 35504
rect 15785 35388 16093 35397
rect 15785 35386 15791 35388
rect 15847 35386 15871 35388
rect 15927 35386 15951 35388
rect 16007 35386 16031 35388
rect 16087 35386 16093 35388
rect 15847 35334 15849 35386
rect 16029 35334 16031 35386
rect 15785 35332 15791 35334
rect 15847 35332 15871 35334
rect 15927 35332 15951 35334
rect 16007 35332 16031 35334
rect 16087 35332 16093 35334
rect 15785 35323 16093 35332
rect 15476 35012 15528 35018
rect 15476 34954 15528 34960
rect 15488 34746 15516 34954
rect 15476 34740 15528 34746
rect 15476 34682 15528 34688
rect 15488 34066 15516 34682
rect 16120 34672 16172 34678
rect 16118 34640 16120 34649
rect 16172 34640 16174 34649
rect 16118 34575 16174 34584
rect 16408 34542 16436 41670
rect 16684 40712 16712 41754
rect 16500 40684 16712 40712
rect 16500 37262 16528 40684
rect 16580 40588 16632 40594
rect 16580 40530 16632 40536
rect 16488 37256 16540 37262
rect 16488 37198 16540 37204
rect 16396 34536 16448 34542
rect 16396 34478 16448 34484
rect 16304 34400 16356 34406
rect 16304 34342 16356 34348
rect 15785 34300 16093 34309
rect 15785 34298 15791 34300
rect 15847 34298 15871 34300
rect 15927 34298 15951 34300
rect 16007 34298 16031 34300
rect 16087 34298 16093 34300
rect 15847 34246 15849 34298
rect 16029 34246 16031 34298
rect 15785 34244 15791 34246
rect 15847 34244 15871 34246
rect 15927 34244 15951 34246
rect 16007 34244 16031 34246
rect 16087 34244 16093 34246
rect 15785 34235 16093 34244
rect 16316 34202 16344 34342
rect 16304 34196 16356 34202
rect 16304 34138 16356 34144
rect 15476 34060 15528 34066
rect 15476 34002 15528 34008
rect 15384 33992 15436 33998
rect 15384 33934 15436 33940
rect 16500 33946 16528 37198
rect 16592 36378 16620 40530
rect 16670 38720 16726 38729
rect 16670 38655 16726 38664
rect 16580 36372 16632 36378
rect 16580 36314 16632 36320
rect 16684 34746 16712 38655
rect 16776 36650 16804 42502
rect 17236 42362 17264 42502
rect 17328 42362 17356 42502
rect 17224 42356 17276 42362
rect 17224 42298 17276 42304
rect 17316 42356 17368 42362
rect 17316 42298 17368 42304
rect 17604 42265 17632 43046
rect 17696 42362 17724 43386
rect 17880 42702 17908 43386
rect 17972 43246 18000 44764
rect 18064 44554 18092 44934
rect 18142 44840 18198 44934
rect 18340 44934 18474 44962
rect 18524 44946 18750 44962
rect 18340 44690 18368 44934
rect 18418 44840 18474 44934
rect 18512 44940 18750 44946
rect 18564 44934 18750 44940
rect 18512 44882 18564 44888
rect 18694 44840 18750 44934
rect 18970 44840 19026 45000
rect 19246 44840 19302 45000
rect 19522 44840 19578 45000
rect 19798 44840 19854 45000
rect 20074 44962 20130 45000
rect 20350 44962 20406 45000
rect 20074 44934 20300 44962
rect 20074 44840 20130 44934
rect 18248 44662 18368 44690
rect 18064 44526 18184 44554
rect 18052 43784 18104 43790
rect 18052 43726 18104 43732
rect 18064 43314 18092 43726
rect 18052 43308 18104 43314
rect 18052 43250 18104 43256
rect 17960 43240 18012 43246
rect 17960 43182 18012 43188
rect 18052 43104 18104 43110
rect 18052 43046 18104 43052
rect 18064 42702 18092 43046
rect 18156 42786 18184 44526
rect 18248 43382 18276 44662
rect 18984 43738 19012 44840
rect 18604 43716 18656 43722
rect 18984 43710 19196 43738
rect 18604 43658 18656 43664
rect 18328 43648 18380 43654
rect 18328 43590 18380 43596
rect 18236 43376 18288 43382
rect 18236 43318 18288 43324
rect 18340 43314 18368 43590
rect 18616 43314 18644 43658
rect 18752 43548 19060 43557
rect 18752 43546 18758 43548
rect 18814 43546 18838 43548
rect 18894 43546 18918 43548
rect 18974 43546 18998 43548
rect 19054 43546 19060 43548
rect 18814 43494 18816 43546
rect 18996 43494 18998 43546
rect 18752 43492 18758 43494
rect 18814 43492 18838 43494
rect 18894 43492 18918 43494
rect 18974 43492 18998 43494
rect 19054 43492 19060 43494
rect 18752 43483 19060 43492
rect 18328 43308 18380 43314
rect 18328 43250 18380 43256
rect 18604 43308 18656 43314
rect 18604 43250 18656 43256
rect 18512 43240 18564 43246
rect 18512 43182 18564 43188
rect 18418 42800 18474 42809
rect 18156 42758 18418 42786
rect 18418 42735 18474 42744
rect 17868 42696 17920 42702
rect 17868 42638 17920 42644
rect 18052 42696 18104 42702
rect 18052 42638 18104 42644
rect 17776 42560 17828 42566
rect 17776 42502 17828 42508
rect 18052 42560 18104 42566
rect 18052 42502 18104 42508
rect 18328 42560 18380 42566
rect 18328 42502 18380 42508
rect 18420 42560 18472 42566
rect 18420 42502 18472 42508
rect 17788 42362 17816 42502
rect 18064 42362 18092 42502
rect 18340 42362 18368 42502
rect 17684 42356 17736 42362
rect 17684 42298 17736 42304
rect 17776 42356 17828 42362
rect 17776 42298 17828 42304
rect 18052 42356 18104 42362
rect 18052 42298 18104 42304
rect 18328 42356 18380 42362
rect 18328 42298 18380 42304
rect 18432 42294 18460 42502
rect 18420 42288 18472 42294
rect 17590 42256 17646 42265
rect 18420 42230 18472 42236
rect 17590 42191 17646 42200
rect 16948 42084 17000 42090
rect 16948 42026 17000 42032
rect 17316 42084 17368 42090
rect 17316 42026 17368 42032
rect 18420 42084 18472 42090
rect 18420 42026 18472 42032
rect 16960 41414 16988 42026
rect 17328 41857 17356 42026
rect 17592 42016 17644 42022
rect 17592 41958 17644 41964
rect 17960 42016 18012 42022
rect 17960 41958 18012 41964
rect 17314 41848 17370 41857
rect 17314 41783 17370 41792
rect 17604 41721 17632 41958
rect 17972 41721 18000 41958
rect 17590 41712 17646 41721
rect 17590 41647 17646 41656
rect 17958 41712 18014 41721
rect 17958 41647 18014 41656
rect 18328 41472 18380 41478
rect 18328 41414 18380 41420
rect 16960 41386 17080 41414
rect 16856 40112 16908 40118
rect 16854 40080 16856 40089
rect 16908 40080 16910 40089
rect 16854 40015 16910 40024
rect 16764 36644 16816 36650
rect 16764 36586 16816 36592
rect 16672 34740 16724 34746
rect 16672 34682 16724 34688
rect 16684 34610 16712 34682
rect 16672 34604 16724 34610
rect 16672 34546 16724 34552
rect 15396 33436 15424 33934
rect 16500 33918 16620 33946
rect 16488 33856 16540 33862
rect 16488 33798 16540 33804
rect 15396 33408 15700 33436
rect 15568 33040 15620 33046
rect 15568 32982 15620 32988
rect 15580 32910 15608 32982
rect 15384 32904 15436 32910
rect 15568 32904 15620 32910
rect 15436 32864 15516 32892
rect 15384 32846 15436 32852
rect 15382 32464 15438 32473
rect 15382 32399 15438 32408
rect 15396 32178 15424 32399
rect 15304 32150 15424 32178
rect 15304 31754 15332 32150
rect 15304 31726 15424 31754
rect 15292 30728 15344 30734
rect 15292 30670 15344 30676
rect 15200 29844 15252 29850
rect 15200 29786 15252 29792
rect 14922 29135 14978 29144
rect 15028 29158 15148 29186
rect 14832 28960 14884 28966
rect 14832 28902 14884 28908
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 14752 27713 14780 28018
rect 14844 28014 14872 28902
rect 14832 28008 14884 28014
rect 14832 27950 14884 27956
rect 14738 27704 14794 27713
rect 14738 27639 14794 27648
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 14740 27328 14792 27334
rect 14740 27270 14792 27276
rect 14752 26994 14780 27270
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 14752 25838 14780 26726
rect 14844 26042 14872 27406
rect 14832 26036 14884 26042
rect 14832 25978 14884 25984
rect 14740 25832 14792 25838
rect 14740 25774 14792 25780
rect 14648 25356 14700 25362
rect 14648 25298 14700 25304
rect 14476 25214 14596 25242
rect 14372 24268 14424 24274
rect 14372 24210 14424 24216
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14384 19922 14412 20402
rect 14372 19916 14424 19922
rect 14372 19858 14424 19864
rect 14384 18630 14412 19858
rect 14476 19417 14504 25214
rect 14556 24676 14608 24682
rect 14556 24618 14608 24624
rect 14568 21010 14596 24618
rect 14660 24342 14688 25298
rect 14648 24336 14700 24342
rect 14648 24278 14700 24284
rect 14648 23656 14700 23662
rect 14752 23644 14780 25774
rect 14844 24818 14872 25978
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14936 24682 14964 29135
rect 15028 28393 15056 29158
rect 15108 29028 15160 29034
rect 15108 28970 15160 28976
rect 15014 28384 15070 28393
rect 15014 28319 15070 28328
rect 15120 26466 15148 28970
rect 15304 28558 15332 30670
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 15304 28121 15332 28494
rect 15290 28112 15346 28121
rect 15290 28047 15346 28056
rect 15292 26580 15344 26586
rect 15292 26522 15344 26528
rect 15120 26438 15240 26466
rect 15304 26450 15332 26522
rect 15108 26376 15160 26382
rect 15108 26318 15160 26324
rect 15120 26246 15148 26318
rect 15108 26240 15160 26246
rect 15108 26182 15160 26188
rect 15212 26194 15240 26438
rect 15292 26444 15344 26450
rect 15292 26386 15344 26392
rect 15120 25362 15148 26182
rect 15212 26166 15332 26194
rect 15200 25968 15252 25974
rect 15200 25910 15252 25916
rect 15212 25498 15240 25910
rect 15200 25492 15252 25498
rect 15200 25434 15252 25440
rect 15304 25362 15332 26166
rect 15396 25974 15424 31726
rect 15488 30734 15516 32864
rect 15568 32846 15620 32852
rect 15580 32502 15608 32846
rect 15568 32496 15620 32502
rect 15672 32473 15700 33408
rect 15785 33212 16093 33221
rect 15785 33210 15791 33212
rect 15847 33210 15871 33212
rect 15927 33210 15951 33212
rect 16007 33210 16031 33212
rect 16087 33210 16093 33212
rect 15847 33158 15849 33210
rect 16029 33158 16031 33210
rect 15785 33156 15791 33158
rect 15847 33156 15871 33158
rect 15927 33156 15951 33158
rect 16007 33156 16031 33158
rect 16087 33156 16093 33158
rect 15785 33147 16093 33156
rect 16500 33114 16528 33798
rect 16488 33108 16540 33114
rect 16408 33068 16488 33096
rect 16304 32904 16356 32910
rect 16304 32846 16356 32852
rect 15568 32438 15620 32444
rect 15658 32464 15714 32473
rect 15658 32399 15714 32408
rect 16120 32428 16172 32434
rect 16120 32370 16172 32376
rect 15568 32224 15620 32230
rect 15568 32166 15620 32172
rect 15580 32065 15608 32166
rect 15785 32124 16093 32133
rect 15785 32122 15791 32124
rect 15847 32122 15871 32124
rect 15927 32122 15951 32124
rect 16007 32122 16031 32124
rect 16087 32122 16093 32124
rect 15847 32070 15849 32122
rect 16029 32070 16031 32122
rect 15785 32068 15791 32070
rect 15847 32068 15871 32070
rect 15927 32068 15951 32070
rect 16007 32068 16031 32070
rect 16087 32068 16093 32070
rect 15566 32056 15622 32065
rect 15785 32059 16093 32068
rect 15566 31991 15622 32000
rect 16026 31920 16082 31929
rect 16026 31855 16082 31864
rect 15568 31816 15620 31822
rect 15568 31758 15620 31764
rect 15580 30802 15608 31758
rect 16040 31346 16068 31855
rect 16028 31340 16080 31346
rect 16028 31282 16080 31288
rect 15785 31036 16093 31045
rect 15785 31034 15791 31036
rect 15847 31034 15871 31036
rect 15927 31034 15951 31036
rect 16007 31034 16031 31036
rect 16087 31034 16093 31036
rect 15847 30982 15849 31034
rect 16029 30982 16031 31034
rect 15785 30980 15791 30982
rect 15847 30980 15871 30982
rect 15927 30980 15951 30982
rect 16007 30980 16031 30982
rect 16087 30980 16093 30982
rect 15785 30971 16093 30980
rect 15568 30796 15620 30802
rect 15568 30738 15620 30744
rect 15936 30796 15988 30802
rect 15936 30738 15988 30744
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15476 30048 15528 30054
rect 15476 29990 15528 29996
rect 15488 29782 15516 29990
rect 15476 29776 15528 29782
rect 15476 29718 15528 29724
rect 15476 28688 15528 28694
rect 15474 28656 15476 28665
rect 15528 28656 15530 28665
rect 15474 28591 15530 28600
rect 15488 26586 15516 28591
rect 15476 26580 15528 26586
rect 15476 26522 15528 26528
rect 15476 26444 15528 26450
rect 15476 26386 15528 26392
rect 15488 26353 15516 26386
rect 15474 26344 15530 26353
rect 15474 26279 15530 26288
rect 15384 25968 15436 25974
rect 15384 25910 15436 25916
rect 15108 25356 15160 25362
rect 15108 25298 15160 25304
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 14924 24676 14976 24682
rect 14924 24618 14976 24624
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 15120 24274 15148 24550
rect 15304 24274 15332 25298
rect 14832 24268 14884 24274
rect 14832 24210 14884 24216
rect 15108 24268 15160 24274
rect 15108 24210 15160 24216
rect 15292 24268 15344 24274
rect 15292 24210 15344 24216
rect 14700 23616 14780 23644
rect 14648 23598 14700 23604
rect 14660 22438 14688 23598
rect 14844 23118 14872 24210
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 14660 21468 14688 22374
rect 14936 21554 14964 23802
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15304 23633 15332 23666
rect 15290 23624 15346 23633
rect 15290 23559 15346 23568
rect 15198 23488 15254 23497
rect 15198 23423 15254 23432
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 15028 21706 15056 23054
rect 15212 23050 15240 23423
rect 15200 23044 15252 23050
rect 15200 22986 15252 22992
rect 15396 22794 15424 25910
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15304 22766 15424 22794
rect 15108 22432 15160 22438
rect 15304 22409 15332 22766
rect 15384 22432 15436 22438
rect 15108 22374 15160 22380
rect 15290 22400 15346 22409
rect 15120 22166 15148 22374
rect 15384 22374 15436 22380
rect 15290 22335 15346 22344
rect 15108 22160 15160 22166
rect 15108 22102 15160 22108
rect 15106 21720 15162 21729
rect 15028 21678 15106 21706
rect 15106 21655 15162 21664
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 14740 21480 14792 21486
rect 14660 21440 14740 21468
rect 14740 21422 14792 21428
rect 14752 21146 14780 21422
rect 14936 21321 14964 21490
rect 15108 21344 15160 21350
rect 14922 21312 14978 21321
rect 15108 21286 15160 21292
rect 14922 21247 14978 21256
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 15028 20466 15056 20946
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 14556 20324 14608 20330
rect 14556 20266 14608 20272
rect 14568 20058 14596 20266
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14462 19408 14518 19417
rect 14462 19343 14518 19352
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14384 17066 14412 18566
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 14372 16584 14424 16590
rect 14568 16572 14596 19994
rect 14752 19854 14780 19994
rect 14922 19952 14978 19961
rect 14922 19887 14978 19896
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14936 19786 14964 19887
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 14832 19304 14884 19310
rect 14832 19246 14884 19252
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14752 18873 14780 19110
rect 14738 18864 14794 18873
rect 14738 18799 14794 18808
rect 14752 18766 14780 18799
rect 14844 18766 14872 19246
rect 14924 19236 14976 19242
rect 14924 19178 14976 19184
rect 14936 18970 14964 19178
rect 14924 18964 14976 18970
rect 14924 18906 14976 18912
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15028 18290 15056 18566
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 14648 18148 14700 18154
rect 14648 18090 14700 18096
rect 14660 17542 14688 18090
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14648 17060 14700 17066
rect 14648 17002 14700 17008
rect 14424 16544 14596 16572
rect 14372 16526 14424 16532
rect 14280 15088 14332 15094
rect 14280 15030 14332 15036
rect 14292 14958 14320 15030
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13780 10696 13860 10724
rect 13912 10736 13964 10742
rect 13728 10678 13780 10684
rect 13912 10678 13964 10684
rect 13450 8800 13506 8809
rect 13450 8735 13506 8744
rect 13464 8362 13492 8735
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13452 8016 13504 8022
rect 13452 7958 13504 7964
rect 13464 7410 13492 7958
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13464 4282 13492 6666
rect 13556 5370 13584 10662
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13648 10266 13676 10542
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13740 9674 13768 10678
rect 13924 10010 13952 10678
rect 14016 10130 14044 11698
rect 14200 10810 14228 14214
rect 14384 13802 14412 16526
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14568 16182 14596 16390
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14464 15496 14516 15502
rect 14556 15496 14608 15502
rect 14464 15438 14516 15444
rect 14554 15464 14556 15473
rect 14608 15464 14610 15473
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14384 12889 14412 13738
rect 14476 12918 14504 15438
rect 14554 15399 14610 15408
rect 14464 12912 14516 12918
rect 14370 12880 14426 12889
rect 14464 12854 14516 12860
rect 14568 12850 14596 15399
rect 14660 14822 14688 17002
rect 14740 16176 14792 16182
rect 14740 16118 14792 16124
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14646 13968 14702 13977
rect 14646 13903 14702 13912
rect 14660 12918 14688 13903
rect 14648 12912 14700 12918
rect 14648 12854 14700 12860
rect 14370 12815 14426 12824
rect 14556 12844 14608 12850
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14292 11898 14320 12242
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14292 11286 14320 11698
rect 14280 11280 14332 11286
rect 14280 11222 14332 11228
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14108 10266 14136 10610
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14384 10062 14412 12815
rect 14556 12786 14608 12792
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14476 11830 14504 12106
rect 14568 12084 14596 12582
rect 14752 12102 14780 16118
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 14936 14958 14964 15098
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14844 14618 14872 14826
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14936 13444 14964 14758
rect 14844 13416 14964 13444
rect 14648 12096 14700 12102
rect 14568 12056 14648 12084
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14464 10668 14516 10674
rect 14568 10656 14596 12056
rect 14648 12038 14700 12044
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14660 11218 14688 11630
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14660 10674 14688 11154
rect 14844 10962 14872 13416
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14752 10934 14872 10962
rect 14516 10628 14596 10656
rect 14648 10668 14700 10674
rect 14464 10610 14516 10616
rect 14648 10610 14700 10616
rect 14372 10056 14424 10062
rect 13924 9982 14136 10010
rect 14372 9998 14424 10004
rect 13648 9646 13768 9674
rect 13648 8566 13676 9646
rect 14108 8838 14136 9982
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13648 8294 13676 8502
rect 14108 8498 14136 8774
rect 14476 8634 14504 10610
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13542 5264 13598 5273
rect 13648 5234 13676 8230
rect 13832 7546 13860 8230
rect 13912 7812 13964 7818
rect 13912 7754 13964 7760
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13726 7304 13782 7313
rect 13726 7239 13782 7248
rect 13542 5199 13598 5208
rect 13636 5228 13688 5234
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13464 3398 13492 4218
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13004 2746 13216 2774
rect 13280 2746 13400 2774
rect 11980 2440 12032 2446
rect 12440 2440 12492 2446
rect 11980 2382 12032 2388
rect 12268 2400 12440 2428
rect 11520 2372 11572 2378
rect 11520 2314 11572 2320
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 11716 2038 11744 2246
rect 11704 2032 11756 2038
rect 11704 1974 11756 1980
rect 11704 1896 11756 1902
rect 11704 1838 11756 1844
rect 11716 1494 11744 1838
rect 11704 1488 11756 1494
rect 11704 1430 11756 1436
rect 11808 1358 11836 2246
rect 11888 1828 11940 1834
rect 11888 1770 11940 1776
rect 11796 1352 11848 1358
rect 11796 1294 11848 1300
rect 11520 1216 11572 1222
rect 11520 1158 11572 1164
rect 11704 1216 11756 1222
rect 11704 1158 11756 1164
rect 11532 814 11560 1158
rect 11520 808 11572 814
rect 11520 750 11572 756
rect 11716 626 11744 1158
rect 11532 598 11744 626
rect 11428 400 11480 406
rect 11428 342 11480 348
rect 11532 160 11560 598
rect 11242 82 11298 160
rect 11164 54 11298 82
rect 11242 0 11298 54
rect 11518 0 11574 160
rect 11794 82 11850 160
rect 11900 82 11928 1770
rect 12084 1494 12112 2246
rect 12268 1766 12296 2400
rect 12440 2382 12492 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 12440 2304 12492 2310
rect 13004 2292 13032 2746
rect 13280 2446 13308 2746
rect 13556 2446 13584 5199
rect 13636 5170 13688 5176
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13544 2440 13596 2446
rect 13648 2417 13676 4150
rect 13740 3058 13768 7239
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5953 13860 6054
rect 13818 5944 13874 5953
rect 13924 5914 13952 7754
rect 13818 5879 13874 5888
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 14016 5166 14044 8434
rect 14200 7546 14228 8434
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13924 3670 13952 3946
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13544 2382 13596 2388
rect 13634 2408 13690 2417
rect 13634 2343 13690 2352
rect 12440 2246 12492 2252
rect 12728 2264 13032 2292
rect 13176 2304 13228 2310
rect 12348 1964 12400 1970
rect 12348 1906 12400 1912
rect 12256 1760 12308 1766
rect 12256 1702 12308 1708
rect 12360 1544 12388 1906
rect 12452 1562 12480 2246
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 12268 1516 12388 1544
rect 12440 1556 12492 1562
rect 11980 1488 12032 1494
rect 11980 1430 12032 1436
rect 12072 1488 12124 1494
rect 12072 1430 12124 1436
rect 11992 898 12020 1430
rect 12268 1426 12296 1516
rect 12440 1498 12492 1504
rect 12532 1556 12584 1562
rect 12532 1498 12584 1504
rect 12544 1442 12572 1498
rect 12256 1420 12308 1426
rect 12256 1362 12308 1368
rect 12360 1414 12572 1442
rect 11992 870 12112 898
rect 12084 160 12112 870
rect 12360 160 12388 1414
rect 12636 160 12664 1702
rect 12728 678 12756 2264
rect 13176 2246 13228 2252
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 12818 2204 13126 2213
rect 12818 2202 12824 2204
rect 12880 2202 12904 2204
rect 12960 2202 12984 2204
rect 13040 2202 13064 2204
rect 13120 2202 13126 2204
rect 12880 2150 12882 2202
rect 13062 2150 13064 2202
rect 12818 2148 12824 2150
rect 12880 2148 12904 2150
rect 12960 2148 12984 2150
rect 13040 2148 13064 2150
rect 13120 2148 13126 2150
rect 12818 2139 13126 2148
rect 13188 1358 13216 2246
rect 13372 2106 13400 2246
rect 13648 2106 13676 2246
rect 13360 2100 13412 2106
rect 13360 2042 13412 2048
rect 13636 2100 13688 2106
rect 13636 2042 13688 2048
rect 13726 2000 13782 2009
rect 13832 1970 13860 3334
rect 13924 2582 13952 3334
rect 14016 2650 14044 5102
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 13912 2576 13964 2582
rect 13912 2518 13964 2524
rect 13726 1935 13728 1944
rect 13780 1935 13782 1944
rect 13820 1964 13872 1970
rect 13728 1906 13780 1912
rect 13820 1906 13872 1912
rect 13360 1760 13412 1766
rect 13360 1702 13412 1708
rect 13636 1760 13688 1766
rect 13636 1702 13688 1708
rect 14096 1760 14148 1766
rect 14096 1702 14148 1708
rect 13372 1562 13400 1702
rect 13360 1556 13412 1562
rect 13360 1498 13412 1504
rect 13648 1358 13676 1702
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 13176 1352 13228 1358
rect 13636 1352 13688 1358
rect 13176 1294 13228 1300
rect 13372 1278 13584 1306
rect 13636 1294 13688 1300
rect 12818 1116 13126 1125
rect 12818 1114 12824 1116
rect 12880 1114 12904 1116
rect 12960 1114 12984 1116
rect 13040 1114 13064 1116
rect 13120 1114 13126 1116
rect 12880 1062 12882 1114
rect 13062 1062 13064 1114
rect 12818 1060 12824 1062
rect 12880 1060 12904 1062
rect 12960 1060 12984 1062
rect 13040 1060 13064 1062
rect 13120 1060 13126 1062
rect 12818 1051 13126 1060
rect 12900 1012 12952 1018
rect 12900 954 12952 960
rect 12716 672 12768 678
rect 12716 614 12768 620
rect 12912 160 12940 954
rect 11794 54 11928 82
rect 11794 0 11850 54
rect 12070 0 12126 160
rect 12346 0 12402 160
rect 12622 0 12678 160
rect 12898 0 12954 160
rect 13174 82 13230 160
rect 13372 82 13400 1278
rect 13452 1216 13504 1222
rect 13556 1204 13584 1278
rect 13636 1216 13688 1222
rect 13556 1176 13636 1204
rect 13452 1158 13504 1164
rect 13636 1158 13688 1164
rect 13464 160 13492 1158
rect 13740 160 13768 1498
rect 14108 1494 14136 1702
rect 14200 1494 14228 7142
rect 14646 5808 14702 5817
rect 14646 5743 14702 5752
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14370 5264 14426 5273
rect 14370 5199 14426 5208
rect 14384 4622 14412 5199
rect 14568 5166 14596 5306
rect 14660 5166 14688 5743
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14384 3194 14412 4558
rect 14568 4078 14596 5102
rect 14752 4672 14780 10934
rect 14832 10736 14884 10742
rect 14936 10724 14964 12038
rect 15016 11144 15068 11150
rect 15014 11112 15016 11121
rect 15068 11112 15070 11121
rect 15014 11047 15070 11056
rect 14884 10696 14964 10724
rect 14832 10678 14884 10684
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14844 8974 14872 10542
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14844 7342 14872 8910
rect 14936 8566 14964 10696
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 15028 8412 15056 8774
rect 14936 8384 15056 8412
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14844 4826 14872 5170
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14832 4684 14884 4690
rect 14752 4644 14832 4672
rect 14832 4626 14884 4632
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14476 3738 14504 3878
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14936 3534 14964 8384
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 15028 4146 15056 8230
rect 15016 4140 15068 4146
rect 15016 4082 15068 4088
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 14280 1964 14332 1970
rect 14280 1906 14332 1912
rect 14292 1873 14320 1906
rect 14278 1864 14334 1873
rect 14278 1799 14334 1808
rect 14280 1760 14332 1766
rect 14280 1702 14332 1708
rect 14096 1488 14148 1494
rect 14096 1430 14148 1436
rect 14188 1488 14240 1494
rect 14188 1430 14240 1436
rect 14004 1216 14056 1222
rect 14004 1158 14056 1164
rect 14016 160 14044 1158
rect 14292 160 14320 1702
rect 14384 1018 14412 2790
rect 14830 2680 14886 2689
rect 14830 2615 14886 2624
rect 14738 2544 14794 2553
rect 14738 2479 14794 2488
rect 14752 2446 14780 2479
rect 14844 2446 14872 2615
rect 15120 2446 15148 21286
rect 15304 20534 15332 22335
rect 15396 22098 15424 22374
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15382 21720 15438 21729
rect 15382 21655 15438 21664
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 15304 19666 15332 20334
rect 15212 19638 15332 19666
rect 15212 19310 15240 19638
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15212 17882 15240 19246
rect 15304 18834 15332 19246
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15212 17678 15240 17818
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15212 15570 15240 17614
rect 15396 16998 15424 21655
rect 15488 20777 15516 24754
rect 15580 20874 15608 30738
rect 15660 30728 15712 30734
rect 15660 30670 15712 30676
rect 15672 28558 15700 30670
rect 15948 30394 15976 30738
rect 15936 30388 15988 30394
rect 15936 30330 15988 30336
rect 15785 29948 16093 29957
rect 15785 29946 15791 29948
rect 15847 29946 15871 29948
rect 15927 29946 15951 29948
rect 16007 29946 16031 29948
rect 16087 29946 16093 29948
rect 15847 29894 15849 29946
rect 16029 29894 16031 29946
rect 15785 29892 15791 29894
rect 15847 29892 15871 29894
rect 15927 29892 15951 29894
rect 16007 29892 16031 29894
rect 16087 29892 16093 29894
rect 15785 29883 16093 29892
rect 15752 29844 15804 29850
rect 15752 29786 15804 29792
rect 15764 29646 15792 29786
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15785 28860 16093 28869
rect 15785 28858 15791 28860
rect 15847 28858 15871 28860
rect 15927 28858 15951 28860
rect 16007 28858 16031 28860
rect 16087 28858 16093 28860
rect 15847 28806 15849 28858
rect 16029 28806 16031 28858
rect 15785 28804 15791 28806
rect 15847 28804 15871 28806
rect 15927 28804 15951 28806
rect 16007 28804 16031 28806
rect 16087 28804 16093 28806
rect 15785 28795 16093 28804
rect 15936 28620 15988 28626
rect 15936 28562 15988 28568
rect 15660 28552 15712 28558
rect 15660 28494 15712 28500
rect 15672 25809 15700 28494
rect 15752 28212 15804 28218
rect 15752 28154 15804 28160
rect 15764 28121 15792 28154
rect 15750 28112 15806 28121
rect 15948 28082 15976 28562
rect 15750 28047 15806 28056
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 15785 27772 16093 27781
rect 15785 27770 15791 27772
rect 15847 27770 15871 27772
rect 15927 27770 15951 27772
rect 16007 27770 16031 27772
rect 16087 27770 16093 27772
rect 15847 27718 15849 27770
rect 16029 27718 16031 27770
rect 15785 27716 15791 27718
rect 15847 27716 15871 27718
rect 15927 27716 15951 27718
rect 16007 27716 16031 27718
rect 16087 27716 16093 27718
rect 15785 27707 16093 27716
rect 15785 26684 16093 26693
rect 15785 26682 15791 26684
rect 15847 26682 15871 26684
rect 15927 26682 15951 26684
rect 16007 26682 16031 26684
rect 16087 26682 16093 26684
rect 15847 26630 15849 26682
rect 16029 26630 16031 26682
rect 15785 26628 15791 26630
rect 15847 26628 15871 26630
rect 15927 26628 15951 26630
rect 16007 26628 16031 26630
rect 16087 26628 16093 26630
rect 15785 26619 16093 26628
rect 15844 26580 15896 26586
rect 15844 26522 15896 26528
rect 15856 26330 15884 26522
rect 16132 26450 16160 32370
rect 16316 31754 16344 32846
rect 16408 31958 16436 33068
rect 16488 33050 16540 33056
rect 16592 32994 16620 33918
rect 16500 32966 16620 32994
rect 16396 31952 16448 31958
rect 16396 31894 16448 31900
rect 16500 31754 16528 32966
rect 16684 32434 16712 34546
rect 16868 33590 16896 40015
rect 16948 39840 17000 39846
rect 16948 39782 17000 39788
rect 16856 33584 16908 33590
rect 16856 33526 16908 33532
rect 16764 32972 16816 32978
rect 16816 32932 16896 32960
rect 16764 32914 16816 32920
rect 16762 32600 16818 32609
rect 16762 32535 16818 32544
rect 16776 32502 16804 32535
rect 16764 32496 16816 32502
rect 16764 32438 16816 32444
rect 16672 32428 16724 32434
rect 16672 32370 16724 32376
rect 16868 32212 16896 32932
rect 16960 32314 16988 39782
rect 17052 32994 17080 41386
rect 17316 40996 17368 41002
rect 17316 40938 17368 40944
rect 17224 34672 17276 34678
rect 17224 34614 17276 34620
rect 17132 33992 17184 33998
rect 17132 33934 17184 33940
rect 17144 33114 17172 33934
rect 17132 33108 17184 33114
rect 17132 33050 17184 33056
rect 17236 33017 17264 34614
rect 17328 33674 17356 40938
rect 17958 40624 18014 40633
rect 17958 40559 18014 40568
rect 17972 39302 18000 40559
rect 17960 39296 18012 39302
rect 17960 39238 18012 39244
rect 18340 39030 18368 41414
rect 18328 39024 18380 39030
rect 18328 38966 18380 38972
rect 18144 38344 18196 38350
rect 18144 38286 18196 38292
rect 18156 38010 18184 38286
rect 18144 38004 18196 38010
rect 18144 37946 18196 37952
rect 17776 36644 17828 36650
rect 17776 36586 17828 36592
rect 18144 36644 18196 36650
rect 18144 36586 18196 36592
rect 17684 35624 17736 35630
rect 17684 35566 17736 35572
rect 17408 34740 17460 34746
rect 17408 34682 17460 34688
rect 17420 33998 17448 34682
rect 17500 34400 17552 34406
rect 17500 34342 17552 34348
rect 17512 34202 17540 34342
rect 17500 34196 17552 34202
rect 17500 34138 17552 34144
rect 17408 33992 17460 33998
rect 17408 33934 17460 33940
rect 17592 33992 17644 33998
rect 17592 33934 17644 33940
rect 17328 33646 17540 33674
rect 17604 33658 17632 33934
rect 17408 33584 17460 33590
rect 17408 33526 17460 33532
rect 17316 33516 17368 33522
rect 17316 33458 17368 33464
rect 17222 33008 17278 33017
rect 17052 32966 17172 32994
rect 17038 32464 17094 32473
rect 17038 32399 17040 32408
rect 17092 32399 17094 32408
rect 17040 32370 17092 32376
rect 16960 32286 17080 32314
rect 16948 32224 17000 32230
rect 16868 32184 16948 32212
rect 16672 32020 16724 32026
rect 16672 31962 16724 31968
rect 16684 31822 16712 31962
rect 16868 31890 16896 32184
rect 16948 32166 17000 32172
rect 16856 31884 16908 31890
rect 16856 31826 16908 31832
rect 16672 31816 16724 31822
rect 17052 31770 17080 32286
rect 17144 32008 17172 32966
rect 17222 32943 17278 32952
rect 17328 32026 17356 33458
rect 17316 32020 17368 32026
rect 17144 31980 17264 32008
rect 16672 31758 16724 31764
rect 16224 31726 16344 31754
rect 16408 31726 16528 31754
rect 16224 28558 16252 31726
rect 16304 30932 16356 30938
rect 16304 30874 16356 30880
rect 16316 30802 16344 30874
rect 16304 30796 16356 30802
rect 16304 30738 16356 30744
rect 16304 29640 16356 29646
rect 16304 29582 16356 29588
rect 16212 28552 16264 28558
rect 16212 28494 16264 28500
rect 16224 28422 16252 28494
rect 16212 28416 16264 28422
rect 16212 28358 16264 28364
rect 16316 28200 16344 29582
rect 16224 28172 16344 28200
rect 16120 26444 16172 26450
rect 16120 26386 16172 26392
rect 15856 26302 16160 26330
rect 15658 25800 15714 25809
rect 15658 25735 15714 25744
rect 15660 25696 15712 25702
rect 15660 25638 15712 25644
rect 15672 22642 15700 25638
rect 15785 25596 16093 25605
rect 15785 25594 15791 25596
rect 15847 25594 15871 25596
rect 15927 25594 15951 25596
rect 16007 25594 16031 25596
rect 16087 25594 16093 25596
rect 15847 25542 15849 25594
rect 16029 25542 16031 25594
rect 15785 25540 15791 25542
rect 15847 25540 15871 25542
rect 15927 25540 15951 25542
rect 16007 25540 16031 25542
rect 16087 25540 16093 25542
rect 15785 25531 16093 25540
rect 16132 25242 16160 26302
rect 16224 25344 16252 28172
rect 16304 26444 16356 26450
rect 16304 26386 16356 26392
rect 16316 26058 16344 26386
rect 16408 26217 16436 31726
rect 16488 31136 16540 31142
rect 16488 31078 16540 31084
rect 16500 30802 16528 31078
rect 16488 30796 16540 30802
rect 16488 30738 16540 30744
rect 16488 29776 16540 29782
rect 16488 29718 16540 29724
rect 16500 28626 16528 29718
rect 16488 28620 16540 28626
rect 16488 28562 16540 28568
rect 16488 28416 16540 28422
rect 16488 28358 16540 28364
rect 16580 28416 16632 28422
rect 16580 28358 16632 28364
rect 16394 26208 16450 26217
rect 16394 26143 16450 26152
rect 16316 26030 16436 26058
rect 16304 25356 16356 25362
rect 16224 25316 16304 25344
rect 16304 25298 16356 25304
rect 16132 25214 16344 25242
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 15948 24954 15976 25094
rect 15936 24948 15988 24954
rect 15936 24890 15988 24896
rect 16120 24744 16172 24750
rect 16120 24686 16172 24692
rect 15785 24508 16093 24517
rect 15785 24506 15791 24508
rect 15847 24506 15871 24508
rect 15927 24506 15951 24508
rect 16007 24506 16031 24508
rect 16087 24506 16093 24508
rect 15847 24454 15849 24506
rect 16029 24454 16031 24506
rect 15785 24452 15791 24454
rect 15847 24452 15871 24454
rect 15927 24452 15951 24454
rect 16007 24452 16031 24454
rect 16087 24452 16093 24454
rect 15785 24443 16093 24452
rect 16132 24410 16160 24686
rect 16212 24608 16264 24614
rect 16212 24550 16264 24556
rect 16224 24410 16252 24550
rect 16120 24404 16172 24410
rect 16120 24346 16172 24352
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 16316 24290 16344 25214
rect 16224 24262 16344 24290
rect 16120 23520 16172 23526
rect 16120 23462 16172 23468
rect 15785 23420 16093 23429
rect 15785 23418 15791 23420
rect 15847 23418 15871 23420
rect 15927 23418 15951 23420
rect 16007 23418 16031 23420
rect 16087 23418 16093 23420
rect 15847 23366 15849 23418
rect 16029 23366 16031 23418
rect 15785 23364 15791 23366
rect 15847 23364 15871 23366
rect 15927 23364 15951 23366
rect 16007 23364 16031 23366
rect 16087 23364 16093 23366
rect 15785 23355 16093 23364
rect 16132 23254 16160 23462
rect 16120 23248 16172 23254
rect 16120 23190 16172 23196
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15785 22332 16093 22341
rect 15785 22330 15791 22332
rect 15847 22330 15871 22332
rect 15927 22330 15951 22332
rect 16007 22330 16031 22332
rect 16087 22330 16093 22332
rect 15847 22278 15849 22330
rect 16029 22278 16031 22330
rect 15785 22276 15791 22278
rect 15847 22276 15871 22278
rect 15927 22276 15951 22278
rect 16007 22276 16031 22278
rect 16087 22276 16093 22278
rect 15785 22267 16093 22276
rect 16028 22092 16080 22098
rect 16080 22052 16160 22080
rect 16028 22034 16080 22040
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 15672 21690 15700 21966
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 16132 21457 16160 22052
rect 16118 21448 16174 21457
rect 16118 21383 16174 21392
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15474 20768 15530 20777
rect 15474 20703 15530 20712
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15488 19378 15516 19654
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15488 18426 15516 18906
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15488 16810 15516 18362
rect 15396 16782 15516 16810
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 15212 14958 15240 15370
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15212 14521 15240 14758
rect 15198 14512 15254 14521
rect 15198 14447 15254 14456
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15200 13796 15252 13802
rect 15304 13784 15332 13942
rect 15252 13756 15332 13784
rect 15200 13738 15252 13744
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15212 11150 15240 12106
rect 15304 11218 15332 13466
rect 15396 13308 15424 16782
rect 15580 15434 15608 20810
rect 15672 16794 15700 21286
rect 15785 21244 16093 21253
rect 15785 21242 15791 21244
rect 15847 21242 15871 21244
rect 15927 21242 15951 21244
rect 16007 21242 16031 21244
rect 16087 21242 16093 21244
rect 15847 21190 15849 21242
rect 16029 21190 16031 21242
rect 15785 21188 15791 21190
rect 15847 21188 15871 21190
rect 15927 21188 15951 21190
rect 16007 21188 16031 21190
rect 16087 21188 16093 21190
rect 15785 21179 16093 21188
rect 16132 20913 16160 21383
rect 16118 20904 16174 20913
rect 16118 20839 16174 20848
rect 15785 20156 16093 20165
rect 15785 20154 15791 20156
rect 15847 20154 15871 20156
rect 15927 20154 15951 20156
rect 16007 20154 16031 20156
rect 16087 20154 16093 20156
rect 15847 20102 15849 20154
rect 16029 20102 16031 20154
rect 15785 20100 15791 20102
rect 15847 20100 15871 20102
rect 15927 20100 15951 20102
rect 16007 20100 16031 20102
rect 16087 20100 16093 20102
rect 15785 20091 16093 20100
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15764 19281 15792 19654
rect 15750 19272 15806 19281
rect 15750 19207 15806 19216
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 15785 19068 16093 19077
rect 15785 19066 15791 19068
rect 15847 19066 15871 19068
rect 15927 19066 15951 19068
rect 16007 19066 16031 19068
rect 16087 19066 16093 19068
rect 15847 19014 15849 19066
rect 16029 19014 16031 19066
rect 15785 19012 15791 19014
rect 15847 19012 15871 19014
rect 15927 19012 15951 19014
rect 16007 19012 16031 19014
rect 16087 19012 16093 19014
rect 15785 19003 16093 19012
rect 16132 18193 16160 19110
rect 15934 18184 15990 18193
rect 15934 18119 15990 18128
rect 16118 18184 16174 18193
rect 16118 18119 16174 18128
rect 15948 18086 15976 18119
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 15785 17980 16093 17989
rect 15785 17978 15791 17980
rect 15847 17978 15871 17980
rect 15927 17978 15951 17980
rect 16007 17978 16031 17980
rect 16087 17978 16093 17980
rect 15847 17926 15849 17978
rect 16029 17926 16031 17978
rect 15785 17924 15791 17926
rect 15847 17924 15871 17926
rect 15927 17924 15951 17926
rect 16007 17924 16031 17926
rect 16087 17924 16093 17926
rect 15785 17915 16093 17924
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 15785 16892 16093 16901
rect 15785 16890 15791 16892
rect 15847 16890 15871 16892
rect 15927 16890 15951 16892
rect 16007 16890 16031 16892
rect 16087 16890 16093 16892
rect 15847 16838 15849 16890
rect 16029 16838 16031 16890
rect 15785 16836 15791 16838
rect 15847 16836 15871 16838
rect 15927 16836 15951 16838
rect 16007 16836 16031 16838
rect 16087 16836 16093 16838
rect 15785 16827 16093 16836
rect 16132 16794 16160 16934
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15488 13462 15516 15302
rect 15580 13530 15608 15370
rect 15568 13524 15620 13530
rect 15672 13512 15700 16730
rect 16028 16652 16080 16658
rect 16080 16612 16160 16640
rect 16028 16594 16080 16600
rect 15785 15804 16093 15813
rect 15785 15802 15791 15804
rect 15847 15802 15871 15804
rect 15927 15802 15951 15804
rect 16007 15802 16031 15804
rect 16087 15802 16093 15804
rect 15847 15750 15849 15802
rect 16029 15750 16031 15802
rect 15785 15748 15791 15750
rect 15847 15748 15871 15750
rect 15927 15748 15951 15750
rect 16007 15748 16031 15750
rect 16087 15748 16093 15750
rect 15785 15739 16093 15748
rect 15785 14716 16093 14725
rect 15785 14714 15791 14716
rect 15847 14714 15871 14716
rect 15927 14714 15951 14716
rect 16007 14714 16031 14716
rect 16087 14714 16093 14716
rect 15847 14662 15849 14714
rect 16029 14662 16031 14714
rect 15785 14660 15791 14662
rect 15847 14660 15871 14662
rect 15927 14660 15951 14662
rect 16007 14660 16031 14662
rect 16087 14660 16093 14662
rect 15785 14651 16093 14660
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15856 13938 15884 14214
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15785 13628 16093 13637
rect 15785 13626 15791 13628
rect 15847 13626 15871 13628
rect 15927 13626 15951 13628
rect 16007 13626 16031 13628
rect 16087 13626 16093 13628
rect 15847 13574 15849 13626
rect 16029 13574 16031 13626
rect 15785 13572 15791 13574
rect 15847 13572 15871 13574
rect 15927 13572 15951 13574
rect 16007 13572 16031 13574
rect 16087 13572 16093 13574
rect 15785 13563 16093 13572
rect 15672 13484 16068 13512
rect 15568 13466 15620 13472
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15396 13280 15516 13308
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15396 12918 15424 13126
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15212 9330 15240 11086
rect 15304 10810 15332 11154
rect 15396 11150 15424 12242
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15290 10568 15346 10577
rect 15290 10503 15346 10512
rect 15304 10470 15332 10503
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15212 9302 15332 9330
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15212 5710 15240 7822
rect 15304 7206 15332 9302
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15304 6390 15332 6734
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15292 5704 15344 5710
rect 15396 5692 15424 11086
rect 15488 9674 15516 13280
rect 15672 12646 15700 13330
rect 16040 13172 16068 13484
rect 16132 13274 16160 16612
rect 16224 16114 16252 24262
rect 16304 24200 16356 24206
rect 16304 24142 16356 24148
rect 16316 23118 16344 24142
rect 16304 23112 16356 23118
rect 16304 23054 16356 23060
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 16316 17202 16344 22578
rect 16408 21486 16436 26030
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 16500 21350 16528 28358
rect 16592 26518 16620 28358
rect 16684 26790 16712 31758
rect 16868 31742 17080 31770
rect 16764 31680 16816 31686
rect 16764 31622 16816 31628
rect 16776 28801 16804 31622
rect 16762 28792 16818 28801
rect 16762 28727 16818 28736
rect 16672 26784 16724 26790
rect 16672 26726 16724 26732
rect 16776 26738 16804 28727
rect 16868 28082 16896 31742
rect 17040 29572 17092 29578
rect 17040 29514 17092 29520
rect 16948 29164 17000 29170
rect 16948 29106 17000 29112
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 16868 26897 16896 28018
rect 16854 26888 16910 26897
rect 16854 26823 16910 26832
rect 16684 26602 16712 26726
rect 16776 26710 16896 26738
rect 16684 26574 16804 26602
rect 16580 26512 16632 26518
rect 16580 26454 16632 26460
rect 16776 26450 16804 26574
rect 16672 26444 16724 26450
rect 16672 26386 16724 26392
rect 16764 26444 16816 26450
rect 16764 26386 16816 26392
rect 16684 26042 16712 26386
rect 16868 26330 16896 26710
rect 16776 26302 16896 26330
rect 16672 26036 16724 26042
rect 16672 25978 16724 25984
rect 16580 25356 16632 25362
rect 16580 25298 16632 25304
rect 16592 25158 16620 25298
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16592 23866 16620 25094
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 16580 23520 16632 23526
rect 16580 23462 16632 23468
rect 16670 23488 16726 23497
rect 16592 23118 16620 23462
rect 16670 23423 16726 23432
rect 16580 23112 16632 23118
rect 16580 23054 16632 23060
rect 16684 22930 16712 23423
rect 16592 22902 16712 22930
rect 16488 21344 16540 21350
rect 16488 21286 16540 21292
rect 16394 21040 16450 21049
rect 16394 20975 16450 20984
rect 16408 18970 16436 20975
rect 16488 20596 16540 20602
rect 16488 20538 16540 20544
rect 16500 19854 16528 20538
rect 16488 19848 16540 19854
rect 16592 19825 16620 22902
rect 16672 22772 16724 22778
rect 16672 22714 16724 22720
rect 16684 21554 16712 22714
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16488 19790 16540 19796
rect 16578 19816 16634 19825
rect 16500 19446 16528 19790
rect 16578 19751 16634 19760
rect 16488 19440 16540 19446
rect 16488 19382 16540 19388
rect 16684 19310 16712 21082
rect 16776 20942 16804 26302
rect 16856 24676 16908 24682
rect 16856 24618 16908 24624
rect 16868 24274 16896 24618
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16868 23866 16896 24006
rect 16856 23860 16908 23866
rect 16856 23802 16908 23808
rect 16856 21480 16908 21486
rect 16856 21422 16908 21428
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16500 18970 16528 19110
rect 16396 18964 16448 18970
rect 16396 18906 16448 18912
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16396 18828 16448 18834
rect 16396 18770 16448 18776
rect 16408 18426 16436 18770
rect 16684 18630 16712 19246
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16396 18420 16448 18426
rect 16396 18362 16448 18368
rect 16776 17954 16804 20878
rect 16868 19514 16896 21422
rect 16960 20330 16988 29106
rect 17052 29102 17080 29514
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 17052 28150 17080 29038
rect 17236 28994 17264 31980
rect 17316 31962 17368 31968
rect 17316 30320 17368 30326
rect 17316 30262 17368 30268
rect 17144 28966 17264 28994
rect 17040 28144 17092 28150
rect 17040 28086 17092 28092
rect 17040 27532 17092 27538
rect 17040 27474 17092 27480
rect 17052 26382 17080 27474
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 17052 22778 17080 26318
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 17052 21078 17080 21286
rect 17040 21072 17092 21078
rect 17040 21014 17092 21020
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 17052 19922 17080 20402
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16868 19394 16896 19450
rect 16868 19366 16988 19394
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16684 17926 16804 17954
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16304 17196 16356 17202
rect 16356 17156 16528 17184
rect 16304 17138 16356 17144
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16224 14618 16252 14894
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16316 14074 16344 16934
rect 16408 16590 16436 17002
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16316 13938 16344 14010
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 13462 16252 13670
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16408 13274 16436 15506
rect 16132 13246 16252 13274
rect 16040 13144 16160 13172
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15580 12238 15608 12582
rect 15672 12442 15700 12582
rect 15785 12540 16093 12549
rect 15785 12538 15791 12540
rect 15847 12538 15871 12540
rect 15927 12538 15951 12540
rect 16007 12538 16031 12540
rect 16087 12538 16093 12540
rect 15847 12486 15849 12538
rect 16029 12486 16031 12538
rect 15785 12484 15791 12486
rect 15847 12484 15871 12486
rect 15927 12484 15951 12486
rect 16007 12484 16031 12486
rect 16087 12484 16093 12486
rect 15785 12475 16093 12484
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15785 11452 16093 11461
rect 15785 11450 15791 11452
rect 15847 11450 15871 11452
rect 15927 11450 15951 11452
rect 16007 11450 16031 11452
rect 16087 11450 16093 11452
rect 15847 11398 15849 11450
rect 16029 11398 16031 11450
rect 15785 11396 15791 11398
rect 15847 11396 15871 11398
rect 15927 11396 15951 11398
rect 16007 11396 16031 11398
rect 16087 11396 16093 11398
rect 15785 11387 16093 11396
rect 16132 11268 16160 13144
rect 16224 11370 16252 13246
rect 16316 13246 16436 13274
rect 16316 12442 16344 13246
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16408 12322 16436 13126
rect 16316 12306 16436 12322
rect 16304 12300 16436 12306
rect 16356 12294 16436 12300
rect 16304 12242 16356 12248
rect 16500 11762 16528 17156
rect 16592 15094 16620 17478
rect 16684 16794 16712 17926
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16684 15366 16712 16730
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16580 15088 16632 15094
rect 16580 15030 16632 15036
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16592 13326 16620 13466
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16592 12918 16620 13262
rect 16580 12912 16632 12918
rect 16580 12854 16632 12860
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16224 11342 16528 11370
rect 16026 11248 16082 11257
rect 15844 11212 15896 11218
rect 16132 11240 16436 11268
rect 16026 11183 16082 11192
rect 15844 11154 15896 11160
rect 15856 10810 15884 11154
rect 16040 11132 16068 11183
rect 16120 11144 16172 11150
rect 16040 11104 16120 11132
rect 16172 11104 16344 11132
rect 16120 11086 16172 11092
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15568 10668 15620 10674
rect 15620 10628 15700 10656
rect 15568 10610 15620 10616
rect 15488 9646 15608 9674
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15488 7886 15516 8910
rect 15580 8906 15608 9646
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15580 6458 15608 7142
rect 15672 6798 15700 10628
rect 15785 10364 16093 10373
rect 15785 10362 15791 10364
rect 15847 10362 15871 10364
rect 15927 10362 15951 10364
rect 16007 10362 16031 10364
rect 16087 10362 16093 10364
rect 15847 10310 15849 10362
rect 16029 10310 16031 10362
rect 15785 10308 15791 10310
rect 15847 10308 15871 10310
rect 15927 10308 15951 10310
rect 16007 10308 16031 10310
rect 16087 10308 16093 10310
rect 15785 10299 16093 10308
rect 15785 9276 16093 9285
rect 15785 9274 15791 9276
rect 15847 9274 15871 9276
rect 15927 9274 15951 9276
rect 16007 9274 16031 9276
rect 16087 9274 16093 9276
rect 15847 9222 15849 9274
rect 16029 9222 16031 9274
rect 15785 9220 15791 9222
rect 15847 9220 15871 9222
rect 15927 9220 15951 9222
rect 16007 9220 16031 9222
rect 16087 9220 16093 9222
rect 15785 9211 16093 9220
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 15785 8188 16093 8197
rect 15785 8186 15791 8188
rect 15847 8186 15871 8188
rect 15927 8186 15951 8188
rect 16007 8186 16031 8188
rect 16087 8186 16093 8188
rect 15847 8134 15849 8186
rect 16029 8134 16031 8186
rect 15785 8132 15791 8134
rect 15847 8132 15871 8134
rect 15927 8132 15951 8134
rect 16007 8132 16031 8134
rect 16087 8132 16093 8134
rect 15785 8123 16093 8132
rect 16132 8022 16160 8774
rect 16120 8016 16172 8022
rect 16120 7958 16172 7964
rect 16316 7954 16344 11104
rect 16408 8362 16436 11240
rect 16500 9110 16528 11342
rect 16684 10810 16712 11630
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16670 10160 16726 10169
rect 16670 10095 16726 10104
rect 16578 10024 16634 10033
rect 16578 9959 16634 9968
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16408 7954 16436 8298
rect 16500 8090 16528 9046
rect 16592 8634 16620 9959
rect 16684 9654 16712 10095
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16684 8498 16712 9454
rect 16776 8634 16804 17478
rect 16868 13530 16896 18702
rect 16960 16182 16988 19366
rect 17144 17626 17172 28966
rect 17328 27606 17356 30262
rect 17420 29170 17448 33526
rect 17512 31822 17540 33646
rect 17592 33652 17644 33658
rect 17592 33594 17644 33600
rect 17592 32904 17644 32910
rect 17696 32892 17724 35566
rect 17644 32864 17724 32892
rect 17592 32846 17644 32852
rect 17500 31816 17552 31822
rect 17500 31758 17552 31764
rect 17500 30796 17552 30802
rect 17604 30784 17632 32846
rect 17788 31906 17816 36586
rect 17960 36032 18012 36038
rect 17960 35974 18012 35980
rect 17972 35698 18000 35974
rect 18156 35834 18184 36586
rect 18328 36304 18380 36310
rect 18328 36246 18380 36252
rect 18144 35828 18196 35834
rect 18144 35770 18196 35776
rect 17960 35692 18012 35698
rect 17960 35634 18012 35640
rect 17972 35034 18000 35634
rect 17880 35006 18000 35034
rect 18052 35080 18104 35086
rect 18052 35022 18104 35028
rect 17880 34950 17908 35006
rect 17868 34944 17920 34950
rect 17868 34886 17920 34892
rect 17866 34640 17922 34649
rect 17866 34575 17868 34584
rect 17920 34575 17922 34584
rect 17868 34546 17920 34552
rect 17960 33516 18012 33522
rect 17960 33458 18012 33464
rect 17972 32842 18000 33458
rect 18064 33114 18092 35022
rect 18156 34762 18184 35770
rect 18236 35012 18288 35018
rect 18236 34954 18288 34960
rect 18248 34921 18276 34954
rect 18234 34912 18290 34921
rect 18234 34847 18290 34856
rect 18156 34734 18276 34762
rect 18052 33108 18104 33114
rect 18052 33050 18104 33056
rect 17960 32836 18012 32842
rect 17960 32778 18012 32784
rect 18064 32502 18092 33050
rect 18142 32872 18198 32881
rect 18142 32807 18198 32816
rect 18052 32496 18104 32502
rect 18052 32438 18104 32444
rect 17868 32360 17920 32366
rect 17868 32302 17920 32308
rect 17552 30756 17632 30784
rect 17696 31878 17816 31906
rect 17500 30738 17552 30744
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 17500 28620 17552 28626
rect 17420 28580 17500 28608
rect 17316 27600 17368 27606
rect 17316 27542 17368 27548
rect 17420 27538 17448 28580
rect 17500 28562 17552 28568
rect 17498 28384 17554 28393
rect 17498 28319 17554 28328
rect 17408 27532 17460 27538
rect 17408 27474 17460 27480
rect 17512 27418 17540 28319
rect 17696 27674 17724 31878
rect 17776 31816 17828 31822
rect 17776 31758 17828 31764
rect 17788 31396 17816 31758
rect 17880 31498 17908 32302
rect 18156 31958 18184 32807
rect 18144 31952 18196 31958
rect 18144 31894 18196 31900
rect 17880 31470 18000 31498
rect 17788 31368 17908 31396
rect 17880 30580 17908 31368
rect 17788 30552 17908 30580
rect 17788 27713 17816 30552
rect 17972 30258 18000 31470
rect 18052 31476 18104 31482
rect 18052 31418 18104 31424
rect 17960 30252 18012 30258
rect 17960 30194 18012 30200
rect 17960 30048 18012 30054
rect 17960 29990 18012 29996
rect 17866 29200 17922 29209
rect 17866 29135 17868 29144
rect 17920 29135 17922 29144
rect 17868 29106 17920 29112
rect 17868 28688 17920 28694
rect 17868 28630 17920 28636
rect 17880 28218 17908 28630
rect 17868 28212 17920 28218
rect 17868 28154 17920 28160
rect 17868 27940 17920 27946
rect 17868 27882 17920 27888
rect 17774 27704 17830 27713
rect 17684 27668 17736 27674
rect 17774 27639 17830 27648
rect 17684 27610 17736 27616
rect 17592 27532 17644 27538
rect 17592 27474 17644 27480
rect 17328 27390 17540 27418
rect 17222 26888 17278 26897
rect 17222 26823 17278 26832
rect 17236 22001 17264 26823
rect 17328 22030 17356 27390
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 17420 26897 17448 26930
rect 17406 26888 17462 26897
rect 17406 26823 17462 26832
rect 17408 26784 17460 26790
rect 17408 26726 17460 26732
rect 17316 22024 17368 22030
rect 17222 21992 17278 22001
rect 17316 21966 17368 21972
rect 17222 21927 17278 21936
rect 17420 20942 17448 26726
rect 17500 25288 17552 25294
rect 17500 25230 17552 25236
rect 17512 24682 17540 25230
rect 17500 24676 17552 24682
rect 17500 24618 17552 24624
rect 17604 24426 17632 27474
rect 17880 27146 17908 27882
rect 17972 27282 18000 29990
rect 18064 27384 18092 31418
rect 18144 31340 18196 31346
rect 18144 31282 18196 31288
rect 18156 30734 18184 31282
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 18248 30258 18276 34734
rect 18340 31906 18368 36246
rect 18432 32026 18460 42026
rect 18524 41138 18552 43182
rect 18604 42832 18656 42838
rect 18604 42774 18656 42780
rect 18616 42226 18644 42774
rect 18752 42460 19060 42469
rect 18752 42458 18758 42460
rect 18814 42458 18838 42460
rect 18894 42458 18918 42460
rect 18974 42458 18998 42460
rect 19054 42458 19060 42460
rect 18814 42406 18816 42458
rect 18996 42406 18998 42458
rect 18752 42404 18758 42406
rect 18814 42404 18838 42406
rect 18894 42404 18918 42406
rect 18974 42404 18998 42406
rect 19054 42404 19060 42406
rect 18752 42395 19060 42404
rect 19168 42226 19196 43710
rect 19260 43246 19288 44840
rect 19432 43308 19484 43314
rect 19432 43250 19484 43256
rect 19248 43240 19300 43246
rect 19248 43182 19300 43188
rect 19340 43104 19392 43110
rect 19340 43046 19392 43052
rect 19248 42628 19300 42634
rect 19248 42570 19300 42576
rect 18604 42220 18656 42226
rect 18604 42162 18656 42168
rect 18880 42220 18932 42226
rect 18880 42162 18932 42168
rect 19156 42220 19208 42226
rect 19156 42162 19208 42168
rect 18696 42016 18748 42022
rect 18696 41958 18748 41964
rect 18708 41698 18736 41958
rect 18892 41818 18920 42162
rect 19064 42016 19116 42022
rect 19064 41958 19116 41964
rect 19076 41857 19104 41958
rect 19062 41848 19118 41857
rect 18880 41812 18932 41818
rect 19062 41783 19118 41792
rect 18880 41754 18932 41760
rect 18616 41670 18736 41698
rect 18512 41132 18564 41138
rect 18512 41074 18564 41080
rect 18616 38654 18644 41670
rect 18696 41608 18748 41614
rect 18694 41576 18696 41585
rect 18748 41576 18750 41585
rect 18694 41511 18750 41520
rect 19156 41472 19208 41478
rect 19156 41414 19208 41420
rect 18752 41372 19060 41381
rect 18752 41370 18758 41372
rect 18814 41370 18838 41372
rect 18894 41370 18918 41372
rect 18974 41370 18998 41372
rect 19054 41370 19060 41372
rect 18814 41318 18816 41370
rect 18996 41318 18998 41370
rect 18752 41316 18758 41318
rect 18814 41316 18838 41318
rect 18894 41316 18918 41318
rect 18974 41316 18998 41318
rect 19054 41316 19060 41318
rect 18752 41307 19060 41316
rect 19168 41206 19196 41414
rect 19156 41200 19208 41206
rect 19156 41142 19208 41148
rect 19156 40996 19208 41002
rect 19156 40938 19208 40944
rect 18752 40284 19060 40293
rect 18752 40282 18758 40284
rect 18814 40282 18838 40284
rect 18894 40282 18918 40284
rect 18974 40282 18998 40284
rect 19054 40282 19060 40284
rect 18814 40230 18816 40282
rect 18996 40230 18998 40282
rect 18752 40228 18758 40230
rect 18814 40228 18838 40230
rect 18894 40228 18918 40230
rect 18974 40228 18998 40230
rect 19054 40228 19060 40230
rect 18752 40219 19060 40228
rect 18752 39196 19060 39205
rect 18752 39194 18758 39196
rect 18814 39194 18838 39196
rect 18894 39194 18918 39196
rect 18974 39194 18998 39196
rect 19054 39194 19060 39196
rect 18814 39142 18816 39194
rect 18996 39142 18998 39194
rect 18752 39140 18758 39142
rect 18814 39140 18838 39142
rect 18894 39140 18918 39142
rect 18974 39140 18998 39142
rect 19054 39140 19060 39142
rect 18752 39131 19060 39140
rect 18524 38626 18644 38654
rect 18420 32020 18472 32026
rect 18420 31962 18472 31968
rect 18340 31878 18460 31906
rect 18326 31648 18382 31657
rect 18326 31583 18382 31592
rect 18236 30252 18288 30258
rect 18236 30194 18288 30200
rect 18236 30048 18288 30054
rect 18236 29990 18288 29996
rect 18248 28937 18276 29990
rect 18234 28928 18290 28937
rect 18234 28863 18290 28872
rect 18142 28792 18198 28801
rect 18142 28727 18198 28736
rect 18156 28626 18184 28727
rect 18144 28620 18196 28626
rect 18144 28562 18196 28568
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 18248 28393 18276 28494
rect 18234 28384 18290 28393
rect 18234 28319 18290 28328
rect 18340 28200 18368 31583
rect 18432 29209 18460 31878
rect 18418 29200 18474 29209
rect 18418 29135 18474 29144
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 18432 28558 18460 28902
rect 18420 28552 18472 28558
rect 18420 28494 18472 28500
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18432 28218 18460 28358
rect 18309 28172 18368 28200
rect 18420 28212 18472 28218
rect 18309 28064 18337 28172
rect 18420 28154 18472 28160
rect 18309 28036 18368 28064
rect 18234 27976 18290 27985
rect 18234 27911 18290 27920
rect 18248 27606 18276 27911
rect 18236 27600 18288 27606
rect 18236 27542 18288 27548
rect 18064 27356 18184 27384
rect 17972 27254 18092 27282
rect 17880 27118 18000 27146
rect 17684 26784 17736 26790
rect 17684 26726 17736 26732
rect 17696 26586 17724 26726
rect 17684 26580 17736 26586
rect 17684 26522 17736 26528
rect 17868 26376 17920 26382
rect 17868 26318 17920 26324
rect 17880 25974 17908 26318
rect 17868 25968 17920 25974
rect 17868 25910 17920 25916
rect 17972 25702 18000 27118
rect 17960 25696 18012 25702
rect 17960 25638 18012 25644
rect 18064 25378 18092 27254
rect 17880 25350 18092 25378
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17512 24410 17724 24426
rect 17500 24404 17724 24410
rect 17552 24398 17724 24404
rect 17500 24346 17552 24352
rect 17500 23656 17552 23662
rect 17500 23598 17552 23604
rect 17316 20936 17368 20942
rect 17316 20878 17368 20884
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17222 20768 17278 20777
rect 17222 20703 17278 20712
rect 17052 17598 17172 17626
rect 17052 17542 17080 17598
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17144 17241 17172 17478
rect 17130 17232 17186 17241
rect 17130 17167 17186 17176
rect 17040 16992 17092 16998
rect 17236 16980 17264 20703
rect 17328 17882 17356 20878
rect 17316 17876 17368 17882
rect 17316 17818 17368 17824
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17092 16952 17264 16980
rect 17040 16934 17092 16940
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 17052 16028 17080 16934
rect 17328 16794 17356 17614
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 16960 16000 17080 16028
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16868 10062 16896 12378
rect 16960 11898 16988 16000
rect 17328 15502 17356 16526
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17420 15162 17448 20878
rect 17512 20602 17540 23598
rect 17696 22094 17724 24398
rect 17788 23118 17816 24550
rect 17776 23112 17828 23118
rect 17776 23054 17828 23060
rect 17880 22166 17908 25350
rect 17960 25220 18012 25226
rect 17960 25162 18012 25168
rect 17972 24886 18000 25162
rect 17960 24880 18012 24886
rect 17960 24822 18012 24828
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17696 22066 17816 22094
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17696 21554 17724 21966
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17684 21344 17736 21350
rect 17684 21286 17736 21292
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17604 20602 17632 20878
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17592 20596 17644 20602
rect 17592 20538 17644 20544
rect 17498 20496 17554 20505
rect 17498 20431 17554 20440
rect 17512 19786 17540 20431
rect 17696 20369 17724 21286
rect 17682 20360 17738 20369
rect 17682 20295 17738 20304
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17590 19544 17646 19553
rect 17590 19479 17646 19488
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17512 17270 17540 18566
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17512 16522 17540 17070
rect 17500 16516 17552 16522
rect 17500 16458 17552 16464
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17040 14408 17092 14414
rect 17092 14368 17172 14396
rect 17040 14350 17092 14356
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 17052 11762 17080 12310
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16960 10810 16988 11018
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 17052 9738 17080 10746
rect 16868 9710 17080 9738
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16488 8084 16540 8090
rect 16868 8072 16896 9710
rect 17144 9674 17172 14368
rect 17316 13932 17368 13938
rect 17236 13892 17316 13920
rect 17236 11121 17264 13892
rect 17316 13874 17368 13880
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17328 11830 17356 12378
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 17222 11112 17278 11121
rect 17222 11047 17224 11056
rect 17276 11047 17278 11056
rect 17224 11018 17276 11024
rect 17236 9761 17264 11018
rect 17420 10146 17448 15098
rect 17512 13530 17540 15642
rect 17604 13938 17632 19479
rect 17788 19334 17816 22066
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 17880 20602 17908 21422
rect 17868 20596 17920 20602
rect 17868 20538 17920 20544
rect 17788 19306 17908 19334
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17696 18834 17724 19110
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17696 18329 17724 18634
rect 17682 18320 17738 18329
rect 17682 18255 17738 18264
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17696 16794 17724 16934
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17880 16454 17908 19306
rect 17972 18154 18000 24142
rect 18052 24064 18104 24070
rect 18052 24006 18104 24012
rect 18064 23730 18092 24006
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 18064 23118 18092 23666
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 18064 18714 18092 21422
rect 18156 18850 18184 27356
rect 18236 27124 18288 27130
rect 18236 27066 18288 27072
rect 18248 22710 18276 27066
rect 18340 24206 18368 28036
rect 18524 26874 18552 38626
rect 18752 38108 19060 38117
rect 18752 38106 18758 38108
rect 18814 38106 18838 38108
rect 18894 38106 18918 38108
rect 18974 38106 18998 38108
rect 19054 38106 19060 38108
rect 18814 38054 18816 38106
rect 18996 38054 18998 38106
rect 18752 38052 18758 38054
rect 18814 38052 18838 38054
rect 18894 38052 18918 38054
rect 18974 38052 18998 38054
rect 19054 38052 19060 38054
rect 18752 38043 19060 38052
rect 19168 37398 19196 40938
rect 19260 38418 19288 42570
rect 19352 42294 19380 43046
rect 19340 42288 19392 42294
rect 19340 42230 19392 42236
rect 19340 42016 19392 42022
rect 19338 41984 19340 41993
rect 19392 41984 19394 41993
rect 19338 41919 19394 41928
rect 19340 41812 19392 41818
rect 19340 41754 19392 41760
rect 19352 41614 19380 41754
rect 19340 41608 19392 41614
rect 19340 41550 19392 41556
rect 19444 41414 19472 43250
rect 19536 41614 19564 44840
rect 19708 42832 19760 42838
rect 19708 42774 19760 42780
rect 19616 42696 19668 42702
rect 19616 42638 19668 42644
rect 19628 42362 19656 42638
rect 19616 42356 19668 42362
rect 19616 42298 19668 42304
rect 19720 41818 19748 42774
rect 19708 41812 19760 41818
rect 19708 41754 19760 41760
rect 19812 41682 19840 44840
rect 19984 43648 20036 43654
rect 19984 43590 20036 43596
rect 19996 42362 20024 43590
rect 20076 43172 20128 43178
rect 20076 43114 20128 43120
rect 20088 42770 20116 43114
rect 20272 42906 20300 44934
rect 20350 44934 20484 44962
rect 20350 44840 20406 44934
rect 20456 43450 20484 44934
rect 20626 44840 20682 45000
rect 20902 44840 20958 45000
rect 21178 44840 21234 45000
rect 21454 44840 21510 45000
rect 21730 44962 21786 45000
rect 21730 44934 21956 44962
rect 21730 44840 21786 44934
rect 20640 43450 20668 44840
rect 20916 43466 20944 44840
rect 21192 44146 21220 44840
rect 21192 44118 21404 44146
rect 20444 43444 20496 43450
rect 20444 43386 20496 43392
rect 20628 43444 20680 43450
rect 20916 43438 21036 43466
rect 21376 43450 21404 44118
rect 20628 43386 20680 43392
rect 20352 43308 20404 43314
rect 20352 43250 20404 43256
rect 20904 43308 20956 43314
rect 20904 43250 20956 43256
rect 20260 42900 20312 42906
rect 20260 42842 20312 42848
rect 20076 42764 20128 42770
rect 20076 42706 20128 42712
rect 20168 42764 20220 42770
rect 20168 42706 20220 42712
rect 19984 42356 20036 42362
rect 19984 42298 20036 42304
rect 19984 42220 20036 42226
rect 19984 42162 20036 42168
rect 19892 42016 19944 42022
rect 19892 41958 19944 41964
rect 19800 41676 19852 41682
rect 19800 41618 19852 41624
rect 19904 41614 19932 41958
rect 19996 41818 20024 42162
rect 19984 41812 20036 41818
rect 19984 41754 20036 41760
rect 19524 41608 19576 41614
rect 19524 41550 19576 41556
rect 19892 41608 19944 41614
rect 19892 41550 19944 41556
rect 19444 41386 19656 41414
rect 19628 41274 19656 41386
rect 19616 41268 19668 41274
rect 19616 41210 19668 41216
rect 19432 40928 19484 40934
rect 19432 40870 19484 40876
rect 19444 40526 19472 40870
rect 20180 40730 20208 42706
rect 20364 42362 20392 43250
rect 20720 42560 20772 42566
rect 20720 42502 20772 42508
rect 20352 42356 20404 42362
rect 20352 42298 20404 42304
rect 20260 42288 20312 42294
rect 20260 42230 20312 42236
rect 20272 41478 20300 42230
rect 20444 42220 20496 42226
rect 20444 42162 20496 42168
rect 20456 41818 20484 42162
rect 20444 41812 20496 41818
rect 20444 41754 20496 41760
rect 20628 41608 20680 41614
rect 20628 41550 20680 41556
rect 20260 41472 20312 41478
rect 20260 41414 20312 41420
rect 20352 41472 20404 41478
rect 20352 41414 20404 41420
rect 20444 41472 20496 41478
rect 20444 41414 20496 41420
rect 20364 41274 20392 41414
rect 20352 41268 20404 41274
rect 20352 41210 20404 41216
rect 20352 41132 20404 41138
rect 20352 41074 20404 41080
rect 20168 40724 20220 40730
rect 20168 40666 20220 40672
rect 20258 40624 20314 40633
rect 20258 40559 20314 40568
rect 19432 40520 19484 40526
rect 19432 40462 19484 40468
rect 20076 40520 20128 40526
rect 20076 40462 20128 40468
rect 19432 40384 19484 40390
rect 19432 40326 19484 40332
rect 19892 40384 19944 40390
rect 19892 40326 19944 40332
rect 19444 40089 19472 40326
rect 19904 40225 19932 40326
rect 19890 40216 19946 40225
rect 19890 40151 19946 40160
rect 19430 40080 19486 40089
rect 19430 40015 19486 40024
rect 20088 39545 20116 40462
rect 20272 40186 20300 40559
rect 20260 40180 20312 40186
rect 20260 40122 20312 40128
rect 20168 40044 20220 40050
rect 20168 39986 20220 39992
rect 20180 39953 20208 39986
rect 20166 39944 20222 39953
rect 20166 39879 20222 39888
rect 20074 39536 20130 39545
rect 20074 39471 20130 39480
rect 20168 39432 20220 39438
rect 20168 39374 20220 39380
rect 19340 39364 19392 39370
rect 19340 39306 19392 39312
rect 19248 38412 19300 38418
rect 19248 38354 19300 38360
rect 19156 37392 19208 37398
rect 19156 37334 19208 37340
rect 19352 37330 19380 39306
rect 20180 39098 20208 39374
rect 20364 39114 20392 41074
rect 20456 40050 20484 41414
rect 20534 41304 20590 41313
rect 20640 41274 20668 41550
rect 20534 41239 20590 41248
rect 20628 41268 20680 41274
rect 20548 40934 20576 41239
rect 20628 41210 20680 41216
rect 20732 41154 20760 42502
rect 20916 42362 20944 43250
rect 21008 43110 21036 43438
rect 21364 43444 21416 43450
rect 21364 43386 21416 43392
rect 21468 43382 21496 44840
rect 21272 43376 21324 43382
rect 21272 43318 21324 43324
rect 21456 43376 21508 43382
rect 21456 43318 21508 43324
rect 21088 43308 21140 43314
rect 21088 43250 21140 43256
rect 20996 43104 21048 43110
rect 20996 43046 21048 43052
rect 20996 42628 21048 42634
rect 20996 42570 21048 42576
rect 20904 42356 20956 42362
rect 20904 42298 20956 42304
rect 21008 41818 21036 42570
rect 20996 41812 21048 41818
rect 20996 41754 21048 41760
rect 20994 41440 21050 41449
rect 20994 41375 21050 41384
rect 20640 41126 20760 41154
rect 20812 41132 20864 41138
rect 20536 40928 20588 40934
rect 20536 40870 20588 40876
rect 20534 40760 20590 40769
rect 20534 40695 20590 40704
rect 20548 40594 20576 40695
rect 20536 40588 20588 40594
rect 20536 40530 20588 40536
rect 20640 40118 20668 41126
rect 20812 41074 20864 41080
rect 20824 40610 20852 41074
rect 20902 41032 20958 41041
rect 20902 40967 20958 40976
rect 20916 40662 20944 40967
rect 21008 40662 21036 41375
rect 21100 40730 21128 43250
rect 21180 41608 21232 41614
rect 21180 41550 21232 41556
rect 21192 40934 21220 41550
rect 21284 41274 21312 43318
rect 21548 43308 21600 43314
rect 21548 43250 21600 43256
rect 21560 43058 21588 43250
rect 21928 43110 21956 44934
rect 22006 44840 22062 45000
rect 22282 44840 22338 45000
rect 22558 44840 22614 45000
rect 22834 44840 22890 45000
rect 23110 44840 23166 45000
rect 23386 44840 23442 45000
rect 23662 44840 23718 45000
rect 23938 44840 23994 45000
rect 24214 44840 24270 45000
rect 24490 44962 24546 45000
rect 24766 44962 24822 45000
rect 24320 44934 24546 44962
rect 21468 43030 21588 43058
rect 21916 43104 21968 43110
rect 22020 43092 22048 44840
rect 22100 43308 22152 43314
rect 22100 43250 22152 43256
rect 22112 43217 22140 43250
rect 22098 43208 22154 43217
rect 22098 43143 22154 43152
rect 22020 43064 22140 43092
rect 21916 43046 21968 43052
rect 21364 42696 21416 42702
rect 21364 42638 21416 42644
rect 21376 42129 21404 42638
rect 21362 42120 21418 42129
rect 21362 42055 21418 42064
rect 21468 41818 21496 43030
rect 21719 43004 22027 43013
rect 21719 43002 21725 43004
rect 21781 43002 21805 43004
rect 21861 43002 21885 43004
rect 21941 43002 21965 43004
rect 22021 43002 22027 43004
rect 21781 42950 21783 43002
rect 21963 42950 21965 43002
rect 21719 42948 21725 42950
rect 21781 42948 21805 42950
rect 21861 42948 21885 42950
rect 21941 42948 21965 42950
rect 22021 42948 22027 42950
rect 21719 42939 22027 42948
rect 21548 42900 21600 42906
rect 21548 42842 21600 42848
rect 21560 41834 21588 42842
rect 22112 42786 22140 43064
rect 22112 42758 22232 42786
rect 22296 42770 22324 44840
rect 22572 43314 22600 44840
rect 22652 43648 22704 43654
rect 22652 43590 22704 43596
rect 22664 43450 22692 43590
rect 22652 43444 22704 43450
rect 22652 43386 22704 43392
rect 22560 43308 22612 43314
rect 22560 43250 22612 43256
rect 22848 42786 22876 44840
rect 23018 43888 23074 43897
rect 23018 43823 23074 43832
rect 22928 42900 22980 42906
rect 22928 42842 22980 42848
rect 22940 42786 22968 42842
rect 22100 42288 22152 42294
rect 22100 42230 22152 42236
rect 21719 41916 22027 41925
rect 21719 41914 21725 41916
rect 21781 41914 21805 41916
rect 21861 41914 21885 41916
rect 21941 41914 21965 41916
rect 22021 41914 22027 41916
rect 21781 41862 21783 41914
rect 21963 41862 21965 41914
rect 21719 41860 21725 41862
rect 21781 41860 21805 41862
rect 21861 41860 21885 41862
rect 21941 41860 21965 41862
rect 22021 41860 22027 41862
rect 21719 41851 22027 41860
rect 21456 41812 21508 41818
rect 21560 41806 21680 41834
rect 21652 41800 21680 41806
rect 21732 41812 21784 41818
rect 21652 41772 21732 41800
rect 21456 41754 21508 41760
rect 21732 41754 21784 41760
rect 21548 41744 21600 41750
rect 21548 41686 21600 41692
rect 21272 41268 21324 41274
rect 21272 41210 21324 41216
rect 21456 41132 21508 41138
rect 21284 41092 21456 41120
rect 21180 40928 21232 40934
rect 21180 40870 21232 40876
rect 21284 40746 21312 41092
rect 21456 41074 21508 41080
rect 21364 40996 21416 41002
rect 21364 40938 21416 40944
rect 21088 40724 21140 40730
rect 21088 40666 21140 40672
rect 21192 40718 21312 40746
rect 20732 40582 20852 40610
rect 20904 40656 20956 40662
rect 20904 40598 20956 40604
rect 20996 40656 21048 40662
rect 20996 40598 21048 40604
rect 20732 40458 20760 40582
rect 20812 40520 20864 40526
rect 20812 40462 20864 40468
rect 20904 40520 20956 40526
rect 20904 40462 20956 40468
rect 21086 40488 21142 40497
rect 20720 40452 20772 40458
rect 20720 40394 20772 40400
rect 20824 40118 20852 40462
rect 20916 40186 20944 40462
rect 21086 40423 21142 40432
rect 20904 40180 20956 40186
rect 20904 40122 20956 40128
rect 20628 40112 20680 40118
rect 20628 40054 20680 40060
rect 20812 40112 20864 40118
rect 20812 40054 20864 40060
rect 20902 40080 20958 40089
rect 20444 40044 20496 40050
rect 20444 39986 20496 39992
rect 20720 40044 20772 40050
rect 21100 40050 21128 40423
rect 20902 40015 20958 40024
rect 21088 40044 21140 40050
rect 20720 39986 20772 39992
rect 20168 39092 20220 39098
rect 20168 39034 20220 39040
rect 20272 39086 20392 39114
rect 20732 39098 20760 39986
rect 20916 39914 20944 40015
rect 21088 39986 21140 39992
rect 20904 39908 20956 39914
rect 20904 39850 20956 39856
rect 20812 39568 20864 39574
rect 20812 39510 20864 39516
rect 20824 39273 20852 39510
rect 20810 39264 20866 39273
rect 20810 39199 20866 39208
rect 20720 39092 20772 39098
rect 19432 38956 19484 38962
rect 19432 38898 19484 38904
rect 19444 38554 19472 38898
rect 20272 38654 20300 39086
rect 20720 39034 20772 39040
rect 20352 38956 20404 38962
rect 20352 38898 20404 38904
rect 19996 38626 20300 38654
rect 19432 38548 19484 38554
rect 19432 38490 19484 38496
rect 19708 38412 19760 38418
rect 19708 38354 19760 38360
rect 19616 38344 19668 38350
rect 19616 38286 19668 38292
rect 19628 37466 19656 38286
rect 19616 37460 19668 37466
rect 19616 37402 19668 37408
rect 19340 37324 19392 37330
rect 19340 37266 19392 37272
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 18752 37020 19060 37029
rect 18752 37018 18758 37020
rect 18814 37018 18838 37020
rect 18894 37018 18918 37020
rect 18974 37018 18998 37020
rect 19054 37018 19060 37020
rect 18814 36966 18816 37018
rect 18996 36966 18998 37018
rect 18752 36964 18758 36966
rect 18814 36964 18838 36966
rect 18894 36964 18918 36966
rect 18974 36964 18998 36966
rect 19054 36964 19060 36966
rect 18752 36955 19060 36964
rect 19444 36922 19472 37198
rect 19432 36916 19484 36922
rect 19432 36858 19484 36864
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 19432 36168 19484 36174
rect 19432 36110 19484 36116
rect 18752 35932 19060 35941
rect 18752 35930 18758 35932
rect 18814 35930 18838 35932
rect 18894 35930 18918 35932
rect 18974 35930 18998 35932
rect 19054 35930 19060 35932
rect 18814 35878 18816 35930
rect 18996 35878 18998 35930
rect 18752 35876 18758 35878
rect 18814 35876 18838 35878
rect 18894 35876 18918 35878
rect 18974 35876 18998 35878
rect 19054 35876 19060 35878
rect 18752 35867 19060 35876
rect 19260 35698 19288 36110
rect 19340 36032 19392 36038
rect 19340 35974 19392 35980
rect 19156 35692 19208 35698
rect 19156 35634 19208 35640
rect 19248 35692 19300 35698
rect 19248 35634 19300 35640
rect 19168 35222 19196 35634
rect 19156 35216 19208 35222
rect 19156 35158 19208 35164
rect 19168 35086 19196 35158
rect 19352 35154 19380 35974
rect 19444 35834 19472 36110
rect 19720 35834 19748 38354
rect 19996 36310 20024 38626
rect 20364 38214 20392 38898
rect 20352 38208 20404 38214
rect 20352 38150 20404 38156
rect 21088 37868 21140 37874
rect 21088 37810 21140 37816
rect 20260 37800 20312 37806
rect 20260 37742 20312 37748
rect 20536 37800 20588 37806
rect 20536 37742 20588 37748
rect 19984 36304 20036 36310
rect 19984 36246 20036 36252
rect 19892 36032 19944 36038
rect 19892 35974 19944 35980
rect 19432 35828 19484 35834
rect 19432 35770 19484 35776
rect 19708 35828 19760 35834
rect 19708 35770 19760 35776
rect 19904 35766 19932 35974
rect 19892 35760 19944 35766
rect 19892 35702 19944 35708
rect 19432 35624 19484 35630
rect 19432 35566 19484 35572
rect 19444 35290 19472 35566
rect 19432 35284 19484 35290
rect 19432 35226 19484 35232
rect 19340 35148 19392 35154
rect 19340 35090 19392 35096
rect 19156 35080 19208 35086
rect 19156 35022 19208 35028
rect 19708 34944 19760 34950
rect 19708 34886 19760 34892
rect 18752 34844 19060 34853
rect 18752 34842 18758 34844
rect 18814 34842 18838 34844
rect 18894 34842 18918 34844
rect 18974 34842 18998 34844
rect 19054 34842 19060 34844
rect 18814 34790 18816 34842
rect 18996 34790 18998 34842
rect 18752 34788 18758 34790
rect 18814 34788 18838 34790
rect 18894 34788 18918 34790
rect 18974 34788 18998 34790
rect 19054 34788 19060 34790
rect 18752 34779 19060 34788
rect 19340 34672 19392 34678
rect 19340 34614 19392 34620
rect 19352 33998 19380 34614
rect 19432 34536 19484 34542
rect 19432 34478 19484 34484
rect 19340 33992 19392 33998
rect 19340 33934 19392 33940
rect 18752 33756 19060 33765
rect 18752 33754 18758 33756
rect 18814 33754 18838 33756
rect 18894 33754 18918 33756
rect 18974 33754 18998 33756
rect 19054 33754 19060 33756
rect 18814 33702 18816 33754
rect 18996 33702 18998 33754
rect 18752 33700 18758 33702
rect 18814 33700 18838 33702
rect 18894 33700 18918 33702
rect 18974 33700 18998 33702
rect 19054 33700 19060 33702
rect 18752 33691 19060 33700
rect 19156 33448 19208 33454
rect 19156 33390 19208 33396
rect 18604 33380 18656 33386
rect 18604 33322 18656 33328
rect 18616 31482 18644 33322
rect 18752 32668 19060 32677
rect 18752 32666 18758 32668
rect 18814 32666 18838 32668
rect 18894 32666 18918 32668
rect 18974 32666 18998 32668
rect 19054 32666 19060 32668
rect 18814 32614 18816 32666
rect 18996 32614 18998 32666
rect 18752 32612 18758 32614
rect 18814 32612 18838 32614
rect 18894 32612 18918 32614
rect 18974 32612 18998 32614
rect 19054 32612 19060 32614
rect 18752 32603 19060 32612
rect 19168 32570 19196 33390
rect 19340 33312 19392 33318
rect 19260 33272 19340 33300
rect 19260 33114 19288 33272
rect 19340 33254 19392 33260
rect 19248 33108 19300 33114
rect 19248 33050 19300 33056
rect 19340 32768 19392 32774
rect 19340 32710 19392 32716
rect 19156 32564 19208 32570
rect 19156 32506 19208 32512
rect 19352 32434 19380 32710
rect 19340 32428 19392 32434
rect 19340 32370 19392 32376
rect 19444 32366 19472 34478
rect 19524 33584 19576 33590
rect 19524 33526 19576 33532
rect 19536 32842 19564 33526
rect 19616 33516 19668 33522
rect 19616 33458 19668 33464
rect 19524 32836 19576 32842
rect 19524 32778 19576 32784
rect 19628 32570 19656 33458
rect 19616 32564 19668 32570
rect 19616 32506 19668 32512
rect 19720 32434 19748 34886
rect 20168 34604 20220 34610
rect 20168 34546 20220 34552
rect 19708 32428 19760 32434
rect 19708 32370 19760 32376
rect 20076 32428 20128 32434
rect 20076 32370 20128 32376
rect 19432 32360 19484 32366
rect 19432 32302 19484 32308
rect 19156 32020 19208 32026
rect 19156 31962 19208 31968
rect 18752 31580 19060 31589
rect 18752 31578 18758 31580
rect 18814 31578 18838 31580
rect 18894 31578 18918 31580
rect 18974 31578 18998 31580
rect 19054 31578 19060 31580
rect 18814 31526 18816 31578
rect 18996 31526 18998 31578
rect 18752 31524 18758 31526
rect 18814 31524 18838 31526
rect 18894 31524 18918 31526
rect 18974 31524 18998 31526
rect 19054 31524 19060 31526
rect 18752 31515 19060 31524
rect 18604 31476 18656 31482
rect 18604 31418 18656 31424
rect 18696 31204 18748 31210
rect 18696 31146 18748 31152
rect 18604 31136 18656 31142
rect 18604 31078 18656 31084
rect 18616 30938 18644 31078
rect 18604 30932 18656 30938
rect 18604 30874 18656 30880
rect 18708 30580 18736 31146
rect 18972 30864 19024 30870
rect 18972 30806 19024 30812
rect 18984 30666 19012 30806
rect 18972 30660 19024 30666
rect 18972 30602 19024 30608
rect 18616 30552 18736 30580
rect 18616 29288 18644 30552
rect 18752 30492 19060 30501
rect 18752 30490 18758 30492
rect 18814 30490 18838 30492
rect 18894 30490 18918 30492
rect 18974 30490 18998 30492
rect 19054 30490 19060 30492
rect 18814 30438 18816 30490
rect 18996 30438 18998 30490
rect 18752 30436 18758 30438
rect 18814 30436 18838 30438
rect 18894 30436 18918 30438
rect 18974 30436 18998 30438
rect 19054 30436 19060 30438
rect 18752 30427 19060 30436
rect 19064 30252 19116 30258
rect 19064 30194 19116 30200
rect 19076 29578 19104 30194
rect 19064 29572 19116 29578
rect 19064 29514 19116 29520
rect 18752 29404 19060 29413
rect 18752 29402 18758 29404
rect 18814 29402 18838 29404
rect 18894 29402 18918 29404
rect 18974 29402 18998 29404
rect 19054 29402 19060 29404
rect 18814 29350 18816 29402
rect 18996 29350 18998 29402
rect 18752 29348 18758 29350
rect 18814 29348 18838 29350
rect 18894 29348 18918 29350
rect 18974 29348 18998 29350
rect 19054 29348 19060 29350
rect 18752 29339 19060 29348
rect 18616 29260 18920 29288
rect 18694 29064 18750 29073
rect 18694 28999 18750 29008
rect 18604 28960 18656 28966
rect 18604 28902 18656 28908
rect 18616 28762 18644 28902
rect 18604 28756 18656 28762
rect 18604 28698 18656 28704
rect 18602 28656 18658 28665
rect 18602 28591 18604 28600
rect 18656 28591 18658 28600
rect 18604 28562 18656 28568
rect 18708 28472 18736 28999
rect 18432 26846 18552 26874
rect 18616 28444 18736 28472
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 18328 23588 18380 23594
rect 18328 23530 18380 23536
rect 18236 22704 18288 22710
rect 18236 22646 18288 22652
rect 18248 22030 18276 22646
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18248 20913 18276 20946
rect 18234 20904 18290 20913
rect 18234 20839 18290 20848
rect 18156 18822 18276 18850
rect 18064 18686 18184 18714
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 18064 18290 18092 18566
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 18064 17882 18092 18226
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17696 13394 17724 13670
rect 17880 13530 17908 16390
rect 17972 16114 18000 17614
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 18064 15910 18092 16390
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 18050 15192 18106 15201
rect 18050 15127 18106 15136
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17972 12782 18000 14962
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17500 12640 17552 12646
rect 18064 12628 18092 15127
rect 17500 12582 17552 12588
rect 17880 12600 18092 12628
rect 17512 12238 17540 12582
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17774 11792 17830 11801
rect 17684 11756 17736 11762
rect 17774 11727 17830 11736
rect 17684 11698 17736 11704
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17512 10742 17540 11630
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17420 10118 17632 10146
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17222 9752 17278 9761
rect 17222 9687 17278 9696
rect 17052 9646 17172 9674
rect 17224 9648 17276 9654
rect 17052 9586 17080 9646
rect 17224 9590 17276 9596
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17144 9178 17172 9318
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 17144 8634 17172 8978
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 16488 8026 16540 8032
rect 16776 8044 16896 8072
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 15785 7100 16093 7109
rect 15785 7098 15791 7100
rect 15847 7098 15871 7100
rect 15927 7098 15951 7100
rect 16007 7098 16031 7100
rect 16087 7098 16093 7100
rect 15847 7046 15849 7098
rect 16029 7046 16031 7098
rect 15785 7044 15791 7046
rect 15847 7044 15871 7046
rect 15927 7044 15951 7046
rect 16007 7044 16031 7046
rect 16087 7044 16093 7046
rect 15785 7035 16093 7044
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 16316 6361 16344 7890
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16592 7546 16620 7822
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16302 6352 16358 6361
rect 16302 6287 16358 6296
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15672 5914 15700 6054
rect 15785 6012 16093 6021
rect 15785 6010 15791 6012
rect 15847 6010 15871 6012
rect 15927 6010 15951 6012
rect 16007 6010 16031 6012
rect 16087 6010 16093 6012
rect 15847 5958 15849 6010
rect 16029 5958 16031 6010
rect 15785 5956 15791 5958
rect 15847 5956 15871 5958
rect 15927 5956 15951 5958
rect 16007 5956 16031 5958
rect 16087 5956 16093 5958
rect 15785 5947 16093 5956
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15344 5664 15424 5692
rect 15568 5704 15620 5710
rect 15292 5646 15344 5652
rect 15568 5646 15620 5652
rect 15212 4282 15240 5646
rect 15304 5370 15332 5646
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15580 4078 15608 5646
rect 15764 5012 15792 5850
rect 15672 4984 15792 5012
rect 15672 4146 15700 4984
rect 15785 4924 16093 4933
rect 15785 4922 15791 4924
rect 15847 4922 15871 4924
rect 15927 4922 15951 4924
rect 16007 4922 16031 4924
rect 16087 4922 16093 4924
rect 15847 4870 15849 4922
rect 16029 4870 16031 4922
rect 15785 4868 15791 4870
rect 15847 4868 15871 4870
rect 15927 4868 15951 4870
rect 16007 4868 16031 4870
rect 16087 4868 16093 4870
rect 15785 4859 16093 4868
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15396 3738 15424 3946
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15580 3466 15608 4014
rect 15785 3836 16093 3845
rect 15785 3834 15791 3836
rect 15847 3834 15871 3836
rect 15927 3834 15951 3836
rect 16007 3834 16031 3836
rect 16087 3834 16093 3836
rect 15847 3782 15849 3834
rect 16029 3782 16031 3834
rect 15785 3780 15791 3782
rect 15847 3780 15871 3782
rect 15927 3780 15951 3782
rect 16007 3780 16031 3782
rect 16087 3780 16093 3782
rect 15785 3771 16093 3780
rect 16132 3738 16160 6122
rect 16316 5914 16344 6287
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16316 5778 16344 5850
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 16302 4584 16358 4593
rect 16302 4519 16358 4528
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 16316 3058 16344 4519
rect 16408 3534 16436 7346
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16684 7177 16712 7278
rect 16670 7168 16726 7177
rect 16670 7103 16726 7112
rect 16486 6760 16542 6769
rect 16486 6695 16542 6704
rect 16500 6118 16528 6695
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16592 2854 16620 5306
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 15785 2748 16093 2757
rect 15785 2746 15791 2748
rect 15847 2746 15871 2748
rect 15927 2746 15951 2748
rect 16007 2746 16031 2748
rect 16087 2746 16093 2748
rect 15847 2694 15849 2746
rect 16029 2694 16031 2746
rect 15785 2692 15791 2694
rect 15847 2692 15871 2694
rect 15927 2692 15951 2694
rect 16007 2692 16031 2694
rect 16087 2692 16093 2694
rect 15474 2680 15530 2689
rect 15785 2683 16093 2692
rect 16776 2650 16804 8044
rect 16854 7984 16910 7993
rect 16854 7919 16910 7928
rect 16868 3058 16896 7919
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16960 4758 16988 4966
rect 16948 4752 17000 4758
rect 16948 4694 17000 4700
rect 17052 4604 17080 8570
rect 17236 6254 17264 9590
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17132 5772 17184 5778
rect 17236 5760 17264 6190
rect 17184 5732 17264 5760
rect 17132 5714 17184 5720
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17236 4622 17264 5102
rect 16960 4576 17080 4604
rect 17224 4616 17276 4622
rect 16960 3108 16988 4576
rect 17224 4558 17276 4564
rect 17328 4486 17356 9862
rect 17420 8974 17448 9998
rect 17604 9466 17632 10118
rect 17696 9994 17724 11698
rect 17788 11150 17816 11727
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17604 9438 17816 9466
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 9194 17724 9318
rect 17678 9166 17724 9194
rect 17678 9160 17706 9166
rect 17604 9132 17706 9160
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17500 8968 17552 8974
rect 17604 8956 17632 9132
rect 17684 8968 17736 8974
rect 17604 8928 17684 8956
rect 17500 8910 17552 8916
rect 17684 8910 17736 8916
rect 17420 8480 17448 8910
rect 17512 8820 17540 8910
rect 17788 8820 17816 9438
rect 17512 8809 17816 8820
rect 17498 8800 17816 8809
rect 17554 8792 17816 8800
rect 17498 8735 17554 8744
rect 17420 8452 17540 8480
rect 17406 8392 17462 8401
rect 17406 8327 17462 8336
rect 17420 5710 17448 8327
rect 17512 6662 17540 8452
rect 17880 7970 17908 12600
rect 18156 12434 18184 18686
rect 18248 16250 18276 18822
rect 18340 17241 18368 23530
rect 18432 22250 18460 26846
rect 18512 26240 18564 26246
rect 18512 26182 18564 26188
rect 18524 25974 18552 26182
rect 18512 25968 18564 25974
rect 18512 25910 18564 25916
rect 18616 25786 18644 28444
rect 18892 28422 18920 29260
rect 18880 28416 18932 28422
rect 18880 28358 18932 28364
rect 18752 28316 19060 28325
rect 18752 28314 18758 28316
rect 18814 28314 18838 28316
rect 18894 28314 18918 28316
rect 18974 28314 18998 28316
rect 19054 28314 19060 28316
rect 18814 28262 18816 28314
rect 18996 28262 18998 28314
rect 18752 28260 18758 28262
rect 18814 28260 18838 28262
rect 18894 28260 18918 28262
rect 18974 28260 18998 28262
rect 19054 28260 19060 28262
rect 18752 28251 19060 28260
rect 18696 28144 18748 28150
rect 18788 28144 18840 28150
rect 18696 28086 18748 28092
rect 18786 28112 18788 28121
rect 18840 28112 18842 28121
rect 18708 27538 18736 28086
rect 18786 28047 18842 28056
rect 18696 27532 18748 27538
rect 18696 27474 18748 27480
rect 18752 27228 19060 27237
rect 18752 27226 18758 27228
rect 18814 27226 18838 27228
rect 18894 27226 18918 27228
rect 18974 27226 18998 27228
rect 19054 27226 19060 27228
rect 18814 27174 18816 27226
rect 18996 27174 18998 27226
rect 18752 27172 18758 27174
rect 18814 27172 18838 27174
rect 18894 27172 18918 27174
rect 18974 27172 18998 27174
rect 19054 27172 19060 27174
rect 18752 27163 19060 27172
rect 18752 26140 19060 26149
rect 18752 26138 18758 26140
rect 18814 26138 18838 26140
rect 18894 26138 18918 26140
rect 18974 26138 18998 26140
rect 19054 26138 19060 26140
rect 18814 26086 18816 26138
rect 18996 26086 18998 26138
rect 18752 26084 18758 26086
rect 18814 26084 18838 26086
rect 18894 26084 18918 26086
rect 18974 26084 18998 26086
rect 19054 26084 19060 26086
rect 18752 26075 19060 26084
rect 18616 25758 18736 25786
rect 18512 25696 18564 25702
rect 18512 25638 18564 25644
rect 18604 25696 18656 25702
rect 18604 25638 18656 25644
rect 18524 24750 18552 25638
rect 18616 25498 18644 25638
rect 18604 25492 18656 25498
rect 18604 25434 18656 25440
rect 18708 25242 18736 25758
rect 18616 25214 18736 25242
rect 18512 24744 18564 24750
rect 18512 24686 18564 24692
rect 18524 22438 18552 24686
rect 18616 23848 18644 25214
rect 18752 25052 19060 25061
rect 18752 25050 18758 25052
rect 18814 25050 18838 25052
rect 18894 25050 18918 25052
rect 18974 25050 18998 25052
rect 19054 25050 19060 25052
rect 18814 24998 18816 25050
rect 18996 24998 18998 25050
rect 18752 24996 18758 24998
rect 18814 24996 18838 24998
rect 18894 24996 18918 24998
rect 18974 24996 18998 24998
rect 19054 24996 19060 24998
rect 18752 24987 19060 24996
rect 18788 24812 18840 24818
rect 18788 24754 18840 24760
rect 18800 24206 18828 24754
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18752 23964 19060 23973
rect 18752 23962 18758 23964
rect 18814 23962 18838 23964
rect 18894 23962 18918 23964
rect 18974 23962 18998 23964
rect 19054 23962 19060 23964
rect 18814 23910 18816 23962
rect 18996 23910 18998 23962
rect 18752 23908 18758 23910
rect 18814 23908 18838 23910
rect 18894 23908 18918 23910
rect 18974 23908 18998 23910
rect 19054 23908 19060 23910
rect 18752 23899 19060 23908
rect 18616 23820 18736 23848
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18616 23322 18644 23666
rect 18708 23497 18736 23820
rect 18786 23624 18842 23633
rect 18786 23559 18842 23568
rect 18800 23526 18828 23559
rect 18788 23520 18840 23526
rect 18694 23488 18750 23497
rect 18788 23462 18840 23468
rect 18694 23423 18750 23432
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 18752 22876 19060 22885
rect 18752 22874 18758 22876
rect 18814 22874 18838 22876
rect 18894 22874 18918 22876
rect 18974 22874 18998 22876
rect 19054 22874 19060 22876
rect 18814 22822 18816 22874
rect 18996 22822 18998 22874
rect 18752 22820 18758 22822
rect 18814 22820 18838 22822
rect 18894 22820 18918 22822
rect 18974 22820 18998 22822
rect 19054 22820 19060 22822
rect 18752 22811 19060 22820
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 18432 22222 18552 22250
rect 18420 22160 18472 22166
rect 18420 22102 18472 22108
rect 18432 17252 18460 22102
rect 18524 22094 18552 22222
rect 18524 22066 18644 22094
rect 18616 21486 18644 22066
rect 18752 21788 19060 21797
rect 18752 21786 18758 21788
rect 18814 21786 18838 21788
rect 18894 21786 18918 21788
rect 18974 21786 18998 21788
rect 19054 21786 19060 21788
rect 18814 21734 18816 21786
rect 18996 21734 18998 21786
rect 18752 21732 18758 21734
rect 18814 21732 18838 21734
rect 18894 21732 18918 21734
rect 18974 21732 18998 21734
rect 19054 21732 19060 21734
rect 18752 21723 19060 21732
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18524 20942 18552 21286
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18524 20602 18552 20742
rect 18512 20596 18564 20602
rect 18512 20538 18564 20544
rect 18616 20466 18644 21082
rect 18970 21040 19026 21049
rect 18970 20975 18972 20984
rect 19024 20975 19026 20984
rect 18972 20946 19024 20952
rect 19076 20913 19104 21082
rect 19062 20904 19118 20913
rect 19062 20839 19118 20848
rect 18752 20700 19060 20709
rect 18752 20698 18758 20700
rect 18814 20698 18838 20700
rect 18894 20698 18918 20700
rect 18974 20698 18998 20700
rect 19054 20698 19060 20700
rect 18814 20646 18816 20698
rect 18996 20646 18998 20698
rect 18752 20644 18758 20646
rect 18814 20644 18838 20646
rect 18894 20644 18918 20646
rect 18974 20644 18998 20646
rect 19054 20644 19060 20646
rect 18752 20635 19060 20644
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18524 20058 18552 20402
rect 19064 20324 19116 20330
rect 19064 20266 19116 20272
rect 19076 20058 19104 20266
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 18752 19612 19060 19621
rect 18752 19610 18758 19612
rect 18814 19610 18838 19612
rect 18894 19610 18918 19612
rect 18974 19610 18998 19612
rect 19054 19610 19060 19612
rect 18814 19558 18816 19610
rect 18996 19558 18998 19610
rect 18752 19556 18758 19558
rect 18814 19556 18838 19558
rect 18894 19556 18918 19558
rect 18974 19556 18998 19558
rect 19054 19556 19060 19558
rect 18752 19547 19060 19556
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18326 17232 18382 17241
rect 18432 17224 18552 17252
rect 18326 17167 18382 17176
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18248 13938 18276 14554
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 17604 7942 17908 7970
rect 17972 12406 18184 12434
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17512 5710 17540 6054
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17420 5234 17448 5646
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 17052 3738 17080 4014
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 17604 3534 17632 7942
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17880 5166 17908 6734
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17682 4040 17738 4049
rect 17682 3975 17738 3984
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17132 3460 17184 3466
rect 17132 3402 17184 3408
rect 17040 3120 17092 3126
rect 16960 3080 17040 3108
rect 17040 3062 17092 3068
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 15474 2615 15530 2624
rect 16764 2644 16816 2650
rect 15488 2446 15516 2615
rect 16764 2586 16816 2592
rect 16026 2544 16082 2553
rect 16026 2479 16082 2488
rect 16040 2446 16068 2479
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 14568 1290 14596 2246
rect 14936 2106 14964 2246
rect 15856 2106 15884 2246
rect 14924 2100 14976 2106
rect 14924 2042 14976 2048
rect 15844 2100 15896 2106
rect 15844 2042 15896 2048
rect 16120 1964 16172 1970
rect 16120 1906 16172 1912
rect 15384 1828 15436 1834
rect 15384 1770 15436 1776
rect 14740 1760 14792 1766
rect 14740 1702 14792 1708
rect 14556 1284 14608 1290
rect 14556 1226 14608 1232
rect 14372 1012 14424 1018
rect 14372 954 14424 960
rect 13174 54 13400 82
rect 13174 0 13230 54
rect 13450 0 13506 160
rect 13726 0 13782 160
rect 14002 0 14058 160
rect 14278 0 14334 160
rect 14554 82 14610 160
rect 14752 82 14780 1702
rect 14924 1556 14976 1562
rect 14924 1498 14976 1504
rect 14936 626 14964 1498
rect 15200 1488 15252 1494
rect 14844 598 14964 626
rect 15120 1436 15200 1442
rect 15120 1430 15252 1436
rect 15120 1414 15240 1430
rect 14844 160 14872 598
rect 15120 160 15148 1414
rect 15396 160 15424 1770
rect 15752 1760 15804 1766
rect 15672 1720 15752 1748
rect 15672 160 15700 1720
rect 15752 1702 15804 1708
rect 15785 1660 16093 1669
rect 15785 1658 15791 1660
rect 15847 1658 15871 1660
rect 15927 1658 15951 1660
rect 16007 1658 16031 1660
rect 16087 1658 16093 1660
rect 15847 1606 15849 1658
rect 16029 1606 16031 1658
rect 15785 1604 15791 1606
rect 15847 1604 15871 1606
rect 15927 1604 15951 1606
rect 16007 1604 16031 1606
rect 16087 1604 16093 1606
rect 15785 1595 16093 1604
rect 16132 1562 16160 1906
rect 16120 1556 16172 1562
rect 16120 1498 16172 1504
rect 16028 1488 16080 1494
rect 16028 1430 16080 1436
rect 14554 54 14780 82
rect 14554 0 14610 54
rect 14830 0 14886 160
rect 15106 0 15162 160
rect 15382 0 15438 160
rect 15658 0 15714 160
rect 15934 82 15990 160
rect 16040 82 16068 1430
rect 16212 1420 16264 1426
rect 16212 1362 16264 1368
rect 16224 160 16252 1362
rect 16684 1358 16712 2246
rect 16868 1970 16896 2790
rect 16946 2544 17002 2553
rect 16946 2479 16948 2488
rect 17000 2479 17002 2488
rect 16948 2450 17000 2456
rect 17144 2310 17172 3402
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17316 2916 17368 2922
rect 17316 2858 17368 2864
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 16856 1964 16908 1970
rect 16856 1906 16908 1912
rect 17132 1828 17184 1834
rect 17052 1788 17132 1816
rect 16856 1760 16908 1766
rect 16856 1702 16908 1708
rect 16488 1352 16540 1358
rect 16486 1320 16488 1329
rect 16672 1352 16724 1358
rect 16540 1320 16542 1329
rect 16672 1294 16724 1300
rect 16486 1255 16542 1264
rect 16488 1216 16540 1222
rect 16488 1158 16540 1164
rect 16500 160 16528 1158
rect 15934 54 16068 82
rect 15934 0 15990 54
rect 16210 0 16266 160
rect 16486 0 16542 160
rect 16762 82 16818 160
rect 16868 82 16896 1702
rect 17052 160 17080 1788
rect 17132 1770 17184 1776
rect 17236 1358 17264 2790
rect 17328 2446 17356 2858
rect 17512 2774 17540 3334
rect 17696 3058 17724 3975
rect 17866 3496 17922 3505
rect 17866 3431 17868 3440
rect 17920 3431 17922 3440
rect 17868 3402 17920 3408
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 17880 2802 17908 2994
rect 17972 2922 18000 12406
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 18064 10742 18092 12038
rect 18156 11898 18184 12242
rect 18248 12186 18276 13466
rect 18340 12374 18368 16662
rect 18432 16046 18460 16934
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 18432 12986 18460 13194
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18328 12368 18380 12374
rect 18326 12336 18328 12345
rect 18380 12336 18382 12345
rect 18326 12271 18382 12280
rect 18248 12158 18368 12186
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18248 11082 18276 12038
rect 18340 11898 18368 12158
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 8498 18092 9454
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 18326 9072 18382 9081
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 17960 2916 18012 2922
rect 17960 2858 18012 2864
rect 18064 2802 18092 5510
rect 18156 5302 18184 9046
rect 18326 9007 18328 9016
rect 18380 9007 18382 9016
rect 18328 8978 18380 8984
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18248 7002 18276 7346
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18340 6662 18368 7278
rect 18420 7200 18472 7206
rect 18418 7168 18420 7177
rect 18472 7168 18474 7177
rect 18418 7103 18474 7112
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18248 4214 18276 4422
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18156 3602 18184 4014
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 18248 3534 18276 4150
rect 18524 4146 18552 17224
rect 18616 13920 18644 19110
rect 18752 18524 19060 18533
rect 18752 18522 18758 18524
rect 18814 18522 18838 18524
rect 18894 18522 18918 18524
rect 18974 18522 18998 18524
rect 19054 18522 19060 18524
rect 18814 18470 18816 18522
rect 18996 18470 18998 18522
rect 18752 18468 18758 18470
rect 18814 18468 18838 18470
rect 18894 18468 18918 18470
rect 18974 18468 18998 18470
rect 19054 18468 19060 18470
rect 18752 18459 19060 18468
rect 19064 17808 19116 17814
rect 19064 17750 19116 17756
rect 19076 17542 19104 17750
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 18752 17436 19060 17445
rect 18752 17434 18758 17436
rect 18814 17434 18838 17436
rect 18894 17434 18918 17436
rect 18974 17434 18998 17436
rect 19054 17434 19060 17436
rect 18814 17382 18816 17434
rect 18996 17382 18998 17434
rect 18752 17380 18758 17382
rect 18814 17380 18838 17382
rect 18894 17380 18918 17382
rect 18974 17380 18998 17382
rect 19054 17380 19060 17382
rect 18752 17371 19060 17380
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18708 16726 18736 17138
rect 18696 16720 18748 16726
rect 18696 16662 18748 16668
rect 18752 16348 19060 16357
rect 18752 16346 18758 16348
rect 18814 16346 18838 16348
rect 18894 16346 18918 16348
rect 18974 16346 18998 16348
rect 19054 16346 19060 16348
rect 18814 16294 18816 16346
rect 18996 16294 18998 16346
rect 18752 16292 18758 16294
rect 18814 16292 18838 16294
rect 18894 16292 18918 16294
rect 18974 16292 18998 16294
rect 19054 16292 19060 16294
rect 18752 16283 19060 16292
rect 18752 15260 19060 15269
rect 18752 15258 18758 15260
rect 18814 15258 18838 15260
rect 18894 15258 18918 15260
rect 18974 15258 18998 15260
rect 19054 15258 19060 15260
rect 18814 15206 18816 15258
rect 18996 15206 18998 15258
rect 18752 15204 18758 15206
rect 18814 15204 18838 15206
rect 18894 15204 18918 15206
rect 18974 15204 18998 15206
rect 19054 15204 19060 15206
rect 18752 15195 19060 15204
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18800 14482 18828 14962
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 19168 14362 19196 31962
rect 19720 31754 19748 32370
rect 19720 31726 19840 31754
rect 19708 31272 19760 31278
rect 19708 31214 19760 31220
rect 19248 30592 19300 30598
rect 19248 30534 19300 30540
rect 19340 30592 19392 30598
rect 19340 30534 19392 30540
rect 19616 30592 19668 30598
rect 19616 30534 19668 30540
rect 19260 30394 19288 30534
rect 19248 30388 19300 30394
rect 19248 30330 19300 30336
rect 19260 29646 19288 30330
rect 19352 29850 19380 30534
rect 19628 29850 19656 30534
rect 19340 29844 19392 29850
rect 19340 29786 19392 29792
rect 19616 29844 19668 29850
rect 19616 29786 19668 29792
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19432 29640 19484 29646
rect 19432 29582 19484 29588
rect 19248 29504 19300 29510
rect 19248 29446 19300 29452
rect 19260 28762 19288 29446
rect 19248 28756 19300 28762
rect 19248 28698 19300 28704
rect 19340 28756 19392 28762
rect 19340 28698 19392 28704
rect 19248 28416 19300 28422
rect 19248 28358 19300 28364
rect 19260 26858 19288 28358
rect 19352 27878 19380 28698
rect 19444 28014 19472 29582
rect 19524 29504 19576 29510
rect 19524 29446 19576 29452
rect 19432 28008 19484 28014
rect 19432 27950 19484 27956
rect 19340 27872 19392 27878
rect 19340 27814 19392 27820
rect 19248 26852 19300 26858
rect 19248 26794 19300 26800
rect 19352 26194 19380 27814
rect 19352 26166 19472 26194
rect 19248 25696 19300 25702
rect 19248 25638 19300 25644
rect 19260 25498 19288 25638
rect 19248 25492 19300 25498
rect 19248 25434 19300 25440
rect 19338 25256 19394 25265
rect 19338 25191 19394 25200
rect 19248 24880 19300 24886
rect 19248 24822 19300 24828
rect 19260 22642 19288 24822
rect 19352 23322 19380 25191
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 19260 22094 19288 22374
rect 19260 22066 19380 22094
rect 19352 20482 19380 22066
rect 19444 20890 19472 26166
rect 19536 23050 19564 29446
rect 19614 28248 19670 28257
rect 19614 28183 19670 28192
rect 19628 28150 19656 28183
rect 19616 28144 19668 28150
rect 19616 28086 19668 28092
rect 19720 24018 19748 31214
rect 19812 29782 19840 31726
rect 20088 30870 20116 32370
rect 20076 30864 20128 30870
rect 20076 30806 20128 30812
rect 19800 29776 19852 29782
rect 19800 29718 19852 29724
rect 20180 29646 20208 34546
rect 20272 34406 20300 37742
rect 20352 37256 20404 37262
rect 20352 37198 20404 37204
rect 20364 36922 20392 37198
rect 20352 36916 20404 36922
rect 20352 36858 20404 36864
rect 20352 36236 20404 36242
rect 20352 36178 20404 36184
rect 20260 34400 20312 34406
rect 20260 34342 20312 34348
rect 20260 33992 20312 33998
rect 20260 33934 20312 33940
rect 20168 29640 20220 29646
rect 20168 29582 20220 29588
rect 20180 28994 20208 29582
rect 19996 28966 20208 28994
rect 19800 28552 19852 28558
rect 19800 28494 19852 28500
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 19812 27878 19840 28494
rect 19904 28218 19932 28494
rect 19892 28212 19944 28218
rect 19892 28154 19944 28160
rect 19800 27872 19852 27878
rect 19800 27814 19852 27820
rect 19812 27470 19840 27814
rect 19800 27464 19852 27470
rect 19800 27406 19852 27412
rect 19996 26994 20024 28966
rect 20076 28416 20128 28422
rect 20076 28358 20128 28364
rect 20088 27538 20116 28358
rect 20272 28082 20300 33934
rect 20364 30598 20392 36178
rect 20444 35080 20496 35086
rect 20444 35022 20496 35028
rect 20456 34950 20484 35022
rect 20444 34944 20496 34950
rect 20444 34886 20496 34892
rect 20548 32434 20576 37742
rect 20904 37732 20956 37738
rect 20904 37674 20956 37680
rect 20916 37262 20944 37674
rect 21100 37262 21128 37810
rect 20904 37256 20956 37262
rect 20904 37198 20956 37204
rect 21088 37256 21140 37262
rect 21088 37198 21140 37204
rect 20628 36168 20680 36174
rect 20628 36110 20680 36116
rect 20640 35086 20668 36110
rect 21192 35578 21220 40718
rect 21272 40656 21324 40662
rect 21270 40624 21272 40633
rect 21324 40624 21326 40633
rect 21270 40559 21326 40568
rect 21376 40526 21404 40938
rect 21456 40928 21508 40934
rect 21456 40870 21508 40876
rect 21468 40769 21496 40870
rect 21454 40760 21510 40769
rect 21454 40695 21510 40704
rect 21364 40520 21416 40526
rect 21270 40488 21326 40497
rect 21364 40462 21416 40468
rect 21456 40520 21508 40526
rect 21456 40462 21508 40468
rect 21270 40423 21326 40432
rect 21284 39914 21312 40423
rect 21272 39908 21324 39914
rect 21272 39850 21324 39856
rect 21364 39840 21416 39846
rect 21364 39782 21416 39788
rect 21272 39432 21324 39438
rect 21376 39409 21404 39782
rect 21468 39642 21496 40462
rect 21560 40050 21588 41686
rect 22008 41608 22060 41614
rect 22006 41576 22008 41585
rect 22060 41576 22062 41585
rect 21640 41540 21692 41546
rect 22006 41511 22062 41520
rect 21640 41482 21692 41488
rect 21652 40712 21680 41482
rect 22112 41138 22140 42230
rect 22204 41800 22232 42758
rect 22284 42764 22336 42770
rect 22848 42758 22968 42786
rect 22284 42706 22336 42712
rect 22376 42628 22428 42634
rect 22376 42570 22428 42576
rect 22836 42628 22888 42634
rect 22836 42570 22888 42576
rect 22284 41812 22336 41818
rect 22204 41772 22284 41800
rect 22284 41754 22336 41760
rect 22190 41712 22246 41721
rect 22190 41647 22246 41656
rect 22204 41274 22232 41647
rect 22284 41472 22336 41478
rect 22284 41414 22336 41420
rect 22296 41274 22324 41414
rect 22192 41268 22244 41274
rect 22192 41210 22244 41216
rect 22284 41268 22336 41274
rect 22284 41210 22336 41216
rect 22282 41168 22338 41177
rect 22008 41132 22060 41138
rect 22008 41074 22060 41080
rect 22100 41132 22152 41138
rect 22282 41103 22284 41112
rect 22100 41074 22152 41080
rect 22336 41103 22338 41112
rect 22284 41074 22336 41080
rect 22020 40916 22048 41074
rect 22192 41064 22244 41070
rect 22192 41006 22244 41012
rect 22020 40888 22140 40916
rect 21719 40828 22027 40837
rect 21719 40826 21725 40828
rect 21781 40826 21805 40828
rect 21861 40826 21885 40828
rect 21941 40826 21965 40828
rect 22021 40826 22027 40828
rect 21781 40774 21783 40826
rect 21963 40774 21965 40826
rect 21719 40772 21725 40774
rect 21781 40772 21805 40774
rect 21861 40772 21885 40774
rect 21941 40772 21965 40774
rect 22021 40772 22027 40774
rect 21719 40763 22027 40772
rect 21652 40684 21956 40712
rect 21732 40520 21784 40526
rect 21652 40480 21732 40508
rect 21548 40044 21600 40050
rect 21548 39986 21600 39992
rect 21652 39642 21680 40480
rect 21732 40462 21784 40468
rect 21928 40458 21956 40684
rect 22008 40656 22060 40662
rect 22008 40598 22060 40604
rect 21916 40452 21968 40458
rect 21916 40394 21968 40400
rect 22020 40186 22048 40598
rect 22112 40361 22140 40888
rect 22098 40352 22154 40361
rect 22098 40287 22154 40296
rect 22204 40186 22232 41006
rect 22388 40730 22416 42570
rect 22468 42220 22520 42226
rect 22468 42162 22520 42168
rect 22560 42220 22612 42226
rect 22560 42162 22612 42168
rect 22480 41449 22508 42162
rect 22466 41440 22522 41449
rect 22466 41375 22522 41384
rect 22572 40730 22600 42162
rect 22652 41132 22704 41138
rect 22652 41074 22704 41080
rect 22664 41041 22692 41074
rect 22650 41032 22706 41041
rect 22650 40967 22706 40976
rect 22376 40724 22428 40730
rect 22376 40666 22428 40672
rect 22560 40724 22612 40730
rect 22560 40666 22612 40672
rect 22284 40520 22336 40526
rect 22282 40488 22284 40497
rect 22336 40488 22338 40497
rect 22282 40423 22338 40432
rect 22008 40180 22060 40186
rect 22008 40122 22060 40128
rect 22192 40180 22244 40186
rect 22192 40122 22244 40128
rect 21732 40112 21784 40118
rect 21730 40080 21732 40089
rect 21784 40080 21786 40089
rect 21730 40015 21786 40024
rect 22100 40044 22152 40050
rect 22100 39986 22152 39992
rect 22560 40044 22612 40050
rect 22560 39986 22612 39992
rect 21719 39740 22027 39749
rect 21719 39738 21725 39740
rect 21781 39738 21805 39740
rect 21861 39738 21885 39740
rect 21941 39738 21965 39740
rect 22021 39738 22027 39740
rect 21781 39686 21783 39738
rect 21963 39686 21965 39738
rect 21719 39684 21725 39686
rect 21781 39684 21805 39686
rect 21861 39684 21885 39686
rect 21941 39684 21965 39686
rect 22021 39684 22027 39686
rect 21719 39675 22027 39684
rect 21456 39636 21508 39642
rect 21456 39578 21508 39584
rect 21640 39636 21692 39642
rect 22112 39624 22140 39986
rect 22468 39976 22520 39982
rect 22468 39918 22520 39924
rect 22480 39642 22508 39918
rect 22572 39642 22600 39986
rect 21640 39578 21692 39584
rect 21928 39596 22140 39624
rect 22468 39636 22520 39642
rect 21928 39506 21956 39596
rect 22468 39578 22520 39584
rect 22560 39636 22612 39642
rect 22560 39578 22612 39584
rect 21916 39500 21968 39506
rect 21916 39442 21968 39448
rect 22560 39500 22612 39506
rect 22560 39442 22612 39448
rect 22468 39432 22520 39438
rect 21272 39374 21324 39380
rect 21362 39400 21418 39409
rect 21284 38729 21312 39374
rect 22282 39400 22338 39409
rect 21362 39335 21418 39344
rect 22008 39364 22060 39370
rect 22282 39335 22284 39344
rect 22008 39306 22060 39312
rect 22336 39335 22338 39344
rect 22466 39400 22468 39409
rect 22520 39400 22522 39409
rect 22466 39335 22522 39344
rect 22284 39306 22336 39312
rect 21640 39296 21692 39302
rect 22020 39250 22048 39306
rect 21692 39244 22048 39250
rect 21640 39238 22048 39244
rect 22100 39296 22152 39302
rect 22100 39238 22152 39244
rect 21652 39222 22048 39238
rect 21364 38888 21416 38894
rect 21364 38830 21416 38836
rect 21270 38720 21326 38729
rect 21270 38655 21326 38664
rect 21376 38282 21404 38830
rect 21719 38652 22027 38661
rect 21719 38650 21725 38652
rect 21781 38650 21805 38652
rect 21861 38650 21885 38652
rect 21941 38650 21965 38652
rect 22021 38650 22027 38652
rect 21781 38598 21783 38650
rect 21963 38598 21965 38650
rect 21719 38596 21725 38598
rect 21781 38596 21805 38598
rect 21861 38596 21885 38598
rect 21941 38596 21965 38598
rect 22021 38596 22027 38598
rect 21719 38587 22027 38596
rect 22112 38350 22140 39238
rect 22468 38956 22520 38962
rect 22468 38898 22520 38904
rect 22376 38752 22428 38758
rect 22204 38700 22376 38706
rect 22204 38694 22428 38700
rect 22204 38678 22416 38694
rect 22100 38344 22152 38350
rect 22100 38286 22152 38292
rect 21364 38276 21416 38282
rect 21364 38218 21416 38224
rect 21456 38208 21508 38214
rect 21456 38150 21508 38156
rect 21468 38010 21496 38150
rect 21456 38004 21508 38010
rect 21456 37946 21508 37952
rect 21719 37564 22027 37573
rect 21719 37562 21725 37564
rect 21781 37562 21805 37564
rect 21861 37562 21885 37564
rect 21941 37562 21965 37564
rect 22021 37562 22027 37564
rect 21781 37510 21783 37562
rect 21963 37510 21965 37562
rect 21719 37508 21725 37510
rect 21781 37508 21805 37510
rect 21861 37508 21885 37510
rect 21941 37508 21965 37510
rect 22021 37508 22027 37510
rect 21719 37499 22027 37508
rect 21456 37256 21508 37262
rect 21456 37198 21508 37204
rect 21272 37120 21324 37126
rect 21272 37062 21324 37068
rect 21284 36242 21312 37062
rect 21272 36236 21324 36242
rect 21272 36178 21324 36184
rect 21272 35692 21324 35698
rect 21272 35634 21324 35640
rect 20916 35550 21220 35578
rect 20720 35488 20772 35494
rect 20720 35430 20772 35436
rect 20628 35080 20680 35086
rect 20626 35048 20628 35057
rect 20680 35048 20682 35057
rect 20626 34983 20682 34992
rect 20628 32904 20680 32910
rect 20628 32846 20680 32852
rect 20732 32858 20760 35430
rect 20812 33312 20864 33318
rect 20812 33254 20864 33260
rect 20824 33114 20852 33254
rect 20812 33108 20864 33114
rect 20812 33050 20864 33056
rect 20640 32434 20668 32846
rect 20732 32830 20852 32858
rect 20720 32768 20772 32774
rect 20720 32710 20772 32716
rect 20732 32570 20760 32710
rect 20824 32570 20852 32830
rect 20720 32564 20772 32570
rect 20720 32506 20772 32512
rect 20812 32564 20864 32570
rect 20812 32506 20864 32512
rect 20536 32428 20588 32434
rect 20536 32370 20588 32376
rect 20628 32428 20680 32434
rect 20628 32370 20680 32376
rect 20536 31136 20588 31142
rect 20536 31078 20588 31084
rect 20352 30592 20404 30598
rect 20352 30534 20404 30540
rect 20442 30424 20498 30433
rect 20442 30359 20498 30368
rect 20456 30326 20484 30359
rect 20444 30320 20496 30326
rect 20444 30262 20496 30268
rect 20548 28994 20576 31078
rect 20640 30054 20668 32370
rect 20916 30716 20944 35550
rect 21284 35290 21312 35634
rect 21272 35284 21324 35290
rect 21272 35226 21324 35232
rect 21180 35216 21232 35222
rect 21468 35170 21496 37198
rect 21719 36476 22027 36485
rect 21719 36474 21725 36476
rect 21781 36474 21805 36476
rect 21861 36474 21885 36476
rect 21941 36474 21965 36476
rect 22021 36474 22027 36476
rect 21781 36422 21783 36474
rect 21963 36422 21965 36474
rect 21719 36420 21725 36422
rect 21781 36420 21805 36422
rect 21861 36420 21885 36422
rect 21941 36420 21965 36422
rect 22021 36420 22027 36422
rect 21719 36411 22027 36420
rect 21548 36032 21600 36038
rect 21548 35974 21600 35980
rect 22112 35986 22140 38286
rect 22204 37874 22232 38678
rect 22480 38554 22508 38898
rect 22468 38548 22520 38554
rect 22468 38490 22520 38496
rect 22376 38344 22428 38350
rect 22376 38286 22428 38292
rect 22468 38344 22520 38350
rect 22468 38286 22520 38292
rect 22284 38208 22336 38214
rect 22284 38150 22336 38156
rect 22192 37868 22244 37874
rect 22192 37810 22244 37816
rect 22296 37806 22324 38150
rect 22284 37800 22336 37806
rect 22284 37742 22336 37748
rect 22284 36780 22336 36786
rect 22284 36722 22336 36728
rect 22296 36378 22324 36722
rect 22284 36372 22336 36378
rect 22284 36314 22336 36320
rect 21560 35698 21588 35974
rect 22112 35958 22324 35986
rect 21732 35760 21784 35766
rect 21732 35702 21784 35708
rect 22192 35760 22244 35766
rect 22192 35702 22244 35708
rect 21548 35692 21600 35698
rect 21548 35634 21600 35640
rect 21744 35494 21772 35702
rect 22100 35692 22152 35698
rect 22100 35634 22152 35640
rect 21732 35488 21784 35494
rect 21732 35430 21784 35436
rect 21719 35388 22027 35397
rect 21719 35386 21725 35388
rect 21781 35386 21805 35388
rect 21861 35386 21885 35388
rect 21941 35386 21965 35388
rect 22021 35386 22027 35388
rect 21781 35334 21783 35386
rect 21963 35334 21965 35386
rect 21719 35332 21725 35334
rect 21781 35332 21805 35334
rect 21861 35332 21885 35334
rect 21941 35332 21965 35334
rect 22021 35332 22027 35334
rect 21719 35323 22027 35332
rect 21916 35284 21968 35290
rect 22112 35272 22140 35634
rect 21968 35244 22140 35272
rect 21916 35226 21968 35232
rect 21180 35158 21232 35164
rect 21192 35018 21220 35158
rect 21284 35142 21496 35170
rect 21180 35012 21232 35018
rect 21180 34954 21232 34960
rect 21180 33924 21232 33930
rect 21180 33866 21232 33872
rect 21192 32842 21220 33866
rect 21180 32836 21232 32842
rect 21180 32778 21232 32784
rect 20996 32768 21048 32774
rect 20996 32710 21048 32716
rect 20732 30688 20944 30716
rect 20628 30048 20680 30054
rect 20628 29990 20680 29996
rect 20364 28966 20576 28994
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 20076 27532 20128 27538
rect 20076 27474 20128 27480
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 20076 26920 20128 26926
rect 20076 26862 20128 26868
rect 20088 26382 20116 26862
rect 20076 26376 20128 26382
rect 20076 26318 20128 26324
rect 19892 25424 19944 25430
rect 19892 25366 19944 25372
rect 19904 24206 19932 25366
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 19996 24954 20024 25230
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19996 24206 20024 24550
rect 19892 24200 19944 24206
rect 19892 24142 19944 24148
rect 19984 24200 20036 24206
rect 20088 24188 20116 26318
rect 20260 26308 20312 26314
rect 20260 26250 20312 26256
rect 20272 26042 20300 26250
rect 20260 26036 20312 26042
rect 20260 25978 20312 25984
rect 20168 25424 20220 25430
rect 20168 25366 20220 25372
rect 20180 24818 20208 25366
rect 20364 25242 20392 28966
rect 20444 28688 20496 28694
rect 20444 28630 20496 28636
rect 20456 28558 20484 28630
rect 20640 28558 20668 29990
rect 20732 29170 20760 30688
rect 20812 30592 20864 30598
rect 20812 30534 20864 30540
rect 20904 30592 20956 30598
rect 20904 30534 20956 30540
rect 20720 29164 20772 29170
rect 20720 29106 20772 29112
rect 20444 28552 20496 28558
rect 20444 28494 20496 28500
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20536 28416 20588 28422
rect 20536 28358 20588 28364
rect 20548 28257 20576 28358
rect 20534 28248 20590 28257
rect 20534 28183 20536 28192
rect 20588 28183 20590 28192
rect 20536 28154 20588 28160
rect 20640 26926 20668 28494
rect 20718 27704 20774 27713
rect 20718 27639 20774 27648
rect 20628 26920 20680 26926
rect 20628 26862 20680 26868
rect 20272 25214 20392 25242
rect 20444 25288 20496 25294
rect 20444 25230 20496 25236
rect 20272 24954 20300 25214
rect 20352 25152 20404 25158
rect 20352 25094 20404 25100
rect 20260 24948 20312 24954
rect 20260 24890 20312 24896
rect 20272 24818 20300 24890
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20260 24812 20312 24818
rect 20260 24754 20312 24760
rect 20364 24410 20392 25094
rect 20456 24614 20484 25230
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20352 24404 20404 24410
rect 20352 24346 20404 24352
rect 20168 24336 20220 24342
rect 20220 24284 20576 24290
rect 20168 24278 20576 24284
rect 20180 24262 20576 24278
rect 20168 24200 20220 24206
rect 20088 24160 20168 24188
rect 19984 24142 20036 24148
rect 20168 24142 20220 24148
rect 19720 23990 20024 24018
rect 19800 23588 19852 23594
rect 19800 23530 19852 23536
rect 19524 23044 19576 23050
rect 19524 22986 19576 22992
rect 19616 22636 19668 22642
rect 19616 22578 19668 22584
rect 19524 22024 19576 22030
rect 19524 21966 19576 21972
rect 19536 21078 19564 21966
rect 19628 21894 19656 22578
rect 19708 22432 19760 22438
rect 19708 22374 19760 22380
rect 19720 22234 19748 22374
rect 19708 22228 19760 22234
rect 19708 22170 19760 22176
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19524 21072 19576 21078
rect 19524 21014 19576 21020
rect 19444 20862 19656 20890
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19260 20466 19380 20482
rect 19248 20460 19380 20466
rect 19300 20454 19380 20460
rect 19248 20402 19300 20408
rect 19352 18290 19380 20454
rect 19444 19854 19472 20742
rect 19536 20602 19564 20742
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19628 19854 19656 20862
rect 19708 20800 19760 20806
rect 19708 20742 19760 20748
rect 19720 20466 19748 20742
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19812 19904 19840 23530
rect 19892 22500 19944 22506
rect 19892 22442 19944 22448
rect 19904 22098 19932 22442
rect 19892 22092 19944 22098
rect 19996 22094 20024 23990
rect 20180 22098 20208 24142
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 20456 22710 20484 23054
rect 20444 22704 20496 22710
rect 20444 22646 20496 22652
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 20272 22234 20300 22374
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 19996 22066 20116 22094
rect 19892 22034 19944 22040
rect 19904 21690 19932 22034
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19996 21690 20024 21830
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 19892 21344 19944 21350
rect 19892 21286 19944 21292
rect 19904 20058 19932 21286
rect 19984 21072 20036 21078
rect 19984 21014 20036 21020
rect 19892 20052 19944 20058
rect 19892 19994 19944 20000
rect 19812 19876 19932 19904
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19628 19378 19656 19790
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19340 18284 19392 18290
rect 19260 18244 19340 18272
rect 19260 16590 19288 18244
rect 19340 18226 19392 18232
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19444 17898 19472 18226
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19352 17882 19472 17898
rect 19340 17876 19472 17882
rect 19392 17870 19472 17876
rect 19340 17818 19392 17824
rect 19430 17368 19486 17377
rect 19430 17303 19486 17312
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19260 15910 19288 16526
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 19260 15026 19288 15846
rect 19352 15706 19380 16118
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 19260 14482 19288 14962
rect 19444 14929 19472 17303
rect 19536 17202 19564 18022
rect 19628 17882 19656 18702
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19628 17270 19656 17818
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19720 17134 19748 18566
rect 19812 18426 19840 18702
rect 19800 18420 19852 18426
rect 19800 18362 19852 18368
rect 19904 17678 19932 19876
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19708 17128 19760 17134
rect 19708 17070 19760 17076
rect 19800 16244 19852 16250
rect 19800 16186 19852 16192
rect 19812 15570 19840 16186
rect 19996 15910 20024 21014
rect 20088 19718 20116 22066
rect 20168 22092 20220 22098
rect 20168 22034 20220 22040
rect 20548 21962 20576 24262
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 20640 23866 20668 24074
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20628 23044 20680 23050
rect 20628 22986 20680 22992
rect 20640 22506 20668 22986
rect 20628 22500 20680 22506
rect 20628 22442 20680 22448
rect 20732 22094 20760 27639
rect 20824 23118 20852 30534
rect 20916 30258 20944 30534
rect 21008 30297 21036 32710
rect 21088 30592 21140 30598
rect 21088 30534 21140 30540
rect 20994 30288 21050 30297
rect 20904 30252 20956 30258
rect 21100 30256 21128 30534
rect 20994 30223 21050 30232
rect 21088 30250 21140 30256
rect 20904 30194 20956 30200
rect 20916 29850 20944 30194
rect 21088 30192 21140 30198
rect 21180 30252 21232 30258
rect 21180 30194 21232 30200
rect 20996 30048 21048 30054
rect 20996 29990 21048 29996
rect 20904 29844 20956 29850
rect 20904 29786 20956 29792
rect 20904 27396 20956 27402
rect 20904 27338 20956 27344
rect 20916 27062 20944 27338
rect 20904 27056 20956 27062
rect 20904 26998 20956 27004
rect 21008 24818 21036 29990
rect 21088 29708 21140 29714
rect 21088 29650 21140 29656
rect 21100 26450 21128 29650
rect 21192 29646 21220 30194
rect 21180 29640 21232 29646
rect 21180 29582 21232 29588
rect 21088 26444 21140 26450
rect 21088 26386 21140 26392
rect 21100 25430 21128 26386
rect 21284 26194 21312 35142
rect 21456 35080 21508 35086
rect 22204 35034 22232 35702
rect 21456 35022 21508 35028
rect 21468 34746 21496 35022
rect 22112 35006 22232 35034
rect 22112 34950 22140 35006
rect 22100 34944 22152 34950
rect 22100 34886 22152 34892
rect 22296 34762 22324 35958
rect 21456 34740 21508 34746
rect 21456 34682 21508 34688
rect 22112 34734 22324 34762
rect 21719 34300 22027 34309
rect 21719 34298 21725 34300
rect 21781 34298 21805 34300
rect 21861 34298 21885 34300
rect 21941 34298 21965 34300
rect 22021 34298 22027 34300
rect 21781 34246 21783 34298
rect 21963 34246 21965 34298
rect 21719 34244 21725 34246
rect 21781 34244 21805 34246
rect 21861 34244 21885 34246
rect 21941 34244 21965 34246
rect 22021 34244 22027 34246
rect 21719 34235 22027 34244
rect 22112 34202 22140 34734
rect 22100 34196 22152 34202
rect 22100 34138 22152 34144
rect 21364 33992 21416 33998
rect 21364 33934 21416 33940
rect 21376 31958 21404 33934
rect 22112 33538 22140 34138
rect 22192 33856 22244 33862
rect 22192 33798 22244 33804
rect 22204 33658 22232 33798
rect 22192 33652 22244 33658
rect 22192 33594 22244 33600
rect 22112 33510 22232 33538
rect 22100 33312 22152 33318
rect 22100 33254 22152 33260
rect 21719 33212 22027 33221
rect 21719 33210 21725 33212
rect 21781 33210 21805 33212
rect 21861 33210 21885 33212
rect 21941 33210 21965 33212
rect 22021 33210 22027 33212
rect 21781 33158 21783 33210
rect 21963 33158 21965 33210
rect 21719 33156 21725 33158
rect 21781 33156 21805 33158
rect 21861 33156 21885 33158
rect 21941 33156 21965 33158
rect 22021 33156 22027 33158
rect 21546 33144 21602 33153
rect 21719 33147 22027 33156
rect 22112 33114 22140 33254
rect 21546 33079 21602 33088
rect 22100 33108 22152 33114
rect 21456 32224 21508 32230
rect 21456 32166 21508 32172
rect 21468 32026 21496 32166
rect 21456 32020 21508 32026
rect 21456 31962 21508 31968
rect 21364 31952 21416 31958
rect 21364 31894 21416 31900
rect 21376 29322 21404 31894
rect 21456 30728 21508 30734
rect 21456 30670 21508 30676
rect 21468 30394 21496 30670
rect 21456 30388 21508 30394
rect 21456 30330 21508 30336
rect 21376 29294 21496 29322
rect 21364 29164 21416 29170
rect 21364 29106 21416 29112
rect 21376 28762 21404 29106
rect 21364 28756 21416 28762
rect 21364 28698 21416 28704
rect 21364 26988 21416 26994
rect 21364 26930 21416 26936
rect 21376 26586 21404 26930
rect 21364 26580 21416 26586
rect 21364 26522 21416 26528
rect 21364 26308 21416 26314
rect 21468 26296 21496 29294
rect 21416 26268 21496 26296
rect 21364 26250 21416 26256
rect 21284 26166 21496 26194
rect 21088 25424 21140 25430
rect 21088 25366 21140 25372
rect 21180 25220 21232 25226
rect 21180 25162 21232 25168
rect 20996 24812 21048 24818
rect 20996 24754 21048 24760
rect 21192 24138 21220 25162
rect 21362 24712 21418 24721
rect 21362 24647 21418 24656
rect 21376 24410 21404 24647
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 21180 24132 21232 24138
rect 21180 24074 21232 24080
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 20640 22066 20760 22094
rect 20536 21956 20588 21962
rect 20536 21898 20588 21904
rect 20548 21554 20576 21898
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20088 16250 20116 19654
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19430 14920 19486 14929
rect 19430 14855 19486 14864
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19168 14334 19288 14362
rect 18752 14172 19060 14181
rect 18752 14170 18758 14172
rect 18814 14170 18838 14172
rect 18894 14170 18918 14172
rect 18974 14170 18998 14172
rect 19054 14170 19060 14172
rect 18814 14118 18816 14170
rect 18996 14118 18998 14170
rect 18752 14116 18758 14118
rect 18814 14116 18838 14118
rect 18894 14116 18918 14118
rect 18974 14116 18998 14118
rect 19054 14116 19060 14118
rect 18752 14107 19060 14116
rect 18696 13932 18748 13938
rect 18616 13892 18696 13920
rect 18696 13874 18748 13880
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 19076 13462 19104 13670
rect 19064 13456 19116 13462
rect 19064 13398 19116 13404
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18616 12986 18644 13262
rect 18752 13084 19060 13093
rect 18752 13082 18758 13084
rect 18814 13082 18838 13084
rect 18894 13082 18918 13084
rect 18974 13082 18998 13084
rect 19054 13082 19060 13084
rect 18814 13030 18816 13082
rect 18996 13030 18998 13082
rect 18752 13028 18758 13030
rect 18814 13028 18838 13030
rect 18894 13028 18918 13030
rect 18974 13028 18998 13030
rect 19054 13028 19060 13030
rect 18752 13019 19060 13028
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 19260 12434 19288 14334
rect 19352 13938 19380 14486
rect 19536 14346 19564 15506
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19628 14414 19656 14758
rect 19800 14544 19852 14550
rect 19800 14486 19852 14492
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19524 14340 19576 14346
rect 19524 14282 19576 14288
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19432 13864 19484 13870
rect 19536 13818 19564 14282
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19484 13812 19564 13818
rect 19432 13806 19564 13812
rect 19444 13790 19564 13806
rect 19720 13530 19748 14214
rect 19812 13938 19840 14486
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19444 12986 19472 13262
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19812 12434 19840 13874
rect 19168 12406 19288 12434
rect 19720 12406 19840 12434
rect 18752 11996 19060 12005
rect 18752 11994 18758 11996
rect 18814 11994 18838 11996
rect 18894 11994 18918 11996
rect 18974 11994 18998 11996
rect 19054 11994 19060 11996
rect 18814 11942 18816 11994
rect 18996 11942 18998 11994
rect 18752 11940 18758 11942
rect 18814 11940 18838 11942
rect 18894 11940 18918 11942
rect 18974 11940 18998 11942
rect 19054 11940 19060 11942
rect 18752 11931 19060 11940
rect 18752 10908 19060 10917
rect 18752 10906 18758 10908
rect 18814 10906 18838 10908
rect 18894 10906 18918 10908
rect 18974 10906 18998 10908
rect 19054 10906 19060 10908
rect 18814 10854 18816 10906
rect 18996 10854 18998 10906
rect 18752 10852 18758 10854
rect 18814 10852 18838 10854
rect 18894 10852 18918 10854
rect 18974 10852 18998 10854
rect 19054 10852 19060 10854
rect 18752 10843 19060 10852
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18892 10266 18920 10610
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 18752 9820 19060 9829
rect 18752 9818 18758 9820
rect 18814 9818 18838 9820
rect 18894 9818 18918 9820
rect 18974 9818 18998 9820
rect 19054 9818 19060 9820
rect 18814 9766 18816 9818
rect 18996 9766 18998 9818
rect 18752 9764 18758 9766
rect 18814 9764 18838 9766
rect 18894 9764 18918 9766
rect 18974 9764 18998 9766
rect 19054 9764 19060 9766
rect 18752 9755 19060 9764
rect 18752 8732 19060 8741
rect 18752 8730 18758 8732
rect 18814 8730 18838 8732
rect 18894 8730 18918 8732
rect 18974 8730 18998 8732
rect 19054 8730 19060 8732
rect 18814 8678 18816 8730
rect 18996 8678 18998 8730
rect 18752 8676 18758 8678
rect 18814 8676 18838 8678
rect 18894 8676 18918 8678
rect 18974 8676 18998 8678
rect 19054 8676 19060 8678
rect 18752 8667 19060 8676
rect 18752 7644 19060 7653
rect 18752 7642 18758 7644
rect 18814 7642 18838 7644
rect 18894 7642 18918 7644
rect 18974 7642 18998 7644
rect 19054 7642 19060 7644
rect 18814 7590 18816 7642
rect 18996 7590 18998 7642
rect 18752 7588 18758 7590
rect 18814 7588 18838 7590
rect 18894 7588 18918 7590
rect 18974 7588 18998 7590
rect 19054 7588 19060 7590
rect 18752 7579 19060 7588
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18800 7002 18828 7346
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 19168 6882 19196 12406
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19260 11694 19288 12310
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19248 11144 19300 11150
rect 19444 11132 19472 12174
rect 19300 11104 19472 11132
rect 19248 11086 19300 11092
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19352 10674 19380 10950
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19248 9648 19300 9654
rect 19352 9636 19380 9930
rect 19300 9608 19380 9636
rect 19248 9590 19300 9596
rect 19444 9450 19472 11104
rect 19720 10742 19748 12406
rect 19904 10826 19932 14010
rect 20088 13512 20116 15982
rect 20180 15162 20208 19654
rect 20272 16402 20300 20198
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20364 18358 20392 18634
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20272 16374 20392 16402
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 19996 13484 20116 13512
rect 19996 13172 20024 13484
rect 20180 13410 20208 13670
rect 20088 13382 20208 13410
rect 20088 13326 20116 13382
rect 20272 13326 20300 14214
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20168 13184 20220 13190
rect 19996 13144 20116 13172
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19812 10798 19932 10826
rect 19708 10736 19760 10742
rect 19628 10696 19708 10724
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 19536 10266 19564 10610
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19260 7410 19288 8434
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19260 7018 19288 7346
rect 19260 6990 19380 7018
rect 19168 6854 19288 6882
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 18616 6458 18644 6734
rect 18752 6556 19060 6565
rect 18752 6554 18758 6556
rect 18814 6554 18838 6556
rect 18894 6554 18918 6556
rect 18974 6554 18998 6556
rect 19054 6554 19060 6556
rect 18814 6502 18816 6554
rect 18996 6502 18998 6554
rect 18752 6500 18758 6502
rect 18814 6500 18838 6502
rect 18894 6500 18918 6502
rect 18974 6500 18998 6502
rect 19054 6500 19060 6502
rect 18752 6491 19060 6500
rect 19168 6458 19196 6734
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19064 6180 19116 6186
rect 19064 6122 19116 6128
rect 19076 5574 19104 6122
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 18752 5468 19060 5477
rect 18752 5466 18758 5468
rect 18814 5466 18838 5468
rect 18894 5466 18918 5468
rect 18974 5466 18998 5468
rect 19054 5466 19060 5468
rect 18814 5414 18816 5466
rect 18996 5414 18998 5466
rect 18752 5412 18758 5414
rect 18814 5412 18838 5414
rect 18894 5412 18918 5414
rect 18974 5412 18998 5414
rect 19054 5412 19060 5414
rect 18752 5403 19060 5412
rect 18696 5296 18748 5302
rect 18696 5238 18748 5244
rect 18708 4826 18736 5238
rect 18696 4820 18748 4826
rect 18696 4762 18748 4768
rect 18696 4616 18748 4622
rect 18616 4576 18696 4604
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18340 3738 18368 3878
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18524 3194 18552 3470
rect 18616 3398 18644 4576
rect 18696 4558 18748 4564
rect 18752 4380 19060 4389
rect 18752 4378 18758 4380
rect 18814 4378 18838 4380
rect 18894 4378 18918 4380
rect 18974 4378 18998 4380
rect 19054 4378 19060 4380
rect 18814 4326 18816 4378
rect 18996 4326 18998 4378
rect 18752 4324 18758 4326
rect 18814 4324 18838 4326
rect 18894 4324 18918 4326
rect 18974 4324 18998 4326
rect 19054 4324 19060 4326
rect 18752 4315 19060 4324
rect 19260 4162 19288 6854
rect 19352 6390 19380 6990
rect 19444 6798 19472 8502
rect 19628 7002 19656 10696
rect 19708 10678 19760 10684
rect 19812 10554 19840 10798
rect 19892 10736 19944 10742
rect 19996 10724 20024 12922
rect 20088 11064 20116 13144
rect 20168 13126 20220 13132
rect 20180 12238 20208 13126
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20088 11036 20300 11064
rect 20168 10804 20220 10810
rect 19944 10696 20024 10724
rect 20088 10764 20168 10792
rect 19892 10678 19944 10684
rect 19812 10526 19932 10554
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19720 9722 19748 9998
rect 19708 9716 19760 9722
rect 19708 9658 19760 9664
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19720 7546 19748 7822
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19616 6996 19668 7002
rect 19616 6938 19668 6944
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19352 4622 19380 6326
rect 19628 4706 19656 6938
rect 19706 5264 19762 5273
rect 19706 5199 19762 5208
rect 19800 5228 19852 5234
rect 19720 4826 19748 5199
rect 19800 5170 19852 5176
rect 19812 4826 19840 5170
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19628 4678 19748 4706
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19352 4282 19380 4558
rect 19524 4548 19576 4554
rect 19524 4490 19576 4496
rect 19536 4321 19564 4490
rect 19522 4312 19578 4321
rect 19340 4276 19392 4282
rect 19392 4236 19463 4264
rect 19628 4282 19656 4558
rect 19522 4247 19578 4256
rect 19616 4276 19668 4282
rect 19340 4218 19392 4224
rect 19435 4196 19463 4236
rect 19616 4218 19668 4224
rect 19338 4176 19394 4185
rect 19260 4134 19338 4162
rect 19435 4168 19564 4196
rect 19338 4111 19394 4120
rect 19536 3992 19564 4168
rect 19352 3964 19564 3992
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 18892 3602 18920 3878
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18236 3120 18288 3126
rect 18236 3062 18288 3068
rect 18248 2854 18276 3062
rect 17512 2746 17632 2774
rect 17498 2680 17554 2689
rect 17408 2644 17460 2650
rect 17498 2615 17554 2624
rect 17408 2586 17460 2592
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17328 2106 17356 2246
rect 17316 2100 17368 2106
rect 17316 2042 17368 2048
rect 17224 1352 17276 1358
rect 17224 1294 17276 1300
rect 16762 54 16896 82
rect 16762 0 16818 54
rect 17038 0 17094 160
rect 17314 82 17370 160
rect 17420 82 17448 2586
rect 17512 2446 17540 2615
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 17604 2038 17632 2746
rect 17592 2032 17644 2038
rect 17592 1974 17644 1980
rect 17696 1358 17724 2790
rect 17880 2774 18092 2802
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17684 1352 17736 1358
rect 17684 1294 17736 1300
rect 17314 54 17448 82
rect 17590 82 17646 160
rect 17788 82 17816 2246
rect 17960 1760 18012 1766
rect 17880 1720 17960 1748
rect 17880 160 17908 1720
rect 17960 1702 18012 1708
rect 18144 1760 18196 1766
rect 18144 1702 18196 1708
rect 18156 160 18184 1702
rect 18340 1562 18368 2450
rect 18328 1556 18380 1562
rect 18328 1498 18380 1504
rect 18432 160 18460 2790
rect 18510 2544 18566 2553
rect 18616 2514 18644 3334
rect 18752 3292 19060 3301
rect 18752 3290 18758 3292
rect 18814 3290 18838 3292
rect 18894 3290 18918 3292
rect 18974 3290 18998 3292
rect 19054 3290 19060 3292
rect 18814 3238 18816 3290
rect 18996 3238 18998 3290
rect 18752 3236 18758 3238
rect 18814 3236 18838 3238
rect 18894 3236 18918 3238
rect 18974 3236 18998 3238
rect 19054 3236 19060 3238
rect 18752 3227 19060 3236
rect 19168 3040 19196 3878
rect 19246 3768 19302 3777
rect 19246 3703 19302 3712
rect 19260 3534 19288 3703
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19076 3012 19196 3040
rect 18878 2680 18934 2689
rect 19076 2650 19104 3012
rect 19156 2916 19208 2922
rect 19156 2858 19208 2864
rect 18878 2615 18934 2624
rect 19064 2644 19116 2650
rect 18510 2479 18566 2488
rect 18604 2508 18656 2514
rect 18524 2038 18552 2479
rect 18604 2450 18656 2456
rect 18892 2446 18920 2615
rect 19064 2586 19116 2592
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18616 2106 18644 2246
rect 18752 2204 19060 2213
rect 18752 2202 18758 2204
rect 18814 2202 18838 2204
rect 18894 2202 18918 2204
rect 18974 2202 18998 2204
rect 19054 2202 19060 2204
rect 18814 2150 18816 2202
rect 18996 2150 18998 2202
rect 18752 2148 18758 2150
rect 18814 2148 18838 2150
rect 18894 2148 18918 2150
rect 18974 2148 18998 2150
rect 19054 2148 19060 2150
rect 18752 2139 19060 2148
rect 18604 2100 18656 2106
rect 18604 2042 18656 2048
rect 18512 2032 18564 2038
rect 18512 1974 18564 1980
rect 18604 1964 18656 1970
rect 18604 1906 18656 1912
rect 18512 1352 18564 1358
rect 18510 1320 18512 1329
rect 18564 1320 18566 1329
rect 18510 1255 18566 1264
rect 17590 54 17816 82
rect 17314 0 17370 54
rect 17590 0 17646 54
rect 17866 0 17922 160
rect 18142 0 18198 160
rect 18418 0 18474 160
rect 18616 82 18644 1906
rect 18752 1116 19060 1125
rect 18752 1114 18758 1116
rect 18814 1114 18838 1116
rect 18894 1114 18918 1116
rect 18974 1114 18998 1116
rect 19054 1114 19060 1116
rect 18814 1062 18816 1114
rect 18996 1062 18998 1114
rect 18752 1060 18758 1062
rect 18814 1060 18838 1062
rect 18894 1060 18918 1062
rect 18974 1060 18998 1062
rect 19054 1060 19060 1062
rect 18752 1051 19060 1060
rect 18694 82 18750 160
rect 18616 54 18750 82
rect 18694 0 18750 54
rect 18970 82 19026 160
rect 19168 82 19196 2858
rect 19260 2689 19288 3334
rect 19352 3194 19380 3964
rect 19720 3913 19748 4678
rect 19904 4468 19932 10526
rect 19984 9988 20036 9994
rect 19984 9930 20036 9936
rect 19996 6798 20024 9930
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19996 4622 20024 5034
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19904 4440 20024 4468
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 19522 3904 19578 3913
rect 19706 3904 19762 3913
rect 19578 3862 19656 3890
rect 19522 3839 19578 3848
rect 19628 3754 19656 3862
rect 19706 3839 19762 3848
rect 19628 3726 19748 3754
rect 19720 3466 19748 3726
rect 19708 3460 19760 3466
rect 19708 3402 19760 3408
rect 19524 3392 19576 3398
rect 19522 3360 19524 3369
rect 19576 3360 19578 3369
rect 19522 3295 19578 3304
rect 19812 3210 19840 4082
rect 19890 4040 19946 4049
rect 19890 3975 19946 3984
rect 19904 3602 19932 3975
rect 19892 3596 19944 3602
rect 19892 3538 19944 3544
rect 19892 3460 19944 3466
rect 19892 3402 19944 3408
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19432 3188 19484 3194
rect 19536 3182 19840 3210
rect 19536 3176 19564 3182
rect 19484 3148 19564 3176
rect 19432 3130 19484 3136
rect 19616 3120 19668 3126
rect 19522 3088 19578 3097
rect 19340 3052 19392 3058
rect 19444 3046 19522 3074
rect 19444 3040 19472 3046
rect 19392 3012 19472 3040
rect 19668 3080 19748 3108
rect 19616 3062 19668 3068
rect 19522 3023 19578 3032
rect 19340 2994 19392 3000
rect 19720 2990 19748 3080
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 19524 2848 19576 2854
rect 19338 2816 19394 2825
rect 19394 2774 19463 2802
rect 19800 2848 19852 2854
rect 19576 2796 19800 2802
rect 19524 2790 19852 2796
rect 19534 2774 19840 2790
rect 19338 2751 19394 2760
rect 19435 2746 19472 2774
rect 19246 2680 19302 2689
rect 19444 2632 19472 2746
rect 19246 2615 19302 2624
rect 19352 2604 19472 2632
rect 19522 2680 19578 2689
rect 19522 2615 19578 2624
rect 19352 2530 19380 2604
rect 19260 2502 19380 2530
rect 19260 160 19288 2502
rect 19340 2372 19392 2378
rect 19340 2314 19392 2320
rect 19352 2106 19380 2314
rect 19340 2100 19392 2106
rect 19340 2042 19392 2048
rect 19536 1970 19564 2615
rect 19614 2408 19670 2417
rect 19614 2343 19670 2352
rect 19524 1964 19576 1970
rect 19524 1906 19576 1912
rect 19524 1760 19576 1766
rect 19524 1702 19576 1708
rect 19432 1352 19484 1358
rect 19432 1294 19484 1300
rect 19444 950 19472 1294
rect 19432 944 19484 950
rect 19432 886 19484 892
rect 19536 160 19564 1702
rect 19628 1290 19656 2343
rect 19800 2304 19852 2310
rect 19800 2246 19852 2252
rect 19812 2106 19840 2246
rect 19800 2100 19852 2106
rect 19800 2042 19852 2048
rect 19800 1896 19852 1902
rect 19800 1838 19852 1844
rect 19812 1426 19840 1838
rect 19800 1420 19852 1426
rect 19800 1362 19852 1368
rect 19616 1284 19668 1290
rect 19616 1226 19668 1232
rect 18970 54 19196 82
rect 18970 0 19026 54
rect 19246 0 19302 160
rect 19522 0 19578 160
rect 19798 82 19854 160
rect 19904 82 19932 3402
rect 19996 2922 20024 4440
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 20088 2650 20116 10764
rect 20168 10746 20220 10752
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 20180 7002 20208 7754
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 20168 4752 20220 4758
rect 20168 4694 20220 4700
rect 20180 4622 20208 4694
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 20168 4480 20220 4486
rect 20166 4448 20168 4457
rect 20220 4448 20222 4457
rect 20166 4383 20222 4392
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 20180 3602 20208 3946
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20074 2408 20130 2417
rect 20074 2343 20130 2352
rect 20088 160 20116 2343
rect 20180 1766 20208 3334
rect 20272 1970 20300 11036
rect 20364 2106 20392 16374
rect 20456 15434 20484 19314
rect 20640 18737 20668 22066
rect 20810 21992 20866 22001
rect 20810 21927 20866 21936
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20732 20058 20760 20198
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20626 18728 20682 18737
rect 20626 18663 20682 18672
rect 20732 17678 20760 19858
rect 20824 19514 20852 21927
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20732 17542 20760 17614
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20732 17134 20760 17478
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20548 15706 20576 16050
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20640 15706 20668 15846
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20732 15586 20760 15846
rect 20548 15558 20760 15586
rect 20444 15428 20496 15434
rect 20444 15370 20496 15376
rect 20456 12986 20484 15370
rect 20548 13190 20576 15558
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20640 12889 20668 15098
rect 20720 14476 20772 14482
rect 20772 14436 20852 14464
rect 20720 14418 20772 14424
rect 20626 12880 20682 12889
rect 20536 12844 20588 12850
rect 20626 12815 20682 12824
rect 20536 12786 20588 12792
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20456 8974 20484 9318
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20548 7834 20576 12786
rect 20640 8090 20668 12815
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20732 11762 20760 12378
rect 20824 12306 20852 14436
rect 20916 14346 20944 22918
rect 21272 22704 21324 22710
rect 21272 22646 21324 22652
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 21008 18970 21036 21626
rect 21180 21412 21232 21418
rect 21180 21354 21232 21360
rect 21192 21010 21220 21354
rect 21180 21004 21232 21010
rect 21180 20946 21232 20952
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 17338 21036 17614
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 20916 13938 20944 14282
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20996 12640 21048 12646
rect 20996 12582 21048 12588
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20824 9518 20852 12242
rect 21008 11762 21036 12582
rect 21100 12322 21128 19314
rect 21284 17202 21312 22646
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21376 20058 21404 20198
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21362 18048 21418 18057
rect 21468 18034 21496 26166
rect 21560 20058 21588 33079
rect 22100 33050 22152 33056
rect 21640 32836 21692 32842
rect 21640 32778 21692 32784
rect 21652 29646 21680 32778
rect 21719 32124 22027 32133
rect 21719 32122 21725 32124
rect 21781 32122 21805 32124
rect 21861 32122 21885 32124
rect 21941 32122 21965 32124
rect 22021 32122 22027 32124
rect 21781 32070 21783 32122
rect 21963 32070 21965 32122
rect 21719 32068 21725 32070
rect 21781 32068 21805 32070
rect 21861 32068 21885 32070
rect 21941 32068 21965 32070
rect 22021 32068 22027 32070
rect 21719 32059 22027 32068
rect 22204 31498 22232 33510
rect 22388 31754 22416 38286
rect 22480 37466 22508 38286
rect 22572 37738 22600 39442
rect 22744 39432 22796 39438
rect 22744 39374 22796 39380
rect 22652 39024 22704 39030
rect 22756 39012 22784 39374
rect 22704 38984 22784 39012
rect 22652 38966 22704 38972
rect 22652 38752 22704 38758
rect 22652 38694 22704 38700
rect 22664 37942 22692 38694
rect 22652 37936 22704 37942
rect 22652 37878 22704 37884
rect 22560 37732 22612 37738
rect 22560 37674 22612 37680
rect 22468 37460 22520 37466
rect 22468 37402 22520 37408
rect 22848 36378 22876 42570
rect 23032 42362 23060 43823
rect 23124 43432 23152 44840
rect 23400 43602 23428 44840
rect 23400 43574 23520 43602
rect 23388 43444 23440 43450
rect 23124 43404 23388 43432
rect 23388 43386 23440 43392
rect 23388 43308 23440 43314
rect 23388 43250 23440 43256
rect 23112 43240 23164 43246
rect 23112 43182 23164 43188
rect 23124 42809 23152 43182
rect 23110 42800 23166 42809
rect 23110 42735 23166 42744
rect 23400 42684 23428 43250
rect 23492 42786 23520 43574
rect 23676 43466 23704 44840
rect 23676 43438 23796 43466
rect 23662 43344 23718 43353
rect 23662 43279 23718 43288
rect 23492 42770 23612 42786
rect 23492 42764 23624 42770
rect 23492 42758 23572 42764
rect 23572 42706 23624 42712
rect 23400 42656 23520 42684
rect 23020 42356 23072 42362
rect 23020 42298 23072 42304
rect 23202 41712 23258 41721
rect 23202 41647 23258 41656
rect 23216 41274 23244 41647
rect 23296 41540 23348 41546
rect 23296 41482 23348 41488
rect 23204 41268 23256 41274
rect 23204 41210 23256 41216
rect 23112 41132 23164 41138
rect 23112 41074 23164 41080
rect 22928 40520 22980 40526
rect 22928 40462 22980 40468
rect 22940 39098 22968 40462
rect 23020 40452 23072 40458
rect 23020 40394 23072 40400
rect 23032 39386 23060 40394
rect 23124 40186 23152 41074
rect 23308 40730 23336 41482
rect 23388 40996 23440 41002
rect 23388 40938 23440 40944
rect 23296 40724 23348 40730
rect 23296 40666 23348 40672
rect 23204 40452 23256 40458
rect 23204 40394 23256 40400
rect 23112 40180 23164 40186
rect 23112 40122 23164 40128
rect 23032 39358 23152 39386
rect 23020 39296 23072 39302
rect 23020 39238 23072 39244
rect 23032 39098 23060 39238
rect 23124 39098 23152 39358
rect 22928 39092 22980 39098
rect 22928 39034 22980 39040
rect 23020 39092 23072 39098
rect 23020 39034 23072 39040
rect 23112 39092 23164 39098
rect 23112 39034 23164 39040
rect 22928 38888 22980 38894
rect 22928 38830 22980 38836
rect 22940 38214 22968 38830
rect 22928 38208 22980 38214
rect 22928 38150 22980 38156
rect 23020 38004 23072 38010
rect 23020 37946 23072 37952
rect 23032 37874 23060 37946
rect 23020 37868 23072 37874
rect 23020 37810 23072 37816
rect 22928 36576 22980 36582
rect 22928 36518 22980 36524
rect 23020 36576 23072 36582
rect 23020 36518 23072 36524
rect 22836 36372 22888 36378
rect 22836 36314 22888 36320
rect 22744 36168 22796 36174
rect 22744 36110 22796 36116
rect 22756 35834 22784 36110
rect 22744 35828 22796 35834
rect 22744 35770 22796 35776
rect 22560 35692 22612 35698
rect 22560 35634 22612 35640
rect 22572 35290 22600 35634
rect 22940 35562 22968 36518
rect 23032 36145 23060 36518
rect 23018 36136 23074 36145
rect 23018 36071 23074 36080
rect 22928 35556 22980 35562
rect 22928 35498 22980 35504
rect 22560 35284 22612 35290
rect 22560 35226 22612 35232
rect 22744 35148 22796 35154
rect 22744 35090 22796 35096
rect 22756 33658 22784 35090
rect 22744 33652 22796 33658
rect 22744 33594 22796 33600
rect 22652 33516 22704 33522
rect 22652 33458 22704 33464
rect 22388 31726 22508 31754
rect 21836 31470 22232 31498
rect 21836 31278 21864 31470
rect 22192 31340 22244 31346
rect 22192 31282 22244 31288
rect 21824 31272 21876 31278
rect 21824 31214 21876 31220
rect 21719 31036 22027 31045
rect 21719 31034 21725 31036
rect 21781 31034 21805 31036
rect 21861 31034 21885 31036
rect 21941 31034 21965 31036
rect 22021 31034 22027 31036
rect 21781 30982 21783 31034
rect 21963 30982 21965 31034
rect 21719 30980 21725 30982
rect 21781 30980 21805 30982
rect 21861 30980 21885 30982
rect 21941 30980 21965 30982
rect 22021 30980 22027 30982
rect 21719 30971 22027 30980
rect 21719 29948 22027 29957
rect 21719 29946 21725 29948
rect 21781 29946 21805 29948
rect 21861 29946 21885 29948
rect 21941 29946 21965 29948
rect 22021 29946 22027 29948
rect 21781 29894 21783 29946
rect 21963 29894 21965 29946
rect 21719 29892 21725 29894
rect 21781 29892 21805 29894
rect 21861 29892 21885 29894
rect 21941 29892 21965 29894
rect 22021 29892 22027 29894
rect 21719 29883 22027 29892
rect 21640 29640 21692 29646
rect 21640 29582 21692 29588
rect 21824 29572 21876 29578
rect 21824 29514 21876 29520
rect 21730 29200 21786 29209
rect 21836 29170 21864 29514
rect 21730 29135 21786 29144
rect 21824 29164 21876 29170
rect 21638 29064 21694 29073
rect 21638 28999 21694 29008
rect 21652 28218 21680 28999
rect 21744 28966 21772 29135
rect 21824 29106 21876 29112
rect 22100 29028 22152 29034
rect 22100 28970 22152 28976
rect 21732 28960 21784 28966
rect 21732 28902 21784 28908
rect 21719 28860 22027 28869
rect 21719 28858 21725 28860
rect 21781 28858 21805 28860
rect 21861 28858 21885 28860
rect 21941 28858 21965 28860
rect 22021 28858 22027 28860
rect 21781 28806 21783 28858
rect 21963 28806 21965 28858
rect 21719 28804 21725 28806
rect 21781 28804 21805 28806
rect 21861 28804 21885 28806
rect 21941 28804 21965 28806
rect 22021 28804 22027 28806
rect 21719 28795 22027 28804
rect 21640 28212 21692 28218
rect 21640 28154 21692 28160
rect 22112 28082 22140 28970
rect 22204 28694 22232 31282
rect 22284 29708 22336 29714
rect 22284 29650 22336 29656
rect 22296 29238 22324 29650
rect 22376 29504 22428 29510
rect 22376 29446 22428 29452
rect 22284 29232 22336 29238
rect 22284 29174 22336 29180
rect 22388 29170 22416 29446
rect 22480 29209 22508 31726
rect 22560 30048 22612 30054
rect 22560 29990 22612 29996
rect 22572 29850 22600 29990
rect 22560 29844 22612 29850
rect 22560 29786 22612 29792
rect 22466 29200 22522 29209
rect 22376 29164 22428 29170
rect 22466 29135 22522 29144
rect 22560 29164 22612 29170
rect 22376 29106 22428 29112
rect 22560 29106 22612 29112
rect 22192 28688 22244 28694
rect 22192 28630 22244 28636
rect 22204 28218 22232 28630
rect 22388 28558 22416 29106
rect 22468 28960 22520 28966
rect 22468 28902 22520 28908
rect 22480 28626 22508 28902
rect 22572 28762 22600 29106
rect 22560 28756 22612 28762
rect 22560 28698 22612 28704
rect 22468 28620 22520 28626
rect 22468 28562 22520 28568
rect 22376 28552 22428 28558
rect 22376 28494 22428 28500
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22192 28212 22244 28218
rect 22192 28154 22244 28160
rect 22572 28082 22600 28494
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 22560 28076 22612 28082
rect 22560 28018 22612 28024
rect 21719 27772 22027 27781
rect 21719 27770 21725 27772
rect 21781 27770 21805 27772
rect 21861 27770 21885 27772
rect 21941 27770 21965 27772
rect 22021 27770 22027 27772
rect 21781 27718 21783 27770
rect 21963 27718 21965 27770
rect 21719 27716 21725 27718
rect 21781 27716 21805 27718
rect 21861 27716 21885 27718
rect 21941 27716 21965 27718
rect 22021 27716 22027 27718
rect 21719 27707 22027 27716
rect 22100 27668 22152 27674
rect 22100 27610 22152 27616
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 21928 27130 21956 27270
rect 21916 27124 21968 27130
rect 21916 27066 21968 27072
rect 21719 26684 22027 26693
rect 21719 26682 21725 26684
rect 21781 26682 21805 26684
rect 21861 26682 21885 26684
rect 21941 26682 21965 26684
rect 22021 26682 22027 26684
rect 21781 26630 21783 26682
rect 21963 26630 21965 26682
rect 21719 26628 21725 26630
rect 21781 26628 21805 26630
rect 21861 26628 21885 26630
rect 21941 26628 21965 26630
rect 22021 26628 22027 26630
rect 21719 26619 22027 26628
rect 21719 25596 22027 25605
rect 21719 25594 21725 25596
rect 21781 25594 21805 25596
rect 21861 25594 21885 25596
rect 21941 25594 21965 25596
rect 22021 25594 22027 25596
rect 21781 25542 21783 25594
rect 21963 25542 21965 25594
rect 21719 25540 21725 25542
rect 21781 25540 21805 25542
rect 21861 25540 21885 25542
rect 21941 25540 21965 25542
rect 22021 25540 22027 25542
rect 21719 25531 22027 25540
rect 21640 24812 21692 24818
rect 21640 24754 21692 24760
rect 21652 24410 21680 24754
rect 21719 24508 22027 24517
rect 21719 24506 21725 24508
rect 21781 24506 21805 24508
rect 21861 24506 21885 24508
rect 21941 24506 21965 24508
rect 22021 24506 22027 24508
rect 21781 24454 21783 24506
rect 21963 24454 21965 24506
rect 21719 24452 21725 24454
rect 21781 24452 21805 24454
rect 21861 24452 21885 24454
rect 21941 24452 21965 24454
rect 22021 24452 22027 24454
rect 21719 24443 22027 24452
rect 21640 24404 21692 24410
rect 21640 24346 21692 24352
rect 21640 23588 21692 23594
rect 21640 23530 21692 23536
rect 21652 23322 21680 23530
rect 21719 23420 22027 23429
rect 21719 23418 21725 23420
rect 21781 23418 21805 23420
rect 21861 23418 21885 23420
rect 21941 23418 21965 23420
rect 22021 23418 22027 23420
rect 21781 23366 21783 23418
rect 21963 23366 21965 23418
rect 21719 23364 21725 23366
rect 21781 23364 21805 23366
rect 21861 23364 21885 23366
rect 21941 23364 21965 23366
rect 22021 23364 22027 23366
rect 21719 23355 22027 23364
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 21719 22332 22027 22341
rect 21719 22330 21725 22332
rect 21781 22330 21805 22332
rect 21861 22330 21885 22332
rect 21941 22330 21965 22332
rect 22021 22330 22027 22332
rect 21781 22278 21783 22330
rect 21963 22278 21965 22330
rect 21719 22276 21725 22278
rect 21781 22276 21805 22278
rect 21861 22276 21885 22278
rect 21941 22276 21965 22278
rect 22021 22276 22027 22278
rect 21719 22267 22027 22276
rect 21824 22160 21876 22166
rect 21876 22108 21956 22114
rect 21824 22102 21956 22108
rect 21836 22086 21956 22102
rect 21928 21622 21956 22086
rect 22112 22094 22140 27610
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 22204 26874 22232 26930
rect 22204 26846 22324 26874
rect 22192 26784 22244 26790
rect 22192 26726 22244 26732
rect 22204 25838 22232 26726
rect 22296 26586 22324 26846
rect 22284 26580 22336 26586
rect 22284 26522 22336 26528
rect 22296 25906 22324 26522
rect 22468 26444 22520 26450
rect 22468 26386 22520 26392
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 22192 25832 22244 25838
rect 22192 25774 22244 25780
rect 22284 24676 22336 24682
rect 22284 24618 22336 24624
rect 22296 24206 22324 24618
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22388 23730 22416 24550
rect 22480 23730 22508 26386
rect 22560 25696 22612 25702
rect 22560 25638 22612 25644
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22480 23186 22508 23666
rect 22468 23180 22520 23186
rect 22468 23122 22520 23128
rect 22112 22066 22232 22094
rect 21916 21616 21968 21622
rect 21916 21558 21968 21564
rect 22008 21548 22060 21554
rect 22060 21508 22140 21536
rect 22008 21490 22060 21496
rect 21719 21244 22027 21253
rect 21719 21242 21725 21244
rect 21781 21242 21805 21244
rect 21861 21242 21885 21244
rect 21941 21242 21965 21244
rect 22021 21242 22027 21244
rect 21781 21190 21783 21242
rect 21963 21190 21965 21242
rect 21719 21188 21725 21190
rect 21781 21188 21805 21190
rect 21861 21188 21885 21190
rect 21941 21188 21965 21190
rect 22021 21188 22027 21190
rect 21719 21179 22027 21188
rect 22112 21146 22140 21508
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 21719 20156 22027 20165
rect 21719 20154 21725 20156
rect 21781 20154 21805 20156
rect 21861 20154 21885 20156
rect 21941 20154 21965 20156
rect 22021 20154 22027 20156
rect 21781 20102 21783 20154
rect 21963 20102 21965 20154
rect 21719 20100 21725 20102
rect 21781 20100 21805 20102
rect 21861 20100 21885 20102
rect 21941 20100 21965 20102
rect 22021 20100 22027 20102
rect 21719 20091 22027 20100
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21836 19378 21864 19790
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 21719 19068 22027 19077
rect 21719 19066 21725 19068
rect 21781 19066 21805 19068
rect 21861 19066 21885 19068
rect 21941 19066 21965 19068
rect 22021 19066 22027 19068
rect 21781 19014 21783 19066
rect 21963 19014 21965 19066
rect 21719 19012 21725 19014
rect 21781 19012 21805 19014
rect 21861 19012 21885 19014
rect 21941 19012 21965 19014
rect 22021 19012 22027 19014
rect 21719 19003 22027 19012
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21928 18290 21956 18566
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 21640 18284 21692 18290
rect 21640 18226 21692 18232
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 21418 18006 21496 18034
rect 21362 17983 21418 17992
rect 21652 17882 21680 18226
rect 21719 17980 22027 17989
rect 21719 17978 21725 17980
rect 21781 17978 21805 17980
rect 21861 17978 21885 17980
rect 21941 17978 21965 17980
rect 22021 17978 22027 17980
rect 21781 17926 21783 17978
rect 21963 17926 21965 17978
rect 21719 17924 21725 17926
rect 21781 17924 21805 17926
rect 21861 17924 21885 17926
rect 21941 17924 21965 17926
rect 22021 17924 22027 17926
rect 21719 17915 22027 17924
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 22112 17338 22140 18294
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21284 16590 21312 17138
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21272 16584 21324 16590
rect 21272 16526 21324 16532
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21376 15706 21404 15846
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21376 13274 21404 14214
rect 21560 13682 21588 16934
rect 21652 16046 21680 17070
rect 21719 16892 22027 16901
rect 21719 16890 21725 16892
rect 21781 16890 21805 16892
rect 21861 16890 21885 16892
rect 21941 16890 21965 16892
rect 22021 16890 22027 16892
rect 21781 16838 21783 16890
rect 21963 16838 21965 16890
rect 21719 16836 21725 16838
rect 21781 16836 21805 16838
rect 21861 16836 21885 16838
rect 21941 16836 21965 16838
rect 22021 16836 22027 16838
rect 21719 16827 22027 16836
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 21652 14958 21680 15982
rect 21719 15804 22027 15813
rect 21719 15802 21725 15804
rect 21781 15802 21805 15804
rect 21861 15802 21885 15804
rect 21941 15802 21965 15804
rect 22021 15802 22027 15804
rect 21781 15750 21783 15802
rect 21963 15750 21965 15802
rect 21719 15748 21725 15750
rect 21781 15748 21805 15750
rect 21861 15748 21885 15750
rect 21941 15748 21965 15750
rect 22021 15748 22027 15750
rect 21719 15739 22027 15748
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 21652 13870 21680 14894
rect 21719 14716 22027 14725
rect 21719 14714 21725 14716
rect 21781 14714 21805 14716
rect 21861 14714 21885 14716
rect 21941 14714 21965 14716
rect 22021 14714 22027 14716
rect 21781 14662 21783 14714
rect 21963 14662 21965 14714
rect 21719 14660 21725 14662
rect 21781 14660 21805 14662
rect 21861 14660 21885 14662
rect 21941 14660 21965 14662
rect 22021 14660 22027 14662
rect 21719 14651 22027 14660
rect 22204 14498 22232 22066
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22296 19854 22324 21966
rect 22480 21554 22508 23122
rect 22572 23050 22600 25638
rect 22560 23044 22612 23050
rect 22560 22986 22612 22992
rect 22664 22094 22692 33458
rect 22836 31680 22888 31686
rect 22836 31622 22888 31628
rect 22848 31482 22876 31622
rect 22836 31476 22888 31482
rect 22836 31418 22888 31424
rect 22836 30592 22888 30598
rect 22836 30534 22888 30540
rect 22848 30326 22876 30534
rect 22836 30320 22888 30326
rect 22836 30262 22888 30268
rect 22940 29730 22968 35498
rect 23216 35290 23244 40394
rect 23296 40044 23348 40050
rect 23296 39986 23348 39992
rect 23308 39098 23336 39986
rect 23400 39914 23428 40938
rect 23492 40633 23520 42656
rect 23572 42220 23624 42226
rect 23572 42162 23624 42168
rect 23478 40624 23534 40633
rect 23478 40559 23534 40568
rect 23478 40216 23534 40225
rect 23478 40151 23534 40160
rect 23492 40118 23520 40151
rect 23480 40112 23532 40118
rect 23480 40054 23532 40060
rect 23388 39908 23440 39914
rect 23388 39850 23440 39856
rect 23584 39642 23612 42162
rect 23676 41818 23704 43279
rect 23768 42294 23796 43438
rect 23848 42628 23900 42634
rect 23848 42570 23900 42576
rect 23756 42288 23808 42294
rect 23756 42230 23808 42236
rect 23756 42152 23808 42158
rect 23756 42094 23808 42100
rect 23664 41812 23716 41818
rect 23664 41754 23716 41760
rect 23664 40928 23716 40934
rect 23664 40870 23716 40876
rect 23676 40633 23704 40870
rect 23662 40624 23718 40633
rect 23662 40559 23718 40568
rect 23768 40372 23796 42094
rect 23860 41664 23888 42570
rect 23952 41818 23980 44840
rect 24122 42800 24178 42809
rect 24122 42735 24178 42744
rect 24136 42702 24164 42735
rect 24124 42696 24176 42702
rect 24124 42638 24176 42644
rect 24228 42362 24256 44840
rect 24216 42356 24268 42362
rect 24216 42298 24268 42304
rect 24030 42256 24086 42265
rect 24030 42191 24032 42200
rect 24084 42191 24086 42200
rect 24124 42220 24176 42226
rect 24032 42162 24084 42168
rect 24124 42162 24176 42168
rect 23940 41812 23992 41818
rect 23940 41754 23992 41760
rect 23860 41636 23980 41664
rect 23848 41540 23900 41546
rect 23848 41482 23900 41488
rect 23860 41313 23888 41482
rect 23846 41304 23902 41313
rect 23846 41239 23902 41248
rect 23952 40662 23980 41636
rect 24136 40662 24164 42162
rect 24320 41274 24348 44934
rect 24490 44840 24546 44934
rect 24596 44934 24822 44962
rect 24596 41818 24624 44934
rect 24766 44840 24822 44934
rect 25042 44840 25098 45000
rect 25318 44840 25374 45000
rect 25594 44840 25650 45000
rect 24686 43548 24994 43557
rect 24686 43546 24692 43548
rect 24748 43546 24772 43548
rect 24828 43546 24852 43548
rect 24908 43546 24932 43548
rect 24988 43546 24994 43548
rect 24748 43494 24750 43546
rect 24930 43494 24932 43546
rect 24686 43492 24692 43494
rect 24748 43492 24772 43494
rect 24828 43492 24852 43494
rect 24908 43492 24932 43494
rect 24988 43492 24994 43494
rect 24686 43483 24994 43492
rect 25056 42566 25084 44840
rect 25044 42560 25096 42566
rect 25044 42502 25096 42508
rect 24686 42460 24994 42469
rect 24686 42458 24692 42460
rect 24748 42458 24772 42460
rect 24828 42458 24852 42460
rect 24908 42458 24932 42460
rect 24988 42458 24994 42460
rect 24748 42406 24750 42458
rect 24930 42406 24932 42458
rect 24686 42404 24692 42406
rect 24748 42404 24772 42406
rect 24828 42404 24852 42406
rect 24908 42404 24932 42406
rect 24988 42404 24994 42406
rect 24686 42395 24994 42404
rect 25044 42220 25096 42226
rect 25044 42162 25096 42168
rect 24584 41812 24636 41818
rect 24584 41754 24636 41760
rect 24492 41472 24544 41478
rect 24492 41414 24544 41420
rect 24308 41268 24360 41274
rect 24308 41210 24360 41216
rect 23940 40656 23992 40662
rect 23940 40598 23992 40604
rect 24124 40656 24176 40662
rect 24124 40598 24176 40604
rect 23848 40452 23900 40458
rect 23848 40394 23900 40400
rect 24216 40452 24268 40458
rect 24216 40394 24268 40400
rect 23676 40344 23796 40372
rect 23676 40186 23704 40344
rect 23664 40180 23716 40186
rect 23664 40122 23716 40128
rect 23756 40180 23808 40186
rect 23756 40122 23808 40128
rect 23664 40044 23716 40050
rect 23664 39986 23716 39992
rect 23572 39636 23624 39642
rect 23572 39578 23624 39584
rect 23478 39536 23534 39545
rect 23478 39471 23534 39480
rect 23296 39092 23348 39098
rect 23296 39034 23348 39040
rect 23388 38956 23440 38962
rect 23388 38898 23440 38904
rect 23400 38010 23428 38898
rect 23492 38826 23520 39471
rect 23572 38888 23624 38894
rect 23572 38830 23624 38836
rect 23480 38820 23532 38826
rect 23480 38762 23532 38768
rect 23388 38004 23440 38010
rect 23388 37946 23440 37952
rect 23296 37868 23348 37874
rect 23296 37810 23348 37816
rect 23308 37466 23336 37810
rect 23388 37664 23440 37670
rect 23388 37606 23440 37612
rect 23296 37460 23348 37466
rect 23296 37402 23348 37408
rect 23308 37330 23336 37402
rect 23296 37324 23348 37330
rect 23296 37266 23348 37272
rect 23296 36236 23348 36242
rect 23296 36178 23348 36184
rect 23308 35834 23336 36178
rect 23296 35828 23348 35834
rect 23296 35770 23348 35776
rect 23204 35284 23256 35290
rect 23204 35226 23256 35232
rect 23204 34944 23256 34950
rect 23204 34886 23256 34892
rect 23216 34610 23244 34886
rect 23020 34604 23072 34610
rect 23020 34546 23072 34552
rect 23204 34604 23256 34610
rect 23204 34546 23256 34552
rect 23032 34474 23060 34546
rect 23400 34474 23428 37606
rect 23480 37256 23532 37262
rect 23480 37198 23532 37204
rect 23492 36310 23520 37198
rect 23584 36922 23612 38830
rect 23676 37262 23704 39986
rect 23768 39953 23796 40122
rect 23754 39944 23810 39953
rect 23754 39879 23810 39888
rect 23860 39273 23888 40394
rect 24228 40089 24256 40394
rect 24214 40080 24270 40089
rect 24032 40044 24084 40050
rect 24214 40015 24270 40024
rect 24032 39986 24084 39992
rect 23846 39264 23902 39273
rect 23846 39199 23902 39208
rect 24044 39114 24072 39986
rect 24400 39840 24452 39846
rect 24400 39782 24452 39788
rect 24412 39545 24440 39782
rect 24398 39536 24454 39545
rect 24398 39471 24454 39480
rect 24124 39296 24176 39302
rect 24124 39238 24176 39244
rect 23952 39086 24072 39114
rect 23952 38826 23980 39086
rect 24136 39001 24164 39238
rect 24122 38992 24178 39001
rect 24032 38956 24084 38962
rect 24122 38927 24178 38936
rect 24032 38898 24084 38904
rect 23940 38820 23992 38826
rect 23940 38762 23992 38768
rect 24044 38554 24072 38898
rect 24400 38752 24452 38758
rect 24400 38694 24452 38700
rect 24412 38593 24440 38694
rect 24398 38584 24454 38593
rect 24032 38548 24084 38554
rect 24398 38519 24454 38528
rect 24032 38490 24084 38496
rect 24124 38208 24176 38214
rect 24124 38150 24176 38156
rect 24136 37913 24164 38150
rect 24122 37904 24178 37913
rect 23848 37868 23900 37874
rect 24122 37839 24178 37848
rect 23848 37810 23900 37816
rect 23860 37466 23888 37810
rect 24032 37664 24084 37670
rect 24032 37606 24084 37612
rect 24400 37664 24452 37670
rect 24400 37606 24452 37612
rect 23848 37460 23900 37466
rect 23848 37402 23900 37408
rect 23756 37392 23808 37398
rect 23756 37334 23808 37340
rect 23664 37256 23716 37262
rect 23664 37198 23716 37204
rect 23572 36916 23624 36922
rect 23572 36858 23624 36864
rect 23480 36304 23532 36310
rect 23480 36246 23532 36252
rect 23768 35714 23796 37334
rect 23848 37256 23900 37262
rect 23848 37198 23900 37204
rect 23940 37256 23992 37262
rect 23940 37198 23992 37204
rect 23860 35834 23888 37198
rect 23952 36922 23980 37198
rect 23940 36916 23992 36922
rect 23940 36858 23992 36864
rect 24044 36854 24072 37606
rect 24412 37369 24440 37606
rect 24398 37360 24454 37369
rect 24398 37295 24454 37304
rect 24124 37120 24176 37126
rect 24124 37062 24176 37068
rect 24032 36848 24084 36854
rect 24136 36825 24164 37062
rect 24032 36790 24084 36796
rect 24122 36816 24178 36825
rect 24122 36751 24178 36760
rect 24400 36576 24452 36582
rect 24400 36518 24452 36524
rect 24308 36304 24360 36310
rect 24412 36281 24440 36518
rect 24308 36246 24360 36252
rect 24398 36272 24454 36281
rect 24124 36032 24176 36038
rect 24124 35974 24176 35980
rect 24136 35873 24164 35974
rect 24122 35864 24178 35873
rect 23848 35828 23900 35834
rect 24122 35799 24178 35808
rect 23848 35770 23900 35776
rect 23768 35686 24072 35714
rect 23572 35012 23624 35018
rect 23572 34954 23624 34960
rect 23584 34746 23612 34954
rect 23572 34740 23624 34746
rect 23572 34682 23624 34688
rect 23020 34468 23072 34474
rect 23020 34410 23072 34416
rect 23388 34468 23440 34474
rect 23388 34410 23440 34416
rect 23296 33992 23348 33998
rect 23296 33934 23348 33940
rect 23664 33992 23716 33998
rect 23664 33934 23716 33940
rect 23308 33658 23336 33934
rect 23388 33856 23440 33862
rect 23388 33798 23440 33804
rect 23400 33658 23428 33798
rect 23676 33658 23704 33934
rect 23296 33652 23348 33658
rect 23296 33594 23348 33600
rect 23388 33652 23440 33658
rect 23388 33594 23440 33600
rect 23664 33652 23716 33658
rect 23664 33594 23716 33600
rect 23296 33516 23348 33522
rect 23296 33458 23348 33464
rect 23940 33516 23992 33522
rect 23940 33458 23992 33464
rect 23308 33114 23336 33458
rect 23848 33312 23900 33318
rect 23848 33254 23900 33260
rect 23296 33108 23348 33114
rect 23296 33050 23348 33056
rect 23860 32910 23888 33254
rect 23480 32904 23532 32910
rect 23480 32846 23532 32852
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23296 32768 23348 32774
rect 23296 32710 23348 32716
rect 23112 32292 23164 32298
rect 23112 32234 23164 32240
rect 23020 31408 23072 31414
rect 23020 31350 23072 31356
rect 23032 30938 23060 31350
rect 23020 30932 23072 30938
rect 23020 30874 23072 30880
rect 23124 30818 23152 32234
rect 23308 31754 23336 32710
rect 23492 32570 23520 32846
rect 23572 32768 23624 32774
rect 23572 32710 23624 32716
rect 23584 32570 23612 32710
rect 23480 32564 23532 32570
rect 23480 32506 23532 32512
rect 23572 32564 23624 32570
rect 23572 32506 23624 32512
rect 23756 32496 23808 32502
rect 23756 32438 23808 32444
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 23296 31748 23348 31754
rect 23296 31690 23348 31696
rect 23204 31136 23256 31142
rect 23204 31078 23256 31084
rect 23216 30938 23244 31078
rect 23400 30938 23428 32370
rect 23572 32360 23624 32366
rect 23572 32302 23624 32308
rect 23480 32224 23532 32230
rect 23480 32166 23532 32172
rect 23492 31890 23520 32166
rect 23480 31884 23532 31890
rect 23480 31826 23532 31832
rect 23584 31822 23612 32302
rect 23662 31920 23718 31929
rect 23662 31855 23718 31864
rect 23676 31822 23704 31855
rect 23572 31816 23624 31822
rect 23572 31758 23624 31764
rect 23664 31816 23716 31822
rect 23664 31758 23716 31764
rect 23480 31476 23532 31482
rect 23480 31418 23532 31424
rect 23204 30932 23256 30938
rect 23204 30874 23256 30880
rect 23388 30932 23440 30938
rect 23388 30874 23440 30880
rect 23124 30790 23244 30818
rect 23216 30734 23244 30790
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23018 30424 23074 30433
rect 23018 30359 23074 30368
rect 23032 30258 23060 30359
rect 23202 30288 23258 30297
rect 23020 30252 23072 30258
rect 23202 30223 23258 30232
rect 23388 30252 23440 30258
rect 23020 30194 23072 30200
rect 22940 29702 23152 29730
rect 22928 29572 22980 29578
rect 22928 29514 22980 29520
rect 22940 29034 22968 29514
rect 22928 29028 22980 29034
rect 22928 28970 22980 28976
rect 22744 27464 22796 27470
rect 22744 27406 22796 27412
rect 22756 27062 22784 27406
rect 22836 27328 22888 27334
rect 22836 27270 22888 27276
rect 22744 27056 22796 27062
rect 22744 26998 22796 27004
rect 22848 26042 22876 27270
rect 23020 26784 23072 26790
rect 23020 26726 23072 26732
rect 22836 26036 22888 26042
rect 22836 25978 22888 25984
rect 22928 24608 22980 24614
rect 22928 24550 22980 24556
rect 22940 24410 22968 24550
rect 22928 24404 22980 24410
rect 22928 24346 22980 24352
rect 22836 23724 22888 23730
rect 22836 23666 22888 23672
rect 22744 23248 22796 23254
rect 22744 23190 22796 23196
rect 22572 22066 22692 22094
rect 22468 21548 22520 21554
rect 22388 21508 22468 21536
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22388 19378 22416 21508
rect 22468 21490 22520 21496
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22480 21146 22508 21286
rect 22468 21140 22520 21146
rect 22468 21082 22520 21088
rect 22572 20618 22600 22066
rect 22652 21956 22704 21962
rect 22652 21898 22704 21904
rect 22664 21690 22692 21898
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22652 21412 22704 21418
rect 22652 21354 22704 21360
rect 22664 21146 22692 21354
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22480 20590 22600 20618
rect 22756 20602 22784 23190
rect 22848 20874 22876 23666
rect 23032 22094 23060 26726
rect 23124 26382 23152 29702
rect 23216 28370 23244 30223
rect 23388 30194 23440 30200
rect 23400 29782 23428 30194
rect 23388 29776 23440 29782
rect 23388 29718 23440 29724
rect 23294 29200 23350 29209
rect 23294 29135 23350 29144
rect 23308 28558 23336 29135
rect 23388 29028 23440 29034
rect 23388 28970 23440 28976
rect 23400 28762 23428 28970
rect 23388 28756 23440 28762
rect 23388 28698 23440 28704
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23216 28342 23336 28370
rect 23112 26376 23164 26382
rect 23112 26318 23164 26324
rect 23124 23798 23152 26318
rect 23204 24812 23256 24818
rect 23204 24754 23256 24760
rect 23216 24410 23244 24754
rect 23204 24404 23256 24410
rect 23204 24346 23256 24352
rect 23112 23792 23164 23798
rect 23112 23734 23164 23740
rect 23110 23488 23166 23497
rect 23110 23423 23166 23432
rect 22940 22066 23060 22094
rect 22836 20868 22888 20874
rect 22836 20810 22888 20816
rect 22744 20596 22796 20602
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 22296 17882 22324 18362
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 22480 17626 22508 20590
rect 22744 20538 22796 20544
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22572 19786 22600 20402
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22560 19780 22612 19786
rect 22560 19722 22612 19728
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22664 17678 22692 19654
rect 22756 18766 22784 20198
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22756 17678 22784 18022
rect 22296 17598 22508 17626
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22744 17672 22796 17678
rect 22744 17614 22796 17620
rect 22296 16250 22324 17598
rect 22376 17536 22428 17542
rect 22376 17478 22428 17484
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22388 16726 22416 17478
rect 22572 17202 22600 17478
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 22376 16720 22428 16726
rect 22376 16662 22428 16668
rect 22480 16590 22508 16934
rect 22572 16674 22600 17138
rect 22664 16794 22692 17614
rect 22744 17060 22796 17066
rect 22744 17002 22796 17008
rect 22756 16794 22784 17002
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22572 16646 22784 16674
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22572 15706 22600 16390
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22112 14470 22232 14498
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21560 13654 21680 13682
rect 21376 13246 21588 13274
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21192 12442 21220 12786
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 21100 12294 21220 12322
rect 21088 12164 21140 12170
rect 21088 12106 21140 12112
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20720 7880 20772 7886
rect 20548 7806 20668 7834
rect 20720 7822 20772 7828
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20548 7546 20576 7686
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20640 6458 20668 7806
rect 20732 7546 20760 7822
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20824 7206 20852 8774
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20718 6760 20774 6769
rect 20718 6695 20720 6704
rect 20772 6695 20774 6704
rect 20720 6666 20772 6672
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20640 5914 20668 6258
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20732 5545 20760 6054
rect 20916 5778 20944 10406
rect 20996 9988 21048 9994
rect 20996 9930 21048 9936
rect 21008 9450 21036 9930
rect 21100 9874 21128 12106
rect 21192 11064 21220 12294
rect 21284 11744 21312 12582
rect 21376 11898 21404 12786
rect 21468 12170 21496 12786
rect 21560 12442 21588 13246
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21364 11756 21416 11762
rect 21284 11716 21364 11744
rect 21364 11698 21416 11704
rect 21192 11036 21312 11064
rect 21178 10976 21234 10985
rect 21178 10911 21234 10920
rect 21192 10062 21220 10911
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21100 9846 21220 9874
rect 20996 9444 21048 9450
rect 20996 9386 21048 9392
rect 21008 8090 21036 9386
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21100 7342 21128 8434
rect 21088 7336 21140 7342
rect 21086 7304 21088 7313
rect 21140 7304 21142 7313
rect 21086 7239 21142 7248
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 20812 5568 20864 5574
rect 20718 5536 20774 5545
rect 20812 5510 20864 5516
rect 20718 5471 20774 5480
rect 20718 5400 20774 5409
rect 20718 5335 20720 5344
rect 20772 5335 20774 5344
rect 20720 5306 20772 5312
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20732 4826 20760 5170
rect 20824 5166 20852 5510
rect 20916 5370 20944 5714
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20536 4684 20588 4690
rect 20588 4644 20852 4672
rect 20536 4626 20588 4632
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20456 4214 20484 4558
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20718 4448 20774 4457
rect 20444 4208 20496 4214
rect 20444 4150 20496 4156
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20456 3913 20484 4014
rect 20442 3904 20498 3913
rect 20442 3839 20498 3848
rect 20352 2100 20404 2106
rect 20352 2042 20404 2048
rect 20456 1986 20484 3839
rect 20548 3097 20576 4422
rect 20718 4383 20774 4392
rect 20732 3754 20760 4383
rect 20640 3726 20760 3754
rect 20640 3482 20668 3726
rect 20718 3632 20774 3641
rect 20718 3567 20720 3576
rect 20772 3567 20774 3576
rect 20720 3538 20772 3544
rect 20640 3454 20760 3482
rect 20534 3088 20590 3097
rect 20534 3023 20590 3032
rect 20732 2922 20760 3454
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20824 2514 20852 4644
rect 21008 4554 21036 5714
rect 21100 5250 21128 7142
rect 21192 6118 21220 9846
rect 21284 9722 21312 11036
rect 21560 9994 21588 12106
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21272 9716 21324 9722
rect 21324 9676 21404 9704
rect 21272 9658 21324 9664
rect 21376 9382 21404 9676
rect 21548 9512 21600 9518
rect 21652 9489 21680 13654
rect 21719 13628 22027 13637
rect 21719 13626 21725 13628
rect 21781 13626 21805 13628
rect 21861 13626 21885 13628
rect 21941 13626 21965 13628
rect 22021 13626 22027 13628
rect 21781 13574 21783 13626
rect 21963 13574 21965 13626
rect 21719 13572 21725 13574
rect 21781 13572 21805 13574
rect 21861 13572 21885 13574
rect 21941 13572 21965 13574
rect 22021 13572 22027 13574
rect 21719 13563 22027 13572
rect 22112 13274 22140 14470
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22204 14074 22232 14350
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22020 13246 22140 13274
rect 22020 12866 22048 13246
rect 22020 12838 22140 12866
rect 21719 12540 22027 12549
rect 21719 12538 21725 12540
rect 21781 12538 21805 12540
rect 21861 12538 21885 12540
rect 21941 12538 21965 12540
rect 22021 12538 22027 12540
rect 21781 12486 21783 12538
rect 21963 12486 21965 12538
rect 21719 12484 21725 12486
rect 21781 12484 21805 12486
rect 21861 12484 21885 12486
rect 21941 12484 21965 12486
rect 22021 12484 22027 12486
rect 21719 12475 22027 12484
rect 22112 12322 22140 12838
rect 22020 12306 22140 12322
rect 22008 12300 22140 12306
rect 22060 12294 22140 12300
rect 22008 12242 22060 12248
rect 22204 12186 22232 13874
rect 22296 13530 22324 14214
rect 22480 13938 22508 15302
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22572 14618 22600 14962
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22664 13394 22692 15438
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22468 13184 22520 13190
rect 22756 13138 22784 16646
rect 22468 13126 22520 13132
rect 22388 12850 22416 13126
rect 22480 12986 22508 13126
rect 22572 13110 22784 13138
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22112 12158 22232 12186
rect 21916 11824 21968 11830
rect 21914 11792 21916 11801
rect 21968 11792 21970 11801
rect 21914 11727 21970 11736
rect 21719 11452 22027 11461
rect 21719 11450 21725 11452
rect 21781 11450 21805 11452
rect 21861 11450 21885 11452
rect 21941 11450 21965 11452
rect 22021 11450 22027 11452
rect 21781 11398 21783 11450
rect 21963 11398 21965 11450
rect 21719 11396 21725 11398
rect 21781 11396 21805 11398
rect 21861 11396 21885 11398
rect 21941 11396 21965 11398
rect 22021 11396 22027 11398
rect 21719 11387 22027 11396
rect 22112 11150 22140 12158
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 22204 11898 22232 12038
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22374 11792 22430 11801
rect 22374 11727 22430 11736
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 22388 11064 22416 11727
rect 22480 11694 22508 12038
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22480 11354 22508 11494
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22388 11036 22508 11064
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 22100 10600 22152 10606
rect 22100 10542 22152 10548
rect 21719 10364 22027 10373
rect 21719 10362 21725 10364
rect 21781 10362 21805 10364
rect 21861 10362 21885 10364
rect 21941 10362 21965 10364
rect 22021 10362 22027 10364
rect 21781 10310 21783 10362
rect 21963 10310 21965 10362
rect 21719 10308 21725 10310
rect 21781 10308 21805 10310
rect 21861 10308 21885 10310
rect 21941 10308 21965 10310
rect 22021 10308 22027 10310
rect 21719 10299 22027 10308
rect 22112 10198 22140 10542
rect 22388 10266 22416 10610
rect 22376 10260 22428 10266
rect 22376 10202 22428 10208
rect 22100 10192 22152 10198
rect 22100 10134 22152 10140
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 21744 9722 21772 9998
rect 21732 9716 21784 9722
rect 21732 9658 21784 9664
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 21548 9454 21600 9460
rect 21638 9480 21694 9489
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21560 8430 21588 9454
rect 21638 9415 21694 9424
rect 21719 9276 22027 9285
rect 21719 9274 21725 9276
rect 21781 9274 21805 9276
rect 21861 9274 21885 9276
rect 21941 9274 21965 9276
rect 22021 9274 22027 9276
rect 21781 9222 21783 9274
rect 21963 9222 21965 9274
rect 21719 9220 21725 9222
rect 21781 9220 21805 9222
rect 21861 9220 21885 9222
rect 21941 9220 21965 9222
rect 22021 9220 22027 9222
rect 21719 9211 22027 9220
rect 21640 9036 21692 9042
rect 21640 8978 21692 8984
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21284 7002 21312 7278
rect 21468 7002 21496 7482
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21560 6866 21588 8366
rect 21652 8362 21680 8978
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 21836 8634 21864 8910
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21640 8356 21692 8362
rect 21640 8298 21692 8304
rect 22100 8288 22152 8294
rect 22100 8230 22152 8236
rect 21719 8188 22027 8197
rect 21719 8186 21725 8188
rect 21781 8186 21805 8188
rect 21861 8186 21885 8188
rect 21941 8186 21965 8188
rect 22021 8186 22027 8188
rect 21781 8134 21783 8186
rect 21963 8134 21965 8186
rect 21719 8132 21725 8134
rect 21781 8132 21805 8134
rect 21861 8132 21885 8134
rect 21941 8132 21965 8134
rect 22021 8132 22027 8134
rect 21719 8123 22027 8132
rect 22112 7834 22140 8230
rect 22020 7806 22140 7834
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 22020 7478 22048 7806
rect 22204 7750 22232 7822
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22008 7472 22060 7478
rect 22008 7414 22060 7420
rect 22112 7410 22140 7686
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 21719 7100 22027 7109
rect 21719 7098 21725 7100
rect 21781 7098 21805 7100
rect 21861 7098 21885 7100
rect 21941 7098 21965 7100
rect 22021 7098 22027 7100
rect 21781 7046 21783 7098
rect 21963 7046 21965 7098
rect 21719 7044 21725 7046
rect 21781 7044 21805 7046
rect 21861 7044 21885 7046
rect 21941 7044 21965 7046
rect 22021 7044 22027 7046
rect 21719 7035 22027 7044
rect 21916 6996 21968 7002
rect 21916 6938 21968 6944
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21376 6458 21404 6598
rect 21364 6452 21416 6458
rect 21364 6394 21416 6400
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 21192 5370 21220 5850
rect 21284 5817 21312 6258
rect 21270 5808 21326 5817
rect 21270 5743 21326 5752
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21284 5370 21312 5646
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 21100 5222 21312 5250
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 21088 4548 21140 4554
rect 21088 4490 21140 4496
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 21008 3466 21036 3878
rect 20996 3460 21048 3466
rect 20996 3402 21048 3408
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 20824 2417 20852 2450
rect 20810 2408 20866 2417
rect 20628 2372 20680 2378
rect 20810 2343 20866 2352
rect 20628 2314 20680 2320
rect 20640 2122 20668 2314
rect 20640 2094 20852 2122
rect 20260 1964 20312 1970
rect 20260 1906 20312 1912
rect 20364 1958 20484 1986
rect 20720 1964 20772 1970
rect 20168 1760 20220 1766
rect 20168 1702 20220 1708
rect 20364 1358 20392 1958
rect 20720 1906 20772 1912
rect 20732 1442 20760 1906
rect 20640 1414 20760 1442
rect 20352 1352 20404 1358
rect 20352 1294 20404 1300
rect 20444 1352 20496 1358
rect 20444 1294 20496 1300
rect 19798 54 19932 82
rect 19798 0 19854 54
rect 20074 0 20130 160
rect 20350 82 20406 160
rect 20456 82 20484 1294
rect 20640 160 20668 1414
rect 20350 54 20484 82
rect 20350 0 20406 54
rect 20626 0 20682 160
rect 20824 82 20852 2094
rect 20916 1222 20944 2926
rect 20996 1352 21048 1358
rect 20994 1320 20996 1329
rect 21048 1320 21050 1329
rect 20994 1255 21050 1264
rect 20904 1216 20956 1222
rect 20904 1158 20956 1164
rect 21100 921 21128 4490
rect 21284 4298 21312 5222
rect 21376 4457 21404 6258
rect 21468 5846 21496 6394
rect 21560 6254 21588 6802
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21560 5914 21588 6054
rect 21652 5914 21680 6666
rect 21928 6186 21956 6938
rect 22112 6322 22140 7346
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 22204 6322 22232 7142
rect 22296 6322 22324 7142
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 21916 6180 21968 6186
rect 21916 6122 21968 6128
rect 22192 6180 22244 6186
rect 22192 6122 22244 6128
rect 21719 6012 22027 6021
rect 21719 6010 21725 6012
rect 21781 6010 21805 6012
rect 21861 6010 21885 6012
rect 21941 6010 21965 6012
rect 22021 6010 22027 6012
rect 21781 5958 21783 6010
rect 21963 5958 21965 6010
rect 21719 5956 21725 5958
rect 21781 5956 21805 5958
rect 21861 5956 21885 5958
rect 21941 5956 21965 5958
rect 22021 5956 22027 5958
rect 21719 5947 22027 5956
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 21456 5840 21508 5846
rect 21456 5782 21508 5788
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 21640 5704 21692 5710
rect 21638 5672 21640 5681
rect 21692 5672 21694 5681
rect 21638 5607 21694 5616
rect 21548 5160 21600 5166
rect 21548 5102 21600 5108
rect 21560 4826 21588 5102
rect 21744 5012 21772 5782
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 21928 5273 21956 5646
rect 22112 5273 22140 5646
rect 21914 5264 21970 5273
rect 21914 5199 21970 5208
rect 22098 5264 22154 5273
rect 22098 5199 22154 5208
rect 21652 4984 21772 5012
rect 21548 4820 21600 4826
rect 21548 4762 21600 4768
rect 21362 4448 21418 4457
rect 21362 4383 21418 4392
rect 21284 4270 21404 4298
rect 21180 3936 21232 3942
rect 21178 3904 21180 3913
rect 21232 3904 21234 3913
rect 21178 3839 21234 3848
rect 21178 3768 21234 3777
rect 21376 3754 21404 4270
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21456 3936 21508 3942
rect 21454 3904 21456 3913
rect 21508 3904 21510 3913
rect 21454 3839 21510 3848
rect 21376 3726 21496 3754
rect 21178 3703 21234 3712
rect 21192 2009 21220 3703
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 21178 2000 21234 2009
rect 21178 1935 21234 1944
rect 21284 1494 21312 2790
rect 21376 2122 21404 3606
rect 21468 2378 21496 3726
rect 21560 2854 21588 4082
rect 21652 3534 21680 4984
rect 21719 4924 22027 4933
rect 21719 4922 21725 4924
rect 21781 4922 21805 4924
rect 21861 4922 21885 4924
rect 21941 4922 21965 4924
rect 22021 4922 22027 4924
rect 21781 4870 21783 4922
rect 21963 4870 21965 4922
rect 21719 4868 21725 4870
rect 21781 4868 21805 4870
rect 21861 4868 21885 4870
rect 21941 4868 21965 4870
rect 22021 4868 22027 4870
rect 21719 4859 22027 4868
rect 21914 4312 21970 4321
rect 21970 4270 22048 4298
rect 21914 4247 21970 4256
rect 22020 3924 22048 4270
rect 22100 4140 22152 4146
rect 22204 4128 22232 6122
rect 22282 5536 22338 5545
rect 22282 5471 22338 5480
rect 22296 5370 22324 5471
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22152 4100 22232 4128
rect 22100 4082 22152 4088
rect 22296 4060 22324 5170
rect 22388 4826 22416 9658
rect 22480 7002 22508 11036
rect 22572 7886 22600 13110
rect 22652 12436 22704 12442
rect 22848 12434 22876 20198
rect 22940 16028 22968 22066
rect 23018 21584 23074 21593
rect 23018 21519 23020 21528
rect 23072 21519 23074 21528
rect 23020 21490 23072 21496
rect 23124 17649 23152 23423
rect 23204 22976 23256 22982
rect 23204 22918 23256 22924
rect 23216 22778 23244 22918
rect 23204 22772 23256 22778
rect 23204 22714 23256 22720
rect 23308 19854 23336 28342
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23400 25498 23428 25842
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 23492 25362 23520 31418
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23584 30394 23612 30534
rect 23572 30388 23624 30394
rect 23572 30330 23624 30336
rect 23572 30252 23624 30258
rect 23572 30194 23624 30200
rect 23584 29850 23612 30194
rect 23572 29844 23624 29850
rect 23572 29786 23624 29792
rect 23664 28552 23716 28558
rect 23584 28500 23664 28506
rect 23584 28494 23716 28500
rect 23584 28478 23704 28494
rect 23584 28218 23612 28478
rect 23664 28416 23716 28422
rect 23664 28358 23716 28364
rect 23676 28218 23704 28358
rect 23572 28212 23624 28218
rect 23572 28154 23624 28160
rect 23664 28212 23716 28218
rect 23664 28154 23716 28160
rect 23664 27872 23716 27878
rect 23664 27814 23716 27820
rect 23676 27470 23704 27814
rect 23768 27470 23796 32438
rect 23952 31482 23980 33458
rect 23940 31476 23992 31482
rect 23940 31418 23992 31424
rect 23848 30660 23900 30666
rect 23848 30602 23900 30608
rect 23860 30054 23888 30602
rect 23848 30048 23900 30054
rect 23848 29990 23900 29996
rect 23940 28960 23992 28966
rect 23940 28902 23992 28908
rect 23848 28688 23900 28694
rect 23848 28630 23900 28636
rect 23860 28200 23888 28630
rect 23952 28558 23980 28902
rect 23940 28552 23992 28558
rect 23940 28494 23992 28500
rect 23860 28172 23980 28200
rect 23848 28076 23900 28082
rect 23848 28018 23900 28024
rect 23860 27674 23888 28018
rect 23848 27668 23900 27674
rect 23848 27610 23900 27616
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23756 27464 23808 27470
rect 23756 27406 23808 27412
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 23584 27033 23612 27270
rect 23570 27024 23626 27033
rect 23570 26959 23626 26968
rect 23756 26784 23808 26790
rect 23756 26726 23808 26732
rect 23480 25356 23532 25362
rect 23480 25298 23532 25304
rect 23768 25294 23796 26726
rect 23848 26240 23900 26246
rect 23848 26182 23900 26188
rect 23860 26042 23888 26182
rect 23848 26036 23900 26042
rect 23848 25978 23900 25984
rect 23952 25974 23980 28172
rect 23940 25968 23992 25974
rect 23940 25910 23992 25916
rect 23848 25696 23900 25702
rect 23848 25638 23900 25644
rect 23756 25288 23808 25294
rect 23756 25230 23808 25236
rect 23400 24942 23612 24970
rect 23400 24818 23428 24942
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23492 23866 23520 24754
rect 23584 24698 23612 24942
rect 23584 24670 23796 24698
rect 23572 24608 23624 24614
rect 23572 24550 23624 24556
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23584 24410 23612 24550
rect 23572 24404 23624 24410
rect 23572 24346 23624 24352
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 23492 23322 23520 23802
rect 23584 23322 23612 24006
rect 23480 23316 23532 23322
rect 23480 23258 23532 23264
rect 23572 23316 23624 23322
rect 23572 23258 23624 23264
rect 23676 23254 23704 24550
rect 23664 23248 23716 23254
rect 23664 23190 23716 23196
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23400 22681 23428 23054
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23676 22681 23704 22918
rect 23768 22778 23796 24670
rect 23756 22772 23808 22778
rect 23756 22714 23808 22720
rect 23386 22672 23442 22681
rect 23662 22672 23718 22681
rect 23386 22607 23442 22616
rect 23572 22636 23624 22642
rect 23662 22607 23718 22616
rect 23572 22578 23624 22584
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23492 21486 23520 22374
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23584 20602 23612 22578
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 23676 21690 23704 22510
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 23572 20596 23624 20602
rect 23572 20538 23624 20544
rect 23768 20534 23796 21830
rect 23860 20534 23888 25638
rect 23940 25356 23992 25362
rect 23940 25298 23992 25304
rect 23952 24206 23980 25298
rect 23940 24200 23992 24206
rect 24044 24177 24072 35686
rect 24124 35692 24176 35698
rect 24124 35634 24176 35640
rect 24136 35290 24164 35634
rect 24124 35284 24176 35290
rect 24124 35226 24176 35232
rect 24216 35012 24268 35018
rect 24216 34954 24268 34960
rect 24228 34649 24256 34954
rect 24214 34640 24270 34649
rect 24214 34575 24270 34584
rect 24124 33856 24176 33862
rect 24124 33798 24176 33804
rect 24136 33561 24164 33798
rect 24122 33552 24178 33561
rect 24122 33487 24178 33496
rect 24124 32768 24176 32774
rect 24124 32710 24176 32716
rect 24136 32473 24164 32710
rect 24122 32464 24178 32473
rect 24122 32399 24178 32408
rect 24216 31816 24268 31822
rect 24216 31758 24268 31764
rect 24228 31657 24256 31758
rect 24214 31648 24270 31657
rect 24214 31583 24270 31592
rect 24216 30660 24268 30666
rect 24216 30602 24268 30608
rect 24228 30297 24256 30602
rect 24214 30288 24270 30297
rect 24214 30223 24270 30232
rect 24216 29572 24268 29578
rect 24216 29514 24268 29520
rect 24228 29209 24256 29514
rect 24214 29200 24270 29209
rect 24124 29164 24176 29170
rect 24214 29135 24270 29144
rect 24124 29106 24176 29112
rect 24136 29073 24164 29106
rect 24122 29064 24178 29073
rect 24122 28999 24178 29008
rect 24124 28416 24176 28422
rect 24124 28358 24176 28364
rect 24136 28121 24164 28358
rect 24122 28112 24178 28121
rect 24122 28047 24178 28056
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 24228 26489 24256 26726
rect 24214 26480 24270 26489
rect 24214 26415 24270 26424
rect 24124 25152 24176 25158
rect 24124 25094 24176 25100
rect 24136 24857 24164 25094
rect 24122 24848 24178 24857
rect 24122 24783 24178 24792
rect 23940 24142 23992 24148
rect 24030 24168 24086 24177
rect 24030 24103 24086 24112
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24136 23769 24164 24006
rect 24122 23760 24178 23769
rect 24032 23724 24084 23730
rect 24122 23695 24178 23704
rect 24032 23666 24084 23672
rect 23940 23520 23992 23526
rect 23940 23462 23992 23468
rect 23952 22094 23980 23462
rect 24044 23322 24072 23666
rect 24032 23316 24084 23322
rect 24032 23258 24084 23264
rect 23952 22066 24072 22094
rect 23940 20800 23992 20806
rect 23940 20742 23992 20748
rect 23952 20641 23980 20742
rect 23938 20632 23994 20641
rect 23938 20567 23994 20576
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23848 20528 23900 20534
rect 23848 20470 23900 20476
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23768 19961 23796 20198
rect 23848 20052 23900 20058
rect 23848 19994 23900 20000
rect 23754 19952 23810 19961
rect 23754 19887 23810 19896
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23492 18766 23520 19110
rect 23584 18766 23612 19654
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23480 18760 23532 18766
rect 23400 18720 23480 18748
rect 23400 18426 23428 18720
rect 23480 18702 23532 18708
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23492 18426 23520 18566
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23110 17640 23166 17649
rect 23110 17575 23166 17584
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 23032 16250 23060 17274
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 23308 16590 23336 16934
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 23020 16040 23072 16046
rect 22940 16000 23020 16028
rect 23020 15982 23072 15988
rect 23124 15910 23152 16526
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 23124 15586 23152 15846
rect 23400 15706 23428 16390
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23124 15558 23244 15586
rect 23216 15502 23244 15558
rect 23584 15502 23612 18566
rect 23676 18426 23704 18770
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23768 17338 23796 18226
rect 23756 17332 23808 17338
rect 23756 17274 23808 17280
rect 23860 16114 23888 19994
rect 24044 19446 24072 22066
rect 24124 21888 24176 21894
rect 24124 21830 24176 21836
rect 24136 21593 24164 21830
rect 24122 21584 24178 21593
rect 24122 21519 24178 21528
rect 24320 21434 24348 36246
rect 24398 36207 24454 36216
rect 24400 35488 24452 35494
rect 24400 35430 24452 35436
rect 24412 35193 24440 35430
rect 24398 35184 24454 35193
rect 24398 35119 24454 35128
rect 24400 34536 24452 34542
rect 24398 34504 24400 34513
rect 24452 34504 24454 34513
rect 24398 34439 24454 34448
rect 24504 34202 24532 41414
rect 24686 41372 24994 41381
rect 24686 41370 24692 41372
rect 24748 41370 24772 41372
rect 24828 41370 24852 41372
rect 24908 41370 24932 41372
rect 24988 41370 24994 41372
rect 24748 41318 24750 41370
rect 24930 41318 24932 41370
rect 24686 41316 24692 41318
rect 24748 41316 24772 41318
rect 24828 41316 24852 41318
rect 24908 41316 24932 41318
rect 24988 41316 24994 41318
rect 24686 41307 24994 41316
rect 25056 41177 25084 42162
rect 25042 41168 25098 41177
rect 25042 41103 25098 41112
rect 25332 40730 25360 44840
rect 25608 42158 25636 44840
rect 25596 42152 25648 42158
rect 25596 42094 25648 42100
rect 25688 42016 25740 42022
rect 25688 41958 25740 41964
rect 25700 41414 25728 41958
rect 25700 41386 25820 41414
rect 25320 40724 25372 40730
rect 25320 40666 25372 40672
rect 24686 40284 24994 40293
rect 24686 40282 24692 40284
rect 24748 40282 24772 40284
rect 24828 40282 24852 40284
rect 24908 40282 24932 40284
rect 24988 40282 24994 40284
rect 24748 40230 24750 40282
rect 24930 40230 24932 40282
rect 24686 40228 24692 40230
rect 24748 40228 24772 40230
rect 24828 40228 24852 40230
rect 24908 40228 24932 40230
rect 24988 40228 24994 40230
rect 24686 40219 24994 40228
rect 24582 39400 24638 39409
rect 24582 39335 24638 39344
rect 24492 34196 24544 34202
rect 24492 34138 24544 34144
rect 24400 33312 24452 33318
rect 24400 33254 24452 33260
rect 24412 33153 24440 33254
rect 24398 33144 24454 33153
rect 24398 33079 24454 33088
rect 24400 32224 24452 32230
rect 24400 32166 24452 32172
rect 24412 31929 24440 32166
rect 24492 31952 24544 31958
rect 24398 31920 24454 31929
rect 24492 31894 24544 31900
rect 24398 31855 24454 31864
rect 24400 31136 24452 31142
rect 24400 31078 24452 31084
rect 24412 30841 24440 31078
rect 24398 30832 24454 30841
rect 24398 30767 24454 30776
rect 24400 30048 24452 30054
rect 24400 29990 24452 29996
rect 24412 29753 24440 29990
rect 24398 29744 24454 29753
rect 24398 29679 24454 29688
rect 24400 29028 24452 29034
rect 24400 28970 24452 28976
rect 24412 28937 24440 28970
rect 24398 28928 24454 28937
rect 24398 28863 24454 28872
rect 24400 27872 24452 27878
rect 24400 27814 24452 27820
rect 24412 27577 24440 27814
rect 24398 27568 24454 27577
rect 24398 27503 24454 27512
rect 24400 25696 24452 25702
rect 24400 25638 24452 25644
rect 24412 25401 24440 25638
rect 24398 25392 24454 25401
rect 24398 25327 24454 25336
rect 24400 24608 24452 24614
rect 24400 24550 24452 24556
rect 24412 24313 24440 24550
rect 24398 24304 24454 24313
rect 24398 24239 24454 24248
rect 24400 23520 24452 23526
rect 24398 23488 24400 23497
rect 24452 23488 24454 23497
rect 24398 23423 24454 23432
rect 24400 22432 24452 22438
rect 24400 22374 24452 22380
rect 24412 22137 24440 22374
rect 24398 22128 24454 22137
rect 24398 22063 24454 22072
rect 24504 21554 24532 31894
rect 24492 21548 24544 21554
rect 24492 21490 24544 21496
rect 24124 21412 24176 21418
rect 24320 21406 24532 21434
rect 24124 21354 24176 21360
rect 24032 19440 24084 19446
rect 24032 19382 24084 19388
rect 24136 18766 24164 21354
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24228 21146 24256 21286
rect 24306 21176 24362 21185
rect 24216 21140 24268 21146
rect 24306 21111 24362 21120
rect 24216 21082 24268 21088
rect 24216 19780 24268 19786
rect 24216 19722 24268 19728
rect 24228 19417 24256 19722
rect 24214 19408 24270 19417
rect 24214 19343 24270 19352
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 24124 18624 24176 18630
rect 24124 18566 24176 18572
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 23940 18080 23992 18086
rect 23940 18022 23992 18028
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 23952 17134 23980 18022
rect 24044 17241 24072 18022
rect 24136 17921 24164 18566
rect 24228 18290 24256 18566
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 24122 17912 24178 17921
rect 24122 17847 24178 17856
rect 24030 17232 24086 17241
rect 24030 17167 24086 17176
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23952 16561 23980 16594
rect 23938 16552 23994 16561
rect 23938 16487 23994 16496
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 24216 16040 24268 16046
rect 24216 15982 24268 15988
rect 23756 15904 23808 15910
rect 23756 15846 23808 15852
rect 23768 15609 23796 15846
rect 23754 15600 23810 15609
rect 23754 15535 23810 15544
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 23112 15496 23164 15502
rect 23112 15438 23164 15444
rect 23204 15496 23256 15502
rect 23204 15438 23256 15444
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23032 15094 23060 15438
rect 23124 15162 23152 15438
rect 23664 15428 23716 15434
rect 23664 15370 23716 15376
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 22928 15088 22980 15094
rect 22928 15030 22980 15036
rect 23020 15088 23072 15094
rect 23020 15030 23072 15036
rect 22940 14940 22968 15030
rect 23400 14940 23428 15302
rect 23492 15094 23520 15302
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23480 15088 23532 15094
rect 23480 15030 23532 15036
rect 22940 14912 23060 14940
rect 23400 14912 23520 14940
rect 23032 14006 23060 14912
rect 23112 14340 23164 14346
rect 23112 14282 23164 14288
rect 23020 14000 23072 14006
rect 23020 13942 23072 13948
rect 22928 13728 22980 13734
rect 22928 13670 22980 13676
rect 22940 13462 22968 13670
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 22652 12378 22704 12384
rect 22756 12406 22876 12434
rect 22664 12345 22692 12378
rect 22650 12336 22706 12345
rect 22650 12271 22706 12280
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22664 11694 22692 12174
rect 22652 11688 22704 11694
rect 22652 11630 22704 11636
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22664 10266 22692 10610
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22756 10146 22784 12406
rect 22928 12164 22980 12170
rect 22928 12106 22980 12112
rect 22834 11792 22890 11801
rect 22834 11727 22836 11736
rect 22888 11727 22890 11736
rect 22836 11698 22888 11704
rect 22940 11150 22968 12106
rect 23032 11150 23060 13942
rect 23124 13190 23152 14282
rect 23204 14272 23256 14278
rect 23204 14214 23256 14220
rect 23216 13530 23244 14214
rect 23492 14074 23520 14912
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23584 13938 23612 15098
rect 23676 13938 23704 15370
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 24136 15201 24164 15302
rect 24122 15192 24178 15201
rect 24122 15127 24178 15136
rect 23296 13932 23348 13938
rect 23296 13874 23348 13880
rect 23572 13932 23624 13938
rect 23572 13874 23624 13880
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23308 13326 23336 13874
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 24032 13252 24084 13258
rect 24032 13194 24084 13200
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22848 10266 22876 10406
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 22756 10118 22876 10146
rect 22560 7880 22612 7886
rect 22560 7822 22612 7828
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22468 6996 22520 7002
rect 22468 6938 22520 6944
rect 22572 6769 22600 7686
rect 22744 7404 22796 7410
rect 22744 7346 22796 7352
rect 22756 7002 22784 7346
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 22744 6792 22796 6798
rect 22558 6760 22614 6769
rect 22744 6734 22796 6740
rect 22558 6695 22614 6704
rect 22650 6216 22706 6225
rect 22650 6151 22652 6160
rect 22704 6151 22706 6160
rect 22652 6122 22704 6128
rect 22558 5808 22614 5817
rect 22558 5743 22614 5752
rect 22572 5710 22600 5743
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 22756 5574 22784 6734
rect 22744 5568 22796 5574
rect 22558 5536 22614 5545
rect 22744 5510 22796 5516
rect 22558 5471 22614 5480
rect 22572 5370 22600 5471
rect 22560 5364 22612 5370
rect 22560 5306 22612 5312
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22296 4032 22416 4060
rect 22284 3936 22336 3942
rect 22020 3896 22232 3924
rect 21719 3836 22027 3845
rect 21719 3834 21725 3836
rect 21781 3834 21805 3836
rect 21861 3834 21885 3836
rect 21941 3834 21965 3836
rect 22021 3834 22027 3836
rect 21781 3782 21783 3834
rect 21963 3782 21965 3834
rect 21719 3780 21725 3782
rect 21781 3780 21805 3782
rect 21861 3780 21885 3782
rect 21941 3780 21965 3782
rect 22021 3780 22027 3782
rect 21719 3771 22027 3780
rect 21640 3528 21692 3534
rect 22100 3528 22152 3534
rect 21640 3470 21692 3476
rect 22098 3496 22100 3505
rect 22152 3496 22154 3505
rect 22098 3431 22154 3440
rect 21640 3052 21692 3058
rect 21640 2994 21692 3000
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 21376 2094 21588 2122
rect 21364 1964 21416 1970
rect 21364 1906 21416 1912
rect 21272 1488 21324 1494
rect 21272 1430 21324 1436
rect 21272 1284 21324 1290
rect 21272 1226 21324 1232
rect 21284 1018 21312 1226
rect 21272 1012 21324 1018
rect 21272 954 21324 960
rect 21086 912 21142 921
rect 21086 847 21142 856
rect 21272 672 21324 678
rect 21192 632 21272 660
rect 21192 160 21220 632
rect 21272 614 21324 620
rect 20902 82 20958 160
rect 20824 54 20958 82
rect 20902 0 20958 54
rect 21178 0 21234 160
rect 21376 82 21404 1906
rect 21454 82 21510 160
rect 21376 54 21510 82
rect 21560 82 21588 2094
rect 21652 1442 21680 2994
rect 21719 2748 22027 2757
rect 21719 2746 21725 2748
rect 21781 2746 21805 2748
rect 21861 2746 21885 2748
rect 21941 2746 21965 2748
rect 22021 2746 22027 2748
rect 21781 2694 21783 2746
rect 21963 2694 21965 2746
rect 21719 2692 21725 2694
rect 21781 2692 21805 2694
rect 21861 2692 21885 2694
rect 21941 2692 21965 2694
rect 22021 2692 22027 2694
rect 21719 2683 22027 2692
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 21928 2553 21956 2586
rect 21914 2544 21970 2553
rect 21914 2479 21970 2488
rect 21732 2372 21784 2378
rect 21732 2314 21784 2320
rect 21744 2106 21772 2314
rect 21732 2100 21784 2106
rect 21732 2042 21784 2048
rect 21719 1660 22027 1669
rect 21719 1658 21725 1660
rect 21781 1658 21805 1660
rect 21861 1658 21885 1660
rect 21941 1658 21965 1660
rect 22021 1658 22027 1660
rect 21781 1606 21783 1658
rect 21963 1606 21965 1658
rect 21719 1604 21725 1606
rect 21781 1604 21805 1606
rect 21861 1604 21885 1606
rect 21941 1604 21965 1606
rect 22021 1604 22027 1606
rect 21719 1595 22027 1604
rect 21652 1414 22048 1442
rect 22020 160 22048 1414
rect 22204 1290 22232 3896
rect 22284 3878 22336 3884
rect 22296 3602 22324 3878
rect 22284 3596 22336 3602
rect 22284 3538 22336 3544
rect 22388 3097 22416 4032
rect 22480 3738 22508 5170
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22652 4616 22704 4622
rect 22756 4593 22784 5510
rect 22652 4558 22704 4564
rect 22742 4584 22798 4593
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 22374 3088 22430 3097
rect 22284 3052 22336 3058
rect 22374 3023 22430 3032
rect 22284 2994 22336 3000
rect 22192 1284 22244 1290
rect 22192 1226 22244 1232
rect 22296 160 22324 2994
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 22480 2514 22508 2926
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22572 1465 22600 4558
rect 22664 3670 22692 4558
rect 22742 4519 22798 4528
rect 22652 3664 22704 3670
rect 22652 3606 22704 3612
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 22558 1456 22614 1465
rect 22558 1391 22614 1400
rect 22468 1284 22520 1290
rect 22468 1226 22520 1232
rect 22480 678 22508 1226
rect 22468 672 22520 678
rect 22468 614 22520 620
rect 21730 82 21786 160
rect 21560 54 21786 82
rect 21454 0 21510 54
rect 21730 0 21786 54
rect 22006 0 22062 160
rect 22282 0 22338 160
rect 22558 82 22614 160
rect 22664 82 22692 3470
rect 22848 3126 22876 10118
rect 22940 9994 22968 11086
rect 22928 9988 22980 9994
rect 22928 9930 22980 9936
rect 22940 6202 22968 9930
rect 23124 9722 23152 13126
rect 24044 12889 24072 13194
rect 24030 12880 24086 12889
rect 23480 12844 23532 12850
rect 24030 12815 24086 12824
rect 23480 12786 23532 12792
rect 23492 11762 23520 12786
rect 23848 12640 23900 12646
rect 23848 12582 23900 12588
rect 23860 12345 23888 12582
rect 23846 12336 23902 12345
rect 23846 12271 23902 12280
rect 23848 12096 23900 12102
rect 23848 12038 23900 12044
rect 23860 11898 23888 12038
rect 23756 11892 23808 11898
rect 23756 11834 23808 11840
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23492 10742 23520 11494
rect 23676 11354 23704 11494
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23676 10742 23704 10950
rect 23480 10736 23532 10742
rect 23480 10678 23532 10684
rect 23664 10736 23716 10742
rect 23664 10678 23716 10684
rect 23204 10668 23256 10674
rect 23204 10610 23256 10616
rect 23216 9722 23244 10610
rect 23112 9716 23164 9722
rect 23112 9658 23164 9664
rect 23204 9716 23256 9722
rect 23204 9658 23256 9664
rect 23768 9654 23796 11834
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23860 10169 23888 10406
rect 23846 10160 23902 10169
rect 23846 10095 23902 10104
rect 24124 9920 24176 9926
rect 24124 9862 24176 9868
rect 23756 9648 23808 9654
rect 23756 9590 23808 9596
rect 23938 9616 23994 9625
rect 23572 9580 23624 9586
rect 23938 9551 23940 9560
rect 23572 9522 23624 9528
rect 23992 9551 23994 9560
rect 23940 9522 23992 9528
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 23020 7200 23072 7206
rect 23020 7142 23072 7148
rect 23032 6458 23060 7142
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23032 6322 23060 6394
rect 23020 6316 23072 6322
rect 23020 6258 23072 6264
rect 23124 6236 23152 9318
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 23216 8498 23244 8774
rect 23204 8492 23256 8498
rect 23204 8434 23256 8440
rect 23308 8090 23336 8910
rect 23492 8634 23520 8910
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 23584 8090 23612 9522
rect 23846 9072 23902 9081
rect 23846 9007 23902 9016
rect 23664 8560 23716 8566
rect 23664 8502 23716 8508
rect 23296 8084 23348 8090
rect 23296 8026 23348 8032
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23492 7562 23520 8026
rect 23492 7534 23612 7562
rect 23676 7546 23704 8502
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 23584 7410 23612 7534
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23768 7410 23796 8434
rect 23860 7886 23888 9007
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 23940 8900 23992 8906
rect 23940 8842 23992 8848
rect 23952 8537 23980 8842
rect 23938 8528 23994 8537
rect 23938 8463 23994 8472
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 24044 7546 24072 8910
rect 24136 7886 24164 9862
rect 24228 9722 24256 15982
rect 24216 9716 24268 9722
rect 24216 9658 24268 9664
rect 24216 9580 24268 9586
rect 24216 9522 24268 9528
rect 24228 8022 24256 9522
rect 24216 8016 24268 8022
rect 24216 7958 24268 7964
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 24216 7812 24268 7818
rect 24216 7754 24268 7760
rect 24228 7546 24256 7754
rect 24032 7540 24084 7546
rect 24032 7482 24084 7488
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24214 7440 24270 7449
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 23756 7404 23808 7410
rect 24214 7375 24216 7384
rect 23756 7346 23808 7352
rect 24268 7375 24270 7384
rect 24216 7346 24268 7352
rect 23216 6361 23244 7346
rect 23492 6905 23520 7346
rect 24214 7304 24270 7313
rect 24214 7239 24270 7248
rect 23478 6896 23534 6905
rect 23478 6831 23534 6840
rect 23572 6792 23624 6798
rect 23386 6760 23442 6769
rect 23572 6734 23624 6740
rect 23386 6695 23442 6704
rect 23202 6352 23258 6361
rect 23202 6287 23258 6296
rect 23124 6208 23244 6236
rect 22940 6174 23060 6202
rect 22928 5636 22980 5642
rect 22928 5578 22980 5584
rect 22940 5234 22968 5578
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 22928 5024 22980 5030
rect 22928 4966 22980 4972
rect 22940 4690 22968 4966
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 23032 3602 23060 6174
rect 23112 5228 23164 5234
rect 23112 5170 23164 5176
rect 23124 3641 23152 5170
rect 23216 4690 23244 6208
rect 23400 5817 23428 6695
rect 23386 5808 23442 5817
rect 23442 5766 23520 5794
rect 23386 5743 23442 5752
rect 23492 5284 23520 5766
rect 23584 5409 23612 6734
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23570 5400 23626 5409
rect 23570 5335 23626 5344
rect 23664 5364 23716 5370
rect 23664 5306 23716 5312
rect 23492 5256 23612 5284
rect 23478 5128 23534 5137
rect 23388 5092 23440 5098
rect 23478 5063 23480 5072
rect 23388 5034 23440 5040
rect 23532 5063 23534 5072
rect 23480 5034 23532 5040
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 23110 3632 23166 3641
rect 23020 3596 23072 3602
rect 23110 3567 23166 3576
rect 23020 3538 23072 3544
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 22744 3120 22796 3126
rect 22744 3062 22796 3068
rect 22836 3120 22888 3126
rect 22836 3062 22888 3068
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 22756 1834 22784 3062
rect 22744 1828 22796 1834
rect 22744 1770 22796 1776
rect 23032 1358 23060 3062
rect 23020 1352 23072 1358
rect 23020 1294 23072 1300
rect 22836 944 22888 950
rect 22836 886 22888 892
rect 22848 160 22876 886
rect 23124 160 23152 3470
rect 23400 160 23428 5034
rect 23584 3670 23612 5256
rect 23676 4706 23704 5306
rect 23768 5302 23796 6054
rect 24228 5914 24256 7239
rect 24216 5908 24268 5914
rect 24216 5850 24268 5856
rect 23940 5704 23992 5710
rect 23846 5672 23902 5681
rect 23940 5646 23992 5652
rect 23846 5607 23902 5616
rect 23756 5296 23808 5302
rect 23756 5238 23808 5244
rect 23860 5114 23888 5607
rect 23768 5086 23888 5114
rect 23768 4842 23796 5086
rect 23952 5001 23980 5646
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 23938 4992 23994 5001
rect 23938 4927 23994 4936
rect 23768 4814 23980 4842
rect 23676 4678 23796 4706
rect 23664 4548 23716 4554
rect 23664 4490 23716 4496
rect 23572 3664 23624 3670
rect 23572 3606 23624 3612
rect 23480 2372 23532 2378
rect 23480 2314 23532 2320
rect 23492 2106 23520 2314
rect 23480 2100 23532 2106
rect 23480 2042 23532 2048
rect 23676 160 23704 4490
rect 23768 2774 23796 4678
rect 23768 2746 23888 2774
rect 23860 2446 23888 2746
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 23768 1272 23796 2382
rect 23952 2106 23980 4814
rect 24044 2553 24072 5170
rect 24216 5160 24268 5166
rect 24216 5102 24268 5108
rect 24124 5024 24176 5030
rect 24124 4966 24176 4972
rect 24136 3126 24164 4966
rect 24228 4078 24256 5102
rect 24216 4072 24268 4078
rect 24216 4014 24268 4020
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 24216 2848 24268 2854
rect 24216 2790 24268 2796
rect 24030 2544 24086 2553
rect 24030 2479 24086 2488
rect 23940 2100 23992 2106
rect 23940 2042 23992 2048
rect 23768 1244 23980 1272
rect 23952 160 23980 1244
rect 24228 160 24256 2790
rect 24320 1970 24348 21111
rect 24398 21040 24454 21049
rect 24398 20975 24454 20984
rect 24412 20602 24440 20975
rect 24400 20596 24452 20602
rect 24400 20538 24452 20544
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24412 18873 24440 19110
rect 24398 18864 24454 18873
rect 24398 18799 24454 18808
rect 24400 18420 24452 18426
rect 24400 18362 24452 18368
rect 24412 18329 24440 18362
rect 24398 18320 24454 18329
rect 24398 18255 24454 18264
rect 24398 16688 24454 16697
rect 24398 16623 24454 16632
rect 24412 16250 24440 16623
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24412 14521 24440 14758
rect 24398 14512 24454 14521
rect 24398 14447 24454 14456
rect 24504 14362 24532 21406
rect 24412 14334 24532 14362
rect 24412 12434 24440 14334
rect 24490 13968 24546 13977
rect 24490 13903 24546 13912
rect 24504 12986 24532 13903
rect 24492 12980 24544 12986
rect 24492 12922 24544 12928
rect 24412 12406 24532 12434
rect 24400 11892 24452 11898
rect 24400 11834 24452 11840
rect 24412 11801 24440 11834
rect 24398 11792 24454 11801
rect 24398 11727 24454 11736
rect 24504 11642 24532 12406
rect 24412 11614 24532 11642
rect 24412 5370 24440 11614
rect 24490 10704 24546 10713
rect 24490 10639 24492 10648
rect 24544 10639 24546 10648
rect 24492 10610 24544 10616
rect 24490 8936 24546 8945
rect 24490 8871 24546 8880
rect 24504 6934 24532 8871
rect 24492 6928 24544 6934
rect 24492 6870 24544 6876
rect 24400 5364 24452 5370
rect 24400 5306 24452 5312
rect 24400 4276 24452 4282
rect 24400 4218 24452 4224
rect 24308 1964 24360 1970
rect 24308 1906 24360 1912
rect 22558 54 22692 82
rect 22558 0 22614 54
rect 22834 0 22890 160
rect 23110 0 23166 160
rect 23386 0 23442 160
rect 23662 0 23718 160
rect 23938 0 23994 160
rect 24214 0 24270 160
rect 24412 82 24440 4218
rect 24492 2848 24544 2854
rect 24492 2790 24544 2796
rect 24504 2106 24532 2790
rect 24596 2650 24624 39335
rect 24686 39196 24994 39205
rect 24686 39194 24692 39196
rect 24748 39194 24772 39196
rect 24828 39194 24852 39196
rect 24908 39194 24932 39196
rect 24988 39194 24994 39196
rect 24748 39142 24750 39194
rect 24930 39142 24932 39194
rect 24686 39140 24692 39142
rect 24748 39140 24772 39142
rect 24828 39140 24852 39142
rect 24908 39140 24932 39142
rect 24988 39140 24994 39142
rect 24686 39131 24994 39140
rect 25228 39024 25280 39030
rect 25228 38966 25280 38972
rect 24686 38108 24994 38117
rect 24686 38106 24692 38108
rect 24748 38106 24772 38108
rect 24828 38106 24852 38108
rect 24908 38106 24932 38108
rect 24988 38106 24994 38108
rect 24748 38054 24750 38106
rect 24930 38054 24932 38106
rect 24686 38052 24692 38054
rect 24748 38052 24772 38054
rect 24828 38052 24852 38054
rect 24908 38052 24932 38054
rect 24988 38052 24994 38054
rect 24686 38043 24994 38052
rect 24686 37020 24994 37029
rect 24686 37018 24692 37020
rect 24748 37018 24772 37020
rect 24828 37018 24852 37020
rect 24908 37018 24932 37020
rect 24988 37018 24994 37020
rect 24748 36966 24750 37018
rect 24930 36966 24932 37018
rect 24686 36964 24692 36966
rect 24748 36964 24772 36966
rect 24828 36964 24852 36966
rect 24908 36964 24932 36966
rect 24988 36964 24994 36966
rect 24686 36955 24994 36964
rect 24686 35932 24994 35941
rect 24686 35930 24692 35932
rect 24748 35930 24772 35932
rect 24828 35930 24852 35932
rect 24908 35930 24932 35932
rect 24988 35930 24994 35932
rect 24748 35878 24750 35930
rect 24930 35878 24932 35930
rect 24686 35876 24692 35878
rect 24748 35876 24772 35878
rect 24828 35876 24852 35878
rect 24908 35876 24932 35878
rect 24988 35876 24994 35878
rect 24686 35867 24994 35876
rect 24686 34844 24994 34853
rect 24686 34842 24692 34844
rect 24748 34842 24772 34844
rect 24828 34842 24852 34844
rect 24908 34842 24932 34844
rect 24988 34842 24994 34844
rect 24748 34790 24750 34842
rect 24930 34790 24932 34842
rect 24686 34788 24692 34790
rect 24748 34788 24772 34790
rect 24828 34788 24852 34790
rect 24908 34788 24932 34790
rect 24988 34788 24994 34790
rect 24686 34779 24994 34788
rect 24686 33756 24994 33765
rect 24686 33754 24692 33756
rect 24748 33754 24772 33756
rect 24828 33754 24852 33756
rect 24908 33754 24932 33756
rect 24988 33754 24994 33756
rect 24748 33702 24750 33754
rect 24930 33702 24932 33754
rect 24686 33700 24692 33702
rect 24748 33700 24772 33702
rect 24828 33700 24852 33702
rect 24908 33700 24932 33702
rect 24988 33700 24994 33702
rect 24686 33691 24994 33700
rect 24686 32668 24994 32677
rect 24686 32666 24692 32668
rect 24748 32666 24772 32668
rect 24828 32666 24852 32668
rect 24908 32666 24932 32668
rect 24988 32666 24994 32668
rect 24748 32614 24750 32666
rect 24930 32614 24932 32666
rect 24686 32612 24692 32614
rect 24748 32612 24772 32614
rect 24828 32612 24852 32614
rect 24908 32612 24932 32614
rect 24988 32612 24994 32614
rect 24686 32603 24994 32612
rect 24686 31580 24994 31589
rect 24686 31578 24692 31580
rect 24748 31578 24772 31580
rect 24828 31578 24852 31580
rect 24908 31578 24932 31580
rect 24988 31578 24994 31580
rect 24748 31526 24750 31578
rect 24930 31526 24932 31578
rect 24686 31524 24692 31526
rect 24748 31524 24772 31526
rect 24828 31524 24852 31526
rect 24908 31524 24932 31526
rect 24988 31524 24994 31526
rect 24686 31515 24994 31524
rect 25044 31340 25096 31346
rect 25044 31282 25096 31288
rect 24686 30492 24994 30501
rect 24686 30490 24692 30492
rect 24748 30490 24772 30492
rect 24828 30490 24852 30492
rect 24908 30490 24932 30492
rect 24988 30490 24994 30492
rect 24748 30438 24750 30490
rect 24930 30438 24932 30490
rect 24686 30436 24692 30438
rect 24748 30436 24772 30438
rect 24828 30436 24852 30438
rect 24908 30436 24932 30438
rect 24988 30436 24994 30438
rect 24686 30427 24994 30436
rect 24686 29404 24994 29413
rect 24686 29402 24692 29404
rect 24748 29402 24772 29404
rect 24828 29402 24852 29404
rect 24908 29402 24932 29404
rect 24988 29402 24994 29404
rect 24748 29350 24750 29402
rect 24930 29350 24932 29402
rect 24686 29348 24692 29350
rect 24748 29348 24772 29350
rect 24828 29348 24852 29350
rect 24908 29348 24932 29350
rect 24988 29348 24994 29350
rect 24686 29339 24994 29348
rect 24686 28316 24994 28325
rect 24686 28314 24692 28316
rect 24748 28314 24772 28316
rect 24828 28314 24852 28316
rect 24908 28314 24932 28316
rect 24988 28314 24994 28316
rect 24748 28262 24750 28314
rect 24930 28262 24932 28314
rect 24686 28260 24692 28262
rect 24748 28260 24772 28262
rect 24828 28260 24852 28262
rect 24908 28260 24932 28262
rect 24988 28260 24994 28262
rect 24686 28251 24994 28260
rect 24686 27228 24994 27237
rect 24686 27226 24692 27228
rect 24748 27226 24772 27228
rect 24828 27226 24852 27228
rect 24908 27226 24932 27228
rect 24988 27226 24994 27228
rect 24748 27174 24750 27226
rect 24930 27174 24932 27226
rect 24686 27172 24692 27174
rect 24748 27172 24772 27174
rect 24828 27172 24852 27174
rect 24908 27172 24932 27174
rect 24988 27172 24994 27174
rect 24686 27163 24994 27172
rect 24686 26140 24994 26149
rect 24686 26138 24692 26140
rect 24748 26138 24772 26140
rect 24828 26138 24852 26140
rect 24908 26138 24932 26140
rect 24988 26138 24994 26140
rect 24748 26086 24750 26138
rect 24930 26086 24932 26138
rect 24686 26084 24692 26086
rect 24748 26084 24772 26086
rect 24828 26084 24852 26086
rect 24908 26084 24932 26086
rect 24988 26084 24994 26086
rect 24686 26075 24994 26084
rect 24686 25052 24994 25061
rect 24686 25050 24692 25052
rect 24748 25050 24772 25052
rect 24828 25050 24852 25052
rect 24908 25050 24932 25052
rect 24988 25050 24994 25052
rect 24748 24998 24750 25050
rect 24930 24998 24932 25050
rect 24686 24996 24692 24998
rect 24748 24996 24772 24998
rect 24828 24996 24852 24998
rect 24908 24996 24932 24998
rect 24988 24996 24994 24998
rect 24686 24987 24994 24996
rect 24686 23964 24994 23973
rect 24686 23962 24692 23964
rect 24748 23962 24772 23964
rect 24828 23962 24852 23964
rect 24908 23962 24932 23964
rect 24988 23962 24994 23964
rect 24748 23910 24750 23962
rect 24930 23910 24932 23962
rect 24686 23908 24692 23910
rect 24748 23908 24772 23910
rect 24828 23908 24852 23910
rect 24908 23908 24932 23910
rect 24988 23908 24994 23910
rect 24686 23899 24994 23908
rect 24686 22876 24994 22885
rect 24686 22874 24692 22876
rect 24748 22874 24772 22876
rect 24828 22874 24852 22876
rect 24908 22874 24932 22876
rect 24988 22874 24994 22876
rect 24748 22822 24750 22874
rect 24930 22822 24932 22874
rect 24686 22820 24692 22822
rect 24748 22820 24772 22822
rect 24828 22820 24852 22822
rect 24908 22820 24932 22822
rect 24988 22820 24994 22822
rect 24686 22811 24994 22820
rect 24686 21788 24994 21797
rect 24686 21786 24692 21788
rect 24748 21786 24772 21788
rect 24828 21786 24852 21788
rect 24908 21786 24932 21788
rect 24988 21786 24994 21788
rect 24748 21734 24750 21786
rect 24930 21734 24932 21786
rect 24686 21732 24692 21734
rect 24748 21732 24772 21734
rect 24828 21732 24852 21734
rect 24908 21732 24932 21734
rect 24988 21732 24994 21734
rect 24686 21723 24994 21732
rect 24686 20700 24994 20709
rect 24686 20698 24692 20700
rect 24748 20698 24772 20700
rect 24828 20698 24852 20700
rect 24908 20698 24932 20700
rect 24988 20698 24994 20700
rect 24748 20646 24750 20698
rect 24930 20646 24932 20698
rect 24686 20644 24692 20646
rect 24748 20644 24772 20646
rect 24828 20644 24852 20646
rect 24908 20644 24932 20646
rect 24988 20644 24994 20646
rect 24686 20635 24994 20644
rect 24686 19612 24994 19621
rect 24686 19610 24692 19612
rect 24748 19610 24772 19612
rect 24828 19610 24852 19612
rect 24908 19610 24932 19612
rect 24988 19610 24994 19612
rect 24748 19558 24750 19610
rect 24930 19558 24932 19610
rect 24686 19556 24692 19558
rect 24748 19556 24772 19558
rect 24828 19556 24852 19558
rect 24908 19556 24932 19558
rect 24988 19556 24994 19558
rect 24686 19547 24994 19556
rect 24686 18524 24994 18533
rect 24686 18522 24692 18524
rect 24748 18522 24772 18524
rect 24828 18522 24852 18524
rect 24908 18522 24932 18524
rect 24988 18522 24994 18524
rect 24748 18470 24750 18522
rect 24930 18470 24932 18522
rect 24686 18468 24692 18470
rect 24748 18468 24772 18470
rect 24828 18468 24852 18470
rect 24908 18468 24932 18470
rect 24988 18468 24994 18470
rect 24686 18459 24994 18468
rect 24686 17436 24994 17445
rect 24686 17434 24692 17436
rect 24748 17434 24772 17436
rect 24828 17434 24852 17436
rect 24908 17434 24932 17436
rect 24988 17434 24994 17436
rect 24748 17382 24750 17434
rect 24930 17382 24932 17434
rect 24686 17380 24692 17382
rect 24748 17380 24772 17382
rect 24828 17380 24852 17382
rect 24908 17380 24932 17382
rect 24988 17380 24994 17382
rect 24686 17371 24994 17380
rect 25056 17134 25084 31282
rect 25136 27396 25188 27402
rect 25136 27338 25188 27344
rect 25148 25945 25176 27338
rect 25134 25936 25190 25945
rect 25134 25871 25190 25880
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 25044 17128 25096 17134
rect 25044 17070 25096 17076
rect 24686 16348 24994 16357
rect 24686 16346 24692 16348
rect 24748 16346 24772 16348
rect 24828 16346 24852 16348
rect 24908 16346 24932 16348
rect 24988 16346 24994 16348
rect 24748 16294 24750 16346
rect 24930 16294 24932 16346
rect 24686 16292 24692 16294
rect 24748 16292 24772 16294
rect 24828 16292 24852 16294
rect 24908 16292 24932 16294
rect 24988 16292 24994 16294
rect 24686 16283 24994 16292
rect 24686 15260 24994 15269
rect 24686 15258 24692 15260
rect 24748 15258 24772 15260
rect 24828 15258 24852 15260
rect 24908 15258 24932 15260
rect 24988 15258 24994 15260
rect 24748 15206 24750 15258
rect 24930 15206 24932 15258
rect 24686 15204 24692 15206
rect 24748 15204 24772 15206
rect 24828 15204 24852 15206
rect 24908 15204 24932 15206
rect 24988 15204 24994 15206
rect 24686 15195 24994 15204
rect 24686 14172 24994 14181
rect 24686 14170 24692 14172
rect 24748 14170 24772 14172
rect 24828 14170 24852 14172
rect 24908 14170 24932 14172
rect 24988 14170 24994 14172
rect 24748 14118 24750 14170
rect 24930 14118 24932 14170
rect 24686 14116 24692 14118
rect 24748 14116 24772 14118
rect 24828 14116 24852 14118
rect 24908 14116 24932 14118
rect 24988 14116 24994 14118
rect 24686 14107 24994 14116
rect 24676 13456 24728 13462
rect 24674 13424 24676 13433
rect 24728 13424 24730 13433
rect 24674 13359 24730 13368
rect 24686 13084 24994 13093
rect 24686 13082 24692 13084
rect 24748 13082 24772 13084
rect 24828 13082 24852 13084
rect 24908 13082 24932 13084
rect 24988 13082 24994 13084
rect 24748 13030 24750 13082
rect 24930 13030 24932 13082
rect 24686 13028 24692 13030
rect 24748 13028 24772 13030
rect 24828 13028 24852 13030
rect 24908 13028 24932 13030
rect 24988 13028 24994 13030
rect 24686 13019 24994 13028
rect 24686 11996 24994 12005
rect 24686 11994 24692 11996
rect 24748 11994 24772 11996
rect 24828 11994 24852 11996
rect 24908 11994 24932 11996
rect 24988 11994 24994 11996
rect 24748 11942 24750 11994
rect 24930 11942 24932 11994
rect 24686 11940 24692 11942
rect 24748 11940 24772 11942
rect 24828 11940 24852 11942
rect 24908 11940 24932 11942
rect 24988 11940 24994 11942
rect 24686 11931 24994 11940
rect 25042 11248 25098 11257
rect 25042 11183 25098 11192
rect 24686 10908 24994 10917
rect 24686 10906 24692 10908
rect 24748 10906 24772 10908
rect 24828 10906 24852 10908
rect 24908 10906 24932 10908
rect 24988 10906 24994 10908
rect 24748 10854 24750 10906
rect 24930 10854 24932 10906
rect 24686 10852 24692 10854
rect 24748 10852 24772 10854
rect 24828 10852 24852 10854
rect 24908 10852 24932 10854
rect 24988 10852 24994 10854
rect 24686 10843 24994 10852
rect 24686 9820 24994 9829
rect 24686 9818 24692 9820
rect 24748 9818 24772 9820
rect 24828 9818 24852 9820
rect 24908 9818 24932 9820
rect 24988 9818 24994 9820
rect 24748 9766 24750 9818
rect 24930 9766 24932 9818
rect 24686 9764 24692 9766
rect 24748 9764 24772 9766
rect 24828 9764 24852 9766
rect 24908 9764 24932 9766
rect 24988 9764 24994 9766
rect 24686 9755 24994 9764
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24964 9466 24992 9658
rect 25056 9654 25084 11183
rect 25044 9648 25096 9654
rect 25044 9590 25096 9596
rect 24964 9438 25084 9466
rect 24686 8732 24994 8741
rect 24686 8730 24692 8732
rect 24748 8730 24772 8732
rect 24828 8730 24852 8732
rect 24908 8730 24932 8732
rect 24988 8730 24994 8732
rect 24748 8678 24750 8730
rect 24930 8678 24932 8730
rect 24686 8676 24692 8678
rect 24748 8676 24772 8678
rect 24828 8676 24852 8678
rect 24908 8676 24932 8678
rect 24988 8676 24994 8678
rect 24686 8667 24994 8676
rect 24686 7644 24994 7653
rect 24686 7642 24692 7644
rect 24748 7642 24772 7644
rect 24828 7642 24852 7644
rect 24908 7642 24932 7644
rect 24988 7642 24994 7644
rect 24748 7590 24750 7642
rect 24930 7590 24932 7642
rect 24686 7588 24692 7590
rect 24748 7588 24772 7590
rect 24828 7588 24852 7590
rect 24908 7588 24932 7590
rect 24988 7588 24994 7590
rect 24686 7579 24994 7588
rect 25056 7460 25084 9438
rect 25148 7562 25176 25774
rect 25240 8106 25268 38966
rect 25412 36100 25464 36106
rect 25412 36042 25464 36048
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25332 25838 25360 29582
rect 25320 25832 25372 25838
rect 25320 25774 25372 25780
rect 25320 21548 25372 21554
rect 25320 21490 25372 21496
rect 25332 12850 25360 21490
rect 25424 17354 25452 36042
rect 25688 35556 25740 35562
rect 25688 35498 25740 35504
rect 25596 34468 25648 34474
rect 25596 34410 25648 34416
rect 25504 34400 25556 34406
rect 25504 34342 25556 34348
rect 25516 17474 25544 34342
rect 25608 17626 25636 34410
rect 25700 22030 25728 35498
rect 25792 24410 25820 41386
rect 25872 25492 25924 25498
rect 25872 25434 25924 25440
rect 25780 24404 25832 24410
rect 25780 24346 25832 24352
rect 25688 22024 25740 22030
rect 25688 21966 25740 21972
rect 25884 20466 25912 25434
rect 25872 20460 25924 20466
rect 25872 20402 25924 20408
rect 25778 20224 25834 20233
rect 25778 20159 25834 20168
rect 25608 17598 25728 17626
rect 25504 17468 25556 17474
rect 25504 17410 25556 17416
rect 25424 17326 25636 17354
rect 25504 17264 25556 17270
rect 25504 17206 25556 17212
rect 25412 17128 25464 17134
rect 25412 17070 25464 17076
rect 25320 12844 25372 12850
rect 25320 12786 25372 12792
rect 25320 12708 25372 12714
rect 25320 12650 25372 12656
rect 25332 8242 25360 12650
rect 25424 10538 25452 17070
rect 25412 10532 25464 10538
rect 25412 10474 25464 10480
rect 25516 9042 25544 17206
rect 25608 10606 25636 17326
rect 25700 13326 25728 17598
rect 25688 13320 25740 13326
rect 25688 13262 25740 13268
rect 25792 13138 25820 20159
rect 25872 19372 25924 19378
rect 25872 19314 25924 19320
rect 25700 13110 25820 13138
rect 25700 12714 25728 13110
rect 25688 12708 25740 12714
rect 25688 12650 25740 12656
rect 25688 12096 25740 12102
rect 25688 12038 25740 12044
rect 25596 10600 25648 10606
rect 25596 10542 25648 10548
rect 25504 9036 25556 9042
rect 25504 8978 25556 8984
rect 25332 8214 25544 8242
rect 25240 8078 25452 8106
rect 25318 7984 25374 7993
rect 25318 7919 25374 7928
rect 25148 7534 25268 7562
rect 25056 7432 25176 7460
rect 24686 6556 24994 6565
rect 24686 6554 24692 6556
rect 24748 6554 24772 6556
rect 24828 6554 24852 6556
rect 24908 6554 24932 6556
rect 24988 6554 24994 6556
rect 24748 6502 24750 6554
rect 24930 6502 24932 6554
rect 24686 6500 24692 6502
rect 24748 6500 24772 6502
rect 24828 6500 24852 6502
rect 24908 6500 24932 6502
rect 24988 6500 24994 6502
rect 24686 6491 24994 6500
rect 24686 5468 24994 5477
rect 24686 5466 24692 5468
rect 24748 5466 24772 5468
rect 24828 5466 24852 5468
rect 24908 5466 24932 5468
rect 24988 5466 24994 5468
rect 24748 5414 24750 5466
rect 24930 5414 24932 5466
rect 24686 5412 24692 5414
rect 24748 5412 24772 5414
rect 24828 5412 24852 5414
rect 24908 5412 24932 5414
rect 24988 5412 24994 5414
rect 24686 5403 24994 5412
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 24686 4380 24994 4389
rect 24686 4378 24692 4380
rect 24748 4378 24772 4380
rect 24828 4378 24852 4380
rect 24908 4378 24932 4380
rect 24988 4378 24994 4380
rect 24748 4326 24750 4378
rect 24930 4326 24932 4378
rect 24686 4324 24692 4326
rect 24748 4324 24772 4326
rect 24828 4324 24852 4326
rect 24908 4324 24932 4326
rect 24988 4324 24994 4326
rect 24686 4315 24994 4324
rect 24686 3292 24994 3301
rect 24686 3290 24692 3292
rect 24748 3290 24772 3292
rect 24828 3290 24852 3292
rect 24908 3290 24932 3292
rect 24988 3290 24994 3292
rect 24748 3238 24750 3290
rect 24930 3238 24932 3290
rect 24686 3236 24692 3238
rect 24748 3236 24772 3238
rect 24828 3236 24852 3238
rect 24908 3236 24932 3238
rect 24988 3236 24994 3238
rect 24686 3227 24994 3236
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 24686 2204 24994 2213
rect 24686 2202 24692 2204
rect 24748 2202 24772 2204
rect 24828 2202 24852 2204
rect 24908 2202 24932 2204
rect 24988 2202 24994 2204
rect 24748 2150 24750 2202
rect 24930 2150 24932 2202
rect 24686 2148 24692 2150
rect 24748 2148 24772 2150
rect 24828 2148 24852 2150
rect 24908 2148 24932 2150
rect 24988 2148 24994 2150
rect 24686 2139 24994 2148
rect 24492 2100 24544 2106
rect 24492 2042 24544 2048
rect 24492 1556 24544 1562
rect 24544 1516 24624 1544
rect 24492 1498 24544 1504
rect 24490 82 24546 160
rect 24412 54 24546 82
rect 24596 82 24624 1516
rect 24686 1116 24994 1125
rect 24686 1114 24692 1116
rect 24748 1114 24772 1116
rect 24828 1114 24852 1116
rect 24908 1114 24932 1116
rect 24988 1114 24994 1116
rect 24748 1062 24750 1114
rect 24930 1062 24932 1114
rect 24686 1060 24692 1062
rect 24748 1060 24772 1062
rect 24828 1060 24852 1062
rect 24908 1060 24932 1062
rect 24988 1060 24994 1062
rect 24686 1051 24994 1060
rect 25056 160 25084 5170
rect 25148 2378 25176 7432
rect 25240 2774 25268 7534
rect 25332 5710 25360 7919
rect 25320 5704 25372 5710
rect 25320 5646 25372 5652
rect 25424 4826 25452 8078
rect 25412 4820 25464 4826
rect 25412 4762 25464 4768
rect 25318 4040 25374 4049
rect 25516 4026 25544 8214
rect 25700 4146 25728 12038
rect 25884 5778 25912 19314
rect 25872 5772 25924 5778
rect 25872 5714 25924 5720
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25374 3998 25544 4026
rect 25318 3975 25374 3984
rect 25596 3732 25648 3738
rect 25596 3674 25648 3680
rect 25240 2746 25452 2774
rect 25136 2372 25188 2378
rect 25136 2314 25188 2320
rect 25320 1896 25372 1902
rect 25424 1873 25452 2746
rect 25320 1838 25372 1844
rect 25410 1864 25466 1873
rect 25332 160 25360 1838
rect 25410 1799 25466 1808
rect 25608 160 25636 3674
rect 24766 82 24822 160
rect 24596 54 24822 82
rect 24490 0 24546 54
rect 24766 0 24822 54
rect 25042 0 25098 160
rect 25318 0 25374 160
rect 25594 0 25650 160
<< via2 >>
rect 1030 41656 1086 41712
rect 662 40160 718 40216
rect 478 36080 534 36136
rect 478 26832 534 26888
rect 478 19760 534 19816
rect 18 1808 74 1864
rect 938 40024 994 40080
rect 754 28056 810 28112
rect 662 26016 718 26072
rect 938 25336 994 25392
rect 846 25064 902 25120
rect 662 22752 718 22808
rect 846 24656 902 24712
rect 938 23840 994 23896
rect 1398 39480 1454 39536
rect 1674 40996 1730 41032
rect 1674 40976 1676 40996
rect 1676 40976 1728 40996
rect 1728 40976 1730 40996
rect 1490 39072 1546 39128
rect 1398 38664 1454 38720
rect 1490 38392 1546 38448
rect 1306 38120 1362 38176
rect 1214 37576 1270 37632
rect 1674 38256 1730 38312
rect 2502 42220 2558 42256
rect 2502 42200 2504 42220
rect 2504 42200 2556 42220
rect 2556 42200 2558 42220
rect 2226 42100 2228 42120
rect 2228 42100 2280 42120
rect 2280 42100 2282 42120
rect 2226 42064 2282 42100
rect 2226 40568 2282 40624
rect 2042 40296 2098 40352
rect 1582 37032 1638 37088
rect 2594 40568 2650 40624
rect 2686 40432 2742 40488
rect 2410 39752 2466 39808
rect 2502 39480 2558 39536
rect 2318 39208 2374 39264
rect 1950 38664 2006 38720
rect 1674 36624 1730 36680
rect 1306 35944 1362 36000
rect 1306 34856 1362 34912
rect 1214 34448 1270 34504
rect 1674 35572 1676 35592
rect 1676 35572 1728 35592
rect 1728 35572 1730 35592
rect 1674 35536 1730 35572
rect 1398 34040 1454 34096
rect 1306 32408 1362 32464
rect 1674 33632 1730 33688
rect 1582 33496 1638 33552
rect 1398 32000 1454 32056
rect 1122 30776 1178 30832
rect 1122 29688 1178 29744
rect 1674 32408 1730 32464
rect 1490 31456 1546 31512
rect 1306 30504 1362 30560
rect 1398 30232 1454 30288
rect 1582 30232 1638 30288
rect 1306 29416 1362 29472
rect 1214 28600 1270 28656
rect 1398 28056 1454 28112
rect 1214 27376 1270 27432
rect 1214 26968 1270 27024
rect 1306 26696 1362 26752
rect 1674 28872 1730 28928
rect 1950 32136 2006 32192
rect 2226 33904 2282 33960
rect 2134 32544 2190 32600
rect 2226 31628 2228 31648
rect 2228 31628 2280 31648
rect 2280 31628 2282 31648
rect 2226 31592 2282 31628
rect 2226 30776 2282 30832
rect 2134 30368 2190 30424
rect 2870 37848 2926 37904
rect 2778 37304 2834 37360
rect 2778 35400 2834 35456
rect 2870 34584 2926 34640
rect 2502 32816 2558 32872
rect 2778 32952 2834 33008
rect 2778 32816 2834 32872
rect 2686 32680 2742 32736
rect 2870 32408 2926 32464
rect 2134 29416 2190 29472
rect 1582 27920 1638 27976
rect 1674 27104 1730 27160
rect 1122 23024 1178 23080
rect 1582 26288 1638 26344
rect 1398 25608 1454 25664
rect 1306 24792 1362 24848
rect 1582 25100 1584 25120
rect 1584 25100 1636 25120
rect 1636 25100 1638 25120
rect 1582 25064 1638 25100
rect 1306 24556 1308 24576
rect 1308 24556 1360 24576
rect 1360 24556 1362 24576
rect 1306 24520 1362 24556
rect 1306 23432 1362 23488
rect 1306 22888 1362 22944
rect 846 21800 902 21856
rect 1030 21564 1032 21584
rect 1032 21564 1084 21584
rect 1084 21564 1086 21584
rect 1030 21528 1086 21564
rect 938 21256 994 21312
rect 754 19080 810 19136
rect 754 18536 810 18592
rect 938 19488 994 19544
rect 938 18828 994 18864
rect 938 18808 940 18828
rect 940 18808 992 18828
rect 992 18808 994 18828
rect 938 17448 994 17504
rect 1674 23976 1730 24032
rect 1674 23724 1730 23760
rect 1674 23704 1676 23724
rect 1676 23704 1728 23724
rect 1728 23704 1730 23724
rect 2134 28872 2190 28928
rect 2778 31320 2834 31376
rect 2778 29688 2834 29744
rect 2410 28192 2466 28248
rect 2042 26696 2098 26752
rect 2226 26560 2282 26616
rect 1858 24792 1914 24848
rect 1950 24248 2006 24304
rect 2134 26424 2190 26480
rect 2134 25880 2190 25936
rect 2226 25744 2282 25800
rect 2594 27512 2650 27568
rect 2502 26832 2558 26888
rect 2502 26152 2558 26208
rect 2410 25764 2466 25800
rect 2410 25744 2412 25764
rect 2412 25744 2464 25764
rect 2464 25744 2466 25764
rect 3923 43002 3979 43004
rect 4003 43002 4059 43004
rect 4083 43002 4139 43004
rect 4163 43002 4219 43004
rect 3923 42950 3969 43002
rect 3969 42950 3979 43002
rect 4003 42950 4033 43002
rect 4033 42950 4045 43002
rect 4045 42950 4059 43002
rect 4083 42950 4097 43002
rect 4097 42950 4109 43002
rect 4109 42950 4139 43002
rect 4163 42950 4173 43002
rect 4173 42950 4219 43002
rect 3923 42948 3979 42950
rect 4003 42948 4059 42950
rect 4083 42948 4139 42950
rect 4163 42948 4219 42950
rect 3923 41914 3979 41916
rect 4003 41914 4059 41916
rect 4083 41914 4139 41916
rect 4163 41914 4219 41916
rect 3923 41862 3969 41914
rect 3969 41862 3979 41914
rect 4003 41862 4033 41914
rect 4033 41862 4045 41914
rect 4045 41862 4059 41914
rect 4083 41862 4097 41914
rect 4097 41862 4109 41914
rect 4109 41862 4139 41914
rect 4163 41862 4173 41914
rect 4173 41862 4219 41914
rect 3923 41860 3979 41862
rect 4003 41860 4059 41862
rect 4083 41860 4139 41862
rect 4163 41860 4219 41862
rect 3606 39480 3662 39536
rect 3422 38956 3478 38992
rect 3422 38936 3424 38956
rect 3424 38936 3476 38956
rect 3476 38936 3478 38956
rect 3238 38292 3240 38312
rect 3240 38292 3292 38312
rect 3292 38292 3294 38312
rect 3238 38256 3294 38292
rect 3054 36216 3110 36272
rect 3238 36488 3294 36544
rect 3146 34992 3202 35048
rect 3054 31184 3110 31240
rect 3054 28328 3110 28384
rect 3054 27648 3110 27704
rect 2962 27412 2964 27432
rect 2964 27412 3016 27432
rect 3016 27412 3018 27432
rect 2962 27376 3018 27412
rect 2778 27240 2834 27296
rect 2962 27240 3018 27296
rect 2870 26696 2926 26752
rect 2686 25236 2688 25256
rect 2688 25236 2740 25256
rect 2740 25236 2742 25256
rect 2686 25200 2742 25236
rect 1490 22616 1546 22672
rect 1306 22228 1362 22264
rect 1306 22208 1308 22228
rect 1308 22208 1360 22228
rect 1360 22208 1362 22228
rect 1306 22072 1362 22128
rect 1674 21936 1730 21992
rect 1582 20984 1638 21040
rect 1398 20712 1454 20768
rect 1490 20576 1546 20632
rect 1214 20168 1270 20224
rect 1306 19896 1362 19952
rect 2134 21392 2190 21448
rect 1306 19352 1362 19408
rect 1582 19372 1638 19408
rect 1582 19352 1584 19372
rect 1584 19352 1636 19372
rect 1636 19352 1638 19372
rect 1398 17992 1454 18048
rect 1306 17720 1362 17776
rect 1306 16904 1362 16960
rect 1306 16632 1362 16688
rect 1122 16224 1178 16280
rect 1582 18672 1638 18728
rect 1950 18844 1952 18864
rect 1952 18844 2004 18864
rect 2004 18844 2006 18864
rect 1950 18808 2006 18844
rect 1950 18128 2006 18184
rect 1766 17720 1822 17776
rect 1858 17176 1914 17232
rect 1674 16904 1730 16960
rect 1674 16668 1676 16688
rect 1676 16668 1728 16688
rect 1728 16668 1730 16688
rect 1674 16632 1730 16668
rect 1582 16088 1638 16144
rect 1398 15408 1454 15464
rect 1306 14492 1308 14512
rect 1308 14492 1360 14512
rect 1360 14492 1362 14512
rect 1306 14456 1362 14492
rect 1490 14728 1546 14784
rect 1306 13912 1362 13968
rect 1306 13776 1362 13832
rect 1766 16360 1822 16416
rect 1766 15000 1822 15056
rect 1490 13776 1546 13832
rect 1306 13368 1362 13424
rect 1674 14184 1730 14240
rect 2134 20848 2190 20904
rect 2594 24792 2650 24848
rect 3054 24656 3110 24712
rect 3238 34040 3294 34096
rect 3882 41112 3938 41168
rect 3923 40826 3979 40828
rect 4003 40826 4059 40828
rect 4083 40826 4139 40828
rect 4163 40826 4219 40828
rect 3923 40774 3969 40826
rect 3969 40774 3979 40826
rect 4003 40774 4033 40826
rect 4033 40774 4045 40826
rect 4045 40774 4059 40826
rect 4083 40774 4097 40826
rect 4097 40774 4109 40826
rect 4109 40774 4139 40826
rect 4163 40774 4173 40826
rect 4173 40774 4219 40826
rect 3923 40772 3979 40774
rect 4003 40772 4059 40774
rect 4083 40772 4139 40774
rect 4163 40772 4219 40774
rect 3882 40432 3938 40488
rect 4158 40452 4214 40488
rect 4158 40432 4160 40452
rect 4160 40432 4212 40452
rect 4212 40432 4214 40452
rect 3974 39888 4030 39944
rect 4250 40024 4306 40080
rect 3923 39738 3979 39740
rect 4003 39738 4059 39740
rect 4083 39738 4139 39740
rect 4163 39738 4219 39740
rect 3923 39686 3969 39738
rect 3969 39686 3979 39738
rect 4003 39686 4033 39738
rect 4033 39686 4045 39738
rect 4045 39686 4059 39738
rect 4083 39686 4097 39738
rect 4097 39686 4109 39738
rect 4109 39686 4139 39738
rect 4163 39686 4173 39738
rect 4173 39686 4219 39738
rect 3923 39684 3979 39686
rect 4003 39684 4059 39686
rect 4083 39684 4139 39686
rect 4163 39684 4219 39686
rect 4710 41656 4766 41712
rect 3923 38650 3979 38652
rect 4003 38650 4059 38652
rect 4083 38650 4139 38652
rect 4163 38650 4219 38652
rect 3923 38598 3969 38650
rect 3969 38598 3979 38650
rect 4003 38598 4033 38650
rect 4033 38598 4045 38650
rect 4045 38598 4059 38650
rect 4083 38598 4097 38650
rect 4097 38598 4109 38650
rect 4109 38598 4139 38650
rect 4163 38598 4173 38650
rect 4173 38598 4219 38650
rect 3923 38596 3979 38598
rect 4003 38596 4059 38598
rect 4083 38596 4139 38598
rect 4163 38596 4219 38598
rect 4066 37868 4122 37904
rect 4066 37848 4068 37868
rect 4068 37848 4120 37868
rect 4120 37848 4122 37868
rect 4158 37748 4160 37768
rect 4160 37748 4212 37768
rect 4212 37748 4214 37768
rect 4158 37712 4214 37748
rect 3923 37562 3979 37564
rect 4003 37562 4059 37564
rect 4083 37562 4139 37564
rect 4163 37562 4219 37564
rect 3923 37510 3969 37562
rect 3969 37510 3979 37562
rect 4003 37510 4033 37562
rect 4033 37510 4045 37562
rect 4045 37510 4059 37562
rect 4083 37510 4097 37562
rect 4097 37510 4109 37562
rect 4109 37510 4139 37562
rect 4163 37510 4173 37562
rect 4173 37510 4219 37562
rect 3923 37508 3979 37510
rect 4003 37508 4059 37510
rect 4083 37508 4139 37510
rect 4163 37508 4219 37510
rect 5170 41556 5172 41576
rect 5172 41556 5224 41576
rect 5224 41556 5226 41576
rect 5170 41520 5226 41556
rect 4618 37984 4674 38040
rect 3882 36760 3938 36816
rect 3923 36474 3979 36476
rect 4003 36474 4059 36476
rect 4083 36474 4139 36476
rect 4163 36474 4219 36476
rect 3923 36422 3969 36474
rect 3969 36422 3979 36474
rect 4003 36422 4033 36474
rect 4033 36422 4045 36474
rect 4045 36422 4059 36474
rect 4083 36422 4097 36474
rect 4097 36422 4109 36474
rect 4109 36422 4139 36474
rect 4163 36422 4173 36474
rect 4173 36422 4219 36474
rect 3923 36420 3979 36422
rect 4003 36420 4059 36422
rect 4083 36420 4139 36422
rect 4163 36420 4219 36422
rect 3974 35944 4030 36000
rect 3790 35808 3846 35864
rect 4066 35536 4122 35592
rect 3923 35386 3979 35388
rect 4003 35386 4059 35388
rect 4083 35386 4139 35388
rect 4163 35386 4219 35388
rect 3923 35334 3969 35386
rect 3969 35334 3979 35386
rect 4003 35334 4033 35386
rect 4033 35334 4045 35386
rect 4045 35334 4059 35386
rect 4083 35334 4097 35386
rect 4097 35334 4109 35386
rect 4109 35334 4139 35386
rect 4163 35334 4173 35386
rect 4173 35334 4219 35386
rect 3923 35332 3979 35334
rect 4003 35332 4059 35334
rect 4083 35332 4139 35334
rect 4163 35332 4219 35334
rect 4342 36216 4398 36272
rect 4526 36216 4582 36272
rect 4342 35672 4398 35728
rect 3330 31728 3386 31784
rect 3238 30368 3294 30424
rect 3606 32952 3662 33008
rect 3790 34992 3846 35048
rect 3923 34298 3979 34300
rect 4003 34298 4059 34300
rect 4083 34298 4139 34300
rect 4163 34298 4219 34300
rect 3923 34246 3969 34298
rect 3969 34246 3979 34298
rect 4003 34246 4033 34298
rect 4033 34246 4045 34298
rect 4045 34246 4059 34298
rect 4083 34246 4097 34298
rect 4097 34246 4109 34298
rect 4109 34246 4139 34298
rect 4163 34246 4173 34298
rect 4173 34246 4219 34298
rect 3923 34244 3979 34246
rect 4003 34244 4059 34246
rect 4083 34244 4139 34246
rect 4163 34244 4219 34246
rect 3882 33768 3938 33824
rect 3790 33360 3846 33416
rect 3923 33210 3979 33212
rect 4003 33210 4059 33212
rect 4083 33210 4139 33212
rect 4163 33210 4219 33212
rect 3923 33158 3969 33210
rect 3969 33158 3979 33210
rect 4003 33158 4033 33210
rect 4033 33158 4045 33210
rect 4045 33158 4059 33210
rect 4083 33158 4097 33210
rect 4097 33158 4109 33210
rect 4109 33158 4139 33210
rect 4163 33158 4173 33210
rect 4173 33158 4219 33210
rect 3923 33156 3979 33158
rect 4003 33156 4059 33158
rect 4083 33156 4139 33158
rect 4163 33156 4219 33158
rect 4342 33088 4398 33144
rect 3974 32816 4030 32872
rect 4250 32272 4306 32328
rect 3606 30504 3662 30560
rect 3923 32122 3979 32124
rect 4003 32122 4059 32124
rect 4083 32122 4139 32124
rect 4163 32122 4219 32124
rect 3923 32070 3969 32122
rect 3969 32070 3979 32122
rect 4003 32070 4033 32122
rect 4033 32070 4045 32122
rect 4045 32070 4059 32122
rect 4083 32070 4097 32122
rect 4097 32070 4109 32122
rect 4109 32070 4139 32122
rect 4163 32070 4173 32122
rect 4173 32070 4219 32122
rect 3923 32068 3979 32070
rect 4003 32068 4059 32070
rect 4083 32068 4139 32070
rect 4163 32068 4219 32070
rect 3882 31320 3938 31376
rect 3923 31034 3979 31036
rect 4003 31034 4059 31036
rect 4083 31034 4139 31036
rect 4163 31034 4219 31036
rect 3923 30982 3969 31034
rect 3969 30982 3979 31034
rect 4003 30982 4033 31034
rect 4033 30982 4045 31034
rect 4045 30982 4059 31034
rect 4083 30982 4097 31034
rect 4097 30982 4109 31034
rect 4109 30982 4139 31034
rect 4163 30982 4173 31034
rect 4173 30982 4219 31034
rect 3923 30980 3979 30982
rect 4003 30980 4059 30982
rect 4083 30980 4139 30982
rect 4163 30980 4219 30982
rect 3923 29946 3979 29948
rect 4003 29946 4059 29948
rect 4083 29946 4139 29948
rect 4163 29946 4219 29948
rect 3923 29894 3969 29946
rect 3969 29894 3979 29946
rect 4003 29894 4033 29946
rect 4033 29894 4045 29946
rect 4045 29894 4059 29946
rect 4083 29894 4097 29946
rect 4097 29894 4109 29946
rect 4109 29894 4139 29946
rect 4163 29894 4173 29946
rect 4173 29894 4219 29946
rect 3923 29892 3979 29894
rect 4003 29892 4059 29894
rect 4083 29892 4139 29894
rect 4163 29892 4219 29894
rect 2778 24112 2834 24168
rect 2778 22480 2834 22536
rect 2686 22208 2742 22264
rect 2778 21800 2834 21856
rect 3238 21800 3294 21856
rect 2226 20304 2282 20360
rect 2594 19352 2650 19408
rect 3606 28056 3662 28112
rect 3923 28858 3979 28860
rect 4003 28858 4059 28860
rect 4083 28858 4139 28860
rect 4163 28858 4219 28860
rect 3923 28806 3969 28858
rect 3969 28806 3979 28858
rect 4003 28806 4033 28858
rect 4033 28806 4045 28858
rect 4045 28806 4059 28858
rect 4083 28806 4097 28858
rect 4097 28806 4109 28858
rect 4109 28806 4139 28858
rect 4163 28806 4173 28858
rect 4173 28806 4219 28858
rect 3923 28804 3979 28806
rect 4003 28804 4059 28806
rect 4083 28804 4139 28806
rect 4163 28804 4219 28806
rect 3882 28484 3938 28520
rect 3882 28464 3884 28484
rect 3884 28464 3936 28484
rect 3936 28464 3938 28484
rect 3790 27784 3846 27840
rect 3606 27512 3662 27568
rect 3923 27770 3979 27772
rect 4003 27770 4059 27772
rect 4083 27770 4139 27772
rect 4163 27770 4219 27772
rect 3923 27718 3969 27770
rect 3969 27718 3979 27770
rect 4003 27718 4033 27770
rect 4033 27718 4045 27770
rect 4045 27718 4059 27770
rect 4083 27718 4097 27770
rect 4097 27718 4109 27770
rect 4109 27718 4139 27770
rect 4163 27718 4173 27770
rect 4173 27718 4219 27770
rect 3923 27716 3979 27718
rect 4003 27716 4059 27718
rect 4083 27716 4139 27718
rect 4163 27716 4219 27718
rect 3923 26682 3979 26684
rect 4003 26682 4059 26684
rect 4083 26682 4139 26684
rect 4163 26682 4219 26684
rect 3923 26630 3969 26682
rect 3969 26630 3979 26682
rect 4003 26630 4033 26682
rect 4033 26630 4045 26682
rect 4045 26630 4059 26682
rect 4083 26630 4097 26682
rect 4097 26630 4109 26682
rect 4109 26630 4139 26682
rect 4163 26630 4173 26682
rect 4173 26630 4219 26682
rect 3923 26628 3979 26630
rect 4003 26628 4059 26630
rect 4083 26628 4139 26630
rect 4163 26628 4219 26630
rect 3606 26016 3662 26072
rect 4158 26016 4214 26072
rect 4802 35944 4858 36000
rect 4618 34992 4674 35048
rect 4618 32000 4674 32056
rect 4618 31476 4674 31512
rect 4618 31456 4620 31476
rect 4620 31456 4672 31476
rect 4672 31456 4674 31476
rect 4618 31048 4674 31104
rect 4802 34856 4858 34912
rect 4802 30776 4858 30832
rect 5262 40296 5318 40352
rect 5446 40160 5502 40216
rect 5170 36100 5226 36136
rect 5170 36080 5172 36100
rect 5172 36080 5224 36100
rect 5224 36080 5226 36100
rect 5078 33224 5134 33280
rect 4802 30232 4858 30288
rect 3923 25594 3979 25596
rect 4003 25594 4059 25596
rect 4083 25594 4139 25596
rect 4163 25594 4219 25596
rect 3923 25542 3969 25594
rect 3969 25542 3979 25594
rect 4003 25542 4033 25594
rect 4033 25542 4045 25594
rect 4045 25542 4059 25594
rect 4083 25542 4097 25594
rect 4097 25542 4109 25594
rect 4109 25542 4139 25594
rect 4163 25542 4173 25594
rect 4173 25542 4219 25594
rect 3923 25540 3979 25542
rect 4003 25540 4059 25542
rect 4083 25540 4139 25542
rect 4163 25540 4219 25542
rect 3923 24506 3979 24508
rect 4003 24506 4059 24508
rect 4083 24506 4139 24508
rect 4163 24506 4219 24508
rect 3923 24454 3969 24506
rect 3969 24454 3979 24506
rect 4003 24454 4033 24506
rect 4033 24454 4045 24506
rect 4045 24454 4059 24506
rect 4083 24454 4097 24506
rect 4097 24454 4109 24506
rect 4109 24454 4139 24506
rect 4163 24454 4173 24506
rect 4173 24454 4219 24506
rect 3923 24452 3979 24454
rect 4003 24452 4059 24454
rect 4083 24452 4139 24454
rect 4163 24452 4219 24454
rect 3422 23160 3478 23216
rect 3923 23418 3979 23420
rect 4003 23418 4059 23420
rect 4083 23418 4139 23420
rect 4163 23418 4219 23420
rect 3923 23366 3969 23418
rect 3969 23366 3979 23418
rect 4003 23366 4033 23418
rect 4033 23366 4045 23418
rect 4045 23366 4059 23418
rect 4083 23366 4097 23418
rect 4097 23366 4109 23418
rect 4109 23366 4139 23418
rect 4163 23366 4173 23418
rect 4173 23366 4219 23418
rect 3923 23364 3979 23366
rect 4003 23364 4059 23366
rect 4083 23364 4139 23366
rect 4163 23364 4219 23366
rect 3974 23024 4030 23080
rect 3790 22888 3846 22944
rect 4066 22636 4122 22672
rect 4066 22616 4068 22636
rect 4068 22616 4120 22636
rect 4120 22616 4122 22636
rect 3923 22330 3979 22332
rect 4003 22330 4059 22332
rect 4083 22330 4139 22332
rect 4163 22330 4219 22332
rect 3923 22278 3969 22330
rect 3969 22278 3979 22330
rect 4003 22278 4033 22330
rect 4033 22278 4045 22330
rect 4045 22278 4059 22330
rect 4083 22278 4097 22330
rect 4097 22278 4109 22330
rect 4109 22278 4139 22330
rect 4163 22278 4173 22330
rect 4173 22278 4219 22330
rect 3923 22276 3979 22278
rect 4003 22276 4059 22278
rect 4083 22276 4139 22278
rect 4163 22276 4219 22278
rect 4618 27920 4674 27976
rect 4618 27784 4674 27840
rect 4894 29416 4950 29472
rect 4894 29280 4950 29336
rect 4894 28736 4950 28792
rect 4894 28464 4950 28520
rect 4894 28192 4950 28248
rect 4710 24676 4766 24712
rect 4710 24656 4712 24676
rect 4712 24656 4764 24676
rect 4764 24656 4766 24676
rect 5078 30660 5134 30696
rect 5078 30640 5080 30660
rect 5080 30640 5132 30660
rect 5132 30640 5134 30660
rect 6182 41792 6238 41848
rect 6890 43546 6946 43548
rect 6970 43546 7026 43548
rect 7050 43546 7106 43548
rect 7130 43546 7186 43548
rect 6890 43494 6936 43546
rect 6936 43494 6946 43546
rect 6970 43494 7000 43546
rect 7000 43494 7012 43546
rect 7012 43494 7026 43546
rect 7050 43494 7064 43546
rect 7064 43494 7076 43546
rect 7076 43494 7106 43546
rect 7130 43494 7140 43546
rect 7140 43494 7186 43546
rect 6890 43492 6946 43494
rect 6970 43492 7026 43494
rect 7050 43492 7106 43494
rect 7130 43492 7186 43494
rect 6890 42458 6946 42460
rect 6970 42458 7026 42460
rect 7050 42458 7106 42460
rect 7130 42458 7186 42460
rect 6890 42406 6936 42458
rect 6936 42406 6946 42458
rect 6970 42406 7000 42458
rect 7000 42406 7012 42458
rect 7012 42406 7026 42458
rect 7050 42406 7064 42458
rect 7064 42406 7076 42458
rect 7076 42406 7106 42458
rect 7130 42406 7140 42458
rect 7140 42406 7186 42458
rect 6890 42404 6946 42406
rect 6970 42404 7026 42406
rect 7050 42404 7106 42406
rect 7130 42404 7186 42406
rect 6642 41792 6698 41848
rect 7378 41792 7434 41848
rect 6734 41556 6736 41576
rect 6736 41556 6788 41576
rect 6788 41556 6790 41576
rect 6734 41520 6790 41556
rect 6890 41370 6946 41372
rect 6970 41370 7026 41372
rect 7050 41370 7106 41372
rect 7130 41370 7186 41372
rect 6890 41318 6936 41370
rect 6936 41318 6946 41370
rect 6970 41318 7000 41370
rect 7000 41318 7012 41370
rect 7012 41318 7026 41370
rect 7050 41318 7064 41370
rect 7064 41318 7076 41370
rect 7076 41318 7106 41370
rect 7130 41318 7140 41370
rect 7140 41318 7186 41370
rect 6890 41316 6946 41318
rect 6970 41316 7026 41318
rect 7050 41316 7106 41318
rect 7130 41316 7186 41318
rect 5262 31184 5318 31240
rect 5170 29960 5226 30016
rect 5538 31476 5594 31512
rect 5538 31456 5540 31476
rect 5540 31456 5592 31476
rect 5592 31456 5594 31476
rect 5446 31184 5502 31240
rect 5354 28464 5410 28520
rect 5170 27920 5226 27976
rect 5170 27376 5226 27432
rect 3790 21936 3846 21992
rect 3422 20304 3478 20360
rect 3330 19624 3386 19680
rect 3054 19352 3110 19408
rect 3514 19624 3570 19680
rect 3606 19352 3662 19408
rect 2870 18536 2926 18592
rect 2226 17196 2282 17232
rect 2226 17176 2228 17196
rect 2228 17176 2280 17196
rect 2280 17176 2282 17196
rect 1858 13776 1914 13832
rect 1582 12824 1638 12880
rect 1306 12008 1362 12064
rect 1674 12552 1730 12608
rect 1490 10376 1546 10432
rect 1398 9832 1454 9888
rect 1306 9016 1362 9072
rect 1766 11192 1822 11248
rect 1858 8880 1914 8936
rect 1582 8472 1638 8528
rect 1306 7656 1362 7712
rect 1398 7248 1454 7304
rect 1306 7112 1362 7168
rect 1214 6296 1270 6352
rect 938 6160 994 6216
rect 1122 5480 1178 5536
rect 1766 8064 1822 8120
rect 2226 14456 2282 14512
rect 2318 13912 2374 13968
rect 2686 16108 2742 16144
rect 2686 16088 2688 16108
rect 2688 16088 2740 16108
rect 2740 16088 2742 16108
rect 2594 15544 2650 15600
rect 2318 13504 2374 13560
rect 2318 12280 2374 12336
rect 2318 10104 2374 10160
rect 2134 9424 2190 9480
rect 2134 7828 2136 7848
rect 2136 7828 2188 7848
rect 2188 7828 2190 7848
rect 2134 7792 2190 7828
rect 2318 8880 2374 8936
rect 1582 6024 1638 6080
rect 1674 5652 1676 5672
rect 1676 5652 1728 5672
rect 1728 5652 1730 5672
rect 1674 5616 1730 5652
rect 1582 4276 1638 4312
rect 1582 4256 1584 4276
rect 1584 4256 1636 4276
rect 1636 4256 1638 4276
rect 2134 6568 2190 6624
rect 2594 13368 2650 13424
rect 3054 13776 3110 13832
rect 3514 19216 3570 19272
rect 3923 21242 3979 21244
rect 4003 21242 4059 21244
rect 4083 21242 4139 21244
rect 4163 21242 4219 21244
rect 3923 21190 3969 21242
rect 3969 21190 3979 21242
rect 4003 21190 4033 21242
rect 4033 21190 4045 21242
rect 4045 21190 4059 21242
rect 4083 21190 4097 21242
rect 4097 21190 4109 21242
rect 4109 21190 4139 21242
rect 4163 21190 4173 21242
rect 4173 21190 4219 21242
rect 3923 21188 3979 21190
rect 4003 21188 4059 21190
rect 4083 21188 4139 21190
rect 4163 21188 4219 21190
rect 3790 20440 3846 20496
rect 4250 20304 4306 20360
rect 3923 20154 3979 20156
rect 4003 20154 4059 20156
rect 4083 20154 4139 20156
rect 4163 20154 4219 20156
rect 3923 20102 3969 20154
rect 3969 20102 3979 20154
rect 4003 20102 4033 20154
rect 4033 20102 4045 20154
rect 4045 20102 4059 20154
rect 4083 20102 4097 20154
rect 4097 20102 4109 20154
rect 4109 20102 4139 20154
rect 4163 20102 4173 20154
rect 4173 20102 4219 20154
rect 3923 20100 3979 20102
rect 4003 20100 4059 20102
rect 4083 20100 4139 20102
rect 4163 20100 4219 20102
rect 4250 19488 4306 19544
rect 3923 19066 3979 19068
rect 4003 19066 4059 19068
rect 4083 19066 4139 19068
rect 4163 19066 4219 19068
rect 3923 19014 3969 19066
rect 3969 19014 3979 19066
rect 4003 19014 4033 19066
rect 4033 19014 4045 19066
rect 4045 19014 4059 19066
rect 4083 19014 4097 19066
rect 4097 19014 4109 19066
rect 4109 19014 4139 19066
rect 4163 19014 4173 19066
rect 4173 19014 4219 19066
rect 3923 19012 3979 19014
rect 4003 19012 4059 19014
rect 4083 19012 4139 19014
rect 4163 19012 4219 19014
rect 3514 18264 3570 18320
rect 3238 12960 3294 13016
rect 3514 13640 3570 13696
rect 3514 13096 3570 13152
rect 2778 12144 2834 12200
rect 2686 11192 2742 11248
rect 2870 11600 2926 11656
rect 3422 12552 3478 12608
rect 3330 12144 3386 12200
rect 3238 11464 3294 11520
rect 1766 3576 1822 3632
rect 2502 5480 2558 5536
rect 386 1400 442 1456
rect 2870 9560 2926 9616
rect 2870 8744 2926 8800
rect 3146 10648 3202 10704
rect 3330 10920 3386 10976
rect 4434 21956 4490 21992
rect 4434 21936 4436 21956
rect 4436 21936 4488 21956
rect 4488 21936 4490 21956
rect 4434 19896 4490 19952
rect 3923 17978 3979 17980
rect 4003 17978 4059 17980
rect 4083 17978 4139 17980
rect 4163 17978 4219 17980
rect 3923 17926 3969 17978
rect 3969 17926 3979 17978
rect 4003 17926 4033 17978
rect 4033 17926 4045 17978
rect 4045 17926 4059 17978
rect 4083 17926 4097 17978
rect 4097 17926 4109 17978
rect 4109 17926 4139 17978
rect 4163 17926 4173 17978
rect 4173 17926 4219 17978
rect 3923 17924 3979 17926
rect 4003 17924 4059 17926
rect 4083 17924 4139 17926
rect 4163 17924 4219 17926
rect 4710 22072 4766 22128
rect 4618 18944 4674 19000
rect 4250 17720 4306 17776
rect 3923 16890 3979 16892
rect 4003 16890 4059 16892
rect 4083 16890 4139 16892
rect 4163 16890 4219 16892
rect 3923 16838 3969 16890
rect 3969 16838 3979 16890
rect 4003 16838 4033 16890
rect 4033 16838 4045 16890
rect 4045 16838 4059 16890
rect 4083 16838 4097 16890
rect 4097 16838 4109 16890
rect 4109 16838 4139 16890
rect 4163 16838 4173 16890
rect 4173 16838 4219 16890
rect 3923 16836 3979 16838
rect 4003 16836 4059 16838
rect 4083 16836 4139 16838
rect 4163 16836 4219 16838
rect 4250 16632 4306 16688
rect 3698 15816 3754 15872
rect 3923 15802 3979 15804
rect 4003 15802 4059 15804
rect 4083 15802 4139 15804
rect 4163 15802 4219 15804
rect 3923 15750 3969 15802
rect 3969 15750 3979 15802
rect 4003 15750 4033 15802
rect 4033 15750 4045 15802
rect 4045 15750 4059 15802
rect 4083 15750 4097 15802
rect 4097 15750 4109 15802
rect 4109 15750 4139 15802
rect 4163 15750 4173 15802
rect 4173 15750 4219 15802
rect 3923 15748 3979 15750
rect 4003 15748 4059 15750
rect 4083 15748 4139 15750
rect 4163 15748 4219 15750
rect 4066 15272 4122 15328
rect 3923 14714 3979 14716
rect 4003 14714 4059 14716
rect 4083 14714 4139 14716
rect 4163 14714 4219 14716
rect 3923 14662 3969 14714
rect 3969 14662 3979 14714
rect 4003 14662 4033 14714
rect 4033 14662 4045 14714
rect 4045 14662 4059 14714
rect 4083 14662 4097 14714
rect 4097 14662 4109 14714
rect 4109 14662 4139 14714
rect 4163 14662 4173 14714
rect 4173 14662 4219 14714
rect 3923 14660 3979 14662
rect 4003 14660 4059 14662
rect 4083 14660 4139 14662
rect 4163 14660 4219 14662
rect 4986 20032 5042 20088
rect 4618 15952 4674 16008
rect 4618 15272 4674 15328
rect 3923 13626 3979 13628
rect 4003 13626 4059 13628
rect 4083 13626 4139 13628
rect 4163 13626 4219 13628
rect 3923 13574 3969 13626
rect 3969 13574 3979 13626
rect 4003 13574 4033 13626
rect 4033 13574 4045 13626
rect 4045 13574 4059 13626
rect 4083 13574 4097 13626
rect 4097 13574 4109 13626
rect 4109 13574 4139 13626
rect 4163 13574 4173 13626
rect 4173 13574 4219 13626
rect 3923 13572 3979 13574
rect 4003 13572 4059 13574
rect 4083 13572 4139 13574
rect 4163 13572 4219 13574
rect 3974 12960 4030 13016
rect 3790 12552 3846 12608
rect 3923 12538 3979 12540
rect 4003 12538 4059 12540
rect 4083 12538 4139 12540
rect 4163 12538 4219 12540
rect 3923 12486 3969 12538
rect 3969 12486 3979 12538
rect 4003 12486 4033 12538
rect 4033 12486 4045 12538
rect 4045 12486 4059 12538
rect 4083 12486 4097 12538
rect 4097 12486 4109 12538
rect 4109 12486 4139 12538
rect 4163 12486 4173 12538
rect 4173 12486 4219 12538
rect 3923 12484 3979 12486
rect 4003 12484 4059 12486
rect 4083 12484 4139 12486
rect 4163 12484 4219 12486
rect 3974 11736 4030 11792
rect 4066 11600 4122 11656
rect 3923 11450 3979 11452
rect 4003 11450 4059 11452
rect 4083 11450 4139 11452
rect 4163 11450 4219 11452
rect 3923 11398 3969 11450
rect 3969 11398 3979 11450
rect 4003 11398 4033 11450
rect 4033 11398 4045 11450
rect 4045 11398 4059 11450
rect 4083 11398 4097 11450
rect 4097 11398 4109 11450
rect 4109 11398 4139 11450
rect 4163 11398 4173 11450
rect 4173 11398 4219 11450
rect 3923 11396 3979 11398
rect 4003 11396 4059 11398
rect 4083 11396 4139 11398
rect 4163 11396 4219 11398
rect 3422 8880 3478 8936
rect 3330 8472 3386 8528
rect 3054 7928 3110 7984
rect 2778 5752 2834 5808
rect 2962 4664 3018 4720
rect 2594 3984 2650 4040
rect 2870 3440 2926 3496
rect 1674 1300 1676 1320
rect 1676 1300 1728 1320
rect 1728 1300 1730 1320
rect 1674 1264 1730 1300
rect 2042 1300 2044 1320
rect 2044 1300 2096 1320
rect 2096 1300 2098 1320
rect 2042 1264 2098 1300
rect 3330 6860 3386 6896
rect 3330 6840 3332 6860
rect 3332 6840 3384 6860
rect 3384 6840 3386 6860
rect 3330 6432 3386 6488
rect 3974 10668 4030 10704
rect 3974 10648 3976 10668
rect 3976 10648 4028 10668
rect 4028 10648 4030 10668
rect 3923 10362 3979 10364
rect 4003 10362 4059 10364
rect 4083 10362 4139 10364
rect 4163 10362 4219 10364
rect 3923 10310 3969 10362
rect 3969 10310 3979 10362
rect 4003 10310 4033 10362
rect 4033 10310 4045 10362
rect 4045 10310 4059 10362
rect 4083 10310 4097 10362
rect 4097 10310 4109 10362
rect 4109 10310 4139 10362
rect 4163 10310 4173 10362
rect 4173 10310 4219 10362
rect 3923 10308 3979 10310
rect 4003 10308 4059 10310
rect 4083 10308 4139 10310
rect 4163 10308 4219 10310
rect 3923 9274 3979 9276
rect 4003 9274 4059 9276
rect 4083 9274 4139 9276
rect 4163 9274 4219 9276
rect 3923 9222 3969 9274
rect 3969 9222 3979 9274
rect 4003 9222 4033 9274
rect 4033 9222 4045 9274
rect 4045 9222 4059 9274
rect 4083 9222 4097 9274
rect 4097 9222 4109 9274
rect 4109 9222 4139 9274
rect 4163 9222 4173 9274
rect 4173 9222 4219 9274
rect 3923 9220 3979 9222
rect 4003 9220 4059 9222
rect 4083 9220 4139 9222
rect 4163 9220 4219 9222
rect 3790 8472 3846 8528
rect 3974 8472 4030 8528
rect 3790 8336 3846 8392
rect 3698 6604 3700 6624
rect 3700 6604 3752 6624
rect 3752 6604 3754 6624
rect 3698 6568 3754 6604
rect 3698 6160 3754 6216
rect 3422 4564 3424 4584
rect 3424 4564 3476 4584
rect 3476 4564 3478 4584
rect 3422 4528 3478 4564
rect 3923 8186 3979 8188
rect 4003 8186 4059 8188
rect 4083 8186 4139 8188
rect 4163 8186 4219 8188
rect 3923 8134 3969 8186
rect 3969 8134 3979 8186
rect 4003 8134 4033 8186
rect 4033 8134 4045 8186
rect 4045 8134 4059 8186
rect 4083 8134 4097 8186
rect 4097 8134 4109 8186
rect 4109 8134 4139 8186
rect 4163 8134 4173 8186
rect 4173 8134 4219 8186
rect 3923 8132 3979 8134
rect 4003 8132 4059 8134
rect 4083 8132 4139 8134
rect 4163 8132 4219 8134
rect 4618 12844 4674 12880
rect 4618 12824 4620 12844
rect 4620 12824 4672 12844
rect 4672 12824 4674 12844
rect 4618 12280 4674 12336
rect 4802 11212 4858 11248
rect 4802 11192 4804 11212
rect 4804 11192 4856 11212
rect 4856 11192 4858 11212
rect 4802 10104 4858 10160
rect 3923 7098 3979 7100
rect 4003 7098 4059 7100
rect 4083 7098 4139 7100
rect 4163 7098 4219 7100
rect 3923 7046 3969 7098
rect 3969 7046 3979 7098
rect 4003 7046 4033 7098
rect 4033 7046 4045 7098
rect 4045 7046 4059 7098
rect 4083 7046 4097 7098
rect 4097 7046 4109 7098
rect 4109 7046 4139 7098
rect 4163 7046 4173 7098
rect 4173 7046 4219 7098
rect 3923 7044 3979 7046
rect 4003 7044 4059 7046
rect 4083 7044 4139 7046
rect 4163 7044 4219 7046
rect 3923 6010 3979 6012
rect 4003 6010 4059 6012
rect 4083 6010 4139 6012
rect 4163 6010 4219 6012
rect 3923 5958 3969 6010
rect 3969 5958 3979 6010
rect 4003 5958 4033 6010
rect 4033 5958 4045 6010
rect 4045 5958 4059 6010
rect 4083 5958 4097 6010
rect 4097 5958 4109 6010
rect 4109 5958 4139 6010
rect 4163 5958 4173 6010
rect 4173 5958 4219 6010
rect 3923 5956 3979 5958
rect 4003 5956 4059 5958
rect 4083 5956 4139 5958
rect 4163 5956 4219 5958
rect 3923 4922 3979 4924
rect 4003 4922 4059 4924
rect 4083 4922 4139 4924
rect 4163 4922 4219 4924
rect 3923 4870 3969 4922
rect 3969 4870 3979 4922
rect 4003 4870 4033 4922
rect 4033 4870 4045 4922
rect 4045 4870 4059 4922
rect 4083 4870 4097 4922
rect 4097 4870 4109 4922
rect 4109 4870 4139 4922
rect 4163 4870 4173 4922
rect 4173 4870 4219 4922
rect 3923 4868 3979 4870
rect 4003 4868 4059 4870
rect 4083 4868 4139 4870
rect 4163 4868 4219 4870
rect 4066 4664 4122 4720
rect 3923 3834 3979 3836
rect 4003 3834 4059 3836
rect 4083 3834 4139 3836
rect 4163 3834 4219 3836
rect 3923 3782 3969 3834
rect 3969 3782 3979 3834
rect 4003 3782 4033 3834
rect 4033 3782 4045 3834
rect 4045 3782 4059 3834
rect 4083 3782 4097 3834
rect 4097 3782 4109 3834
rect 4109 3782 4139 3834
rect 4163 3782 4173 3834
rect 4173 3782 4219 3834
rect 3923 3780 3979 3782
rect 4003 3780 4059 3782
rect 4083 3780 4139 3782
rect 4163 3780 4219 3782
rect 3923 2746 3979 2748
rect 4003 2746 4059 2748
rect 4083 2746 4139 2748
rect 4163 2746 4219 2748
rect 3923 2694 3969 2746
rect 3969 2694 3979 2746
rect 4003 2694 4033 2746
rect 4033 2694 4045 2746
rect 4045 2694 4059 2746
rect 4083 2694 4097 2746
rect 4097 2694 4109 2746
rect 4109 2694 4139 2746
rect 4163 2694 4173 2746
rect 4173 2694 4219 2746
rect 3923 2692 3979 2694
rect 4003 2692 4059 2694
rect 4083 2692 4139 2694
rect 4163 2692 4219 2694
rect 3974 2216 4030 2272
rect 4618 6432 4674 6488
rect 4618 6160 4674 6216
rect 5446 27412 5448 27432
rect 5448 27412 5500 27432
rect 5500 27412 5502 27432
rect 5446 27376 5502 27412
rect 5446 25744 5502 25800
rect 6090 37848 6146 37904
rect 5722 32836 5778 32872
rect 5722 32816 5724 32836
rect 5724 32816 5776 32836
rect 5776 32816 5778 32836
rect 5722 32272 5778 32328
rect 5722 31592 5778 31648
rect 5630 26016 5686 26072
rect 5630 25064 5686 25120
rect 5446 23296 5502 23352
rect 5722 22752 5778 22808
rect 5906 30540 5908 30560
rect 5908 30540 5960 30560
rect 5960 30540 5962 30560
rect 5906 30504 5962 30540
rect 5906 29144 5962 29200
rect 5906 28756 5962 28792
rect 5906 28736 5908 28756
rect 5908 28736 5960 28756
rect 5960 28736 5962 28756
rect 5906 27940 5962 27976
rect 5906 27920 5908 27940
rect 5908 27920 5960 27940
rect 5960 27920 5962 27940
rect 5906 27376 5962 27432
rect 5906 27104 5962 27160
rect 5906 24812 5962 24848
rect 5906 24792 5908 24812
rect 5908 24792 5960 24812
rect 5960 24792 5962 24812
rect 6182 31748 6238 31784
rect 6182 31728 6184 31748
rect 6184 31728 6236 31748
rect 6236 31728 6238 31748
rect 6182 31048 6238 31104
rect 6826 40568 6882 40624
rect 6918 40468 6920 40488
rect 6920 40468 6972 40488
rect 6972 40468 6974 40488
rect 6918 40432 6974 40468
rect 6890 40282 6946 40284
rect 6970 40282 7026 40284
rect 7050 40282 7106 40284
rect 7130 40282 7186 40284
rect 6890 40230 6936 40282
rect 6936 40230 6946 40282
rect 6970 40230 7000 40282
rect 7000 40230 7012 40282
rect 7012 40230 7026 40282
rect 7050 40230 7064 40282
rect 7064 40230 7076 40282
rect 7076 40230 7106 40282
rect 7130 40230 7140 40282
rect 7140 40230 7186 40282
rect 6890 40228 6946 40230
rect 6970 40228 7026 40230
rect 7050 40228 7106 40230
rect 7130 40228 7186 40230
rect 6826 39480 6882 39536
rect 7010 39480 7066 39536
rect 6642 38936 6698 38992
rect 6890 39194 6946 39196
rect 6970 39194 7026 39196
rect 7050 39194 7106 39196
rect 7130 39194 7186 39196
rect 6890 39142 6936 39194
rect 6936 39142 6946 39194
rect 6970 39142 7000 39194
rect 7000 39142 7012 39194
rect 7012 39142 7026 39194
rect 7050 39142 7064 39194
rect 7064 39142 7076 39194
rect 7076 39142 7106 39194
rect 7130 39142 7140 39194
rect 7140 39142 7186 39194
rect 6890 39140 6946 39142
rect 6970 39140 7026 39142
rect 7050 39140 7106 39142
rect 7130 39140 7186 39142
rect 7286 38936 7342 38992
rect 7378 38528 7434 38584
rect 6890 38106 6946 38108
rect 6970 38106 7026 38108
rect 7050 38106 7106 38108
rect 7130 38106 7186 38108
rect 6890 38054 6936 38106
rect 6936 38054 6946 38106
rect 6970 38054 7000 38106
rect 7000 38054 7012 38106
rect 7012 38054 7026 38106
rect 7050 38054 7064 38106
rect 7064 38054 7076 38106
rect 7076 38054 7106 38106
rect 7130 38054 7140 38106
rect 7140 38054 7186 38106
rect 6890 38052 6946 38054
rect 6970 38052 7026 38054
rect 7050 38052 7106 38054
rect 7130 38052 7186 38054
rect 6642 35536 6698 35592
rect 6642 34620 6644 34640
rect 6644 34620 6696 34640
rect 6696 34620 6698 34640
rect 6642 34584 6698 34620
rect 6642 34448 6698 34504
rect 6550 34040 6606 34096
rect 6090 30932 6146 30968
rect 6090 30912 6092 30932
rect 6092 30912 6144 30932
rect 6144 30912 6146 30932
rect 6274 30096 6330 30152
rect 6274 28736 6330 28792
rect 6274 25336 6330 25392
rect 5354 19352 5410 19408
rect 5630 19488 5686 19544
rect 5262 15444 5264 15464
rect 5264 15444 5316 15464
rect 5316 15444 5318 15464
rect 5262 15408 5318 15444
rect 5906 21120 5962 21176
rect 6890 37018 6946 37020
rect 6970 37018 7026 37020
rect 7050 37018 7106 37020
rect 7130 37018 7186 37020
rect 6890 36966 6936 37018
rect 6936 36966 6946 37018
rect 6970 36966 7000 37018
rect 7000 36966 7012 37018
rect 7012 36966 7026 37018
rect 7050 36966 7064 37018
rect 7064 36966 7076 37018
rect 7076 36966 7106 37018
rect 7130 36966 7140 37018
rect 7140 36966 7186 37018
rect 6890 36964 6946 36966
rect 6970 36964 7026 36966
rect 7050 36964 7106 36966
rect 7130 36964 7186 36966
rect 6890 35930 6946 35932
rect 6970 35930 7026 35932
rect 7050 35930 7106 35932
rect 7130 35930 7186 35932
rect 6890 35878 6936 35930
rect 6936 35878 6946 35930
rect 6970 35878 7000 35930
rect 7000 35878 7012 35930
rect 7012 35878 7026 35930
rect 7050 35878 7064 35930
rect 7064 35878 7076 35930
rect 7076 35878 7106 35930
rect 7130 35878 7140 35930
rect 7140 35878 7186 35930
rect 6890 35876 6946 35878
rect 6970 35876 7026 35878
rect 7050 35876 7106 35878
rect 7130 35876 7186 35878
rect 6890 34842 6946 34844
rect 6970 34842 7026 34844
rect 7050 34842 7106 34844
rect 7130 34842 7186 34844
rect 6890 34790 6936 34842
rect 6936 34790 6946 34842
rect 6970 34790 7000 34842
rect 7000 34790 7012 34842
rect 7012 34790 7026 34842
rect 7050 34790 7064 34842
rect 7064 34790 7076 34842
rect 7076 34790 7106 34842
rect 7130 34790 7140 34842
rect 7140 34790 7186 34842
rect 6890 34788 6946 34790
rect 6970 34788 7026 34790
rect 7050 34788 7106 34790
rect 7130 34788 7186 34790
rect 6890 33754 6946 33756
rect 6970 33754 7026 33756
rect 7050 33754 7106 33756
rect 7130 33754 7186 33756
rect 6890 33702 6936 33754
rect 6936 33702 6946 33754
rect 6970 33702 7000 33754
rect 7000 33702 7012 33754
rect 7012 33702 7026 33754
rect 7050 33702 7064 33754
rect 7064 33702 7076 33754
rect 7076 33702 7106 33754
rect 7130 33702 7140 33754
rect 7140 33702 7186 33754
rect 6890 33700 6946 33702
rect 6970 33700 7026 33702
rect 7050 33700 7106 33702
rect 7130 33700 7186 33702
rect 7102 32952 7158 33008
rect 6918 32836 6974 32872
rect 6918 32816 6920 32836
rect 6920 32816 6972 32836
rect 6972 32816 6974 32836
rect 6734 32544 6790 32600
rect 6890 32666 6946 32668
rect 6970 32666 7026 32668
rect 7050 32666 7106 32668
rect 7130 32666 7186 32668
rect 6890 32614 6936 32666
rect 6936 32614 6946 32666
rect 6970 32614 7000 32666
rect 7000 32614 7012 32666
rect 7012 32614 7026 32666
rect 7050 32614 7064 32666
rect 7064 32614 7076 32666
rect 7076 32614 7106 32666
rect 7130 32614 7140 32666
rect 7140 32614 7186 32666
rect 6890 32612 6946 32614
rect 6970 32612 7026 32614
rect 7050 32612 7106 32614
rect 7130 32612 7186 32614
rect 6550 28328 6606 28384
rect 6550 28212 6606 28248
rect 6550 28192 6552 28212
rect 6552 28192 6604 28212
rect 6604 28192 6606 28212
rect 6458 26560 6514 26616
rect 6890 31578 6946 31580
rect 6970 31578 7026 31580
rect 7050 31578 7106 31580
rect 7130 31578 7186 31580
rect 6890 31526 6936 31578
rect 6936 31526 6946 31578
rect 6970 31526 7000 31578
rect 7000 31526 7012 31578
rect 7012 31526 7026 31578
rect 7050 31526 7064 31578
rect 7064 31526 7076 31578
rect 7076 31526 7106 31578
rect 7130 31526 7140 31578
rect 7140 31526 7186 31578
rect 6890 31524 6946 31526
rect 6970 31524 7026 31526
rect 7050 31524 7106 31526
rect 7130 31524 7186 31526
rect 7746 37304 7802 37360
rect 7562 32408 7618 32464
rect 7562 31864 7618 31920
rect 6890 30490 6946 30492
rect 6970 30490 7026 30492
rect 7050 30490 7106 30492
rect 7130 30490 7186 30492
rect 6890 30438 6936 30490
rect 6936 30438 6946 30490
rect 6970 30438 7000 30490
rect 7000 30438 7012 30490
rect 7012 30438 7026 30490
rect 7050 30438 7064 30490
rect 7064 30438 7076 30490
rect 7076 30438 7106 30490
rect 7130 30438 7140 30490
rect 7140 30438 7186 30490
rect 6890 30436 6946 30438
rect 6970 30436 7026 30438
rect 7050 30436 7106 30438
rect 7130 30436 7186 30438
rect 7194 29824 7250 29880
rect 6890 29402 6946 29404
rect 6970 29402 7026 29404
rect 7050 29402 7106 29404
rect 7130 29402 7186 29404
rect 6890 29350 6936 29402
rect 6936 29350 6946 29402
rect 6970 29350 7000 29402
rect 7000 29350 7012 29402
rect 7012 29350 7026 29402
rect 7050 29350 7064 29402
rect 7064 29350 7076 29402
rect 7076 29350 7106 29402
rect 7130 29350 7140 29402
rect 7140 29350 7186 29402
rect 6890 29348 6946 29350
rect 6970 29348 7026 29350
rect 7050 29348 7106 29350
rect 7130 29348 7186 29350
rect 6890 28314 6946 28316
rect 6970 28314 7026 28316
rect 7050 28314 7106 28316
rect 7130 28314 7186 28316
rect 6890 28262 6936 28314
rect 6936 28262 6946 28314
rect 6970 28262 7000 28314
rect 7000 28262 7012 28314
rect 7012 28262 7026 28314
rect 7050 28262 7064 28314
rect 7064 28262 7076 28314
rect 7076 28262 7106 28314
rect 7130 28262 7140 28314
rect 7140 28262 7186 28314
rect 6890 28260 6946 28262
rect 6970 28260 7026 28262
rect 7050 28260 7106 28262
rect 7130 28260 7186 28262
rect 6918 28056 6974 28112
rect 7746 31456 7802 31512
rect 9857 43002 9913 43004
rect 9937 43002 9993 43004
rect 10017 43002 10073 43004
rect 10097 43002 10153 43004
rect 9857 42950 9903 43002
rect 9903 42950 9913 43002
rect 9937 42950 9967 43002
rect 9967 42950 9979 43002
rect 9979 42950 9993 43002
rect 10017 42950 10031 43002
rect 10031 42950 10043 43002
rect 10043 42950 10073 43002
rect 10097 42950 10107 43002
rect 10107 42950 10153 43002
rect 9857 42948 9913 42950
rect 9937 42948 9993 42950
rect 10017 42948 10073 42950
rect 10097 42948 10153 42950
rect 8114 42064 8170 42120
rect 8022 37712 8078 37768
rect 8298 40468 8300 40488
rect 8300 40468 8352 40488
rect 8352 40468 8354 40488
rect 8298 40432 8354 40468
rect 8206 40024 8262 40080
rect 8206 38936 8262 38992
rect 8206 38276 8262 38312
rect 8206 38256 8208 38276
rect 8208 38256 8260 38276
rect 8260 38256 8262 38276
rect 8022 36080 8078 36136
rect 7930 35944 7986 36000
rect 8758 35536 8814 35592
rect 7930 33396 7932 33416
rect 7932 33396 7984 33416
rect 7984 33396 7986 33416
rect 7930 33360 7986 33396
rect 7930 32272 7986 32328
rect 7838 30640 7894 30696
rect 7470 28736 7526 28792
rect 7378 27512 7434 27568
rect 6890 27226 6946 27228
rect 6970 27226 7026 27228
rect 7050 27226 7106 27228
rect 7130 27226 7186 27228
rect 6890 27174 6936 27226
rect 6936 27174 6946 27226
rect 6970 27174 7000 27226
rect 7000 27174 7012 27226
rect 7012 27174 7026 27226
rect 7050 27174 7064 27226
rect 7064 27174 7076 27226
rect 7076 27174 7106 27226
rect 7130 27174 7140 27226
rect 7140 27174 7186 27226
rect 6890 27172 6946 27174
rect 6970 27172 7026 27174
rect 7050 27172 7106 27174
rect 7130 27172 7186 27174
rect 6918 26696 6974 26752
rect 6734 26424 6790 26480
rect 6366 23432 6422 23488
rect 6090 19760 6146 19816
rect 6090 19624 6146 19680
rect 5998 17720 6054 17776
rect 6458 21528 6514 21584
rect 6890 26138 6946 26140
rect 6970 26138 7026 26140
rect 7050 26138 7106 26140
rect 7130 26138 7186 26140
rect 6890 26086 6936 26138
rect 6936 26086 6946 26138
rect 6970 26086 7000 26138
rect 7000 26086 7012 26138
rect 7012 26086 7026 26138
rect 7050 26086 7064 26138
rect 7064 26086 7076 26138
rect 7076 26086 7106 26138
rect 7130 26086 7140 26138
rect 7140 26086 7186 26138
rect 6890 26084 6946 26086
rect 6970 26084 7026 26086
rect 7050 26084 7106 26086
rect 7130 26084 7186 26086
rect 7470 26968 7526 27024
rect 7562 26832 7618 26888
rect 8298 33360 8354 33416
rect 7838 29824 7894 29880
rect 7746 26696 7802 26752
rect 7470 25608 7526 25664
rect 7562 25200 7618 25256
rect 6890 25050 6946 25052
rect 6970 25050 7026 25052
rect 7050 25050 7106 25052
rect 7130 25050 7186 25052
rect 6890 24998 6936 25050
rect 6936 24998 6946 25050
rect 6970 24998 7000 25050
rect 7000 24998 7012 25050
rect 7012 24998 7026 25050
rect 7050 24998 7064 25050
rect 7064 24998 7076 25050
rect 7076 24998 7106 25050
rect 7130 24998 7140 25050
rect 7140 24998 7186 25050
rect 6890 24996 6946 24998
rect 6970 24996 7026 24998
rect 7050 24996 7106 24998
rect 7130 24996 7186 24998
rect 6890 23962 6946 23964
rect 6970 23962 7026 23964
rect 7050 23962 7106 23964
rect 7130 23962 7186 23964
rect 6890 23910 6936 23962
rect 6936 23910 6946 23962
rect 6970 23910 7000 23962
rect 7000 23910 7012 23962
rect 7012 23910 7026 23962
rect 7050 23910 7064 23962
rect 7064 23910 7076 23962
rect 7076 23910 7106 23962
rect 7130 23910 7140 23962
rect 7140 23910 7186 23962
rect 6890 23908 6946 23910
rect 6970 23908 7026 23910
rect 7050 23908 7106 23910
rect 7130 23908 7186 23910
rect 7562 23840 7618 23896
rect 6890 22874 6946 22876
rect 6970 22874 7026 22876
rect 7050 22874 7106 22876
rect 7130 22874 7186 22876
rect 6890 22822 6936 22874
rect 6936 22822 6946 22874
rect 6970 22822 7000 22874
rect 7000 22822 7012 22874
rect 7012 22822 7026 22874
rect 7050 22822 7064 22874
rect 7064 22822 7076 22874
rect 7076 22822 7106 22874
rect 7130 22822 7140 22874
rect 7140 22822 7186 22874
rect 6890 22820 6946 22822
rect 6970 22820 7026 22822
rect 7050 22820 7106 22822
rect 7130 22820 7186 22822
rect 7378 22108 7380 22128
rect 7380 22108 7432 22128
rect 7432 22108 7434 22128
rect 7378 22072 7434 22108
rect 6890 21786 6946 21788
rect 6970 21786 7026 21788
rect 7050 21786 7106 21788
rect 7130 21786 7186 21788
rect 6890 21734 6936 21786
rect 6936 21734 6946 21786
rect 6970 21734 7000 21786
rect 7000 21734 7012 21786
rect 7012 21734 7026 21786
rect 7050 21734 7064 21786
rect 7064 21734 7076 21786
rect 7076 21734 7106 21786
rect 7130 21734 7140 21786
rect 7140 21734 7186 21786
rect 6890 21732 6946 21734
rect 6970 21732 7026 21734
rect 7050 21732 7106 21734
rect 7130 21732 7186 21734
rect 7838 23704 7894 23760
rect 7838 23296 7894 23352
rect 7194 21392 7250 21448
rect 7378 21392 7434 21448
rect 7562 21256 7618 21312
rect 6890 20698 6946 20700
rect 6970 20698 7026 20700
rect 7050 20698 7106 20700
rect 7130 20698 7186 20700
rect 6890 20646 6936 20698
rect 6936 20646 6946 20698
rect 6970 20646 7000 20698
rect 7000 20646 7012 20698
rect 7012 20646 7026 20698
rect 7050 20646 7064 20698
rect 7064 20646 7076 20698
rect 7076 20646 7106 20698
rect 7130 20646 7140 20698
rect 7140 20646 7186 20698
rect 6890 20644 6946 20646
rect 6970 20644 7026 20646
rect 7050 20644 7106 20646
rect 7130 20644 7186 20646
rect 6890 19610 6946 19612
rect 6970 19610 7026 19612
rect 7050 19610 7106 19612
rect 7130 19610 7186 19612
rect 6890 19558 6936 19610
rect 6936 19558 6946 19610
rect 6970 19558 7000 19610
rect 7000 19558 7012 19610
rect 7012 19558 7026 19610
rect 7050 19558 7064 19610
rect 7064 19558 7076 19610
rect 7076 19558 7106 19610
rect 7130 19558 7140 19610
rect 7140 19558 7186 19610
rect 6890 19556 6946 19558
rect 6970 19556 7026 19558
rect 7050 19556 7106 19558
rect 7130 19556 7186 19558
rect 7194 19352 7250 19408
rect 7194 18808 7250 18864
rect 6734 18672 6790 18728
rect 6890 18522 6946 18524
rect 6970 18522 7026 18524
rect 7050 18522 7106 18524
rect 7130 18522 7186 18524
rect 6890 18470 6936 18522
rect 6936 18470 6946 18522
rect 6970 18470 7000 18522
rect 7000 18470 7012 18522
rect 7012 18470 7026 18522
rect 7050 18470 7064 18522
rect 7064 18470 7076 18522
rect 7076 18470 7106 18522
rect 7130 18470 7140 18522
rect 7140 18470 7186 18522
rect 6890 18468 6946 18470
rect 6970 18468 7026 18470
rect 7050 18468 7106 18470
rect 7130 18468 7186 18470
rect 5446 13912 5502 13968
rect 5538 12688 5594 12744
rect 5170 12300 5226 12336
rect 5170 12280 5172 12300
rect 5172 12280 5224 12300
rect 5224 12280 5226 12300
rect 5170 9580 5226 9616
rect 5170 9560 5172 9580
rect 5172 9560 5224 9580
rect 5224 9560 5226 9580
rect 5906 12180 5908 12200
rect 5908 12180 5960 12200
rect 5960 12180 5962 12200
rect 5906 12144 5962 12180
rect 5538 9560 5594 9616
rect 4618 3984 4674 4040
rect 4342 2896 4398 2952
rect 4802 2760 4858 2816
rect 4434 2352 4490 2408
rect 3923 1658 3979 1660
rect 4003 1658 4059 1660
rect 4083 1658 4139 1660
rect 4163 1658 4219 1660
rect 3923 1606 3969 1658
rect 3969 1606 3979 1658
rect 4003 1606 4033 1658
rect 4033 1606 4045 1658
rect 4045 1606 4059 1658
rect 4083 1606 4097 1658
rect 4097 1606 4109 1658
rect 4109 1606 4139 1658
rect 4163 1606 4173 1658
rect 4173 1606 4219 1658
rect 3923 1604 3979 1606
rect 4003 1604 4059 1606
rect 4083 1604 4139 1606
rect 4163 1604 4219 1606
rect 4434 1672 4490 1728
rect 4434 1300 4436 1320
rect 4436 1300 4488 1320
rect 4488 1300 4490 1320
rect 4434 1264 4490 1300
rect 4802 1536 4858 1592
rect 5906 9152 5962 9208
rect 5262 6160 5318 6216
rect 5446 6296 5502 6352
rect 6890 17434 6946 17436
rect 6970 17434 7026 17436
rect 7050 17434 7106 17436
rect 7130 17434 7186 17436
rect 6890 17382 6936 17434
rect 6936 17382 6946 17434
rect 6970 17382 7000 17434
rect 7000 17382 7012 17434
rect 7012 17382 7026 17434
rect 7050 17382 7064 17434
rect 7064 17382 7076 17434
rect 7076 17382 7106 17434
rect 7130 17382 7140 17434
rect 7140 17382 7186 17434
rect 6890 17380 6946 17382
rect 6970 17380 7026 17382
rect 7050 17380 7106 17382
rect 7130 17380 7186 17382
rect 6890 16346 6946 16348
rect 6970 16346 7026 16348
rect 7050 16346 7106 16348
rect 7130 16346 7186 16348
rect 6890 16294 6936 16346
rect 6936 16294 6946 16346
rect 6970 16294 7000 16346
rect 7000 16294 7012 16346
rect 7012 16294 7026 16346
rect 7050 16294 7064 16346
rect 7064 16294 7076 16346
rect 7076 16294 7106 16346
rect 7130 16294 7140 16346
rect 7140 16294 7186 16346
rect 6890 16292 6946 16294
rect 6970 16292 7026 16294
rect 7050 16292 7106 16294
rect 7130 16292 7186 16294
rect 6826 15564 6882 15600
rect 6826 15544 6828 15564
rect 6828 15544 6880 15564
rect 6880 15544 6882 15564
rect 6642 15308 6644 15328
rect 6644 15308 6696 15328
rect 6696 15308 6698 15328
rect 6642 15272 6698 15308
rect 6890 15258 6946 15260
rect 6970 15258 7026 15260
rect 7050 15258 7106 15260
rect 7130 15258 7186 15260
rect 6890 15206 6936 15258
rect 6936 15206 6946 15258
rect 6970 15206 7000 15258
rect 7000 15206 7012 15258
rect 7012 15206 7026 15258
rect 7050 15206 7064 15258
rect 7064 15206 7076 15258
rect 7076 15206 7106 15258
rect 7130 15206 7140 15258
rect 7140 15206 7186 15258
rect 6890 15204 6946 15206
rect 6970 15204 7026 15206
rect 7050 15204 7106 15206
rect 7130 15204 7186 15206
rect 8114 29824 8170 29880
rect 8206 27648 8262 27704
rect 8114 26152 8170 26208
rect 6890 14170 6946 14172
rect 6970 14170 7026 14172
rect 7050 14170 7106 14172
rect 7130 14170 7186 14172
rect 6890 14118 6936 14170
rect 6936 14118 6946 14170
rect 6970 14118 7000 14170
rect 7000 14118 7012 14170
rect 7012 14118 7026 14170
rect 7050 14118 7064 14170
rect 7064 14118 7076 14170
rect 7076 14118 7106 14170
rect 7130 14118 7140 14170
rect 7140 14118 7186 14170
rect 6890 14116 6946 14118
rect 6970 14116 7026 14118
rect 7050 14116 7106 14118
rect 7130 14116 7186 14118
rect 6642 12316 6644 12336
rect 6644 12316 6696 12336
rect 6696 12316 6698 12336
rect 6642 12280 6698 12316
rect 6890 13082 6946 13084
rect 6970 13082 7026 13084
rect 7050 13082 7106 13084
rect 7130 13082 7186 13084
rect 6890 13030 6936 13082
rect 6936 13030 6946 13082
rect 6970 13030 7000 13082
rect 7000 13030 7012 13082
rect 7012 13030 7026 13082
rect 7050 13030 7064 13082
rect 7064 13030 7076 13082
rect 7076 13030 7106 13082
rect 7130 13030 7140 13082
rect 7140 13030 7186 13082
rect 6890 13028 6946 13030
rect 6970 13028 7026 13030
rect 7050 13028 7106 13030
rect 7130 13028 7186 13030
rect 6890 11994 6946 11996
rect 6970 11994 7026 11996
rect 7050 11994 7106 11996
rect 7130 11994 7186 11996
rect 6890 11942 6936 11994
rect 6936 11942 6946 11994
rect 6970 11942 7000 11994
rect 7000 11942 7012 11994
rect 7012 11942 7026 11994
rect 7050 11942 7064 11994
rect 7064 11942 7076 11994
rect 7076 11942 7106 11994
rect 7130 11942 7140 11994
rect 7140 11942 7186 11994
rect 6890 11940 6946 11942
rect 6970 11940 7026 11942
rect 7050 11940 7106 11942
rect 7130 11940 7186 11942
rect 6890 10906 6946 10908
rect 6970 10906 7026 10908
rect 7050 10906 7106 10908
rect 7130 10906 7186 10908
rect 6890 10854 6936 10906
rect 6936 10854 6946 10906
rect 6970 10854 7000 10906
rect 7000 10854 7012 10906
rect 7012 10854 7026 10906
rect 7050 10854 7064 10906
rect 7064 10854 7076 10906
rect 7076 10854 7106 10906
rect 7130 10854 7140 10906
rect 7140 10854 7186 10906
rect 6890 10852 6946 10854
rect 6970 10852 7026 10854
rect 7050 10852 7106 10854
rect 7130 10852 7186 10854
rect 7378 12824 7434 12880
rect 7470 12688 7526 12744
rect 7746 13640 7802 13696
rect 6826 10648 6882 10704
rect 7194 10512 7250 10568
rect 6918 10260 6974 10296
rect 6918 10240 6920 10260
rect 6920 10240 6972 10260
rect 6972 10240 6974 10260
rect 6890 9818 6946 9820
rect 6970 9818 7026 9820
rect 7050 9818 7106 9820
rect 7130 9818 7186 9820
rect 6890 9766 6936 9818
rect 6936 9766 6946 9818
rect 6970 9766 7000 9818
rect 7000 9766 7012 9818
rect 7012 9766 7026 9818
rect 7050 9766 7064 9818
rect 7064 9766 7076 9818
rect 7076 9766 7106 9818
rect 7130 9766 7140 9818
rect 7140 9766 7186 9818
rect 6890 9764 6946 9766
rect 6970 9764 7026 9766
rect 7050 9764 7106 9766
rect 7130 9764 7186 9766
rect 6918 9036 6974 9072
rect 6918 9016 6920 9036
rect 6920 9016 6972 9036
rect 6972 9016 6974 9036
rect 6890 8730 6946 8732
rect 6970 8730 7026 8732
rect 7050 8730 7106 8732
rect 7130 8730 7186 8732
rect 6890 8678 6936 8730
rect 6936 8678 6946 8730
rect 6970 8678 7000 8730
rect 7000 8678 7012 8730
rect 7012 8678 7026 8730
rect 7050 8678 7064 8730
rect 7064 8678 7076 8730
rect 7076 8678 7106 8730
rect 7130 8678 7140 8730
rect 7140 8678 7186 8730
rect 6890 8676 6946 8678
rect 6970 8676 7026 8678
rect 7050 8676 7106 8678
rect 7130 8676 7186 8678
rect 7378 9152 7434 9208
rect 7654 10512 7710 10568
rect 7562 10240 7618 10296
rect 6550 8336 6606 8392
rect 6890 7642 6946 7644
rect 6970 7642 7026 7644
rect 7050 7642 7106 7644
rect 7130 7642 7186 7644
rect 6890 7590 6936 7642
rect 6936 7590 6946 7642
rect 6970 7590 7000 7642
rect 7000 7590 7012 7642
rect 7012 7590 7026 7642
rect 7050 7590 7064 7642
rect 7064 7590 7076 7642
rect 7076 7590 7106 7642
rect 7130 7590 7140 7642
rect 7140 7590 7186 7642
rect 6890 7588 6946 7590
rect 6970 7588 7026 7590
rect 7050 7588 7106 7590
rect 7130 7588 7186 7590
rect 7470 9016 7526 9072
rect 7654 8508 7656 8528
rect 7656 8508 7708 8528
rect 7708 8508 7710 8528
rect 7654 8472 7710 8508
rect 7470 7792 7526 7848
rect 6734 6840 6790 6896
rect 5538 3304 5594 3360
rect 6890 6554 6946 6556
rect 6970 6554 7026 6556
rect 7050 6554 7106 6556
rect 7130 6554 7186 6556
rect 6890 6502 6936 6554
rect 6936 6502 6946 6554
rect 6970 6502 7000 6554
rect 7000 6502 7012 6554
rect 7012 6502 7026 6554
rect 7050 6502 7064 6554
rect 7064 6502 7076 6554
rect 7076 6502 7106 6554
rect 7130 6502 7140 6554
rect 7140 6502 7186 6554
rect 6890 6500 6946 6502
rect 6970 6500 7026 6502
rect 7050 6500 7106 6502
rect 7130 6500 7186 6502
rect 6890 5466 6946 5468
rect 6970 5466 7026 5468
rect 7050 5466 7106 5468
rect 7130 5466 7186 5468
rect 6890 5414 6936 5466
rect 6936 5414 6946 5466
rect 6970 5414 7000 5466
rect 7000 5414 7012 5466
rect 7012 5414 7026 5466
rect 7050 5414 7064 5466
rect 7064 5414 7076 5466
rect 7076 5414 7106 5466
rect 7130 5414 7140 5466
rect 7140 5414 7186 5466
rect 6890 5412 6946 5414
rect 6970 5412 7026 5414
rect 7050 5412 7106 5414
rect 7130 5412 7186 5414
rect 6890 4378 6946 4380
rect 6970 4378 7026 4380
rect 7050 4378 7106 4380
rect 7130 4378 7186 4380
rect 6890 4326 6936 4378
rect 6936 4326 6946 4378
rect 6970 4326 7000 4378
rect 7000 4326 7012 4378
rect 7012 4326 7026 4378
rect 7050 4326 7064 4378
rect 7064 4326 7076 4378
rect 7076 4326 7106 4378
rect 7130 4326 7140 4378
rect 7140 4326 7186 4378
rect 6890 4324 6946 4326
rect 6970 4324 7026 4326
rect 7050 4324 7106 4326
rect 7130 4324 7186 4326
rect 6890 3290 6946 3292
rect 6970 3290 7026 3292
rect 7050 3290 7106 3292
rect 7130 3290 7186 3292
rect 6890 3238 6936 3290
rect 6936 3238 6946 3290
rect 6970 3238 7000 3290
rect 7000 3238 7012 3290
rect 7012 3238 7026 3290
rect 7050 3238 7064 3290
rect 7064 3238 7076 3290
rect 7076 3238 7106 3290
rect 7130 3238 7140 3290
rect 7140 3238 7186 3290
rect 6890 3236 6946 3238
rect 6970 3236 7026 3238
rect 7050 3236 7106 3238
rect 7130 3236 7186 3238
rect 5906 2760 5962 2816
rect 5722 2488 5778 2544
rect 5538 1944 5594 2000
rect 5998 1944 6054 2000
rect 6090 720 6146 776
rect 6890 2202 6946 2204
rect 6970 2202 7026 2204
rect 7050 2202 7106 2204
rect 7130 2202 7186 2204
rect 6890 2150 6936 2202
rect 6936 2150 6946 2202
rect 6970 2150 7000 2202
rect 7000 2150 7012 2202
rect 7012 2150 7026 2202
rect 7050 2150 7064 2202
rect 7064 2150 7076 2202
rect 7076 2150 7106 2202
rect 7130 2150 7140 2202
rect 7140 2150 7186 2202
rect 6890 2148 6946 2150
rect 6970 2148 7026 2150
rect 7050 2148 7106 2150
rect 7130 2148 7186 2150
rect 7010 1944 7066 2000
rect 6918 1536 6974 1592
rect 6918 1264 6974 1320
rect 6890 1114 6946 1116
rect 6970 1114 7026 1116
rect 7050 1114 7106 1116
rect 7130 1114 7186 1116
rect 6890 1062 6936 1114
rect 6936 1062 6946 1114
rect 6970 1062 7000 1114
rect 7000 1062 7012 1114
rect 7012 1062 7026 1114
rect 7050 1062 7064 1114
rect 7064 1062 7076 1114
rect 7076 1062 7106 1114
rect 7130 1062 7140 1114
rect 7140 1062 7186 1114
rect 6890 1060 6946 1062
rect 6970 1060 7026 1062
rect 7050 1060 7106 1062
rect 7130 1060 7186 1062
rect 7654 3984 7710 4040
rect 8298 25336 8354 25392
rect 8390 21548 8446 21584
rect 8390 21528 8392 21548
rect 8392 21528 8444 21548
rect 8444 21528 8446 21548
rect 8206 20848 8262 20904
rect 8390 20848 8446 20904
rect 8298 18944 8354 19000
rect 7930 8336 7986 8392
rect 8390 9052 8392 9072
rect 8392 9052 8444 9072
rect 8444 9052 8446 9072
rect 8390 9016 8446 9052
rect 10414 42880 10470 42936
rect 9126 41112 9182 41168
rect 9402 41420 9404 41440
rect 9404 41420 9456 41440
rect 9456 41420 9458 41440
rect 9402 41384 9458 41420
rect 9857 41914 9913 41916
rect 9937 41914 9993 41916
rect 10017 41914 10073 41916
rect 10097 41914 10153 41916
rect 9857 41862 9903 41914
rect 9903 41862 9913 41914
rect 9937 41862 9967 41914
rect 9967 41862 9979 41914
rect 9979 41862 9993 41914
rect 10017 41862 10031 41914
rect 10031 41862 10043 41914
rect 10043 41862 10073 41914
rect 10097 41862 10107 41914
rect 10107 41862 10153 41914
rect 9857 41860 9913 41862
rect 9937 41860 9993 41862
rect 10017 41860 10073 41862
rect 10097 41860 10153 41862
rect 10230 41112 10286 41168
rect 9857 40826 9913 40828
rect 9937 40826 9993 40828
rect 10017 40826 10073 40828
rect 10097 40826 10153 40828
rect 9857 40774 9903 40826
rect 9903 40774 9913 40826
rect 9937 40774 9967 40826
rect 9967 40774 9979 40826
rect 9979 40774 9993 40826
rect 10017 40774 10031 40826
rect 10031 40774 10043 40826
rect 10043 40774 10073 40826
rect 10097 40774 10107 40826
rect 10107 40774 10153 40826
rect 9857 40772 9913 40774
rect 9937 40772 9993 40774
rect 10017 40772 10073 40774
rect 10097 40772 10153 40774
rect 9678 40024 9734 40080
rect 10230 40432 10286 40488
rect 10322 40296 10378 40352
rect 10230 40024 10286 40080
rect 9402 39480 9458 39536
rect 9857 39738 9913 39740
rect 9937 39738 9993 39740
rect 10017 39738 10073 39740
rect 10097 39738 10153 39740
rect 9857 39686 9903 39738
rect 9903 39686 9913 39738
rect 9937 39686 9967 39738
rect 9967 39686 9979 39738
rect 9979 39686 9993 39738
rect 10017 39686 10031 39738
rect 10031 39686 10043 39738
rect 10043 39686 10073 39738
rect 10097 39686 10107 39738
rect 10107 39686 10153 39738
rect 9857 39684 9913 39686
rect 9937 39684 9993 39686
rect 10017 39684 10073 39686
rect 10097 39684 10153 39686
rect 9857 38650 9913 38652
rect 9937 38650 9993 38652
rect 10017 38650 10073 38652
rect 10097 38650 10153 38652
rect 9857 38598 9903 38650
rect 9903 38598 9913 38650
rect 9937 38598 9967 38650
rect 9967 38598 9979 38650
rect 9979 38598 9993 38650
rect 10017 38598 10031 38650
rect 10031 38598 10043 38650
rect 10043 38598 10073 38650
rect 10097 38598 10107 38650
rect 10107 38598 10153 38650
rect 9857 38596 9913 38598
rect 9937 38596 9993 38598
rect 10017 38596 10073 38598
rect 10097 38596 10153 38598
rect 8850 34448 8906 34504
rect 8666 32816 8722 32872
rect 8666 31184 8722 31240
rect 8666 28872 8722 28928
rect 8574 27784 8630 27840
rect 8666 23296 8722 23352
rect 8574 21936 8630 21992
rect 8850 31456 8906 31512
rect 9126 33940 9128 33960
rect 9128 33940 9180 33960
rect 9180 33940 9182 33960
rect 9126 33904 9182 33940
rect 9218 33496 9274 33552
rect 9857 37562 9913 37564
rect 9937 37562 9993 37564
rect 10017 37562 10073 37564
rect 10097 37562 10153 37564
rect 9857 37510 9903 37562
rect 9903 37510 9913 37562
rect 9937 37510 9967 37562
rect 9967 37510 9979 37562
rect 9979 37510 9993 37562
rect 10017 37510 10031 37562
rect 10031 37510 10043 37562
rect 10043 37510 10073 37562
rect 10097 37510 10107 37562
rect 10107 37510 10153 37562
rect 9857 37508 9913 37510
rect 9937 37508 9993 37510
rect 10017 37508 10073 37510
rect 10097 37508 10153 37510
rect 9857 36474 9913 36476
rect 9937 36474 9993 36476
rect 10017 36474 10073 36476
rect 10097 36474 10153 36476
rect 9857 36422 9903 36474
rect 9903 36422 9913 36474
rect 9937 36422 9967 36474
rect 9967 36422 9979 36474
rect 9979 36422 9993 36474
rect 10017 36422 10031 36474
rect 10031 36422 10043 36474
rect 10043 36422 10073 36474
rect 10097 36422 10107 36474
rect 10107 36422 10153 36474
rect 9857 36420 9913 36422
rect 9937 36420 9993 36422
rect 10017 36420 10073 36422
rect 10097 36420 10153 36422
rect 10046 35944 10102 36000
rect 10690 40024 10746 40080
rect 9857 35386 9913 35388
rect 9937 35386 9993 35388
rect 10017 35386 10073 35388
rect 10097 35386 10153 35388
rect 9857 35334 9903 35386
rect 9903 35334 9913 35386
rect 9937 35334 9967 35386
rect 9967 35334 9979 35386
rect 9979 35334 9993 35386
rect 10017 35334 10031 35386
rect 10031 35334 10043 35386
rect 10043 35334 10073 35386
rect 10097 35334 10107 35386
rect 10107 35334 10153 35386
rect 9857 35332 9913 35334
rect 9937 35332 9993 35334
rect 10017 35332 10073 35334
rect 10097 35332 10153 35334
rect 9494 34448 9550 34504
rect 9402 33804 9404 33824
rect 9404 33804 9456 33824
rect 9456 33804 9458 33824
rect 9402 33768 9458 33804
rect 9857 34298 9913 34300
rect 9937 34298 9993 34300
rect 10017 34298 10073 34300
rect 10097 34298 10153 34300
rect 9857 34246 9903 34298
rect 9903 34246 9913 34298
rect 9937 34246 9967 34298
rect 9967 34246 9979 34298
rect 9979 34246 9993 34298
rect 10017 34246 10031 34298
rect 10031 34246 10043 34298
rect 10043 34246 10073 34298
rect 10097 34246 10107 34298
rect 10107 34246 10153 34298
rect 9857 34244 9913 34246
rect 9937 34244 9993 34246
rect 10017 34244 10073 34246
rect 10097 34244 10153 34246
rect 9770 33768 9826 33824
rect 9586 33224 9642 33280
rect 9494 32408 9550 32464
rect 9770 33632 9826 33688
rect 9954 33768 10010 33824
rect 9954 33360 10010 33416
rect 9034 31320 9090 31376
rect 9034 30776 9090 30832
rect 8850 29552 8906 29608
rect 9034 30268 9036 30288
rect 9036 30268 9088 30288
rect 9088 30268 9090 30288
rect 9034 30232 9090 30268
rect 9218 29552 9274 29608
rect 8942 24928 8998 24984
rect 9586 32000 9642 32056
rect 9494 30232 9550 30288
rect 9857 33210 9913 33212
rect 9937 33210 9993 33212
rect 10017 33210 10073 33212
rect 10097 33210 10153 33212
rect 9857 33158 9903 33210
rect 9903 33158 9913 33210
rect 9937 33158 9967 33210
rect 9967 33158 9979 33210
rect 9979 33158 9993 33210
rect 10017 33158 10031 33210
rect 10031 33158 10043 33210
rect 10043 33158 10073 33210
rect 10097 33158 10107 33210
rect 10107 33158 10153 33210
rect 9857 33156 9913 33158
rect 9937 33156 9993 33158
rect 10017 33156 10073 33158
rect 10097 33156 10153 33158
rect 10046 32952 10102 33008
rect 10322 35128 10378 35184
rect 10506 33904 10562 33960
rect 10598 33768 10654 33824
rect 9857 32122 9913 32124
rect 9937 32122 9993 32124
rect 10017 32122 10073 32124
rect 10097 32122 10153 32124
rect 9857 32070 9903 32122
rect 9903 32070 9913 32122
rect 9937 32070 9967 32122
rect 9967 32070 9979 32122
rect 9979 32070 9993 32122
rect 10017 32070 10031 32122
rect 10031 32070 10043 32122
rect 10043 32070 10073 32122
rect 10097 32070 10107 32122
rect 10107 32070 10153 32122
rect 9857 32068 9913 32070
rect 9937 32068 9993 32070
rect 10017 32068 10073 32070
rect 10097 32068 10153 32070
rect 10506 32952 10562 33008
rect 11334 38664 11390 38720
rect 11334 34584 11390 34640
rect 10782 33632 10838 33688
rect 9857 31034 9913 31036
rect 9937 31034 9993 31036
rect 10017 31034 10073 31036
rect 10097 31034 10153 31036
rect 9857 30982 9903 31034
rect 9903 30982 9913 31034
rect 9937 30982 9967 31034
rect 9967 30982 9979 31034
rect 9979 30982 9993 31034
rect 10017 30982 10031 31034
rect 10031 30982 10043 31034
rect 10043 30982 10073 31034
rect 10097 30982 10107 31034
rect 10107 30982 10153 31034
rect 9857 30980 9913 30982
rect 9937 30980 9993 30982
rect 10017 30980 10073 30982
rect 10097 30980 10153 30982
rect 9954 30368 10010 30424
rect 10046 30232 10102 30288
rect 9857 29946 9913 29948
rect 9937 29946 9993 29948
rect 10017 29946 10073 29948
rect 10097 29946 10153 29948
rect 9857 29894 9903 29946
rect 9903 29894 9913 29946
rect 9937 29894 9967 29946
rect 9967 29894 9979 29946
rect 9979 29894 9993 29946
rect 10017 29894 10031 29946
rect 10031 29894 10043 29946
rect 10043 29894 10073 29946
rect 10097 29894 10107 29946
rect 10107 29894 10153 29946
rect 9857 29892 9913 29894
rect 9937 29892 9993 29894
rect 10017 29892 10073 29894
rect 10097 29892 10153 29894
rect 10414 29960 10470 30016
rect 9586 29174 9642 29200
rect 9586 29144 9588 29174
rect 9588 29144 9640 29174
rect 9640 29144 9642 29174
rect 9857 28858 9913 28860
rect 9937 28858 9993 28860
rect 10017 28858 10073 28860
rect 10097 28858 10153 28860
rect 9857 28806 9903 28858
rect 9903 28806 9913 28858
rect 9937 28806 9967 28858
rect 9967 28806 9979 28858
rect 9979 28806 9993 28858
rect 10017 28806 10031 28858
rect 10031 28806 10043 28858
rect 10043 28806 10073 28858
rect 10097 28806 10107 28858
rect 10107 28806 10153 28858
rect 9857 28804 9913 28806
rect 9937 28804 9993 28806
rect 10017 28804 10073 28806
rect 10097 28804 10153 28806
rect 9678 28736 9734 28792
rect 9402 24928 9458 24984
rect 9310 23432 9366 23488
rect 8942 20440 8998 20496
rect 9034 20032 9090 20088
rect 8850 19352 8906 19408
rect 9310 21392 9366 21448
rect 9310 21120 9366 21176
rect 8758 19216 8814 19272
rect 8666 18672 8722 18728
rect 8574 13640 8630 13696
rect 8574 6160 8630 6216
rect 9857 27770 9913 27772
rect 9937 27770 9993 27772
rect 10017 27770 10073 27772
rect 10097 27770 10153 27772
rect 9857 27718 9903 27770
rect 9903 27718 9913 27770
rect 9937 27718 9967 27770
rect 9967 27718 9979 27770
rect 9979 27718 9993 27770
rect 10017 27718 10031 27770
rect 10031 27718 10043 27770
rect 10043 27718 10073 27770
rect 10097 27718 10107 27770
rect 10107 27718 10153 27770
rect 9857 27716 9913 27718
rect 9937 27716 9993 27718
rect 10017 27716 10073 27718
rect 10097 27716 10153 27718
rect 10598 28464 10654 28520
rect 10598 27784 10654 27840
rect 10506 27512 10562 27568
rect 9857 26682 9913 26684
rect 9937 26682 9993 26684
rect 10017 26682 10073 26684
rect 10097 26682 10153 26684
rect 9857 26630 9903 26682
rect 9903 26630 9913 26682
rect 9937 26630 9967 26682
rect 9967 26630 9979 26682
rect 9979 26630 9993 26682
rect 10017 26630 10031 26682
rect 10031 26630 10043 26682
rect 10043 26630 10073 26682
rect 10097 26630 10107 26682
rect 10107 26630 10153 26682
rect 9857 26628 9913 26630
rect 9937 26628 9993 26630
rect 10017 26628 10073 26630
rect 10097 26628 10153 26630
rect 9770 26152 9826 26208
rect 9857 25594 9913 25596
rect 9937 25594 9993 25596
rect 10017 25594 10073 25596
rect 10097 25594 10153 25596
rect 9857 25542 9903 25594
rect 9903 25542 9913 25594
rect 9937 25542 9967 25594
rect 9967 25542 9979 25594
rect 9979 25542 9993 25594
rect 10017 25542 10031 25594
rect 10031 25542 10043 25594
rect 10043 25542 10073 25594
rect 10097 25542 10107 25594
rect 10107 25542 10153 25594
rect 9857 25540 9913 25542
rect 9937 25540 9993 25542
rect 10017 25540 10073 25542
rect 10097 25540 10153 25542
rect 9857 24506 9913 24508
rect 9937 24506 9993 24508
rect 10017 24506 10073 24508
rect 10097 24506 10153 24508
rect 9857 24454 9903 24506
rect 9903 24454 9913 24506
rect 9937 24454 9967 24506
rect 9967 24454 9979 24506
rect 9979 24454 9993 24506
rect 10017 24454 10031 24506
rect 10031 24454 10043 24506
rect 10043 24454 10073 24506
rect 10097 24454 10107 24506
rect 10107 24454 10153 24506
rect 9857 24452 9913 24454
rect 9937 24452 9993 24454
rect 10017 24452 10073 24454
rect 10097 24452 10153 24454
rect 10230 23432 10286 23488
rect 9857 23418 9913 23420
rect 9937 23418 9993 23420
rect 10017 23418 10073 23420
rect 10097 23418 10153 23420
rect 9857 23366 9903 23418
rect 9903 23366 9913 23418
rect 9937 23366 9967 23418
rect 9967 23366 9979 23418
rect 9979 23366 9993 23418
rect 10017 23366 10031 23418
rect 10031 23366 10043 23418
rect 10043 23366 10073 23418
rect 10097 23366 10107 23418
rect 10107 23366 10153 23418
rect 9857 23364 9913 23366
rect 9937 23364 9993 23366
rect 10017 23364 10073 23366
rect 10097 23364 10153 23366
rect 10138 22752 10194 22808
rect 9494 19624 9550 19680
rect 9857 22330 9913 22332
rect 9937 22330 9993 22332
rect 10017 22330 10073 22332
rect 10097 22330 10153 22332
rect 9857 22278 9903 22330
rect 9903 22278 9913 22330
rect 9937 22278 9967 22330
rect 9967 22278 9979 22330
rect 9979 22278 9993 22330
rect 10017 22278 10031 22330
rect 10031 22278 10043 22330
rect 10043 22278 10073 22330
rect 10097 22278 10107 22330
rect 10107 22278 10153 22330
rect 9857 22276 9913 22278
rect 9937 22276 9993 22278
rect 10017 22276 10073 22278
rect 10097 22276 10153 22278
rect 9857 21242 9913 21244
rect 9937 21242 9993 21244
rect 10017 21242 10073 21244
rect 10097 21242 10153 21244
rect 9857 21190 9903 21242
rect 9903 21190 9913 21242
rect 9937 21190 9967 21242
rect 9967 21190 9979 21242
rect 9979 21190 9993 21242
rect 10017 21190 10031 21242
rect 10031 21190 10043 21242
rect 10043 21190 10073 21242
rect 10097 21190 10107 21242
rect 10107 21190 10153 21242
rect 9857 21188 9913 21190
rect 9937 21188 9993 21190
rect 10017 21188 10073 21190
rect 10097 21188 10153 21190
rect 10506 24520 10562 24576
rect 10506 24384 10562 24440
rect 10414 22344 10470 22400
rect 9857 20154 9913 20156
rect 9937 20154 9993 20156
rect 10017 20154 10073 20156
rect 10097 20154 10153 20156
rect 9857 20102 9903 20154
rect 9903 20102 9913 20154
rect 9937 20102 9967 20154
rect 9967 20102 9979 20154
rect 9979 20102 9993 20154
rect 10017 20102 10031 20154
rect 10031 20102 10043 20154
rect 10043 20102 10073 20154
rect 10097 20102 10107 20154
rect 10107 20102 10153 20154
rect 9857 20100 9913 20102
rect 9937 20100 9993 20102
rect 10017 20100 10073 20102
rect 10097 20100 10153 20102
rect 9678 17584 9734 17640
rect 9678 17040 9734 17096
rect 9954 19896 10010 19952
rect 10414 20304 10470 20360
rect 9857 19066 9913 19068
rect 9937 19066 9993 19068
rect 10017 19066 10073 19068
rect 10097 19066 10153 19068
rect 9857 19014 9903 19066
rect 9903 19014 9913 19066
rect 9937 19014 9967 19066
rect 9967 19014 9979 19066
rect 9979 19014 9993 19066
rect 10017 19014 10031 19066
rect 10031 19014 10043 19066
rect 10043 19014 10073 19066
rect 10097 19014 10107 19066
rect 10107 19014 10153 19066
rect 9857 19012 9913 19014
rect 9937 19012 9993 19014
rect 10017 19012 10073 19014
rect 10097 19012 10153 19014
rect 10322 19760 10378 19816
rect 9857 17978 9913 17980
rect 9937 17978 9993 17980
rect 10017 17978 10073 17980
rect 10097 17978 10153 17980
rect 9857 17926 9903 17978
rect 9903 17926 9913 17978
rect 9937 17926 9967 17978
rect 9967 17926 9979 17978
rect 9979 17926 9993 17978
rect 10017 17926 10031 17978
rect 10031 17926 10043 17978
rect 10043 17926 10073 17978
rect 10097 17926 10107 17978
rect 10107 17926 10153 17978
rect 9857 17924 9913 17926
rect 9937 17924 9993 17926
rect 10017 17924 10073 17926
rect 10097 17924 10153 17926
rect 10322 17584 10378 17640
rect 9857 16890 9913 16892
rect 9937 16890 9993 16892
rect 10017 16890 10073 16892
rect 10097 16890 10153 16892
rect 9857 16838 9903 16890
rect 9903 16838 9913 16890
rect 9937 16838 9967 16890
rect 9967 16838 9979 16890
rect 9979 16838 9993 16890
rect 10017 16838 10031 16890
rect 10031 16838 10043 16890
rect 10043 16838 10073 16890
rect 10097 16838 10107 16890
rect 10107 16838 10153 16890
rect 9857 16836 9913 16838
rect 9937 16836 9993 16838
rect 10017 16836 10073 16838
rect 10097 16836 10153 16838
rect 9857 15802 9913 15804
rect 9937 15802 9993 15804
rect 10017 15802 10073 15804
rect 10097 15802 10153 15804
rect 9857 15750 9903 15802
rect 9903 15750 9913 15802
rect 9937 15750 9967 15802
rect 9967 15750 9979 15802
rect 9979 15750 9993 15802
rect 10017 15750 10031 15802
rect 10031 15750 10043 15802
rect 10043 15750 10073 15802
rect 10097 15750 10107 15802
rect 10107 15750 10153 15802
rect 9857 15748 9913 15750
rect 9937 15748 9993 15750
rect 10017 15748 10073 15750
rect 10097 15748 10153 15750
rect 9857 14714 9913 14716
rect 9937 14714 9993 14716
rect 10017 14714 10073 14716
rect 10097 14714 10153 14716
rect 9857 14662 9903 14714
rect 9903 14662 9913 14714
rect 9937 14662 9967 14714
rect 9967 14662 9979 14714
rect 9979 14662 9993 14714
rect 10017 14662 10031 14714
rect 10031 14662 10043 14714
rect 10043 14662 10073 14714
rect 10097 14662 10107 14714
rect 10107 14662 10153 14714
rect 9857 14660 9913 14662
rect 9937 14660 9993 14662
rect 10017 14660 10073 14662
rect 10097 14660 10153 14662
rect 11242 32408 11298 32464
rect 11242 31728 11298 31784
rect 11058 28056 11114 28112
rect 11058 25336 11114 25392
rect 11334 24792 11390 24848
rect 11150 22652 11152 22672
rect 11152 22652 11204 22672
rect 11204 22652 11206 22672
rect 11150 22616 11206 22652
rect 10690 20304 10746 20360
rect 10690 18128 10746 18184
rect 10690 16496 10746 16552
rect 9857 13626 9913 13628
rect 9937 13626 9993 13628
rect 10017 13626 10073 13628
rect 10097 13626 10153 13628
rect 9857 13574 9903 13626
rect 9903 13574 9913 13626
rect 9937 13574 9967 13626
rect 9967 13574 9979 13626
rect 9979 13574 9993 13626
rect 10017 13574 10031 13626
rect 10031 13574 10043 13626
rect 10043 13574 10073 13626
rect 10097 13574 10107 13626
rect 10107 13574 10153 13626
rect 9857 13572 9913 13574
rect 9937 13572 9993 13574
rect 10017 13572 10073 13574
rect 10097 13572 10153 13574
rect 10322 13368 10378 13424
rect 9126 10512 9182 10568
rect 9402 9424 9458 9480
rect 9034 6704 9090 6760
rect 8850 5072 8906 5128
rect 8390 3032 8446 3088
rect 7746 2216 7802 2272
rect 8114 2216 8170 2272
rect 7930 856 7986 912
rect 8482 2216 8538 2272
rect 8850 2216 8906 2272
rect 10414 12724 10416 12744
rect 10416 12724 10468 12744
rect 10468 12724 10470 12744
rect 10414 12688 10470 12724
rect 9857 12538 9913 12540
rect 9937 12538 9993 12540
rect 10017 12538 10073 12540
rect 10097 12538 10153 12540
rect 9857 12486 9903 12538
rect 9903 12486 9913 12538
rect 9937 12486 9967 12538
rect 9967 12486 9979 12538
rect 9979 12486 9993 12538
rect 10017 12486 10031 12538
rect 10031 12486 10043 12538
rect 10043 12486 10073 12538
rect 10097 12486 10107 12538
rect 10107 12486 10153 12538
rect 9857 12484 9913 12486
rect 9937 12484 9993 12486
rect 10017 12484 10073 12486
rect 10097 12484 10153 12486
rect 9857 11450 9913 11452
rect 9937 11450 9993 11452
rect 10017 11450 10073 11452
rect 10097 11450 10153 11452
rect 9857 11398 9903 11450
rect 9903 11398 9913 11450
rect 9937 11398 9967 11450
rect 9967 11398 9979 11450
rect 9979 11398 9993 11450
rect 10017 11398 10031 11450
rect 10031 11398 10043 11450
rect 10043 11398 10073 11450
rect 10097 11398 10107 11450
rect 10107 11398 10153 11450
rect 9857 11396 9913 11398
rect 9937 11396 9993 11398
rect 10017 11396 10073 11398
rect 10097 11396 10153 11398
rect 9857 10362 9913 10364
rect 9937 10362 9993 10364
rect 10017 10362 10073 10364
rect 10097 10362 10153 10364
rect 9857 10310 9903 10362
rect 9903 10310 9913 10362
rect 9937 10310 9967 10362
rect 9967 10310 9979 10362
rect 9979 10310 9993 10362
rect 10017 10310 10031 10362
rect 10031 10310 10043 10362
rect 10043 10310 10073 10362
rect 10097 10310 10107 10362
rect 10107 10310 10153 10362
rect 9857 10308 9913 10310
rect 9937 10308 9993 10310
rect 10017 10308 10073 10310
rect 10097 10308 10153 10310
rect 9857 9274 9913 9276
rect 9937 9274 9993 9276
rect 10017 9274 10073 9276
rect 10097 9274 10153 9276
rect 9857 9222 9903 9274
rect 9903 9222 9913 9274
rect 9937 9222 9967 9274
rect 9967 9222 9979 9274
rect 9979 9222 9993 9274
rect 10017 9222 10031 9274
rect 10031 9222 10043 9274
rect 10043 9222 10073 9274
rect 10097 9222 10107 9274
rect 10107 9222 10153 9274
rect 9857 9220 9913 9222
rect 9937 9220 9993 9222
rect 10017 9220 10073 9222
rect 10097 9220 10153 9222
rect 9857 8186 9913 8188
rect 9937 8186 9993 8188
rect 10017 8186 10073 8188
rect 10097 8186 10153 8188
rect 9857 8134 9903 8186
rect 9903 8134 9913 8186
rect 9937 8134 9967 8186
rect 9967 8134 9979 8186
rect 9979 8134 9993 8186
rect 10017 8134 10031 8186
rect 10031 8134 10043 8186
rect 10043 8134 10073 8186
rect 10097 8134 10107 8186
rect 10107 8134 10153 8186
rect 9857 8132 9913 8134
rect 9937 8132 9993 8134
rect 10017 8132 10073 8134
rect 10097 8132 10153 8134
rect 9586 6840 9642 6896
rect 9857 7098 9913 7100
rect 9937 7098 9993 7100
rect 10017 7098 10073 7100
rect 10097 7098 10153 7100
rect 9857 7046 9903 7098
rect 9903 7046 9913 7098
rect 9937 7046 9967 7098
rect 9967 7046 9979 7098
rect 9979 7046 9993 7098
rect 10017 7046 10031 7098
rect 10031 7046 10043 7098
rect 10043 7046 10073 7098
rect 10097 7046 10107 7098
rect 10107 7046 10153 7098
rect 9857 7044 9913 7046
rect 9937 7044 9993 7046
rect 10017 7044 10073 7046
rect 10097 7044 10153 7046
rect 9770 6704 9826 6760
rect 9586 5364 9642 5400
rect 9586 5344 9588 5364
rect 9588 5344 9640 5364
rect 9640 5344 9642 5364
rect 9402 4528 9458 4584
rect 9857 6010 9913 6012
rect 9937 6010 9993 6012
rect 10017 6010 10073 6012
rect 10097 6010 10153 6012
rect 9857 5958 9903 6010
rect 9903 5958 9913 6010
rect 9937 5958 9967 6010
rect 9967 5958 9979 6010
rect 9979 5958 9993 6010
rect 10017 5958 10031 6010
rect 10031 5958 10043 6010
rect 10043 5958 10073 6010
rect 10097 5958 10107 6010
rect 10107 5958 10153 6010
rect 9857 5956 9913 5958
rect 9937 5956 9993 5958
rect 10017 5956 10073 5958
rect 10097 5956 10153 5958
rect 9857 4922 9913 4924
rect 9937 4922 9993 4924
rect 10017 4922 10073 4924
rect 10097 4922 10153 4924
rect 9857 4870 9903 4922
rect 9903 4870 9913 4922
rect 9937 4870 9967 4922
rect 9967 4870 9979 4922
rect 9979 4870 9993 4922
rect 10017 4870 10031 4922
rect 10031 4870 10043 4922
rect 10043 4870 10073 4922
rect 10097 4870 10107 4922
rect 10107 4870 10153 4922
rect 9857 4868 9913 4870
rect 9937 4868 9993 4870
rect 10017 4868 10073 4870
rect 10097 4868 10153 4870
rect 10046 4700 10048 4720
rect 10048 4700 10100 4720
rect 10100 4700 10102 4720
rect 10046 4664 10102 4700
rect 10414 6024 10470 6080
rect 9857 3834 9913 3836
rect 9937 3834 9993 3836
rect 10017 3834 10073 3836
rect 10097 3834 10153 3836
rect 9857 3782 9903 3834
rect 9903 3782 9913 3834
rect 9937 3782 9967 3834
rect 9967 3782 9979 3834
rect 9979 3782 9993 3834
rect 10017 3782 10031 3834
rect 10031 3782 10043 3834
rect 10043 3782 10073 3834
rect 10097 3782 10107 3834
rect 10107 3782 10153 3834
rect 9857 3780 9913 3782
rect 9937 3780 9993 3782
rect 10017 3780 10073 3782
rect 10097 3780 10153 3782
rect 9678 3440 9734 3496
rect 9402 2896 9458 2952
rect 9126 1400 9182 1456
rect 9402 2644 9458 2680
rect 9402 2624 9404 2644
rect 9404 2624 9456 2644
rect 9456 2624 9458 2644
rect 10138 3440 10194 3496
rect 9857 2746 9913 2748
rect 9937 2746 9993 2748
rect 10017 2746 10073 2748
rect 10097 2746 10153 2748
rect 9857 2694 9903 2746
rect 9903 2694 9913 2746
rect 9937 2694 9967 2746
rect 9967 2694 9979 2746
rect 9979 2694 9993 2746
rect 10017 2694 10031 2746
rect 10031 2694 10043 2746
rect 10043 2694 10073 2746
rect 10097 2694 10107 2746
rect 10107 2694 10153 2746
rect 9857 2692 9913 2694
rect 9937 2692 9993 2694
rect 10017 2692 10073 2694
rect 10097 2692 10153 2694
rect 9402 1672 9458 1728
rect 9770 2488 9826 2544
rect 10138 2352 10194 2408
rect 11242 21392 11298 21448
rect 11058 20304 11114 20360
rect 11150 19216 11206 19272
rect 10966 18128 11022 18184
rect 10966 17040 11022 17096
rect 12254 42880 12310 42936
rect 12824 43546 12880 43548
rect 12904 43546 12960 43548
rect 12984 43546 13040 43548
rect 13064 43546 13120 43548
rect 12824 43494 12870 43546
rect 12870 43494 12880 43546
rect 12904 43494 12934 43546
rect 12934 43494 12946 43546
rect 12946 43494 12960 43546
rect 12984 43494 12998 43546
rect 12998 43494 13010 43546
rect 13010 43494 13040 43546
rect 13064 43494 13074 43546
rect 13074 43494 13120 43546
rect 12824 43492 12880 43494
rect 12904 43492 12960 43494
rect 12984 43492 13040 43494
rect 13064 43492 13120 43494
rect 12898 43052 12900 43072
rect 12900 43052 12952 43072
rect 12952 43052 12954 43072
rect 12898 43016 12954 43052
rect 13082 43016 13138 43072
rect 13818 42880 13874 42936
rect 12824 42458 12880 42460
rect 12904 42458 12960 42460
rect 12984 42458 13040 42460
rect 13064 42458 13120 42460
rect 12824 42406 12870 42458
rect 12870 42406 12880 42458
rect 12904 42406 12934 42458
rect 12934 42406 12946 42458
rect 12946 42406 12960 42458
rect 12984 42406 12998 42458
rect 12998 42406 13010 42458
rect 13010 42406 13040 42458
rect 13064 42406 13074 42458
rect 13074 42406 13120 42458
rect 12824 42404 12880 42406
rect 12904 42404 12960 42406
rect 12984 42404 13040 42406
rect 13064 42404 13120 42406
rect 12530 41656 12586 41712
rect 12824 41370 12880 41372
rect 12904 41370 12960 41372
rect 12984 41370 13040 41372
rect 13064 41370 13120 41372
rect 12824 41318 12870 41370
rect 12870 41318 12880 41370
rect 12904 41318 12934 41370
rect 12934 41318 12946 41370
rect 12946 41318 12960 41370
rect 12984 41318 12998 41370
rect 12998 41318 13010 41370
rect 13010 41318 13040 41370
rect 13064 41318 13074 41370
rect 13074 41318 13120 41370
rect 12824 41316 12880 41318
rect 12904 41316 12960 41318
rect 12984 41316 13040 41318
rect 13064 41316 13120 41318
rect 12824 40282 12880 40284
rect 12904 40282 12960 40284
rect 12984 40282 13040 40284
rect 13064 40282 13120 40284
rect 12824 40230 12870 40282
rect 12870 40230 12880 40282
rect 12904 40230 12934 40282
rect 12934 40230 12946 40282
rect 12946 40230 12960 40282
rect 12984 40230 12998 40282
rect 12998 40230 13010 40282
rect 13010 40230 13040 40282
rect 13064 40230 13074 40282
rect 13074 40230 13120 40282
rect 12824 40228 12880 40230
rect 12904 40228 12960 40230
rect 12984 40228 13040 40230
rect 13064 40228 13120 40230
rect 11794 38800 11850 38856
rect 11978 35536 12034 35592
rect 12824 39194 12880 39196
rect 12904 39194 12960 39196
rect 12984 39194 13040 39196
rect 13064 39194 13120 39196
rect 12824 39142 12870 39194
rect 12870 39142 12880 39194
rect 12904 39142 12934 39194
rect 12934 39142 12946 39194
rect 12946 39142 12960 39194
rect 12984 39142 12998 39194
rect 12998 39142 13010 39194
rect 13010 39142 13040 39194
rect 13064 39142 13074 39194
rect 13074 39142 13120 39194
rect 12824 39140 12880 39142
rect 12904 39140 12960 39142
rect 12984 39140 13040 39142
rect 13064 39140 13120 39142
rect 12824 38106 12880 38108
rect 12904 38106 12960 38108
rect 12984 38106 13040 38108
rect 13064 38106 13120 38108
rect 12824 38054 12870 38106
rect 12870 38054 12880 38106
rect 12904 38054 12934 38106
rect 12934 38054 12946 38106
rect 12946 38054 12960 38106
rect 12984 38054 12998 38106
rect 12998 38054 13010 38106
rect 13010 38054 13040 38106
rect 13064 38054 13074 38106
rect 13074 38054 13120 38106
rect 12824 38052 12880 38054
rect 12904 38052 12960 38054
rect 12984 38052 13040 38054
rect 13064 38052 13120 38054
rect 12438 36216 12494 36272
rect 12070 34448 12126 34504
rect 11702 32952 11758 33008
rect 11794 32408 11850 32464
rect 11886 32292 11942 32328
rect 11886 32272 11888 32292
rect 11888 32272 11940 32292
rect 11940 32272 11942 32292
rect 11886 31728 11942 31784
rect 11886 31184 11942 31240
rect 11610 30368 11666 30424
rect 11610 30232 11666 30288
rect 11886 29688 11942 29744
rect 12824 37018 12880 37020
rect 12904 37018 12960 37020
rect 12984 37018 13040 37020
rect 13064 37018 13120 37020
rect 12824 36966 12870 37018
rect 12870 36966 12880 37018
rect 12904 36966 12934 37018
rect 12934 36966 12946 37018
rect 12946 36966 12960 37018
rect 12984 36966 12998 37018
rect 12998 36966 13010 37018
rect 13010 36966 13040 37018
rect 13064 36966 13074 37018
rect 13074 36966 13120 37018
rect 12824 36964 12880 36966
rect 12904 36964 12960 36966
rect 12984 36964 13040 36966
rect 13064 36964 13120 36966
rect 12824 35930 12880 35932
rect 12904 35930 12960 35932
rect 12984 35930 13040 35932
rect 13064 35930 13120 35932
rect 12824 35878 12870 35930
rect 12870 35878 12880 35930
rect 12904 35878 12934 35930
rect 12934 35878 12946 35930
rect 12946 35878 12960 35930
rect 12984 35878 12998 35930
rect 12998 35878 13010 35930
rect 13010 35878 13040 35930
rect 13064 35878 13074 35930
rect 13074 35878 13120 35930
rect 12824 35876 12880 35878
rect 12904 35876 12960 35878
rect 12984 35876 13040 35878
rect 13064 35876 13120 35878
rect 12824 34842 12880 34844
rect 12904 34842 12960 34844
rect 12984 34842 13040 34844
rect 13064 34842 13120 34844
rect 12824 34790 12870 34842
rect 12870 34790 12880 34842
rect 12904 34790 12934 34842
rect 12934 34790 12946 34842
rect 12946 34790 12960 34842
rect 12984 34790 12998 34842
rect 12998 34790 13010 34842
rect 13010 34790 13040 34842
rect 13064 34790 13074 34842
rect 13074 34790 13120 34842
rect 12824 34788 12880 34790
rect 12904 34788 12960 34790
rect 12984 34788 13040 34790
rect 13064 34788 13120 34790
rect 12824 33754 12880 33756
rect 12904 33754 12960 33756
rect 12984 33754 13040 33756
rect 13064 33754 13120 33756
rect 12824 33702 12870 33754
rect 12870 33702 12880 33754
rect 12904 33702 12934 33754
rect 12934 33702 12946 33754
rect 12946 33702 12960 33754
rect 12984 33702 12998 33754
rect 12998 33702 13010 33754
rect 13010 33702 13040 33754
rect 13064 33702 13074 33754
rect 13074 33702 13120 33754
rect 12824 33700 12880 33702
rect 12904 33700 12960 33702
rect 12984 33700 13040 33702
rect 13064 33700 13120 33702
rect 12162 29008 12218 29064
rect 11978 26424 12034 26480
rect 13082 32836 13138 32872
rect 13082 32816 13084 32836
rect 13084 32816 13136 32836
rect 13136 32816 13138 32836
rect 12824 32666 12880 32668
rect 12904 32666 12960 32668
rect 12984 32666 13040 32668
rect 13064 32666 13120 32668
rect 12824 32614 12870 32666
rect 12870 32614 12880 32666
rect 12904 32614 12934 32666
rect 12934 32614 12946 32666
rect 12946 32614 12960 32666
rect 12984 32614 12998 32666
rect 12998 32614 13010 32666
rect 13010 32614 13040 32666
rect 13064 32614 13074 32666
rect 13074 32614 13120 32666
rect 12824 32612 12880 32614
rect 12904 32612 12960 32614
rect 12984 32612 13040 32614
rect 13064 32612 13120 32614
rect 12824 31578 12880 31580
rect 12904 31578 12960 31580
rect 12984 31578 13040 31580
rect 13064 31578 13120 31580
rect 12824 31526 12870 31578
rect 12870 31526 12880 31578
rect 12904 31526 12934 31578
rect 12934 31526 12946 31578
rect 12946 31526 12960 31578
rect 12984 31526 12998 31578
rect 12998 31526 13010 31578
rect 13010 31526 13040 31578
rect 13064 31526 13074 31578
rect 13074 31526 13120 31578
rect 12824 31524 12880 31526
rect 12904 31524 12960 31526
rect 12984 31524 13040 31526
rect 13064 31524 13120 31526
rect 13082 31184 13138 31240
rect 12824 30490 12880 30492
rect 12904 30490 12960 30492
rect 12984 30490 13040 30492
rect 13064 30490 13120 30492
rect 12824 30438 12870 30490
rect 12870 30438 12880 30490
rect 12904 30438 12934 30490
rect 12934 30438 12946 30490
rect 12946 30438 12960 30490
rect 12984 30438 12998 30490
rect 12998 30438 13010 30490
rect 13010 30438 13040 30490
rect 13064 30438 13074 30490
rect 13074 30438 13120 30490
rect 12824 30436 12880 30438
rect 12904 30436 12960 30438
rect 12984 30436 13040 30438
rect 13064 30436 13120 30438
rect 13174 29552 13230 29608
rect 12824 29402 12880 29404
rect 12904 29402 12960 29404
rect 12984 29402 13040 29404
rect 13064 29402 13120 29404
rect 12824 29350 12870 29402
rect 12870 29350 12880 29402
rect 12904 29350 12934 29402
rect 12934 29350 12946 29402
rect 12946 29350 12960 29402
rect 12984 29350 12998 29402
rect 12998 29350 13010 29402
rect 13010 29350 13040 29402
rect 13064 29350 13074 29402
rect 13074 29350 13120 29402
rect 12824 29348 12880 29350
rect 12904 29348 12960 29350
rect 12984 29348 13040 29350
rect 13064 29348 13120 29350
rect 12990 29164 13046 29200
rect 12990 29144 12992 29164
rect 12992 29144 13044 29164
rect 13044 29144 13046 29164
rect 12530 28464 12586 28520
rect 12346 26988 12402 27024
rect 12346 26968 12348 26988
rect 12348 26968 12400 26988
rect 12400 26968 12402 26988
rect 11610 19760 11666 19816
rect 11518 17604 11574 17640
rect 11518 17584 11520 17604
rect 11520 17584 11572 17604
rect 11572 17584 11574 17604
rect 11426 15408 11482 15464
rect 9857 1658 9913 1660
rect 9937 1658 9993 1660
rect 10017 1658 10073 1660
rect 10097 1658 10153 1660
rect 9857 1606 9903 1658
rect 9903 1606 9913 1658
rect 9937 1606 9967 1658
rect 9967 1606 9979 1658
rect 9979 1606 9993 1658
rect 10017 1606 10031 1658
rect 10031 1606 10043 1658
rect 10043 1606 10073 1658
rect 10097 1606 10107 1658
rect 10107 1606 10153 1658
rect 9857 1604 9913 1606
rect 9937 1604 9993 1606
rect 10017 1604 10073 1606
rect 10097 1604 10153 1606
rect 11886 22208 11942 22264
rect 12530 26424 12586 26480
rect 12824 28314 12880 28316
rect 12904 28314 12960 28316
rect 12984 28314 13040 28316
rect 13064 28314 13120 28316
rect 12824 28262 12870 28314
rect 12870 28262 12880 28314
rect 12904 28262 12934 28314
rect 12934 28262 12946 28314
rect 12946 28262 12960 28314
rect 12984 28262 12998 28314
rect 12998 28262 13010 28314
rect 13010 28262 13040 28314
rect 13064 28262 13074 28314
rect 13074 28262 13120 28314
rect 12824 28260 12880 28262
rect 12904 28260 12960 28262
rect 12984 28260 13040 28262
rect 13064 28260 13120 28262
rect 12824 27226 12880 27228
rect 12904 27226 12960 27228
rect 12984 27226 13040 27228
rect 13064 27226 13120 27228
rect 12824 27174 12870 27226
rect 12870 27174 12880 27226
rect 12904 27174 12934 27226
rect 12934 27174 12946 27226
rect 12946 27174 12960 27226
rect 12984 27174 12998 27226
rect 12998 27174 13010 27226
rect 13010 27174 13040 27226
rect 13064 27174 13074 27226
rect 13074 27174 13120 27226
rect 12824 27172 12880 27174
rect 12904 27172 12960 27174
rect 12984 27172 13040 27174
rect 13064 27172 13120 27174
rect 12824 26138 12880 26140
rect 12904 26138 12960 26140
rect 12984 26138 13040 26140
rect 13064 26138 13120 26140
rect 12824 26086 12870 26138
rect 12870 26086 12880 26138
rect 12904 26086 12934 26138
rect 12934 26086 12946 26138
rect 12946 26086 12960 26138
rect 12984 26086 12998 26138
rect 12998 26086 13010 26138
rect 13010 26086 13040 26138
rect 13064 26086 13074 26138
rect 13074 26086 13120 26138
rect 12824 26084 12880 26086
rect 12904 26084 12960 26086
rect 12984 26084 13040 26086
rect 13064 26084 13120 26086
rect 12824 25050 12880 25052
rect 12904 25050 12960 25052
rect 12984 25050 13040 25052
rect 13064 25050 13120 25052
rect 12824 24998 12870 25050
rect 12870 24998 12880 25050
rect 12904 24998 12934 25050
rect 12934 24998 12946 25050
rect 12946 24998 12960 25050
rect 12984 24998 12998 25050
rect 12998 24998 13010 25050
rect 13010 24998 13040 25050
rect 13064 24998 13074 25050
rect 13074 24998 13120 25050
rect 12824 24996 12880 24998
rect 12904 24996 12960 24998
rect 12984 24996 13040 24998
rect 13064 24996 13120 24998
rect 12346 21936 12402 21992
rect 12530 20984 12586 21040
rect 11978 19624 12034 19680
rect 12070 18264 12126 18320
rect 10874 5888 10930 5944
rect 11242 5752 11298 5808
rect 10782 2352 10838 2408
rect 11334 4664 11390 4720
rect 11978 15444 11980 15464
rect 11980 15444 12032 15464
rect 12032 15444 12034 15464
rect 11978 15408 12034 15444
rect 11702 10104 11758 10160
rect 11794 9968 11850 10024
rect 12070 10104 12126 10160
rect 12824 23962 12880 23964
rect 12904 23962 12960 23964
rect 12984 23962 13040 23964
rect 13064 23962 13120 23964
rect 12824 23910 12870 23962
rect 12870 23910 12880 23962
rect 12904 23910 12934 23962
rect 12934 23910 12946 23962
rect 12946 23910 12960 23962
rect 12984 23910 12998 23962
rect 12998 23910 13010 23962
rect 13010 23910 13040 23962
rect 13064 23910 13074 23962
rect 13074 23910 13120 23962
rect 12824 23908 12880 23910
rect 12904 23908 12960 23910
rect 12984 23908 13040 23910
rect 13064 23908 13120 23910
rect 12824 22874 12880 22876
rect 12904 22874 12960 22876
rect 12984 22874 13040 22876
rect 13064 22874 13120 22876
rect 12824 22822 12870 22874
rect 12870 22822 12880 22874
rect 12904 22822 12934 22874
rect 12934 22822 12946 22874
rect 12946 22822 12960 22874
rect 12984 22822 12998 22874
rect 12998 22822 13010 22874
rect 13010 22822 13040 22874
rect 13064 22822 13074 22874
rect 13074 22822 13120 22874
rect 12824 22820 12880 22822
rect 12904 22820 12960 22822
rect 12984 22820 13040 22822
rect 13064 22820 13120 22822
rect 12824 21786 12880 21788
rect 12904 21786 12960 21788
rect 12984 21786 13040 21788
rect 13064 21786 13120 21788
rect 12824 21734 12870 21786
rect 12870 21734 12880 21786
rect 12904 21734 12934 21786
rect 12934 21734 12946 21786
rect 12946 21734 12960 21786
rect 12984 21734 12998 21786
rect 12998 21734 13010 21786
rect 13010 21734 13040 21786
rect 13064 21734 13074 21786
rect 13074 21734 13120 21786
rect 12824 21732 12880 21734
rect 12904 21732 12960 21734
rect 12984 21732 13040 21734
rect 13064 21732 13120 21734
rect 13450 34856 13506 34912
rect 13450 29144 13506 29200
rect 14278 42880 14334 42936
rect 14922 42880 14978 42936
rect 15290 42880 15346 42936
rect 14094 38664 14150 38720
rect 14002 34992 14058 35048
rect 14186 31728 14242 31784
rect 13910 31592 13966 31648
rect 13910 30504 13966 30560
rect 14094 30368 14150 30424
rect 14002 29144 14058 29200
rect 13818 27648 13874 27704
rect 13266 21664 13322 21720
rect 12824 20698 12880 20700
rect 12904 20698 12960 20700
rect 12984 20698 13040 20700
rect 13064 20698 13120 20700
rect 12824 20646 12870 20698
rect 12870 20646 12880 20698
rect 12904 20646 12934 20698
rect 12934 20646 12946 20698
rect 12946 20646 12960 20698
rect 12984 20646 12998 20698
rect 12998 20646 13010 20698
rect 13010 20646 13040 20698
rect 13064 20646 13074 20698
rect 13074 20646 13120 20698
rect 12824 20644 12880 20646
rect 12904 20644 12960 20646
rect 12984 20644 13040 20646
rect 13064 20644 13120 20646
rect 12898 20440 12954 20496
rect 12824 19610 12880 19612
rect 12904 19610 12960 19612
rect 12984 19610 13040 19612
rect 13064 19610 13120 19612
rect 12824 19558 12870 19610
rect 12870 19558 12880 19610
rect 12904 19558 12934 19610
rect 12934 19558 12946 19610
rect 12946 19558 12960 19610
rect 12984 19558 12998 19610
rect 12998 19558 13010 19610
rect 13010 19558 13040 19610
rect 13064 19558 13074 19610
rect 13074 19558 13120 19610
rect 12824 19556 12880 19558
rect 12904 19556 12960 19558
rect 12984 19556 13040 19558
rect 13064 19556 13120 19558
rect 12346 13640 12402 13696
rect 12346 12280 12402 12336
rect 12824 18522 12880 18524
rect 12904 18522 12960 18524
rect 12984 18522 13040 18524
rect 13064 18522 13120 18524
rect 12824 18470 12870 18522
rect 12870 18470 12880 18522
rect 12904 18470 12934 18522
rect 12934 18470 12946 18522
rect 12946 18470 12960 18522
rect 12984 18470 12998 18522
rect 12998 18470 13010 18522
rect 13010 18470 13040 18522
rect 13064 18470 13074 18522
rect 13074 18470 13120 18522
rect 12824 18468 12880 18470
rect 12904 18468 12960 18470
rect 12984 18468 13040 18470
rect 13064 18468 13120 18470
rect 12824 17434 12880 17436
rect 12904 17434 12960 17436
rect 12984 17434 13040 17436
rect 13064 17434 13120 17436
rect 12824 17382 12870 17434
rect 12870 17382 12880 17434
rect 12904 17382 12934 17434
rect 12934 17382 12946 17434
rect 12946 17382 12960 17434
rect 12984 17382 12998 17434
rect 12998 17382 13010 17434
rect 13010 17382 13040 17434
rect 13064 17382 13074 17434
rect 13074 17382 13120 17434
rect 12824 17380 12880 17382
rect 12904 17380 12960 17382
rect 12984 17380 13040 17382
rect 13064 17380 13120 17382
rect 12824 16346 12880 16348
rect 12904 16346 12960 16348
rect 12984 16346 13040 16348
rect 13064 16346 13120 16348
rect 12824 16294 12870 16346
rect 12870 16294 12880 16346
rect 12904 16294 12934 16346
rect 12934 16294 12946 16346
rect 12946 16294 12960 16346
rect 12984 16294 12998 16346
rect 12998 16294 13010 16346
rect 13010 16294 13040 16346
rect 13064 16294 13074 16346
rect 13074 16294 13120 16346
rect 12824 16292 12880 16294
rect 12904 16292 12960 16294
rect 12984 16292 13040 16294
rect 13064 16292 13120 16294
rect 12714 15408 12770 15464
rect 12824 15258 12880 15260
rect 12904 15258 12960 15260
rect 12984 15258 13040 15260
rect 13064 15258 13120 15260
rect 12824 15206 12870 15258
rect 12870 15206 12880 15258
rect 12904 15206 12934 15258
rect 12934 15206 12946 15258
rect 12946 15206 12960 15258
rect 12984 15206 12998 15258
rect 12998 15206 13010 15258
rect 13010 15206 13040 15258
rect 13064 15206 13074 15258
rect 13074 15206 13120 15258
rect 12824 15204 12880 15206
rect 12904 15204 12960 15206
rect 12984 15204 13040 15206
rect 13064 15204 13120 15206
rect 13910 24112 13966 24168
rect 13358 17720 13414 17776
rect 13726 19488 13782 19544
rect 13358 16496 13414 16552
rect 12824 14170 12880 14172
rect 12904 14170 12960 14172
rect 12984 14170 13040 14172
rect 13064 14170 13120 14172
rect 12824 14118 12870 14170
rect 12870 14118 12880 14170
rect 12904 14118 12934 14170
rect 12934 14118 12946 14170
rect 12946 14118 12960 14170
rect 12984 14118 12998 14170
rect 12998 14118 13010 14170
rect 13010 14118 13040 14170
rect 13064 14118 13074 14170
rect 13074 14118 13120 14170
rect 12824 14116 12880 14118
rect 12904 14116 12960 14118
rect 12984 14116 13040 14118
rect 13064 14116 13120 14118
rect 12824 13082 12880 13084
rect 12904 13082 12960 13084
rect 12984 13082 13040 13084
rect 13064 13082 13120 13084
rect 12824 13030 12870 13082
rect 12870 13030 12880 13082
rect 12904 13030 12934 13082
rect 12934 13030 12946 13082
rect 12946 13030 12960 13082
rect 12984 13030 12998 13082
rect 12998 13030 13010 13082
rect 13010 13030 13040 13082
rect 13064 13030 13074 13082
rect 13074 13030 13120 13082
rect 12824 13028 12880 13030
rect 12904 13028 12960 13030
rect 12984 13028 13040 13030
rect 13064 13028 13120 13030
rect 12824 11994 12880 11996
rect 12904 11994 12960 11996
rect 12984 11994 13040 11996
rect 13064 11994 13120 11996
rect 12824 11942 12870 11994
rect 12870 11942 12880 11994
rect 12904 11942 12934 11994
rect 12934 11942 12946 11994
rect 12946 11942 12960 11994
rect 12984 11942 12998 11994
rect 12998 11942 13010 11994
rect 13010 11942 13040 11994
rect 13064 11942 13074 11994
rect 13074 11942 13120 11994
rect 12824 11940 12880 11942
rect 12904 11940 12960 11942
rect 12984 11940 13040 11942
rect 13064 11940 13120 11942
rect 12824 10906 12880 10908
rect 12904 10906 12960 10908
rect 12984 10906 13040 10908
rect 13064 10906 13120 10908
rect 12824 10854 12870 10906
rect 12870 10854 12880 10906
rect 12904 10854 12934 10906
rect 12934 10854 12946 10906
rect 12946 10854 12960 10906
rect 12984 10854 12998 10906
rect 12998 10854 13010 10906
rect 13010 10854 13040 10906
rect 13064 10854 13074 10906
rect 13074 10854 13120 10906
rect 12824 10852 12880 10854
rect 12904 10852 12960 10854
rect 12984 10852 13040 10854
rect 13064 10852 13120 10854
rect 12806 10376 12862 10432
rect 12162 9016 12218 9072
rect 11886 6840 11942 6896
rect 12254 6704 12310 6760
rect 12346 5616 12402 5672
rect 12824 9818 12880 9820
rect 12904 9818 12960 9820
rect 12984 9818 13040 9820
rect 13064 9818 13120 9820
rect 12824 9766 12870 9818
rect 12870 9766 12880 9818
rect 12904 9766 12934 9818
rect 12934 9766 12946 9818
rect 12946 9766 12960 9818
rect 12984 9766 12998 9818
rect 12998 9766 13010 9818
rect 13010 9766 13040 9818
rect 13064 9766 13074 9818
rect 13074 9766 13120 9818
rect 12824 9764 12880 9766
rect 12904 9764 12960 9766
rect 12984 9764 13040 9766
rect 13064 9764 13120 9766
rect 12824 8730 12880 8732
rect 12904 8730 12960 8732
rect 12984 8730 13040 8732
rect 13064 8730 13120 8732
rect 12824 8678 12870 8730
rect 12870 8678 12880 8730
rect 12904 8678 12934 8730
rect 12934 8678 12946 8730
rect 12946 8678 12960 8730
rect 12984 8678 12998 8730
rect 12998 8678 13010 8730
rect 13010 8678 13040 8730
rect 13064 8678 13074 8730
rect 13074 8678 13120 8730
rect 12824 8676 12880 8678
rect 12904 8676 12960 8678
rect 12984 8676 13040 8678
rect 13064 8676 13120 8678
rect 12824 7642 12880 7644
rect 12904 7642 12960 7644
rect 12984 7642 13040 7644
rect 13064 7642 13120 7644
rect 12824 7590 12870 7642
rect 12870 7590 12880 7642
rect 12904 7590 12934 7642
rect 12934 7590 12946 7642
rect 12946 7590 12960 7642
rect 12984 7590 12998 7642
rect 12998 7590 13010 7642
rect 13010 7590 13040 7642
rect 13064 7590 13074 7642
rect 13074 7590 13120 7642
rect 12824 7588 12880 7590
rect 12904 7588 12960 7590
rect 12984 7588 13040 7590
rect 13064 7588 13120 7590
rect 12824 6554 12880 6556
rect 12904 6554 12960 6556
rect 12984 6554 13040 6556
rect 13064 6554 13120 6556
rect 12824 6502 12870 6554
rect 12870 6502 12880 6554
rect 12904 6502 12934 6554
rect 12934 6502 12946 6554
rect 12946 6502 12960 6554
rect 12984 6502 12998 6554
rect 12998 6502 13010 6554
rect 13010 6502 13040 6554
rect 13064 6502 13074 6554
rect 13074 6502 13120 6554
rect 12824 6500 12880 6502
rect 12904 6500 12960 6502
rect 12984 6500 13040 6502
rect 13064 6500 13120 6502
rect 12346 4700 12348 4720
rect 12348 4700 12400 4720
rect 12400 4700 12402 4720
rect 12346 4664 12402 4700
rect 12162 3984 12218 4040
rect 11794 3032 11850 3088
rect 11978 2624 12034 2680
rect 12622 5344 12678 5400
rect 12824 5466 12880 5468
rect 12904 5466 12960 5468
rect 12984 5466 13040 5468
rect 13064 5466 13120 5468
rect 12824 5414 12870 5466
rect 12870 5414 12880 5466
rect 12904 5414 12934 5466
rect 12934 5414 12946 5466
rect 12946 5414 12960 5466
rect 12984 5414 12998 5466
rect 12998 5414 13010 5466
rect 13010 5414 13040 5466
rect 13064 5414 13074 5466
rect 13074 5414 13120 5466
rect 12824 5412 12880 5414
rect 12904 5412 12960 5414
rect 12984 5412 13040 5414
rect 13064 5412 13120 5414
rect 12824 4378 12880 4380
rect 12904 4378 12960 4380
rect 12984 4378 13040 4380
rect 13064 4378 13120 4380
rect 12824 4326 12870 4378
rect 12870 4326 12880 4378
rect 12904 4326 12934 4378
rect 12934 4326 12946 4378
rect 12946 4326 12960 4378
rect 12984 4326 12998 4378
rect 12998 4326 13010 4378
rect 13010 4326 13040 4378
rect 13064 4326 13074 4378
rect 13074 4326 13120 4378
rect 12824 4324 12880 4326
rect 12904 4324 12960 4326
rect 12984 4324 13040 4326
rect 13064 4324 13120 4326
rect 12622 4140 12678 4176
rect 12622 4120 12624 4140
rect 12624 4120 12676 4140
rect 12676 4120 12678 4140
rect 12824 3290 12880 3292
rect 12904 3290 12960 3292
rect 12984 3290 13040 3292
rect 13064 3290 13120 3292
rect 12824 3238 12870 3290
rect 12870 3238 12880 3290
rect 12904 3238 12934 3290
rect 12934 3238 12946 3290
rect 12946 3238 12960 3290
rect 12984 3238 12998 3290
rect 12998 3238 13010 3290
rect 13010 3238 13040 3290
rect 13064 3238 13074 3290
rect 13074 3238 13120 3290
rect 12824 3236 12880 3238
rect 12904 3236 12960 3238
rect 12984 3236 13040 3238
rect 13064 3236 13120 3238
rect 13266 6160 13322 6216
rect 13266 5344 13322 5400
rect 13634 12688 13690 12744
rect 14186 29008 14242 29064
rect 14186 24556 14188 24576
rect 14188 24556 14240 24576
rect 14240 24556 14242 24576
rect 14186 24520 14242 24556
rect 14002 13640 14058 13696
rect 14370 29960 14426 30016
rect 14922 33496 14978 33552
rect 15290 42200 15346 42256
rect 14554 26152 14610 26208
rect 14922 29144 14978 29200
rect 15791 43002 15847 43004
rect 15871 43002 15927 43004
rect 15951 43002 16007 43004
rect 16031 43002 16087 43004
rect 15791 42950 15837 43002
rect 15837 42950 15847 43002
rect 15871 42950 15901 43002
rect 15901 42950 15913 43002
rect 15913 42950 15927 43002
rect 15951 42950 15965 43002
rect 15965 42950 15977 43002
rect 15977 42950 16007 43002
rect 16031 42950 16041 43002
rect 16041 42950 16087 43002
rect 15791 42948 15847 42950
rect 15871 42948 15927 42950
rect 15951 42948 16007 42950
rect 16031 42948 16087 42950
rect 15791 41914 15847 41916
rect 15871 41914 15927 41916
rect 15951 41914 16007 41916
rect 16031 41914 16087 41916
rect 15791 41862 15837 41914
rect 15837 41862 15847 41914
rect 15871 41862 15901 41914
rect 15901 41862 15913 41914
rect 15913 41862 15927 41914
rect 15951 41862 15965 41914
rect 15965 41862 15977 41914
rect 15977 41862 16007 41914
rect 16031 41862 16041 41914
rect 16041 41862 16087 41914
rect 15791 41860 15847 41862
rect 15871 41860 15927 41862
rect 15951 41860 16007 41862
rect 16031 41860 16087 41862
rect 15791 40826 15847 40828
rect 15871 40826 15927 40828
rect 15951 40826 16007 40828
rect 16031 40826 16087 40828
rect 15791 40774 15837 40826
rect 15837 40774 15847 40826
rect 15871 40774 15901 40826
rect 15901 40774 15913 40826
rect 15913 40774 15927 40826
rect 15951 40774 15965 40826
rect 15965 40774 15977 40826
rect 15977 40774 16007 40826
rect 16031 40774 16041 40826
rect 16041 40774 16087 40826
rect 15791 40772 15847 40774
rect 15871 40772 15927 40774
rect 15951 40772 16007 40774
rect 16031 40772 16087 40774
rect 15791 39738 15847 39740
rect 15871 39738 15927 39740
rect 15951 39738 16007 39740
rect 16031 39738 16087 39740
rect 15791 39686 15837 39738
rect 15837 39686 15847 39738
rect 15871 39686 15901 39738
rect 15901 39686 15913 39738
rect 15913 39686 15927 39738
rect 15951 39686 15965 39738
rect 15965 39686 15977 39738
rect 15977 39686 16007 39738
rect 16031 39686 16041 39738
rect 16041 39686 16087 39738
rect 15791 39684 15847 39686
rect 15871 39684 15927 39686
rect 15951 39684 16007 39686
rect 16031 39684 16087 39686
rect 16302 42200 16358 42256
rect 16210 41420 16212 41440
rect 16212 41420 16264 41440
rect 16264 41420 16266 41440
rect 16210 41384 16266 41420
rect 15791 38650 15847 38652
rect 15871 38650 15927 38652
rect 15951 38650 16007 38652
rect 16031 38650 16087 38652
rect 15791 38598 15837 38650
rect 15837 38598 15847 38650
rect 15871 38598 15901 38650
rect 15901 38598 15913 38650
rect 15913 38598 15927 38650
rect 15951 38598 15965 38650
rect 15965 38598 15977 38650
rect 15977 38598 16007 38650
rect 16031 38598 16041 38650
rect 16041 38598 16087 38650
rect 15791 38596 15847 38598
rect 15871 38596 15927 38598
rect 15951 38596 16007 38598
rect 16031 38596 16087 38598
rect 15791 37562 15847 37564
rect 15871 37562 15927 37564
rect 15951 37562 16007 37564
rect 16031 37562 16087 37564
rect 15791 37510 15837 37562
rect 15837 37510 15847 37562
rect 15871 37510 15901 37562
rect 15901 37510 15913 37562
rect 15913 37510 15927 37562
rect 15951 37510 15965 37562
rect 15965 37510 15977 37562
rect 15977 37510 16007 37562
rect 16031 37510 16041 37562
rect 16041 37510 16087 37562
rect 15791 37508 15847 37510
rect 15871 37508 15927 37510
rect 15951 37508 16007 37510
rect 16031 37508 16087 37510
rect 15791 36474 15847 36476
rect 15871 36474 15927 36476
rect 15951 36474 16007 36476
rect 16031 36474 16087 36476
rect 15791 36422 15837 36474
rect 15837 36422 15847 36474
rect 15871 36422 15901 36474
rect 15901 36422 15913 36474
rect 15913 36422 15927 36474
rect 15951 36422 15965 36474
rect 15965 36422 15977 36474
rect 15977 36422 16007 36474
rect 16031 36422 16041 36474
rect 16041 36422 16087 36474
rect 15791 36420 15847 36422
rect 15871 36420 15927 36422
rect 15951 36420 16007 36422
rect 16031 36420 16087 36422
rect 15290 35556 15346 35592
rect 15290 35536 15292 35556
rect 15292 35536 15344 35556
rect 15344 35536 15346 35556
rect 15791 35386 15847 35388
rect 15871 35386 15927 35388
rect 15951 35386 16007 35388
rect 16031 35386 16087 35388
rect 15791 35334 15837 35386
rect 15837 35334 15847 35386
rect 15871 35334 15901 35386
rect 15901 35334 15913 35386
rect 15913 35334 15927 35386
rect 15951 35334 15965 35386
rect 15965 35334 15977 35386
rect 15977 35334 16007 35386
rect 16031 35334 16041 35386
rect 16041 35334 16087 35386
rect 15791 35332 15847 35334
rect 15871 35332 15927 35334
rect 15951 35332 16007 35334
rect 16031 35332 16087 35334
rect 16118 34620 16120 34640
rect 16120 34620 16172 34640
rect 16172 34620 16174 34640
rect 16118 34584 16174 34620
rect 15791 34298 15847 34300
rect 15871 34298 15927 34300
rect 15951 34298 16007 34300
rect 16031 34298 16087 34300
rect 15791 34246 15837 34298
rect 15837 34246 15847 34298
rect 15871 34246 15901 34298
rect 15901 34246 15913 34298
rect 15913 34246 15927 34298
rect 15951 34246 15965 34298
rect 15965 34246 15977 34298
rect 15977 34246 16007 34298
rect 16031 34246 16041 34298
rect 16041 34246 16087 34298
rect 15791 34244 15847 34246
rect 15871 34244 15927 34246
rect 15951 34244 16007 34246
rect 16031 34244 16087 34246
rect 16670 38664 16726 38720
rect 18758 43546 18814 43548
rect 18838 43546 18894 43548
rect 18918 43546 18974 43548
rect 18998 43546 19054 43548
rect 18758 43494 18804 43546
rect 18804 43494 18814 43546
rect 18838 43494 18868 43546
rect 18868 43494 18880 43546
rect 18880 43494 18894 43546
rect 18918 43494 18932 43546
rect 18932 43494 18944 43546
rect 18944 43494 18974 43546
rect 18998 43494 19008 43546
rect 19008 43494 19054 43546
rect 18758 43492 18814 43494
rect 18838 43492 18894 43494
rect 18918 43492 18974 43494
rect 18998 43492 19054 43494
rect 18418 42744 18474 42800
rect 17590 42200 17646 42256
rect 17314 41792 17370 41848
rect 17590 41656 17646 41712
rect 17958 41656 18014 41712
rect 16854 40060 16856 40080
rect 16856 40060 16908 40080
rect 16908 40060 16910 40080
rect 16854 40024 16910 40060
rect 15382 32408 15438 32464
rect 14738 27648 14794 27704
rect 15014 28328 15070 28384
rect 15290 28056 15346 28112
rect 15791 33210 15847 33212
rect 15871 33210 15927 33212
rect 15951 33210 16007 33212
rect 16031 33210 16087 33212
rect 15791 33158 15837 33210
rect 15837 33158 15847 33210
rect 15871 33158 15901 33210
rect 15901 33158 15913 33210
rect 15913 33158 15927 33210
rect 15951 33158 15965 33210
rect 15965 33158 15977 33210
rect 15977 33158 16007 33210
rect 16031 33158 16041 33210
rect 16041 33158 16087 33210
rect 15791 33156 15847 33158
rect 15871 33156 15927 33158
rect 15951 33156 16007 33158
rect 16031 33156 16087 33158
rect 15658 32408 15714 32464
rect 15791 32122 15847 32124
rect 15871 32122 15927 32124
rect 15951 32122 16007 32124
rect 16031 32122 16087 32124
rect 15791 32070 15837 32122
rect 15837 32070 15847 32122
rect 15871 32070 15901 32122
rect 15901 32070 15913 32122
rect 15913 32070 15927 32122
rect 15951 32070 15965 32122
rect 15965 32070 15977 32122
rect 15977 32070 16007 32122
rect 16031 32070 16041 32122
rect 16041 32070 16087 32122
rect 15791 32068 15847 32070
rect 15871 32068 15927 32070
rect 15951 32068 16007 32070
rect 16031 32068 16087 32070
rect 15566 32000 15622 32056
rect 16026 31864 16082 31920
rect 15791 31034 15847 31036
rect 15871 31034 15927 31036
rect 15951 31034 16007 31036
rect 16031 31034 16087 31036
rect 15791 30982 15837 31034
rect 15837 30982 15847 31034
rect 15871 30982 15901 31034
rect 15901 30982 15913 31034
rect 15913 30982 15927 31034
rect 15951 30982 15965 31034
rect 15965 30982 15977 31034
rect 15977 30982 16007 31034
rect 16031 30982 16041 31034
rect 16041 30982 16087 31034
rect 15791 30980 15847 30982
rect 15871 30980 15927 30982
rect 15951 30980 16007 30982
rect 16031 30980 16087 30982
rect 15474 28636 15476 28656
rect 15476 28636 15528 28656
rect 15528 28636 15530 28656
rect 15474 28600 15530 28636
rect 15474 26288 15530 26344
rect 15290 23568 15346 23624
rect 15198 23432 15254 23488
rect 15290 22344 15346 22400
rect 15106 21664 15162 21720
rect 14922 21256 14978 21312
rect 14462 19352 14518 19408
rect 14922 19896 14978 19952
rect 14738 18808 14794 18864
rect 13450 8744 13506 8800
rect 14554 15444 14556 15464
rect 14556 15444 14608 15464
rect 14608 15444 14610 15464
rect 14554 15408 14610 15444
rect 14370 12824 14426 12880
rect 14646 13912 14702 13968
rect 13542 5208 13598 5264
rect 13726 7248 13782 7304
rect 13818 5888 13874 5944
rect 13634 2352 13690 2408
rect 12824 2202 12880 2204
rect 12904 2202 12960 2204
rect 12984 2202 13040 2204
rect 13064 2202 13120 2204
rect 12824 2150 12870 2202
rect 12870 2150 12880 2202
rect 12904 2150 12934 2202
rect 12934 2150 12946 2202
rect 12946 2150 12960 2202
rect 12984 2150 12998 2202
rect 12998 2150 13010 2202
rect 13010 2150 13040 2202
rect 13064 2150 13074 2202
rect 13074 2150 13120 2202
rect 12824 2148 12880 2150
rect 12904 2148 12960 2150
rect 12984 2148 13040 2150
rect 13064 2148 13120 2150
rect 13726 1964 13782 2000
rect 13726 1944 13728 1964
rect 13728 1944 13780 1964
rect 13780 1944 13782 1964
rect 12824 1114 12880 1116
rect 12904 1114 12960 1116
rect 12984 1114 13040 1116
rect 13064 1114 13120 1116
rect 12824 1062 12870 1114
rect 12870 1062 12880 1114
rect 12904 1062 12934 1114
rect 12934 1062 12946 1114
rect 12946 1062 12960 1114
rect 12984 1062 12998 1114
rect 12998 1062 13010 1114
rect 13010 1062 13040 1114
rect 13064 1062 13074 1114
rect 13074 1062 13120 1114
rect 12824 1060 12880 1062
rect 12904 1060 12960 1062
rect 12984 1060 13040 1062
rect 13064 1060 13120 1062
rect 14646 5752 14702 5808
rect 14370 5208 14426 5264
rect 15014 11092 15016 11112
rect 15016 11092 15068 11112
rect 15068 11092 15070 11112
rect 15014 11056 15070 11092
rect 14278 1808 14334 1864
rect 14830 2624 14886 2680
rect 14738 2488 14794 2544
rect 15382 21664 15438 21720
rect 15791 29946 15847 29948
rect 15871 29946 15927 29948
rect 15951 29946 16007 29948
rect 16031 29946 16087 29948
rect 15791 29894 15837 29946
rect 15837 29894 15847 29946
rect 15871 29894 15901 29946
rect 15901 29894 15913 29946
rect 15913 29894 15927 29946
rect 15951 29894 15965 29946
rect 15965 29894 15977 29946
rect 15977 29894 16007 29946
rect 16031 29894 16041 29946
rect 16041 29894 16087 29946
rect 15791 29892 15847 29894
rect 15871 29892 15927 29894
rect 15951 29892 16007 29894
rect 16031 29892 16087 29894
rect 15791 28858 15847 28860
rect 15871 28858 15927 28860
rect 15951 28858 16007 28860
rect 16031 28858 16087 28860
rect 15791 28806 15837 28858
rect 15837 28806 15847 28858
rect 15871 28806 15901 28858
rect 15901 28806 15913 28858
rect 15913 28806 15927 28858
rect 15951 28806 15965 28858
rect 15965 28806 15977 28858
rect 15977 28806 16007 28858
rect 16031 28806 16041 28858
rect 16041 28806 16087 28858
rect 15791 28804 15847 28806
rect 15871 28804 15927 28806
rect 15951 28804 16007 28806
rect 16031 28804 16087 28806
rect 15750 28056 15806 28112
rect 15791 27770 15847 27772
rect 15871 27770 15927 27772
rect 15951 27770 16007 27772
rect 16031 27770 16087 27772
rect 15791 27718 15837 27770
rect 15837 27718 15847 27770
rect 15871 27718 15901 27770
rect 15901 27718 15913 27770
rect 15913 27718 15927 27770
rect 15951 27718 15965 27770
rect 15965 27718 15977 27770
rect 15977 27718 16007 27770
rect 16031 27718 16041 27770
rect 16041 27718 16087 27770
rect 15791 27716 15847 27718
rect 15871 27716 15927 27718
rect 15951 27716 16007 27718
rect 16031 27716 16087 27718
rect 15791 26682 15847 26684
rect 15871 26682 15927 26684
rect 15951 26682 16007 26684
rect 16031 26682 16087 26684
rect 15791 26630 15837 26682
rect 15837 26630 15847 26682
rect 15871 26630 15901 26682
rect 15901 26630 15913 26682
rect 15913 26630 15927 26682
rect 15951 26630 15965 26682
rect 15965 26630 15977 26682
rect 15977 26630 16007 26682
rect 16031 26630 16041 26682
rect 16041 26630 16087 26682
rect 15791 26628 15847 26630
rect 15871 26628 15927 26630
rect 15951 26628 16007 26630
rect 16031 26628 16087 26630
rect 16762 32544 16818 32600
rect 17958 40568 18014 40624
rect 17038 32428 17094 32464
rect 17038 32408 17040 32428
rect 17040 32408 17092 32428
rect 17092 32408 17094 32428
rect 17222 32952 17278 33008
rect 15658 25744 15714 25800
rect 15791 25594 15847 25596
rect 15871 25594 15927 25596
rect 15951 25594 16007 25596
rect 16031 25594 16087 25596
rect 15791 25542 15837 25594
rect 15837 25542 15847 25594
rect 15871 25542 15901 25594
rect 15901 25542 15913 25594
rect 15913 25542 15927 25594
rect 15951 25542 15965 25594
rect 15965 25542 15977 25594
rect 15977 25542 16007 25594
rect 16031 25542 16041 25594
rect 16041 25542 16087 25594
rect 15791 25540 15847 25542
rect 15871 25540 15927 25542
rect 15951 25540 16007 25542
rect 16031 25540 16087 25542
rect 16394 26152 16450 26208
rect 15791 24506 15847 24508
rect 15871 24506 15927 24508
rect 15951 24506 16007 24508
rect 16031 24506 16087 24508
rect 15791 24454 15837 24506
rect 15837 24454 15847 24506
rect 15871 24454 15901 24506
rect 15901 24454 15913 24506
rect 15913 24454 15927 24506
rect 15951 24454 15965 24506
rect 15965 24454 15977 24506
rect 15977 24454 16007 24506
rect 16031 24454 16041 24506
rect 16041 24454 16087 24506
rect 15791 24452 15847 24454
rect 15871 24452 15927 24454
rect 15951 24452 16007 24454
rect 16031 24452 16087 24454
rect 15791 23418 15847 23420
rect 15871 23418 15927 23420
rect 15951 23418 16007 23420
rect 16031 23418 16087 23420
rect 15791 23366 15837 23418
rect 15837 23366 15847 23418
rect 15871 23366 15901 23418
rect 15901 23366 15913 23418
rect 15913 23366 15927 23418
rect 15951 23366 15965 23418
rect 15965 23366 15977 23418
rect 15977 23366 16007 23418
rect 16031 23366 16041 23418
rect 16041 23366 16087 23418
rect 15791 23364 15847 23366
rect 15871 23364 15927 23366
rect 15951 23364 16007 23366
rect 16031 23364 16087 23366
rect 15791 22330 15847 22332
rect 15871 22330 15927 22332
rect 15951 22330 16007 22332
rect 16031 22330 16087 22332
rect 15791 22278 15837 22330
rect 15837 22278 15847 22330
rect 15871 22278 15901 22330
rect 15901 22278 15913 22330
rect 15913 22278 15927 22330
rect 15951 22278 15965 22330
rect 15965 22278 15977 22330
rect 15977 22278 16007 22330
rect 16031 22278 16041 22330
rect 16041 22278 16087 22330
rect 15791 22276 15847 22278
rect 15871 22276 15927 22278
rect 15951 22276 16007 22278
rect 16031 22276 16087 22278
rect 16118 21392 16174 21448
rect 15474 20712 15530 20768
rect 15198 14456 15254 14512
rect 15791 21242 15847 21244
rect 15871 21242 15927 21244
rect 15951 21242 16007 21244
rect 16031 21242 16087 21244
rect 15791 21190 15837 21242
rect 15837 21190 15847 21242
rect 15871 21190 15901 21242
rect 15901 21190 15913 21242
rect 15913 21190 15927 21242
rect 15951 21190 15965 21242
rect 15965 21190 15977 21242
rect 15977 21190 16007 21242
rect 16031 21190 16041 21242
rect 16041 21190 16087 21242
rect 15791 21188 15847 21190
rect 15871 21188 15927 21190
rect 15951 21188 16007 21190
rect 16031 21188 16087 21190
rect 16118 20848 16174 20904
rect 15791 20154 15847 20156
rect 15871 20154 15927 20156
rect 15951 20154 16007 20156
rect 16031 20154 16087 20156
rect 15791 20102 15837 20154
rect 15837 20102 15847 20154
rect 15871 20102 15901 20154
rect 15901 20102 15913 20154
rect 15913 20102 15927 20154
rect 15951 20102 15965 20154
rect 15965 20102 15977 20154
rect 15977 20102 16007 20154
rect 16031 20102 16041 20154
rect 16041 20102 16087 20154
rect 15791 20100 15847 20102
rect 15871 20100 15927 20102
rect 15951 20100 16007 20102
rect 16031 20100 16087 20102
rect 15750 19216 15806 19272
rect 15791 19066 15847 19068
rect 15871 19066 15927 19068
rect 15951 19066 16007 19068
rect 16031 19066 16087 19068
rect 15791 19014 15837 19066
rect 15837 19014 15847 19066
rect 15871 19014 15901 19066
rect 15901 19014 15913 19066
rect 15913 19014 15927 19066
rect 15951 19014 15965 19066
rect 15965 19014 15977 19066
rect 15977 19014 16007 19066
rect 16031 19014 16041 19066
rect 16041 19014 16087 19066
rect 15791 19012 15847 19014
rect 15871 19012 15927 19014
rect 15951 19012 16007 19014
rect 16031 19012 16087 19014
rect 15934 18128 15990 18184
rect 16118 18128 16174 18184
rect 15791 17978 15847 17980
rect 15871 17978 15927 17980
rect 15951 17978 16007 17980
rect 16031 17978 16087 17980
rect 15791 17926 15837 17978
rect 15837 17926 15847 17978
rect 15871 17926 15901 17978
rect 15901 17926 15913 17978
rect 15913 17926 15927 17978
rect 15951 17926 15965 17978
rect 15965 17926 15977 17978
rect 15977 17926 16007 17978
rect 16031 17926 16041 17978
rect 16041 17926 16087 17978
rect 15791 17924 15847 17926
rect 15871 17924 15927 17926
rect 15951 17924 16007 17926
rect 16031 17924 16087 17926
rect 15791 16890 15847 16892
rect 15871 16890 15927 16892
rect 15951 16890 16007 16892
rect 16031 16890 16087 16892
rect 15791 16838 15837 16890
rect 15837 16838 15847 16890
rect 15871 16838 15901 16890
rect 15901 16838 15913 16890
rect 15913 16838 15927 16890
rect 15951 16838 15965 16890
rect 15965 16838 15977 16890
rect 15977 16838 16007 16890
rect 16031 16838 16041 16890
rect 16041 16838 16087 16890
rect 15791 16836 15847 16838
rect 15871 16836 15927 16838
rect 15951 16836 16007 16838
rect 16031 16836 16087 16838
rect 15791 15802 15847 15804
rect 15871 15802 15927 15804
rect 15951 15802 16007 15804
rect 16031 15802 16087 15804
rect 15791 15750 15837 15802
rect 15837 15750 15847 15802
rect 15871 15750 15901 15802
rect 15901 15750 15913 15802
rect 15913 15750 15927 15802
rect 15951 15750 15965 15802
rect 15965 15750 15977 15802
rect 15977 15750 16007 15802
rect 16031 15750 16041 15802
rect 16041 15750 16087 15802
rect 15791 15748 15847 15750
rect 15871 15748 15927 15750
rect 15951 15748 16007 15750
rect 16031 15748 16087 15750
rect 15791 14714 15847 14716
rect 15871 14714 15927 14716
rect 15951 14714 16007 14716
rect 16031 14714 16087 14716
rect 15791 14662 15837 14714
rect 15837 14662 15847 14714
rect 15871 14662 15901 14714
rect 15901 14662 15913 14714
rect 15913 14662 15927 14714
rect 15951 14662 15965 14714
rect 15965 14662 15977 14714
rect 15977 14662 16007 14714
rect 16031 14662 16041 14714
rect 16041 14662 16087 14714
rect 15791 14660 15847 14662
rect 15871 14660 15927 14662
rect 15951 14660 16007 14662
rect 16031 14660 16087 14662
rect 15791 13626 15847 13628
rect 15871 13626 15927 13628
rect 15951 13626 16007 13628
rect 16031 13626 16087 13628
rect 15791 13574 15837 13626
rect 15837 13574 15847 13626
rect 15871 13574 15901 13626
rect 15901 13574 15913 13626
rect 15913 13574 15927 13626
rect 15951 13574 15965 13626
rect 15965 13574 15977 13626
rect 15977 13574 16007 13626
rect 16031 13574 16041 13626
rect 16041 13574 16087 13626
rect 15791 13572 15847 13574
rect 15871 13572 15927 13574
rect 15951 13572 16007 13574
rect 16031 13572 16087 13574
rect 15290 10512 15346 10568
rect 16762 28736 16818 28792
rect 16854 26832 16910 26888
rect 16670 23432 16726 23488
rect 16394 20984 16450 21040
rect 16578 19760 16634 19816
rect 15791 12538 15847 12540
rect 15871 12538 15927 12540
rect 15951 12538 16007 12540
rect 16031 12538 16087 12540
rect 15791 12486 15837 12538
rect 15837 12486 15847 12538
rect 15871 12486 15901 12538
rect 15901 12486 15913 12538
rect 15913 12486 15927 12538
rect 15951 12486 15965 12538
rect 15965 12486 15977 12538
rect 15977 12486 16007 12538
rect 16031 12486 16041 12538
rect 16041 12486 16087 12538
rect 15791 12484 15847 12486
rect 15871 12484 15927 12486
rect 15951 12484 16007 12486
rect 16031 12484 16087 12486
rect 15791 11450 15847 11452
rect 15871 11450 15927 11452
rect 15951 11450 16007 11452
rect 16031 11450 16087 11452
rect 15791 11398 15837 11450
rect 15837 11398 15847 11450
rect 15871 11398 15901 11450
rect 15901 11398 15913 11450
rect 15913 11398 15927 11450
rect 15951 11398 15965 11450
rect 15965 11398 15977 11450
rect 15977 11398 16007 11450
rect 16031 11398 16041 11450
rect 16041 11398 16087 11450
rect 15791 11396 15847 11398
rect 15871 11396 15927 11398
rect 15951 11396 16007 11398
rect 16031 11396 16087 11398
rect 16026 11192 16082 11248
rect 15791 10362 15847 10364
rect 15871 10362 15927 10364
rect 15951 10362 16007 10364
rect 16031 10362 16087 10364
rect 15791 10310 15837 10362
rect 15837 10310 15847 10362
rect 15871 10310 15901 10362
rect 15901 10310 15913 10362
rect 15913 10310 15927 10362
rect 15951 10310 15965 10362
rect 15965 10310 15977 10362
rect 15977 10310 16007 10362
rect 16031 10310 16041 10362
rect 16041 10310 16087 10362
rect 15791 10308 15847 10310
rect 15871 10308 15927 10310
rect 15951 10308 16007 10310
rect 16031 10308 16087 10310
rect 15791 9274 15847 9276
rect 15871 9274 15927 9276
rect 15951 9274 16007 9276
rect 16031 9274 16087 9276
rect 15791 9222 15837 9274
rect 15837 9222 15847 9274
rect 15871 9222 15901 9274
rect 15901 9222 15913 9274
rect 15913 9222 15927 9274
rect 15951 9222 15965 9274
rect 15965 9222 15977 9274
rect 15977 9222 16007 9274
rect 16031 9222 16041 9274
rect 16041 9222 16087 9274
rect 15791 9220 15847 9222
rect 15871 9220 15927 9222
rect 15951 9220 16007 9222
rect 16031 9220 16087 9222
rect 15791 8186 15847 8188
rect 15871 8186 15927 8188
rect 15951 8186 16007 8188
rect 16031 8186 16087 8188
rect 15791 8134 15837 8186
rect 15837 8134 15847 8186
rect 15871 8134 15901 8186
rect 15901 8134 15913 8186
rect 15913 8134 15927 8186
rect 15951 8134 15965 8186
rect 15965 8134 15977 8186
rect 15977 8134 16007 8186
rect 16031 8134 16041 8186
rect 16041 8134 16087 8186
rect 15791 8132 15847 8134
rect 15871 8132 15927 8134
rect 15951 8132 16007 8134
rect 16031 8132 16087 8134
rect 16670 10104 16726 10160
rect 16578 9968 16634 10024
rect 17866 34604 17922 34640
rect 17866 34584 17868 34604
rect 17868 34584 17920 34604
rect 17920 34584 17922 34604
rect 18234 34856 18290 34912
rect 18142 32816 18198 32872
rect 17498 28328 17554 28384
rect 17866 29164 17922 29200
rect 17866 29144 17868 29164
rect 17868 29144 17920 29164
rect 17920 29144 17922 29164
rect 17774 27648 17830 27704
rect 17222 26832 17278 26888
rect 17406 26832 17462 26888
rect 17222 21936 17278 21992
rect 18758 42458 18814 42460
rect 18838 42458 18894 42460
rect 18918 42458 18974 42460
rect 18998 42458 19054 42460
rect 18758 42406 18804 42458
rect 18804 42406 18814 42458
rect 18838 42406 18868 42458
rect 18868 42406 18880 42458
rect 18880 42406 18894 42458
rect 18918 42406 18932 42458
rect 18932 42406 18944 42458
rect 18944 42406 18974 42458
rect 18998 42406 19008 42458
rect 19008 42406 19054 42458
rect 18758 42404 18814 42406
rect 18838 42404 18894 42406
rect 18918 42404 18974 42406
rect 18998 42404 19054 42406
rect 19062 41792 19118 41848
rect 18694 41556 18696 41576
rect 18696 41556 18748 41576
rect 18748 41556 18750 41576
rect 18694 41520 18750 41556
rect 18758 41370 18814 41372
rect 18838 41370 18894 41372
rect 18918 41370 18974 41372
rect 18998 41370 19054 41372
rect 18758 41318 18804 41370
rect 18804 41318 18814 41370
rect 18838 41318 18868 41370
rect 18868 41318 18880 41370
rect 18880 41318 18894 41370
rect 18918 41318 18932 41370
rect 18932 41318 18944 41370
rect 18944 41318 18974 41370
rect 18998 41318 19008 41370
rect 19008 41318 19054 41370
rect 18758 41316 18814 41318
rect 18838 41316 18894 41318
rect 18918 41316 18974 41318
rect 18998 41316 19054 41318
rect 18758 40282 18814 40284
rect 18838 40282 18894 40284
rect 18918 40282 18974 40284
rect 18998 40282 19054 40284
rect 18758 40230 18804 40282
rect 18804 40230 18814 40282
rect 18838 40230 18868 40282
rect 18868 40230 18880 40282
rect 18880 40230 18894 40282
rect 18918 40230 18932 40282
rect 18932 40230 18944 40282
rect 18944 40230 18974 40282
rect 18998 40230 19008 40282
rect 19008 40230 19054 40282
rect 18758 40228 18814 40230
rect 18838 40228 18894 40230
rect 18918 40228 18974 40230
rect 18998 40228 19054 40230
rect 18758 39194 18814 39196
rect 18838 39194 18894 39196
rect 18918 39194 18974 39196
rect 18998 39194 19054 39196
rect 18758 39142 18804 39194
rect 18804 39142 18814 39194
rect 18838 39142 18868 39194
rect 18868 39142 18880 39194
rect 18880 39142 18894 39194
rect 18918 39142 18932 39194
rect 18932 39142 18944 39194
rect 18944 39142 18974 39194
rect 18998 39142 19008 39194
rect 19008 39142 19054 39194
rect 18758 39140 18814 39142
rect 18838 39140 18894 39142
rect 18918 39140 18974 39142
rect 18998 39140 19054 39142
rect 18326 31592 18382 31648
rect 18234 28872 18290 28928
rect 18142 28736 18198 28792
rect 18234 28328 18290 28384
rect 18418 29144 18474 29200
rect 18234 27920 18290 27976
rect 17222 20712 17278 20768
rect 17130 17176 17186 17232
rect 17498 20440 17554 20496
rect 17682 20304 17738 20360
rect 17590 19488 17646 19544
rect 17222 11076 17278 11112
rect 17222 11056 17224 11076
rect 17224 11056 17276 11076
rect 17276 11056 17278 11076
rect 17682 18264 17738 18320
rect 18758 38106 18814 38108
rect 18838 38106 18894 38108
rect 18918 38106 18974 38108
rect 18998 38106 19054 38108
rect 18758 38054 18804 38106
rect 18804 38054 18814 38106
rect 18838 38054 18868 38106
rect 18868 38054 18880 38106
rect 18880 38054 18894 38106
rect 18918 38054 18932 38106
rect 18932 38054 18944 38106
rect 18944 38054 18974 38106
rect 18998 38054 19008 38106
rect 19008 38054 19054 38106
rect 18758 38052 18814 38054
rect 18838 38052 18894 38054
rect 18918 38052 18974 38054
rect 18998 38052 19054 38054
rect 19338 41964 19340 41984
rect 19340 41964 19392 41984
rect 19392 41964 19394 41984
rect 19338 41928 19394 41964
rect 20258 40568 20314 40624
rect 19890 40160 19946 40216
rect 19430 40024 19486 40080
rect 20166 39888 20222 39944
rect 20074 39480 20130 39536
rect 20534 41248 20590 41304
rect 20994 41384 21050 41440
rect 20534 40704 20590 40760
rect 20902 40976 20958 41032
rect 22098 43152 22154 43208
rect 21362 42064 21418 42120
rect 21725 43002 21781 43004
rect 21805 43002 21861 43004
rect 21885 43002 21941 43004
rect 21965 43002 22021 43004
rect 21725 42950 21771 43002
rect 21771 42950 21781 43002
rect 21805 42950 21835 43002
rect 21835 42950 21847 43002
rect 21847 42950 21861 43002
rect 21885 42950 21899 43002
rect 21899 42950 21911 43002
rect 21911 42950 21941 43002
rect 21965 42950 21975 43002
rect 21975 42950 22021 43002
rect 21725 42948 21781 42950
rect 21805 42948 21861 42950
rect 21885 42948 21941 42950
rect 21965 42948 22021 42950
rect 23018 43832 23074 43888
rect 21725 41914 21781 41916
rect 21805 41914 21861 41916
rect 21885 41914 21941 41916
rect 21965 41914 22021 41916
rect 21725 41862 21771 41914
rect 21771 41862 21781 41914
rect 21805 41862 21835 41914
rect 21835 41862 21847 41914
rect 21847 41862 21861 41914
rect 21885 41862 21899 41914
rect 21899 41862 21911 41914
rect 21911 41862 21941 41914
rect 21965 41862 21975 41914
rect 21975 41862 22021 41914
rect 21725 41860 21781 41862
rect 21805 41860 21861 41862
rect 21885 41860 21941 41862
rect 21965 41860 22021 41862
rect 21086 40432 21142 40488
rect 20902 40024 20958 40080
rect 20810 39208 20866 39264
rect 18758 37018 18814 37020
rect 18838 37018 18894 37020
rect 18918 37018 18974 37020
rect 18998 37018 19054 37020
rect 18758 36966 18804 37018
rect 18804 36966 18814 37018
rect 18838 36966 18868 37018
rect 18868 36966 18880 37018
rect 18880 36966 18894 37018
rect 18918 36966 18932 37018
rect 18932 36966 18944 37018
rect 18944 36966 18974 37018
rect 18998 36966 19008 37018
rect 19008 36966 19054 37018
rect 18758 36964 18814 36966
rect 18838 36964 18894 36966
rect 18918 36964 18974 36966
rect 18998 36964 19054 36966
rect 18758 35930 18814 35932
rect 18838 35930 18894 35932
rect 18918 35930 18974 35932
rect 18998 35930 19054 35932
rect 18758 35878 18804 35930
rect 18804 35878 18814 35930
rect 18838 35878 18868 35930
rect 18868 35878 18880 35930
rect 18880 35878 18894 35930
rect 18918 35878 18932 35930
rect 18932 35878 18944 35930
rect 18944 35878 18974 35930
rect 18998 35878 19008 35930
rect 19008 35878 19054 35930
rect 18758 35876 18814 35878
rect 18838 35876 18894 35878
rect 18918 35876 18974 35878
rect 18998 35876 19054 35878
rect 18758 34842 18814 34844
rect 18838 34842 18894 34844
rect 18918 34842 18974 34844
rect 18998 34842 19054 34844
rect 18758 34790 18804 34842
rect 18804 34790 18814 34842
rect 18838 34790 18868 34842
rect 18868 34790 18880 34842
rect 18880 34790 18894 34842
rect 18918 34790 18932 34842
rect 18932 34790 18944 34842
rect 18944 34790 18974 34842
rect 18998 34790 19008 34842
rect 19008 34790 19054 34842
rect 18758 34788 18814 34790
rect 18838 34788 18894 34790
rect 18918 34788 18974 34790
rect 18998 34788 19054 34790
rect 18758 33754 18814 33756
rect 18838 33754 18894 33756
rect 18918 33754 18974 33756
rect 18998 33754 19054 33756
rect 18758 33702 18804 33754
rect 18804 33702 18814 33754
rect 18838 33702 18868 33754
rect 18868 33702 18880 33754
rect 18880 33702 18894 33754
rect 18918 33702 18932 33754
rect 18932 33702 18944 33754
rect 18944 33702 18974 33754
rect 18998 33702 19008 33754
rect 19008 33702 19054 33754
rect 18758 33700 18814 33702
rect 18838 33700 18894 33702
rect 18918 33700 18974 33702
rect 18998 33700 19054 33702
rect 18758 32666 18814 32668
rect 18838 32666 18894 32668
rect 18918 32666 18974 32668
rect 18998 32666 19054 32668
rect 18758 32614 18804 32666
rect 18804 32614 18814 32666
rect 18838 32614 18868 32666
rect 18868 32614 18880 32666
rect 18880 32614 18894 32666
rect 18918 32614 18932 32666
rect 18932 32614 18944 32666
rect 18944 32614 18974 32666
rect 18998 32614 19008 32666
rect 19008 32614 19054 32666
rect 18758 32612 18814 32614
rect 18838 32612 18894 32614
rect 18918 32612 18974 32614
rect 18998 32612 19054 32614
rect 18758 31578 18814 31580
rect 18838 31578 18894 31580
rect 18918 31578 18974 31580
rect 18998 31578 19054 31580
rect 18758 31526 18804 31578
rect 18804 31526 18814 31578
rect 18838 31526 18868 31578
rect 18868 31526 18880 31578
rect 18880 31526 18894 31578
rect 18918 31526 18932 31578
rect 18932 31526 18944 31578
rect 18944 31526 18974 31578
rect 18998 31526 19008 31578
rect 19008 31526 19054 31578
rect 18758 31524 18814 31526
rect 18838 31524 18894 31526
rect 18918 31524 18974 31526
rect 18998 31524 19054 31526
rect 18758 30490 18814 30492
rect 18838 30490 18894 30492
rect 18918 30490 18974 30492
rect 18998 30490 19054 30492
rect 18758 30438 18804 30490
rect 18804 30438 18814 30490
rect 18838 30438 18868 30490
rect 18868 30438 18880 30490
rect 18880 30438 18894 30490
rect 18918 30438 18932 30490
rect 18932 30438 18944 30490
rect 18944 30438 18974 30490
rect 18998 30438 19008 30490
rect 19008 30438 19054 30490
rect 18758 30436 18814 30438
rect 18838 30436 18894 30438
rect 18918 30436 18974 30438
rect 18998 30436 19054 30438
rect 18758 29402 18814 29404
rect 18838 29402 18894 29404
rect 18918 29402 18974 29404
rect 18998 29402 19054 29404
rect 18758 29350 18804 29402
rect 18804 29350 18814 29402
rect 18838 29350 18868 29402
rect 18868 29350 18880 29402
rect 18880 29350 18894 29402
rect 18918 29350 18932 29402
rect 18932 29350 18944 29402
rect 18944 29350 18974 29402
rect 18998 29350 19008 29402
rect 19008 29350 19054 29402
rect 18758 29348 18814 29350
rect 18838 29348 18894 29350
rect 18918 29348 18974 29350
rect 18998 29348 19054 29350
rect 18694 29008 18750 29064
rect 18602 28620 18658 28656
rect 18602 28600 18604 28620
rect 18604 28600 18656 28620
rect 18656 28600 18658 28620
rect 18234 20848 18290 20904
rect 18050 15136 18106 15192
rect 17774 11736 17830 11792
rect 17222 9696 17278 9752
rect 15791 7098 15847 7100
rect 15871 7098 15927 7100
rect 15951 7098 16007 7100
rect 16031 7098 16087 7100
rect 15791 7046 15837 7098
rect 15837 7046 15847 7098
rect 15871 7046 15901 7098
rect 15901 7046 15913 7098
rect 15913 7046 15927 7098
rect 15951 7046 15965 7098
rect 15965 7046 15977 7098
rect 15977 7046 16007 7098
rect 16031 7046 16041 7098
rect 16041 7046 16087 7098
rect 15791 7044 15847 7046
rect 15871 7044 15927 7046
rect 15951 7044 16007 7046
rect 16031 7044 16087 7046
rect 16302 6296 16358 6352
rect 15791 6010 15847 6012
rect 15871 6010 15927 6012
rect 15951 6010 16007 6012
rect 16031 6010 16087 6012
rect 15791 5958 15837 6010
rect 15837 5958 15847 6010
rect 15871 5958 15901 6010
rect 15901 5958 15913 6010
rect 15913 5958 15927 6010
rect 15951 5958 15965 6010
rect 15965 5958 15977 6010
rect 15977 5958 16007 6010
rect 16031 5958 16041 6010
rect 16041 5958 16087 6010
rect 15791 5956 15847 5958
rect 15871 5956 15927 5958
rect 15951 5956 16007 5958
rect 16031 5956 16087 5958
rect 15791 4922 15847 4924
rect 15871 4922 15927 4924
rect 15951 4922 16007 4924
rect 16031 4922 16087 4924
rect 15791 4870 15837 4922
rect 15837 4870 15847 4922
rect 15871 4870 15901 4922
rect 15901 4870 15913 4922
rect 15913 4870 15927 4922
rect 15951 4870 15965 4922
rect 15965 4870 15977 4922
rect 15977 4870 16007 4922
rect 16031 4870 16041 4922
rect 16041 4870 16087 4922
rect 15791 4868 15847 4870
rect 15871 4868 15927 4870
rect 15951 4868 16007 4870
rect 16031 4868 16087 4870
rect 15791 3834 15847 3836
rect 15871 3834 15927 3836
rect 15951 3834 16007 3836
rect 16031 3834 16087 3836
rect 15791 3782 15837 3834
rect 15837 3782 15847 3834
rect 15871 3782 15901 3834
rect 15901 3782 15913 3834
rect 15913 3782 15927 3834
rect 15951 3782 15965 3834
rect 15965 3782 15977 3834
rect 15977 3782 16007 3834
rect 16031 3782 16041 3834
rect 16041 3782 16087 3834
rect 15791 3780 15847 3782
rect 15871 3780 15927 3782
rect 15951 3780 16007 3782
rect 16031 3780 16087 3782
rect 16302 4528 16358 4584
rect 16670 7112 16726 7168
rect 16486 6704 16542 6760
rect 15791 2746 15847 2748
rect 15871 2746 15927 2748
rect 15951 2746 16007 2748
rect 16031 2746 16087 2748
rect 15791 2694 15837 2746
rect 15837 2694 15847 2746
rect 15871 2694 15901 2746
rect 15901 2694 15913 2746
rect 15913 2694 15927 2746
rect 15951 2694 15965 2746
rect 15965 2694 15977 2746
rect 15977 2694 16007 2746
rect 16031 2694 16041 2746
rect 16041 2694 16087 2746
rect 15791 2692 15847 2694
rect 15871 2692 15927 2694
rect 15951 2692 16007 2694
rect 16031 2692 16087 2694
rect 15474 2624 15530 2680
rect 16854 7928 16910 7984
rect 17498 8744 17554 8800
rect 17406 8336 17462 8392
rect 18758 28314 18814 28316
rect 18838 28314 18894 28316
rect 18918 28314 18974 28316
rect 18998 28314 19054 28316
rect 18758 28262 18804 28314
rect 18804 28262 18814 28314
rect 18838 28262 18868 28314
rect 18868 28262 18880 28314
rect 18880 28262 18894 28314
rect 18918 28262 18932 28314
rect 18932 28262 18944 28314
rect 18944 28262 18974 28314
rect 18998 28262 19008 28314
rect 19008 28262 19054 28314
rect 18758 28260 18814 28262
rect 18838 28260 18894 28262
rect 18918 28260 18974 28262
rect 18998 28260 19054 28262
rect 18786 28092 18788 28112
rect 18788 28092 18840 28112
rect 18840 28092 18842 28112
rect 18786 28056 18842 28092
rect 18758 27226 18814 27228
rect 18838 27226 18894 27228
rect 18918 27226 18974 27228
rect 18998 27226 19054 27228
rect 18758 27174 18804 27226
rect 18804 27174 18814 27226
rect 18838 27174 18868 27226
rect 18868 27174 18880 27226
rect 18880 27174 18894 27226
rect 18918 27174 18932 27226
rect 18932 27174 18944 27226
rect 18944 27174 18974 27226
rect 18998 27174 19008 27226
rect 19008 27174 19054 27226
rect 18758 27172 18814 27174
rect 18838 27172 18894 27174
rect 18918 27172 18974 27174
rect 18998 27172 19054 27174
rect 18758 26138 18814 26140
rect 18838 26138 18894 26140
rect 18918 26138 18974 26140
rect 18998 26138 19054 26140
rect 18758 26086 18804 26138
rect 18804 26086 18814 26138
rect 18838 26086 18868 26138
rect 18868 26086 18880 26138
rect 18880 26086 18894 26138
rect 18918 26086 18932 26138
rect 18932 26086 18944 26138
rect 18944 26086 18974 26138
rect 18998 26086 19008 26138
rect 19008 26086 19054 26138
rect 18758 26084 18814 26086
rect 18838 26084 18894 26086
rect 18918 26084 18974 26086
rect 18998 26084 19054 26086
rect 18758 25050 18814 25052
rect 18838 25050 18894 25052
rect 18918 25050 18974 25052
rect 18998 25050 19054 25052
rect 18758 24998 18804 25050
rect 18804 24998 18814 25050
rect 18838 24998 18868 25050
rect 18868 24998 18880 25050
rect 18880 24998 18894 25050
rect 18918 24998 18932 25050
rect 18932 24998 18944 25050
rect 18944 24998 18974 25050
rect 18998 24998 19008 25050
rect 19008 24998 19054 25050
rect 18758 24996 18814 24998
rect 18838 24996 18894 24998
rect 18918 24996 18974 24998
rect 18998 24996 19054 24998
rect 18758 23962 18814 23964
rect 18838 23962 18894 23964
rect 18918 23962 18974 23964
rect 18998 23962 19054 23964
rect 18758 23910 18804 23962
rect 18804 23910 18814 23962
rect 18838 23910 18868 23962
rect 18868 23910 18880 23962
rect 18880 23910 18894 23962
rect 18918 23910 18932 23962
rect 18932 23910 18944 23962
rect 18944 23910 18974 23962
rect 18998 23910 19008 23962
rect 19008 23910 19054 23962
rect 18758 23908 18814 23910
rect 18838 23908 18894 23910
rect 18918 23908 18974 23910
rect 18998 23908 19054 23910
rect 18786 23568 18842 23624
rect 18694 23432 18750 23488
rect 18758 22874 18814 22876
rect 18838 22874 18894 22876
rect 18918 22874 18974 22876
rect 18998 22874 19054 22876
rect 18758 22822 18804 22874
rect 18804 22822 18814 22874
rect 18838 22822 18868 22874
rect 18868 22822 18880 22874
rect 18880 22822 18894 22874
rect 18918 22822 18932 22874
rect 18932 22822 18944 22874
rect 18944 22822 18974 22874
rect 18998 22822 19008 22874
rect 19008 22822 19054 22874
rect 18758 22820 18814 22822
rect 18838 22820 18894 22822
rect 18918 22820 18974 22822
rect 18998 22820 19054 22822
rect 18758 21786 18814 21788
rect 18838 21786 18894 21788
rect 18918 21786 18974 21788
rect 18998 21786 19054 21788
rect 18758 21734 18804 21786
rect 18804 21734 18814 21786
rect 18838 21734 18868 21786
rect 18868 21734 18880 21786
rect 18880 21734 18894 21786
rect 18918 21734 18932 21786
rect 18932 21734 18944 21786
rect 18944 21734 18974 21786
rect 18998 21734 19008 21786
rect 19008 21734 19054 21786
rect 18758 21732 18814 21734
rect 18838 21732 18894 21734
rect 18918 21732 18974 21734
rect 18998 21732 19054 21734
rect 18970 21004 19026 21040
rect 18970 20984 18972 21004
rect 18972 20984 19024 21004
rect 19024 20984 19026 21004
rect 19062 20848 19118 20904
rect 18758 20698 18814 20700
rect 18838 20698 18894 20700
rect 18918 20698 18974 20700
rect 18998 20698 19054 20700
rect 18758 20646 18804 20698
rect 18804 20646 18814 20698
rect 18838 20646 18868 20698
rect 18868 20646 18880 20698
rect 18880 20646 18894 20698
rect 18918 20646 18932 20698
rect 18932 20646 18944 20698
rect 18944 20646 18974 20698
rect 18998 20646 19008 20698
rect 19008 20646 19054 20698
rect 18758 20644 18814 20646
rect 18838 20644 18894 20646
rect 18918 20644 18974 20646
rect 18998 20644 19054 20646
rect 18758 19610 18814 19612
rect 18838 19610 18894 19612
rect 18918 19610 18974 19612
rect 18998 19610 19054 19612
rect 18758 19558 18804 19610
rect 18804 19558 18814 19610
rect 18838 19558 18868 19610
rect 18868 19558 18880 19610
rect 18880 19558 18894 19610
rect 18918 19558 18932 19610
rect 18932 19558 18944 19610
rect 18944 19558 18974 19610
rect 18998 19558 19008 19610
rect 19008 19558 19054 19610
rect 18758 19556 18814 19558
rect 18838 19556 18894 19558
rect 18918 19556 18974 19558
rect 18998 19556 19054 19558
rect 18326 17176 18382 17232
rect 17682 3984 17738 4040
rect 16026 2488 16082 2544
rect 15791 1658 15847 1660
rect 15871 1658 15927 1660
rect 15951 1658 16007 1660
rect 16031 1658 16087 1660
rect 15791 1606 15837 1658
rect 15837 1606 15847 1658
rect 15871 1606 15901 1658
rect 15901 1606 15913 1658
rect 15913 1606 15927 1658
rect 15951 1606 15965 1658
rect 15965 1606 15977 1658
rect 15977 1606 16007 1658
rect 16031 1606 16041 1658
rect 16041 1606 16087 1658
rect 15791 1604 15847 1606
rect 15871 1604 15927 1606
rect 15951 1604 16007 1606
rect 16031 1604 16087 1606
rect 16946 2508 17002 2544
rect 16946 2488 16948 2508
rect 16948 2488 17000 2508
rect 17000 2488 17002 2508
rect 16486 1300 16488 1320
rect 16488 1300 16540 1320
rect 16540 1300 16542 1320
rect 16486 1264 16542 1300
rect 17866 3460 17922 3496
rect 17866 3440 17868 3460
rect 17868 3440 17920 3460
rect 17920 3440 17922 3460
rect 18326 12316 18328 12336
rect 18328 12316 18380 12336
rect 18380 12316 18382 12336
rect 18326 12280 18382 12316
rect 18326 9036 18382 9072
rect 18326 9016 18328 9036
rect 18328 9016 18380 9036
rect 18380 9016 18382 9036
rect 18418 7148 18420 7168
rect 18420 7148 18472 7168
rect 18472 7148 18474 7168
rect 18418 7112 18474 7148
rect 18758 18522 18814 18524
rect 18838 18522 18894 18524
rect 18918 18522 18974 18524
rect 18998 18522 19054 18524
rect 18758 18470 18804 18522
rect 18804 18470 18814 18522
rect 18838 18470 18868 18522
rect 18868 18470 18880 18522
rect 18880 18470 18894 18522
rect 18918 18470 18932 18522
rect 18932 18470 18944 18522
rect 18944 18470 18974 18522
rect 18998 18470 19008 18522
rect 19008 18470 19054 18522
rect 18758 18468 18814 18470
rect 18838 18468 18894 18470
rect 18918 18468 18974 18470
rect 18998 18468 19054 18470
rect 18758 17434 18814 17436
rect 18838 17434 18894 17436
rect 18918 17434 18974 17436
rect 18998 17434 19054 17436
rect 18758 17382 18804 17434
rect 18804 17382 18814 17434
rect 18838 17382 18868 17434
rect 18868 17382 18880 17434
rect 18880 17382 18894 17434
rect 18918 17382 18932 17434
rect 18932 17382 18944 17434
rect 18944 17382 18974 17434
rect 18998 17382 19008 17434
rect 19008 17382 19054 17434
rect 18758 17380 18814 17382
rect 18838 17380 18894 17382
rect 18918 17380 18974 17382
rect 18998 17380 19054 17382
rect 18758 16346 18814 16348
rect 18838 16346 18894 16348
rect 18918 16346 18974 16348
rect 18998 16346 19054 16348
rect 18758 16294 18804 16346
rect 18804 16294 18814 16346
rect 18838 16294 18868 16346
rect 18868 16294 18880 16346
rect 18880 16294 18894 16346
rect 18918 16294 18932 16346
rect 18932 16294 18944 16346
rect 18944 16294 18974 16346
rect 18998 16294 19008 16346
rect 19008 16294 19054 16346
rect 18758 16292 18814 16294
rect 18838 16292 18894 16294
rect 18918 16292 18974 16294
rect 18998 16292 19054 16294
rect 18758 15258 18814 15260
rect 18838 15258 18894 15260
rect 18918 15258 18974 15260
rect 18998 15258 19054 15260
rect 18758 15206 18804 15258
rect 18804 15206 18814 15258
rect 18838 15206 18868 15258
rect 18868 15206 18880 15258
rect 18880 15206 18894 15258
rect 18918 15206 18932 15258
rect 18932 15206 18944 15258
rect 18944 15206 18974 15258
rect 18998 15206 19008 15258
rect 19008 15206 19054 15258
rect 18758 15204 18814 15206
rect 18838 15204 18894 15206
rect 18918 15204 18974 15206
rect 18998 15204 19054 15206
rect 19338 25200 19394 25256
rect 19614 28192 19670 28248
rect 21270 40604 21272 40624
rect 21272 40604 21324 40624
rect 21324 40604 21326 40624
rect 21270 40568 21326 40604
rect 21454 40704 21510 40760
rect 21270 40432 21326 40488
rect 22006 41556 22008 41576
rect 22008 41556 22060 41576
rect 22060 41556 22062 41576
rect 22006 41520 22062 41556
rect 22190 41656 22246 41712
rect 22282 41132 22338 41168
rect 22282 41112 22284 41132
rect 22284 41112 22336 41132
rect 22336 41112 22338 41132
rect 21725 40826 21781 40828
rect 21805 40826 21861 40828
rect 21885 40826 21941 40828
rect 21965 40826 22021 40828
rect 21725 40774 21771 40826
rect 21771 40774 21781 40826
rect 21805 40774 21835 40826
rect 21835 40774 21847 40826
rect 21847 40774 21861 40826
rect 21885 40774 21899 40826
rect 21899 40774 21911 40826
rect 21911 40774 21941 40826
rect 21965 40774 21975 40826
rect 21975 40774 22021 40826
rect 21725 40772 21781 40774
rect 21805 40772 21861 40774
rect 21885 40772 21941 40774
rect 21965 40772 22021 40774
rect 22098 40296 22154 40352
rect 22466 41384 22522 41440
rect 22650 40976 22706 41032
rect 22282 40468 22284 40488
rect 22284 40468 22336 40488
rect 22336 40468 22338 40488
rect 22282 40432 22338 40468
rect 21730 40060 21732 40080
rect 21732 40060 21784 40080
rect 21784 40060 21786 40080
rect 21730 40024 21786 40060
rect 21725 39738 21781 39740
rect 21805 39738 21861 39740
rect 21885 39738 21941 39740
rect 21965 39738 22021 39740
rect 21725 39686 21771 39738
rect 21771 39686 21781 39738
rect 21805 39686 21835 39738
rect 21835 39686 21847 39738
rect 21847 39686 21861 39738
rect 21885 39686 21899 39738
rect 21899 39686 21911 39738
rect 21911 39686 21941 39738
rect 21965 39686 21975 39738
rect 21975 39686 22021 39738
rect 21725 39684 21781 39686
rect 21805 39684 21861 39686
rect 21885 39684 21941 39686
rect 21965 39684 22021 39686
rect 21362 39344 21418 39400
rect 22282 39364 22338 39400
rect 22282 39344 22284 39364
rect 22284 39344 22336 39364
rect 22336 39344 22338 39364
rect 22466 39380 22468 39400
rect 22468 39380 22520 39400
rect 22520 39380 22522 39400
rect 22466 39344 22522 39380
rect 21270 38664 21326 38720
rect 21725 38650 21781 38652
rect 21805 38650 21861 38652
rect 21885 38650 21941 38652
rect 21965 38650 22021 38652
rect 21725 38598 21771 38650
rect 21771 38598 21781 38650
rect 21805 38598 21835 38650
rect 21835 38598 21847 38650
rect 21847 38598 21861 38650
rect 21885 38598 21899 38650
rect 21899 38598 21911 38650
rect 21911 38598 21941 38650
rect 21965 38598 21975 38650
rect 21975 38598 22021 38650
rect 21725 38596 21781 38598
rect 21805 38596 21861 38598
rect 21885 38596 21941 38598
rect 21965 38596 22021 38598
rect 21725 37562 21781 37564
rect 21805 37562 21861 37564
rect 21885 37562 21941 37564
rect 21965 37562 22021 37564
rect 21725 37510 21771 37562
rect 21771 37510 21781 37562
rect 21805 37510 21835 37562
rect 21835 37510 21847 37562
rect 21847 37510 21861 37562
rect 21885 37510 21899 37562
rect 21899 37510 21911 37562
rect 21911 37510 21941 37562
rect 21965 37510 21975 37562
rect 21975 37510 22021 37562
rect 21725 37508 21781 37510
rect 21805 37508 21861 37510
rect 21885 37508 21941 37510
rect 21965 37508 22021 37510
rect 20626 35028 20628 35048
rect 20628 35028 20680 35048
rect 20680 35028 20682 35048
rect 20626 34992 20682 35028
rect 20442 30368 20498 30424
rect 21725 36474 21781 36476
rect 21805 36474 21861 36476
rect 21885 36474 21941 36476
rect 21965 36474 22021 36476
rect 21725 36422 21771 36474
rect 21771 36422 21781 36474
rect 21805 36422 21835 36474
rect 21835 36422 21847 36474
rect 21847 36422 21861 36474
rect 21885 36422 21899 36474
rect 21899 36422 21911 36474
rect 21911 36422 21941 36474
rect 21965 36422 21975 36474
rect 21975 36422 22021 36474
rect 21725 36420 21781 36422
rect 21805 36420 21861 36422
rect 21885 36420 21941 36422
rect 21965 36420 22021 36422
rect 21725 35386 21781 35388
rect 21805 35386 21861 35388
rect 21885 35386 21941 35388
rect 21965 35386 22021 35388
rect 21725 35334 21771 35386
rect 21771 35334 21781 35386
rect 21805 35334 21835 35386
rect 21835 35334 21847 35386
rect 21847 35334 21861 35386
rect 21885 35334 21899 35386
rect 21899 35334 21911 35386
rect 21911 35334 21941 35386
rect 21965 35334 21975 35386
rect 21975 35334 22021 35386
rect 21725 35332 21781 35334
rect 21805 35332 21861 35334
rect 21885 35332 21941 35334
rect 21965 35332 22021 35334
rect 20534 28212 20590 28248
rect 20534 28192 20536 28212
rect 20536 28192 20588 28212
rect 20588 28192 20590 28212
rect 20718 27648 20774 27704
rect 19430 17312 19486 17368
rect 20994 30232 21050 30288
rect 21725 34298 21781 34300
rect 21805 34298 21861 34300
rect 21885 34298 21941 34300
rect 21965 34298 22021 34300
rect 21725 34246 21771 34298
rect 21771 34246 21781 34298
rect 21805 34246 21835 34298
rect 21835 34246 21847 34298
rect 21847 34246 21861 34298
rect 21885 34246 21899 34298
rect 21899 34246 21911 34298
rect 21911 34246 21941 34298
rect 21965 34246 21975 34298
rect 21975 34246 22021 34298
rect 21725 34244 21781 34246
rect 21805 34244 21861 34246
rect 21885 34244 21941 34246
rect 21965 34244 22021 34246
rect 21725 33210 21781 33212
rect 21805 33210 21861 33212
rect 21885 33210 21941 33212
rect 21965 33210 22021 33212
rect 21725 33158 21771 33210
rect 21771 33158 21781 33210
rect 21805 33158 21835 33210
rect 21835 33158 21847 33210
rect 21847 33158 21861 33210
rect 21885 33158 21899 33210
rect 21899 33158 21911 33210
rect 21911 33158 21941 33210
rect 21965 33158 21975 33210
rect 21975 33158 22021 33210
rect 21725 33156 21781 33158
rect 21805 33156 21861 33158
rect 21885 33156 21941 33158
rect 21965 33156 22021 33158
rect 21546 33088 21602 33144
rect 21362 24656 21418 24712
rect 19430 14864 19486 14920
rect 18758 14170 18814 14172
rect 18838 14170 18894 14172
rect 18918 14170 18974 14172
rect 18998 14170 19054 14172
rect 18758 14118 18804 14170
rect 18804 14118 18814 14170
rect 18838 14118 18868 14170
rect 18868 14118 18880 14170
rect 18880 14118 18894 14170
rect 18918 14118 18932 14170
rect 18932 14118 18944 14170
rect 18944 14118 18974 14170
rect 18998 14118 19008 14170
rect 19008 14118 19054 14170
rect 18758 14116 18814 14118
rect 18838 14116 18894 14118
rect 18918 14116 18974 14118
rect 18998 14116 19054 14118
rect 18758 13082 18814 13084
rect 18838 13082 18894 13084
rect 18918 13082 18974 13084
rect 18998 13082 19054 13084
rect 18758 13030 18804 13082
rect 18804 13030 18814 13082
rect 18838 13030 18868 13082
rect 18868 13030 18880 13082
rect 18880 13030 18894 13082
rect 18918 13030 18932 13082
rect 18932 13030 18944 13082
rect 18944 13030 18974 13082
rect 18998 13030 19008 13082
rect 19008 13030 19054 13082
rect 18758 13028 18814 13030
rect 18838 13028 18894 13030
rect 18918 13028 18974 13030
rect 18998 13028 19054 13030
rect 18758 11994 18814 11996
rect 18838 11994 18894 11996
rect 18918 11994 18974 11996
rect 18998 11994 19054 11996
rect 18758 11942 18804 11994
rect 18804 11942 18814 11994
rect 18838 11942 18868 11994
rect 18868 11942 18880 11994
rect 18880 11942 18894 11994
rect 18918 11942 18932 11994
rect 18932 11942 18944 11994
rect 18944 11942 18974 11994
rect 18998 11942 19008 11994
rect 19008 11942 19054 11994
rect 18758 11940 18814 11942
rect 18838 11940 18894 11942
rect 18918 11940 18974 11942
rect 18998 11940 19054 11942
rect 18758 10906 18814 10908
rect 18838 10906 18894 10908
rect 18918 10906 18974 10908
rect 18998 10906 19054 10908
rect 18758 10854 18804 10906
rect 18804 10854 18814 10906
rect 18838 10854 18868 10906
rect 18868 10854 18880 10906
rect 18880 10854 18894 10906
rect 18918 10854 18932 10906
rect 18932 10854 18944 10906
rect 18944 10854 18974 10906
rect 18998 10854 19008 10906
rect 19008 10854 19054 10906
rect 18758 10852 18814 10854
rect 18838 10852 18894 10854
rect 18918 10852 18974 10854
rect 18998 10852 19054 10854
rect 18758 9818 18814 9820
rect 18838 9818 18894 9820
rect 18918 9818 18974 9820
rect 18998 9818 19054 9820
rect 18758 9766 18804 9818
rect 18804 9766 18814 9818
rect 18838 9766 18868 9818
rect 18868 9766 18880 9818
rect 18880 9766 18894 9818
rect 18918 9766 18932 9818
rect 18932 9766 18944 9818
rect 18944 9766 18974 9818
rect 18998 9766 19008 9818
rect 19008 9766 19054 9818
rect 18758 9764 18814 9766
rect 18838 9764 18894 9766
rect 18918 9764 18974 9766
rect 18998 9764 19054 9766
rect 18758 8730 18814 8732
rect 18838 8730 18894 8732
rect 18918 8730 18974 8732
rect 18998 8730 19054 8732
rect 18758 8678 18804 8730
rect 18804 8678 18814 8730
rect 18838 8678 18868 8730
rect 18868 8678 18880 8730
rect 18880 8678 18894 8730
rect 18918 8678 18932 8730
rect 18932 8678 18944 8730
rect 18944 8678 18974 8730
rect 18998 8678 19008 8730
rect 19008 8678 19054 8730
rect 18758 8676 18814 8678
rect 18838 8676 18894 8678
rect 18918 8676 18974 8678
rect 18998 8676 19054 8678
rect 18758 7642 18814 7644
rect 18838 7642 18894 7644
rect 18918 7642 18974 7644
rect 18998 7642 19054 7644
rect 18758 7590 18804 7642
rect 18804 7590 18814 7642
rect 18838 7590 18868 7642
rect 18868 7590 18880 7642
rect 18880 7590 18894 7642
rect 18918 7590 18932 7642
rect 18932 7590 18944 7642
rect 18944 7590 18974 7642
rect 18998 7590 19008 7642
rect 19008 7590 19054 7642
rect 18758 7588 18814 7590
rect 18838 7588 18894 7590
rect 18918 7588 18974 7590
rect 18998 7588 19054 7590
rect 18758 6554 18814 6556
rect 18838 6554 18894 6556
rect 18918 6554 18974 6556
rect 18998 6554 19054 6556
rect 18758 6502 18804 6554
rect 18804 6502 18814 6554
rect 18838 6502 18868 6554
rect 18868 6502 18880 6554
rect 18880 6502 18894 6554
rect 18918 6502 18932 6554
rect 18932 6502 18944 6554
rect 18944 6502 18974 6554
rect 18998 6502 19008 6554
rect 19008 6502 19054 6554
rect 18758 6500 18814 6502
rect 18838 6500 18894 6502
rect 18918 6500 18974 6502
rect 18998 6500 19054 6502
rect 18758 5466 18814 5468
rect 18838 5466 18894 5468
rect 18918 5466 18974 5468
rect 18998 5466 19054 5468
rect 18758 5414 18804 5466
rect 18804 5414 18814 5466
rect 18838 5414 18868 5466
rect 18868 5414 18880 5466
rect 18880 5414 18894 5466
rect 18918 5414 18932 5466
rect 18932 5414 18944 5466
rect 18944 5414 18974 5466
rect 18998 5414 19008 5466
rect 19008 5414 19054 5466
rect 18758 5412 18814 5414
rect 18838 5412 18894 5414
rect 18918 5412 18974 5414
rect 18998 5412 19054 5414
rect 18758 4378 18814 4380
rect 18838 4378 18894 4380
rect 18918 4378 18974 4380
rect 18998 4378 19054 4380
rect 18758 4326 18804 4378
rect 18804 4326 18814 4378
rect 18838 4326 18868 4378
rect 18868 4326 18880 4378
rect 18880 4326 18894 4378
rect 18918 4326 18932 4378
rect 18932 4326 18944 4378
rect 18944 4326 18974 4378
rect 18998 4326 19008 4378
rect 19008 4326 19054 4378
rect 18758 4324 18814 4326
rect 18838 4324 18894 4326
rect 18918 4324 18974 4326
rect 18998 4324 19054 4326
rect 19706 5208 19762 5264
rect 19522 4256 19578 4312
rect 19338 4120 19394 4176
rect 17498 2624 17554 2680
rect 18510 2488 18566 2544
rect 18758 3290 18814 3292
rect 18838 3290 18894 3292
rect 18918 3290 18974 3292
rect 18998 3290 19054 3292
rect 18758 3238 18804 3290
rect 18804 3238 18814 3290
rect 18838 3238 18868 3290
rect 18868 3238 18880 3290
rect 18880 3238 18894 3290
rect 18918 3238 18932 3290
rect 18932 3238 18944 3290
rect 18944 3238 18974 3290
rect 18998 3238 19008 3290
rect 19008 3238 19054 3290
rect 18758 3236 18814 3238
rect 18838 3236 18894 3238
rect 18918 3236 18974 3238
rect 18998 3236 19054 3238
rect 19246 3712 19302 3768
rect 18878 2624 18934 2680
rect 18758 2202 18814 2204
rect 18838 2202 18894 2204
rect 18918 2202 18974 2204
rect 18998 2202 19054 2204
rect 18758 2150 18804 2202
rect 18804 2150 18814 2202
rect 18838 2150 18868 2202
rect 18868 2150 18880 2202
rect 18880 2150 18894 2202
rect 18918 2150 18932 2202
rect 18932 2150 18944 2202
rect 18944 2150 18974 2202
rect 18998 2150 19008 2202
rect 19008 2150 19054 2202
rect 18758 2148 18814 2150
rect 18838 2148 18894 2150
rect 18918 2148 18974 2150
rect 18998 2148 19054 2150
rect 18510 1300 18512 1320
rect 18512 1300 18564 1320
rect 18564 1300 18566 1320
rect 18510 1264 18566 1300
rect 18758 1114 18814 1116
rect 18838 1114 18894 1116
rect 18918 1114 18974 1116
rect 18998 1114 19054 1116
rect 18758 1062 18804 1114
rect 18804 1062 18814 1114
rect 18838 1062 18868 1114
rect 18868 1062 18880 1114
rect 18880 1062 18894 1114
rect 18918 1062 18932 1114
rect 18932 1062 18944 1114
rect 18944 1062 18974 1114
rect 18998 1062 19008 1114
rect 19008 1062 19054 1114
rect 18758 1060 18814 1062
rect 18838 1060 18894 1062
rect 18918 1060 18974 1062
rect 18998 1060 19054 1062
rect 19522 3848 19578 3904
rect 19706 3848 19762 3904
rect 19522 3340 19524 3360
rect 19524 3340 19576 3360
rect 19576 3340 19578 3360
rect 19522 3304 19578 3340
rect 19890 3984 19946 4040
rect 19522 3032 19578 3088
rect 19338 2760 19394 2816
rect 19246 2624 19302 2680
rect 19522 2624 19578 2680
rect 19614 2352 19670 2408
rect 20166 4428 20168 4448
rect 20168 4428 20220 4448
rect 20220 4428 20222 4448
rect 20166 4392 20222 4428
rect 20074 2352 20130 2408
rect 20810 21936 20866 21992
rect 20626 18672 20682 18728
rect 20626 12824 20682 12880
rect 21362 17992 21418 18048
rect 21725 32122 21781 32124
rect 21805 32122 21861 32124
rect 21885 32122 21941 32124
rect 21965 32122 22021 32124
rect 21725 32070 21771 32122
rect 21771 32070 21781 32122
rect 21805 32070 21835 32122
rect 21835 32070 21847 32122
rect 21847 32070 21861 32122
rect 21885 32070 21899 32122
rect 21899 32070 21911 32122
rect 21911 32070 21941 32122
rect 21965 32070 21975 32122
rect 21975 32070 22021 32122
rect 21725 32068 21781 32070
rect 21805 32068 21861 32070
rect 21885 32068 21941 32070
rect 21965 32068 22021 32070
rect 23110 42744 23166 42800
rect 23662 43288 23718 43344
rect 23202 41656 23258 41712
rect 23018 36080 23074 36136
rect 21725 31034 21781 31036
rect 21805 31034 21861 31036
rect 21885 31034 21941 31036
rect 21965 31034 22021 31036
rect 21725 30982 21771 31034
rect 21771 30982 21781 31034
rect 21805 30982 21835 31034
rect 21835 30982 21847 31034
rect 21847 30982 21861 31034
rect 21885 30982 21899 31034
rect 21899 30982 21911 31034
rect 21911 30982 21941 31034
rect 21965 30982 21975 31034
rect 21975 30982 22021 31034
rect 21725 30980 21781 30982
rect 21805 30980 21861 30982
rect 21885 30980 21941 30982
rect 21965 30980 22021 30982
rect 21725 29946 21781 29948
rect 21805 29946 21861 29948
rect 21885 29946 21941 29948
rect 21965 29946 22021 29948
rect 21725 29894 21771 29946
rect 21771 29894 21781 29946
rect 21805 29894 21835 29946
rect 21835 29894 21847 29946
rect 21847 29894 21861 29946
rect 21885 29894 21899 29946
rect 21899 29894 21911 29946
rect 21911 29894 21941 29946
rect 21965 29894 21975 29946
rect 21975 29894 22021 29946
rect 21725 29892 21781 29894
rect 21805 29892 21861 29894
rect 21885 29892 21941 29894
rect 21965 29892 22021 29894
rect 21730 29144 21786 29200
rect 21638 29008 21694 29064
rect 21725 28858 21781 28860
rect 21805 28858 21861 28860
rect 21885 28858 21941 28860
rect 21965 28858 22021 28860
rect 21725 28806 21771 28858
rect 21771 28806 21781 28858
rect 21805 28806 21835 28858
rect 21835 28806 21847 28858
rect 21847 28806 21861 28858
rect 21885 28806 21899 28858
rect 21899 28806 21911 28858
rect 21911 28806 21941 28858
rect 21965 28806 21975 28858
rect 21975 28806 22021 28858
rect 21725 28804 21781 28806
rect 21805 28804 21861 28806
rect 21885 28804 21941 28806
rect 21965 28804 22021 28806
rect 22466 29144 22522 29200
rect 21725 27770 21781 27772
rect 21805 27770 21861 27772
rect 21885 27770 21941 27772
rect 21965 27770 22021 27772
rect 21725 27718 21771 27770
rect 21771 27718 21781 27770
rect 21805 27718 21835 27770
rect 21835 27718 21847 27770
rect 21847 27718 21861 27770
rect 21885 27718 21899 27770
rect 21899 27718 21911 27770
rect 21911 27718 21941 27770
rect 21965 27718 21975 27770
rect 21975 27718 22021 27770
rect 21725 27716 21781 27718
rect 21805 27716 21861 27718
rect 21885 27716 21941 27718
rect 21965 27716 22021 27718
rect 21725 26682 21781 26684
rect 21805 26682 21861 26684
rect 21885 26682 21941 26684
rect 21965 26682 22021 26684
rect 21725 26630 21771 26682
rect 21771 26630 21781 26682
rect 21805 26630 21835 26682
rect 21835 26630 21847 26682
rect 21847 26630 21861 26682
rect 21885 26630 21899 26682
rect 21899 26630 21911 26682
rect 21911 26630 21941 26682
rect 21965 26630 21975 26682
rect 21975 26630 22021 26682
rect 21725 26628 21781 26630
rect 21805 26628 21861 26630
rect 21885 26628 21941 26630
rect 21965 26628 22021 26630
rect 21725 25594 21781 25596
rect 21805 25594 21861 25596
rect 21885 25594 21941 25596
rect 21965 25594 22021 25596
rect 21725 25542 21771 25594
rect 21771 25542 21781 25594
rect 21805 25542 21835 25594
rect 21835 25542 21847 25594
rect 21847 25542 21861 25594
rect 21885 25542 21899 25594
rect 21899 25542 21911 25594
rect 21911 25542 21941 25594
rect 21965 25542 21975 25594
rect 21975 25542 22021 25594
rect 21725 25540 21781 25542
rect 21805 25540 21861 25542
rect 21885 25540 21941 25542
rect 21965 25540 22021 25542
rect 21725 24506 21781 24508
rect 21805 24506 21861 24508
rect 21885 24506 21941 24508
rect 21965 24506 22021 24508
rect 21725 24454 21771 24506
rect 21771 24454 21781 24506
rect 21805 24454 21835 24506
rect 21835 24454 21847 24506
rect 21847 24454 21861 24506
rect 21885 24454 21899 24506
rect 21899 24454 21911 24506
rect 21911 24454 21941 24506
rect 21965 24454 21975 24506
rect 21975 24454 22021 24506
rect 21725 24452 21781 24454
rect 21805 24452 21861 24454
rect 21885 24452 21941 24454
rect 21965 24452 22021 24454
rect 21725 23418 21781 23420
rect 21805 23418 21861 23420
rect 21885 23418 21941 23420
rect 21965 23418 22021 23420
rect 21725 23366 21771 23418
rect 21771 23366 21781 23418
rect 21805 23366 21835 23418
rect 21835 23366 21847 23418
rect 21847 23366 21861 23418
rect 21885 23366 21899 23418
rect 21899 23366 21911 23418
rect 21911 23366 21941 23418
rect 21965 23366 21975 23418
rect 21975 23366 22021 23418
rect 21725 23364 21781 23366
rect 21805 23364 21861 23366
rect 21885 23364 21941 23366
rect 21965 23364 22021 23366
rect 21725 22330 21781 22332
rect 21805 22330 21861 22332
rect 21885 22330 21941 22332
rect 21965 22330 22021 22332
rect 21725 22278 21771 22330
rect 21771 22278 21781 22330
rect 21805 22278 21835 22330
rect 21835 22278 21847 22330
rect 21847 22278 21861 22330
rect 21885 22278 21899 22330
rect 21899 22278 21911 22330
rect 21911 22278 21941 22330
rect 21965 22278 21975 22330
rect 21975 22278 22021 22330
rect 21725 22276 21781 22278
rect 21805 22276 21861 22278
rect 21885 22276 21941 22278
rect 21965 22276 22021 22278
rect 21725 21242 21781 21244
rect 21805 21242 21861 21244
rect 21885 21242 21941 21244
rect 21965 21242 22021 21244
rect 21725 21190 21771 21242
rect 21771 21190 21781 21242
rect 21805 21190 21835 21242
rect 21835 21190 21847 21242
rect 21847 21190 21861 21242
rect 21885 21190 21899 21242
rect 21899 21190 21911 21242
rect 21911 21190 21941 21242
rect 21965 21190 21975 21242
rect 21975 21190 22021 21242
rect 21725 21188 21781 21190
rect 21805 21188 21861 21190
rect 21885 21188 21941 21190
rect 21965 21188 22021 21190
rect 21725 20154 21781 20156
rect 21805 20154 21861 20156
rect 21885 20154 21941 20156
rect 21965 20154 22021 20156
rect 21725 20102 21771 20154
rect 21771 20102 21781 20154
rect 21805 20102 21835 20154
rect 21835 20102 21847 20154
rect 21847 20102 21861 20154
rect 21885 20102 21899 20154
rect 21899 20102 21911 20154
rect 21911 20102 21941 20154
rect 21965 20102 21975 20154
rect 21975 20102 22021 20154
rect 21725 20100 21781 20102
rect 21805 20100 21861 20102
rect 21885 20100 21941 20102
rect 21965 20100 22021 20102
rect 21725 19066 21781 19068
rect 21805 19066 21861 19068
rect 21885 19066 21941 19068
rect 21965 19066 22021 19068
rect 21725 19014 21771 19066
rect 21771 19014 21781 19066
rect 21805 19014 21835 19066
rect 21835 19014 21847 19066
rect 21847 19014 21861 19066
rect 21885 19014 21899 19066
rect 21899 19014 21911 19066
rect 21911 19014 21941 19066
rect 21965 19014 21975 19066
rect 21975 19014 22021 19066
rect 21725 19012 21781 19014
rect 21805 19012 21861 19014
rect 21885 19012 21941 19014
rect 21965 19012 22021 19014
rect 21725 17978 21781 17980
rect 21805 17978 21861 17980
rect 21885 17978 21941 17980
rect 21965 17978 22021 17980
rect 21725 17926 21771 17978
rect 21771 17926 21781 17978
rect 21805 17926 21835 17978
rect 21835 17926 21847 17978
rect 21847 17926 21861 17978
rect 21885 17926 21899 17978
rect 21899 17926 21911 17978
rect 21911 17926 21941 17978
rect 21965 17926 21975 17978
rect 21975 17926 22021 17978
rect 21725 17924 21781 17926
rect 21805 17924 21861 17926
rect 21885 17924 21941 17926
rect 21965 17924 22021 17926
rect 21725 16890 21781 16892
rect 21805 16890 21861 16892
rect 21885 16890 21941 16892
rect 21965 16890 22021 16892
rect 21725 16838 21771 16890
rect 21771 16838 21781 16890
rect 21805 16838 21835 16890
rect 21835 16838 21847 16890
rect 21847 16838 21861 16890
rect 21885 16838 21899 16890
rect 21899 16838 21911 16890
rect 21911 16838 21941 16890
rect 21965 16838 21975 16890
rect 21975 16838 22021 16890
rect 21725 16836 21781 16838
rect 21805 16836 21861 16838
rect 21885 16836 21941 16838
rect 21965 16836 22021 16838
rect 21725 15802 21781 15804
rect 21805 15802 21861 15804
rect 21885 15802 21941 15804
rect 21965 15802 22021 15804
rect 21725 15750 21771 15802
rect 21771 15750 21781 15802
rect 21805 15750 21835 15802
rect 21835 15750 21847 15802
rect 21847 15750 21861 15802
rect 21885 15750 21899 15802
rect 21899 15750 21911 15802
rect 21911 15750 21941 15802
rect 21965 15750 21975 15802
rect 21975 15750 22021 15802
rect 21725 15748 21781 15750
rect 21805 15748 21861 15750
rect 21885 15748 21941 15750
rect 21965 15748 22021 15750
rect 21725 14714 21781 14716
rect 21805 14714 21861 14716
rect 21885 14714 21941 14716
rect 21965 14714 22021 14716
rect 21725 14662 21771 14714
rect 21771 14662 21781 14714
rect 21805 14662 21835 14714
rect 21835 14662 21847 14714
rect 21847 14662 21861 14714
rect 21885 14662 21899 14714
rect 21899 14662 21911 14714
rect 21911 14662 21941 14714
rect 21965 14662 21975 14714
rect 21975 14662 22021 14714
rect 21725 14660 21781 14662
rect 21805 14660 21861 14662
rect 21885 14660 21941 14662
rect 21965 14660 22021 14662
rect 23478 40568 23534 40624
rect 23478 40160 23534 40216
rect 23662 40568 23718 40624
rect 24122 42744 24178 42800
rect 24030 42220 24086 42256
rect 24030 42200 24032 42220
rect 24032 42200 24084 42220
rect 24084 42200 24086 42220
rect 23846 41248 23902 41304
rect 24692 43546 24748 43548
rect 24772 43546 24828 43548
rect 24852 43546 24908 43548
rect 24932 43546 24988 43548
rect 24692 43494 24738 43546
rect 24738 43494 24748 43546
rect 24772 43494 24802 43546
rect 24802 43494 24814 43546
rect 24814 43494 24828 43546
rect 24852 43494 24866 43546
rect 24866 43494 24878 43546
rect 24878 43494 24908 43546
rect 24932 43494 24942 43546
rect 24942 43494 24988 43546
rect 24692 43492 24748 43494
rect 24772 43492 24828 43494
rect 24852 43492 24908 43494
rect 24932 43492 24988 43494
rect 24692 42458 24748 42460
rect 24772 42458 24828 42460
rect 24852 42458 24908 42460
rect 24932 42458 24988 42460
rect 24692 42406 24738 42458
rect 24738 42406 24748 42458
rect 24772 42406 24802 42458
rect 24802 42406 24814 42458
rect 24814 42406 24828 42458
rect 24852 42406 24866 42458
rect 24866 42406 24878 42458
rect 24878 42406 24908 42458
rect 24932 42406 24942 42458
rect 24942 42406 24988 42458
rect 24692 42404 24748 42406
rect 24772 42404 24828 42406
rect 24852 42404 24908 42406
rect 24932 42404 24988 42406
rect 23478 39480 23534 39536
rect 23754 39888 23810 39944
rect 24214 40024 24270 40080
rect 23846 39208 23902 39264
rect 24398 39480 24454 39536
rect 24122 38936 24178 38992
rect 24398 38528 24454 38584
rect 24122 37848 24178 37904
rect 24398 37304 24454 37360
rect 24122 36760 24178 36816
rect 24122 35808 24178 35864
rect 23662 31864 23718 31920
rect 23018 30368 23074 30424
rect 23202 30232 23258 30288
rect 23294 29144 23350 29200
rect 23110 23432 23166 23488
rect 20718 6724 20774 6760
rect 20718 6704 20720 6724
rect 20720 6704 20772 6724
rect 20772 6704 20774 6724
rect 21178 10920 21234 10976
rect 21086 7284 21088 7304
rect 21088 7284 21140 7304
rect 21140 7284 21142 7304
rect 21086 7248 21142 7284
rect 20718 5480 20774 5536
rect 20718 5364 20774 5400
rect 20718 5344 20720 5364
rect 20720 5344 20772 5364
rect 20772 5344 20774 5364
rect 20442 3848 20498 3904
rect 20718 4392 20774 4448
rect 20718 3596 20774 3632
rect 20718 3576 20720 3596
rect 20720 3576 20772 3596
rect 20772 3576 20774 3596
rect 20534 3032 20590 3088
rect 21725 13626 21781 13628
rect 21805 13626 21861 13628
rect 21885 13626 21941 13628
rect 21965 13626 22021 13628
rect 21725 13574 21771 13626
rect 21771 13574 21781 13626
rect 21805 13574 21835 13626
rect 21835 13574 21847 13626
rect 21847 13574 21861 13626
rect 21885 13574 21899 13626
rect 21899 13574 21911 13626
rect 21911 13574 21941 13626
rect 21965 13574 21975 13626
rect 21975 13574 22021 13626
rect 21725 13572 21781 13574
rect 21805 13572 21861 13574
rect 21885 13572 21941 13574
rect 21965 13572 22021 13574
rect 21725 12538 21781 12540
rect 21805 12538 21861 12540
rect 21885 12538 21941 12540
rect 21965 12538 22021 12540
rect 21725 12486 21771 12538
rect 21771 12486 21781 12538
rect 21805 12486 21835 12538
rect 21835 12486 21847 12538
rect 21847 12486 21861 12538
rect 21885 12486 21899 12538
rect 21899 12486 21911 12538
rect 21911 12486 21941 12538
rect 21965 12486 21975 12538
rect 21975 12486 22021 12538
rect 21725 12484 21781 12486
rect 21805 12484 21861 12486
rect 21885 12484 21941 12486
rect 21965 12484 22021 12486
rect 21914 11772 21916 11792
rect 21916 11772 21968 11792
rect 21968 11772 21970 11792
rect 21914 11736 21970 11772
rect 21725 11450 21781 11452
rect 21805 11450 21861 11452
rect 21885 11450 21941 11452
rect 21965 11450 22021 11452
rect 21725 11398 21771 11450
rect 21771 11398 21781 11450
rect 21805 11398 21835 11450
rect 21835 11398 21847 11450
rect 21847 11398 21861 11450
rect 21885 11398 21899 11450
rect 21899 11398 21911 11450
rect 21911 11398 21941 11450
rect 21965 11398 21975 11450
rect 21975 11398 22021 11450
rect 21725 11396 21781 11398
rect 21805 11396 21861 11398
rect 21885 11396 21941 11398
rect 21965 11396 22021 11398
rect 22374 11736 22430 11792
rect 21725 10362 21781 10364
rect 21805 10362 21861 10364
rect 21885 10362 21941 10364
rect 21965 10362 22021 10364
rect 21725 10310 21771 10362
rect 21771 10310 21781 10362
rect 21805 10310 21835 10362
rect 21835 10310 21847 10362
rect 21847 10310 21861 10362
rect 21885 10310 21899 10362
rect 21899 10310 21911 10362
rect 21911 10310 21941 10362
rect 21965 10310 21975 10362
rect 21975 10310 22021 10362
rect 21725 10308 21781 10310
rect 21805 10308 21861 10310
rect 21885 10308 21941 10310
rect 21965 10308 22021 10310
rect 21638 9424 21694 9480
rect 21725 9274 21781 9276
rect 21805 9274 21861 9276
rect 21885 9274 21941 9276
rect 21965 9274 22021 9276
rect 21725 9222 21771 9274
rect 21771 9222 21781 9274
rect 21805 9222 21835 9274
rect 21835 9222 21847 9274
rect 21847 9222 21861 9274
rect 21885 9222 21899 9274
rect 21899 9222 21911 9274
rect 21911 9222 21941 9274
rect 21965 9222 21975 9274
rect 21975 9222 22021 9274
rect 21725 9220 21781 9222
rect 21805 9220 21861 9222
rect 21885 9220 21941 9222
rect 21965 9220 22021 9222
rect 21725 8186 21781 8188
rect 21805 8186 21861 8188
rect 21885 8186 21941 8188
rect 21965 8186 22021 8188
rect 21725 8134 21771 8186
rect 21771 8134 21781 8186
rect 21805 8134 21835 8186
rect 21835 8134 21847 8186
rect 21847 8134 21861 8186
rect 21885 8134 21899 8186
rect 21899 8134 21911 8186
rect 21911 8134 21941 8186
rect 21965 8134 21975 8186
rect 21975 8134 22021 8186
rect 21725 8132 21781 8134
rect 21805 8132 21861 8134
rect 21885 8132 21941 8134
rect 21965 8132 22021 8134
rect 21725 7098 21781 7100
rect 21805 7098 21861 7100
rect 21885 7098 21941 7100
rect 21965 7098 22021 7100
rect 21725 7046 21771 7098
rect 21771 7046 21781 7098
rect 21805 7046 21835 7098
rect 21835 7046 21847 7098
rect 21847 7046 21861 7098
rect 21885 7046 21899 7098
rect 21899 7046 21911 7098
rect 21911 7046 21941 7098
rect 21965 7046 21975 7098
rect 21975 7046 22021 7098
rect 21725 7044 21781 7046
rect 21805 7044 21861 7046
rect 21885 7044 21941 7046
rect 21965 7044 22021 7046
rect 21270 5752 21326 5808
rect 20810 2352 20866 2408
rect 20994 1300 20996 1320
rect 20996 1300 21048 1320
rect 21048 1300 21050 1320
rect 20994 1264 21050 1300
rect 21725 6010 21781 6012
rect 21805 6010 21861 6012
rect 21885 6010 21941 6012
rect 21965 6010 22021 6012
rect 21725 5958 21771 6010
rect 21771 5958 21781 6010
rect 21805 5958 21835 6010
rect 21835 5958 21847 6010
rect 21847 5958 21861 6010
rect 21885 5958 21899 6010
rect 21899 5958 21911 6010
rect 21911 5958 21941 6010
rect 21965 5958 21975 6010
rect 21975 5958 22021 6010
rect 21725 5956 21781 5958
rect 21805 5956 21861 5958
rect 21885 5956 21941 5958
rect 21965 5956 22021 5958
rect 21638 5652 21640 5672
rect 21640 5652 21692 5672
rect 21692 5652 21694 5672
rect 21638 5616 21694 5652
rect 21914 5208 21970 5264
rect 22098 5208 22154 5264
rect 21362 4392 21418 4448
rect 21178 3884 21180 3904
rect 21180 3884 21232 3904
rect 21232 3884 21234 3904
rect 21178 3848 21234 3884
rect 21178 3712 21234 3768
rect 21454 3884 21456 3904
rect 21456 3884 21508 3904
rect 21508 3884 21510 3904
rect 21454 3848 21510 3884
rect 21178 1944 21234 2000
rect 21725 4922 21781 4924
rect 21805 4922 21861 4924
rect 21885 4922 21941 4924
rect 21965 4922 22021 4924
rect 21725 4870 21771 4922
rect 21771 4870 21781 4922
rect 21805 4870 21835 4922
rect 21835 4870 21847 4922
rect 21847 4870 21861 4922
rect 21885 4870 21899 4922
rect 21899 4870 21911 4922
rect 21911 4870 21941 4922
rect 21965 4870 21975 4922
rect 21975 4870 22021 4922
rect 21725 4868 21781 4870
rect 21805 4868 21861 4870
rect 21885 4868 21941 4870
rect 21965 4868 22021 4870
rect 21914 4256 21970 4312
rect 22282 5480 22338 5536
rect 23018 21548 23074 21584
rect 23018 21528 23020 21548
rect 23020 21528 23072 21548
rect 23072 21528 23074 21548
rect 23570 26968 23626 27024
rect 23386 22616 23442 22672
rect 23662 22616 23718 22672
rect 24214 34584 24270 34640
rect 24122 33496 24178 33552
rect 24122 32408 24178 32464
rect 24214 31592 24270 31648
rect 24214 30232 24270 30288
rect 24214 29144 24270 29200
rect 24122 29008 24178 29064
rect 24122 28056 24178 28112
rect 24214 26424 24270 26480
rect 24122 24792 24178 24848
rect 24030 24112 24086 24168
rect 24122 23704 24178 23760
rect 23938 20576 23994 20632
rect 23754 19896 23810 19952
rect 23110 17584 23166 17640
rect 24122 21528 24178 21584
rect 24398 36216 24454 36272
rect 24398 35128 24454 35184
rect 24398 34484 24400 34504
rect 24400 34484 24452 34504
rect 24452 34484 24454 34504
rect 24398 34448 24454 34484
rect 24692 41370 24748 41372
rect 24772 41370 24828 41372
rect 24852 41370 24908 41372
rect 24932 41370 24988 41372
rect 24692 41318 24738 41370
rect 24738 41318 24748 41370
rect 24772 41318 24802 41370
rect 24802 41318 24814 41370
rect 24814 41318 24828 41370
rect 24852 41318 24866 41370
rect 24866 41318 24878 41370
rect 24878 41318 24908 41370
rect 24932 41318 24942 41370
rect 24942 41318 24988 41370
rect 24692 41316 24748 41318
rect 24772 41316 24828 41318
rect 24852 41316 24908 41318
rect 24932 41316 24988 41318
rect 25042 41112 25098 41168
rect 24692 40282 24748 40284
rect 24772 40282 24828 40284
rect 24852 40282 24908 40284
rect 24932 40282 24988 40284
rect 24692 40230 24738 40282
rect 24738 40230 24748 40282
rect 24772 40230 24802 40282
rect 24802 40230 24814 40282
rect 24814 40230 24828 40282
rect 24852 40230 24866 40282
rect 24866 40230 24878 40282
rect 24878 40230 24908 40282
rect 24932 40230 24942 40282
rect 24942 40230 24988 40282
rect 24692 40228 24748 40230
rect 24772 40228 24828 40230
rect 24852 40228 24908 40230
rect 24932 40228 24988 40230
rect 24582 39344 24638 39400
rect 24398 33088 24454 33144
rect 24398 31864 24454 31920
rect 24398 30776 24454 30832
rect 24398 29688 24454 29744
rect 24398 28872 24454 28928
rect 24398 27512 24454 27568
rect 24398 25336 24454 25392
rect 24398 24248 24454 24304
rect 24398 23468 24400 23488
rect 24400 23468 24452 23488
rect 24452 23468 24454 23488
rect 24398 23432 24454 23468
rect 24398 22072 24454 22128
rect 24306 21120 24362 21176
rect 24214 19352 24270 19408
rect 24122 17856 24178 17912
rect 24030 17176 24086 17232
rect 23938 16496 23994 16552
rect 23754 15544 23810 15600
rect 22650 12280 22706 12336
rect 22834 11756 22890 11792
rect 22834 11736 22836 11756
rect 22836 11736 22888 11756
rect 22888 11736 22890 11756
rect 24122 15136 24178 15192
rect 22558 6704 22614 6760
rect 22650 6180 22706 6216
rect 22650 6160 22652 6180
rect 22652 6160 22704 6180
rect 22704 6160 22706 6180
rect 22558 5752 22614 5808
rect 22558 5480 22614 5536
rect 21725 3834 21781 3836
rect 21805 3834 21861 3836
rect 21885 3834 21941 3836
rect 21965 3834 22021 3836
rect 21725 3782 21771 3834
rect 21771 3782 21781 3834
rect 21805 3782 21835 3834
rect 21835 3782 21847 3834
rect 21847 3782 21861 3834
rect 21885 3782 21899 3834
rect 21899 3782 21911 3834
rect 21911 3782 21941 3834
rect 21965 3782 21975 3834
rect 21975 3782 22021 3834
rect 21725 3780 21781 3782
rect 21805 3780 21861 3782
rect 21885 3780 21941 3782
rect 21965 3780 22021 3782
rect 22098 3476 22100 3496
rect 22100 3476 22152 3496
rect 22152 3476 22154 3496
rect 22098 3440 22154 3476
rect 21086 856 21142 912
rect 21725 2746 21781 2748
rect 21805 2746 21861 2748
rect 21885 2746 21941 2748
rect 21965 2746 22021 2748
rect 21725 2694 21771 2746
rect 21771 2694 21781 2746
rect 21805 2694 21835 2746
rect 21835 2694 21847 2746
rect 21847 2694 21861 2746
rect 21885 2694 21899 2746
rect 21899 2694 21911 2746
rect 21911 2694 21941 2746
rect 21965 2694 21975 2746
rect 21975 2694 22021 2746
rect 21725 2692 21781 2694
rect 21805 2692 21861 2694
rect 21885 2692 21941 2694
rect 21965 2692 22021 2694
rect 21914 2488 21970 2544
rect 21725 1658 21781 1660
rect 21805 1658 21861 1660
rect 21885 1658 21941 1660
rect 21965 1658 22021 1660
rect 21725 1606 21771 1658
rect 21771 1606 21781 1658
rect 21805 1606 21835 1658
rect 21835 1606 21847 1658
rect 21847 1606 21861 1658
rect 21885 1606 21899 1658
rect 21899 1606 21911 1658
rect 21911 1606 21941 1658
rect 21965 1606 21975 1658
rect 21975 1606 22021 1658
rect 21725 1604 21781 1606
rect 21805 1604 21861 1606
rect 21885 1604 21941 1606
rect 21965 1604 22021 1606
rect 22374 3032 22430 3088
rect 22742 4528 22798 4584
rect 22558 1400 22614 1456
rect 24030 12824 24086 12880
rect 23846 12280 23902 12336
rect 23846 10104 23902 10160
rect 23938 9580 23994 9616
rect 23938 9560 23940 9580
rect 23940 9560 23992 9580
rect 23992 9560 23994 9580
rect 23846 9016 23902 9072
rect 23938 8472 23994 8528
rect 24214 7404 24270 7440
rect 24214 7384 24216 7404
rect 24216 7384 24268 7404
rect 24268 7384 24270 7404
rect 24214 7248 24270 7304
rect 23478 6840 23534 6896
rect 23386 6704 23442 6760
rect 23202 6296 23258 6352
rect 23386 5752 23442 5808
rect 23570 5344 23626 5400
rect 23478 5092 23534 5128
rect 23478 5072 23480 5092
rect 23480 5072 23532 5092
rect 23532 5072 23534 5092
rect 23110 3576 23166 3632
rect 23846 5616 23902 5672
rect 23938 4936 23994 4992
rect 24030 2488 24086 2544
rect 24398 20984 24454 21040
rect 24398 18808 24454 18864
rect 24398 18264 24454 18320
rect 24398 16632 24454 16688
rect 24398 14456 24454 14512
rect 24490 13912 24546 13968
rect 24398 11736 24454 11792
rect 24490 10668 24546 10704
rect 24490 10648 24492 10668
rect 24492 10648 24544 10668
rect 24544 10648 24546 10668
rect 24490 8880 24546 8936
rect 24692 39194 24748 39196
rect 24772 39194 24828 39196
rect 24852 39194 24908 39196
rect 24932 39194 24988 39196
rect 24692 39142 24738 39194
rect 24738 39142 24748 39194
rect 24772 39142 24802 39194
rect 24802 39142 24814 39194
rect 24814 39142 24828 39194
rect 24852 39142 24866 39194
rect 24866 39142 24878 39194
rect 24878 39142 24908 39194
rect 24932 39142 24942 39194
rect 24942 39142 24988 39194
rect 24692 39140 24748 39142
rect 24772 39140 24828 39142
rect 24852 39140 24908 39142
rect 24932 39140 24988 39142
rect 24692 38106 24748 38108
rect 24772 38106 24828 38108
rect 24852 38106 24908 38108
rect 24932 38106 24988 38108
rect 24692 38054 24738 38106
rect 24738 38054 24748 38106
rect 24772 38054 24802 38106
rect 24802 38054 24814 38106
rect 24814 38054 24828 38106
rect 24852 38054 24866 38106
rect 24866 38054 24878 38106
rect 24878 38054 24908 38106
rect 24932 38054 24942 38106
rect 24942 38054 24988 38106
rect 24692 38052 24748 38054
rect 24772 38052 24828 38054
rect 24852 38052 24908 38054
rect 24932 38052 24988 38054
rect 24692 37018 24748 37020
rect 24772 37018 24828 37020
rect 24852 37018 24908 37020
rect 24932 37018 24988 37020
rect 24692 36966 24738 37018
rect 24738 36966 24748 37018
rect 24772 36966 24802 37018
rect 24802 36966 24814 37018
rect 24814 36966 24828 37018
rect 24852 36966 24866 37018
rect 24866 36966 24878 37018
rect 24878 36966 24908 37018
rect 24932 36966 24942 37018
rect 24942 36966 24988 37018
rect 24692 36964 24748 36966
rect 24772 36964 24828 36966
rect 24852 36964 24908 36966
rect 24932 36964 24988 36966
rect 24692 35930 24748 35932
rect 24772 35930 24828 35932
rect 24852 35930 24908 35932
rect 24932 35930 24988 35932
rect 24692 35878 24738 35930
rect 24738 35878 24748 35930
rect 24772 35878 24802 35930
rect 24802 35878 24814 35930
rect 24814 35878 24828 35930
rect 24852 35878 24866 35930
rect 24866 35878 24878 35930
rect 24878 35878 24908 35930
rect 24932 35878 24942 35930
rect 24942 35878 24988 35930
rect 24692 35876 24748 35878
rect 24772 35876 24828 35878
rect 24852 35876 24908 35878
rect 24932 35876 24988 35878
rect 24692 34842 24748 34844
rect 24772 34842 24828 34844
rect 24852 34842 24908 34844
rect 24932 34842 24988 34844
rect 24692 34790 24738 34842
rect 24738 34790 24748 34842
rect 24772 34790 24802 34842
rect 24802 34790 24814 34842
rect 24814 34790 24828 34842
rect 24852 34790 24866 34842
rect 24866 34790 24878 34842
rect 24878 34790 24908 34842
rect 24932 34790 24942 34842
rect 24942 34790 24988 34842
rect 24692 34788 24748 34790
rect 24772 34788 24828 34790
rect 24852 34788 24908 34790
rect 24932 34788 24988 34790
rect 24692 33754 24748 33756
rect 24772 33754 24828 33756
rect 24852 33754 24908 33756
rect 24932 33754 24988 33756
rect 24692 33702 24738 33754
rect 24738 33702 24748 33754
rect 24772 33702 24802 33754
rect 24802 33702 24814 33754
rect 24814 33702 24828 33754
rect 24852 33702 24866 33754
rect 24866 33702 24878 33754
rect 24878 33702 24908 33754
rect 24932 33702 24942 33754
rect 24942 33702 24988 33754
rect 24692 33700 24748 33702
rect 24772 33700 24828 33702
rect 24852 33700 24908 33702
rect 24932 33700 24988 33702
rect 24692 32666 24748 32668
rect 24772 32666 24828 32668
rect 24852 32666 24908 32668
rect 24932 32666 24988 32668
rect 24692 32614 24738 32666
rect 24738 32614 24748 32666
rect 24772 32614 24802 32666
rect 24802 32614 24814 32666
rect 24814 32614 24828 32666
rect 24852 32614 24866 32666
rect 24866 32614 24878 32666
rect 24878 32614 24908 32666
rect 24932 32614 24942 32666
rect 24942 32614 24988 32666
rect 24692 32612 24748 32614
rect 24772 32612 24828 32614
rect 24852 32612 24908 32614
rect 24932 32612 24988 32614
rect 24692 31578 24748 31580
rect 24772 31578 24828 31580
rect 24852 31578 24908 31580
rect 24932 31578 24988 31580
rect 24692 31526 24738 31578
rect 24738 31526 24748 31578
rect 24772 31526 24802 31578
rect 24802 31526 24814 31578
rect 24814 31526 24828 31578
rect 24852 31526 24866 31578
rect 24866 31526 24878 31578
rect 24878 31526 24908 31578
rect 24932 31526 24942 31578
rect 24942 31526 24988 31578
rect 24692 31524 24748 31526
rect 24772 31524 24828 31526
rect 24852 31524 24908 31526
rect 24932 31524 24988 31526
rect 24692 30490 24748 30492
rect 24772 30490 24828 30492
rect 24852 30490 24908 30492
rect 24932 30490 24988 30492
rect 24692 30438 24738 30490
rect 24738 30438 24748 30490
rect 24772 30438 24802 30490
rect 24802 30438 24814 30490
rect 24814 30438 24828 30490
rect 24852 30438 24866 30490
rect 24866 30438 24878 30490
rect 24878 30438 24908 30490
rect 24932 30438 24942 30490
rect 24942 30438 24988 30490
rect 24692 30436 24748 30438
rect 24772 30436 24828 30438
rect 24852 30436 24908 30438
rect 24932 30436 24988 30438
rect 24692 29402 24748 29404
rect 24772 29402 24828 29404
rect 24852 29402 24908 29404
rect 24932 29402 24988 29404
rect 24692 29350 24738 29402
rect 24738 29350 24748 29402
rect 24772 29350 24802 29402
rect 24802 29350 24814 29402
rect 24814 29350 24828 29402
rect 24852 29350 24866 29402
rect 24866 29350 24878 29402
rect 24878 29350 24908 29402
rect 24932 29350 24942 29402
rect 24942 29350 24988 29402
rect 24692 29348 24748 29350
rect 24772 29348 24828 29350
rect 24852 29348 24908 29350
rect 24932 29348 24988 29350
rect 24692 28314 24748 28316
rect 24772 28314 24828 28316
rect 24852 28314 24908 28316
rect 24932 28314 24988 28316
rect 24692 28262 24738 28314
rect 24738 28262 24748 28314
rect 24772 28262 24802 28314
rect 24802 28262 24814 28314
rect 24814 28262 24828 28314
rect 24852 28262 24866 28314
rect 24866 28262 24878 28314
rect 24878 28262 24908 28314
rect 24932 28262 24942 28314
rect 24942 28262 24988 28314
rect 24692 28260 24748 28262
rect 24772 28260 24828 28262
rect 24852 28260 24908 28262
rect 24932 28260 24988 28262
rect 24692 27226 24748 27228
rect 24772 27226 24828 27228
rect 24852 27226 24908 27228
rect 24932 27226 24988 27228
rect 24692 27174 24738 27226
rect 24738 27174 24748 27226
rect 24772 27174 24802 27226
rect 24802 27174 24814 27226
rect 24814 27174 24828 27226
rect 24852 27174 24866 27226
rect 24866 27174 24878 27226
rect 24878 27174 24908 27226
rect 24932 27174 24942 27226
rect 24942 27174 24988 27226
rect 24692 27172 24748 27174
rect 24772 27172 24828 27174
rect 24852 27172 24908 27174
rect 24932 27172 24988 27174
rect 24692 26138 24748 26140
rect 24772 26138 24828 26140
rect 24852 26138 24908 26140
rect 24932 26138 24988 26140
rect 24692 26086 24738 26138
rect 24738 26086 24748 26138
rect 24772 26086 24802 26138
rect 24802 26086 24814 26138
rect 24814 26086 24828 26138
rect 24852 26086 24866 26138
rect 24866 26086 24878 26138
rect 24878 26086 24908 26138
rect 24932 26086 24942 26138
rect 24942 26086 24988 26138
rect 24692 26084 24748 26086
rect 24772 26084 24828 26086
rect 24852 26084 24908 26086
rect 24932 26084 24988 26086
rect 24692 25050 24748 25052
rect 24772 25050 24828 25052
rect 24852 25050 24908 25052
rect 24932 25050 24988 25052
rect 24692 24998 24738 25050
rect 24738 24998 24748 25050
rect 24772 24998 24802 25050
rect 24802 24998 24814 25050
rect 24814 24998 24828 25050
rect 24852 24998 24866 25050
rect 24866 24998 24878 25050
rect 24878 24998 24908 25050
rect 24932 24998 24942 25050
rect 24942 24998 24988 25050
rect 24692 24996 24748 24998
rect 24772 24996 24828 24998
rect 24852 24996 24908 24998
rect 24932 24996 24988 24998
rect 24692 23962 24748 23964
rect 24772 23962 24828 23964
rect 24852 23962 24908 23964
rect 24932 23962 24988 23964
rect 24692 23910 24738 23962
rect 24738 23910 24748 23962
rect 24772 23910 24802 23962
rect 24802 23910 24814 23962
rect 24814 23910 24828 23962
rect 24852 23910 24866 23962
rect 24866 23910 24878 23962
rect 24878 23910 24908 23962
rect 24932 23910 24942 23962
rect 24942 23910 24988 23962
rect 24692 23908 24748 23910
rect 24772 23908 24828 23910
rect 24852 23908 24908 23910
rect 24932 23908 24988 23910
rect 24692 22874 24748 22876
rect 24772 22874 24828 22876
rect 24852 22874 24908 22876
rect 24932 22874 24988 22876
rect 24692 22822 24738 22874
rect 24738 22822 24748 22874
rect 24772 22822 24802 22874
rect 24802 22822 24814 22874
rect 24814 22822 24828 22874
rect 24852 22822 24866 22874
rect 24866 22822 24878 22874
rect 24878 22822 24908 22874
rect 24932 22822 24942 22874
rect 24942 22822 24988 22874
rect 24692 22820 24748 22822
rect 24772 22820 24828 22822
rect 24852 22820 24908 22822
rect 24932 22820 24988 22822
rect 24692 21786 24748 21788
rect 24772 21786 24828 21788
rect 24852 21786 24908 21788
rect 24932 21786 24988 21788
rect 24692 21734 24738 21786
rect 24738 21734 24748 21786
rect 24772 21734 24802 21786
rect 24802 21734 24814 21786
rect 24814 21734 24828 21786
rect 24852 21734 24866 21786
rect 24866 21734 24878 21786
rect 24878 21734 24908 21786
rect 24932 21734 24942 21786
rect 24942 21734 24988 21786
rect 24692 21732 24748 21734
rect 24772 21732 24828 21734
rect 24852 21732 24908 21734
rect 24932 21732 24988 21734
rect 24692 20698 24748 20700
rect 24772 20698 24828 20700
rect 24852 20698 24908 20700
rect 24932 20698 24988 20700
rect 24692 20646 24738 20698
rect 24738 20646 24748 20698
rect 24772 20646 24802 20698
rect 24802 20646 24814 20698
rect 24814 20646 24828 20698
rect 24852 20646 24866 20698
rect 24866 20646 24878 20698
rect 24878 20646 24908 20698
rect 24932 20646 24942 20698
rect 24942 20646 24988 20698
rect 24692 20644 24748 20646
rect 24772 20644 24828 20646
rect 24852 20644 24908 20646
rect 24932 20644 24988 20646
rect 24692 19610 24748 19612
rect 24772 19610 24828 19612
rect 24852 19610 24908 19612
rect 24932 19610 24988 19612
rect 24692 19558 24738 19610
rect 24738 19558 24748 19610
rect 24772 19558 24802 19610
rect 24802 19558 24814 19610
rect 24814 19558 24828 19610
rect 24852 19558 24866 19610
rect 24866 19558 24878 19610
rect 24878 19558 24908 19610
rect 24932 19558 24942 19610
rect 24942 19558 24988 19610
rect 24692 19556 24748 19558
rect 24772 19556 24828 19558
rect 24852 19556 24908 19558
rect 24932 19556 24988 19558
rect 24692 18522 24748 18524
rect 24772 18522 24828 18524
rect 24852 18522 24908 18524
rect 24932 18522 24988 18524
rect 24692 18470 24738 18522
rect 24738 18470 24748 18522
rect 24772 18470 24802 18522
rect 24802 18470 24814 18522
rect 24814 18470 24828 18522
rect 24852 18470 24866 18522
rect 24866 18470 24878 18522
rect 24878 18470 24908 18522
rect 24932 18470 24942 18522
rect 24942 18470 24988 18522
rect 24692 18468 24748 18470
rect 24772 18468 24828 18470
rect 24852 18468 24908 18470
rect 24932 18468 24988 18470
rect 24692 17434 24748 17436
rect 24772 17434 24828 17436
rect 24852 17434 24908 17436
rect 24932 17434 24988 17436
rect 24692 17382 24738 17434
rect 24738 17382 24748 17434
rect 24772 17382 24802 17434
rect 24802 17382 24814 17434
rect 24814 17382 24828 17434
rect 24852 17382 24866 17434
rect 24866 17382 24878 17434
rect 24878 17382 24908 17434
rect 24932 17382 24942 17434
rect 24942 17382 24988 17434
rect 24692 17380 24748 17382
rect 24772 17380 24828 17382
rect 24852 17380 24908 17382
rect 24932 17380 24988 17382
rect 25134 25880 25190 25936
rect 24692 16346 24748 16348
rect 24772 16346 24828 16348
rect 24852 16346 24908 16348
rect 24932 16346 24988 16348
rect 24692 16294 24738 16346
rect 24738 16294 24748 16346
rect 24772 16294 24802 16346
rect 24802 16294 24814 16346
rect 24814 16294 24828 16346
rect 24852 16294 24866 16346
rect 24866 16294 24878 16346
rect 24878 16294 24908 16346
rect 24932 16294 24942 16346
rect 24942 16294 24988 16346
rect 24692 16292 24748 16294
rect 24772 16292 24828 16294
rect 24852 16292 24908 16294
rect 24932 16292 24988 16294
rect 24692 15258 24748 15260
rect 24772 15258 24828 15260
rect 24852 15258 24908 15260
rect 24932 15258 24988 15260
rect 24692 15206 24738 15258
rect 24738 15206 24748 15258
rect 24772 15206 24802 15258
rect 24802 15206 24814 15258
rect 24814 15206 24828 15258
rect 24852 15206 24866 15258
rect 24866 15206 24878 15258
rect 24878 15206 24908 15258
rect 24932 15206 24942 15258
rect 24942 15206 24988 15258
rect 24692 15204 24748 15206
rect 24772 15204 24828 15206
rect 24852 15204 24908 15206
rect 24932 15204 24988 15206
rect 24692 14170 24748 14172
rect 24772 14170 24828 14172
rect 24852 14170 24908 14172
rect 24932 14170 24988 14172
rect 24692 14118 24738 14170
rect 24738 14118 24748 14170
rect 24772 14118 24802 14170
rect 24802 14118 24814 14170
rect 24814 14118 24828 14170
rect 24852 14118 24866 14170
rect 24866 14118 24878 14170
rect 24878 14118 24908 14170
rect 24932 14118 24942 14170
rect 24942 14118 24988 14170
rect 24692 14116 24748 14118
rect 24772 14116 24828 14118
rect 24852 14116 24908 14118
rect 24932 14116 24988 14118
rect 24674 13404 24676 13424
rect 24676 13404 24728 13424
rect 24728 13404 24730 13424
rect 24674 13368 24730 13404
rect 24692 13082 24748 13084
rect 24772 13082 24828 13084
rect 24852 13082 24908 13084
rect 24932 13082 24988 13084
rect 24692 13030 24738 13082
rect 24738 13030 24748 13082
rect 24772 13030 24802 13082
rect 24802 13030 24814 13082
rect 24814 13030 24828 13082
rect 24852 13030 24866 13082
rect 24866 13030 24878 13082
rect 24878 13030 24908 13082
rect 24932 13030 24942 13082
rect 24942 13030 24988 13082
rect 24692 13028 24748 13030
rect 24772 13028 24828 13030
rect 24852 13028 24908 13030
rect 24932 13028 24988 13030
rect 24692 11994 24748 11996
rect 24772 11994 24828 11996
rect 24852 11994 24908 11996
rect 24932 11994 24988 11996
rect 24692 11942 24738 11994
rect 24738 11942 24748 11994
rect 24772 11942 24802 11994
rect 24802 11942 24814 11994
rect 24814 11942 24828 11994
rect 24852 11942 24866 11994
rect 24866 11942 24878 11994
rect 24878 11942 24908 11994
rect 24932 11942 24942 11994
rect 24942 11942 24988 11994
rect 24692 11940 24748 11942
rect 24772 11940 24828 11942
rect 24852 11940 24908 11942
rect 24932 11940 24988 11942
rect 25042 11192 25098 11248
rect 24692 10906 24748 10908
rect 24772 10906 24828 10908
rect 24852 10906 24908 10908
rect 24932 10906 24988 10908
rect 24692 10854 24738 10906
rect 24738 10854 24748 10906
rect 24772 10854 24802 10906
rect 24802 10854 24814 10906
rect 24814 10854 24828 10906
rect 24852 10854 24866 10906
rect 24866 10854 24878 10906
rect 24878 10854 24908 10906
rect 24932 10854 24942 10906
rect 24942 10854 24988 10906
rect 24692 10852 24748 10854
rect 24772 10852 24828 10854
rect 24852 10852 24908 10854
rect 24932 10852 24988 10854
rect 24692 9818 24748 9820
rect 24772 9818 24828 9820
rect 24852 9818 24908 9820
rect 24932 9818 24988 9820
rect 24692 9766 24738 9818
rect 24738 9766 24748 9818
rect 24772 9766 24802 9818
rect 24802 9766 24814 9818
rect 24814 9766 24828 9818
rect 24852 9766 24866 9818
rect 24866 9766 24878 9818
rect 24878 9766 24908 9818
rect 24932 9766 24942 9818
rect 24942 9766 24988 9818
rect 24692 9764 24748 9766
rect 24772 9764 24828 9766
rect 24852 9764 24908 9766
rect 24932 9764 24988 9766
rect 24692 8730 24748 8732
rect 24772 8730 24828 8732
rect 24852 8730 24908 8732
rect 24932 8730 24988 8732
rect 24692 8678 24738 8730
rect 24738 8678 24748 8730
rect 24772 8678 24802 8730
rect 24802 8678 24814 8730
rect 24814 8678 24828 8730
rect 24852 8678 24866 8730
rect 24866 8678 24878 8730
rect 24878 8678 24908 8730
rect 24932 8678 24942 8730
rect 24942 8678 24988 8730
rect 24692 8676 24748 8678
rect 24772 8676 24828 8678
rect 24852 8676 24908 8678
rect 24932 8676 24988 8678
rect 24692 7642 24748 7644
rect 24772 7642 24828 7644
rect 24852 7642 24908 7644
rect 24932 7642 24988 7644
rect 24692 7590 24738 7642
rect 24738 7590 24748 7642
rect 24772 7590 24802 7642
rect 24802 7590 24814 7642
rect 24814 7590 24828 7642
rect 24852 7590 24866 7642
rect 24866 7590 24878 7642
rect 24878 7590 24908 7642
rect 24932 7590 24942 7642
rect 24942 7590 24988 7642
rect 24692 7588 24748 7590
rect 24772 7588 24828 7590
rect 24852 7588 24908 7590
rect 24932 7588 24988 7590
rect 25778 20168 25834 20224
rect 25318 7928 25374 7984
rect 24692 6554 24748 6556
rect 24772 6554 24828 6556
rect 24852 6554 24908 6556
rect 24932 6554 24988 6556
rect 24692 6502 24738 6554
rect 24738 6502 24748 6554
rect 24772 6502 24802 6554
rect 24802 6502 24814 6554
rect 24814 6502 24828 6554
rect 24852 6502 24866 6554
rect 24866 6502 24878 6554
rect 24878 6502 24908 6554
rect 24932 6502 24942 6554
rect 24942 6502 24988 6554
rect 24692 6500 24748 6502
rect 24772 6500 24828 6502
rect 24852 6500 24908 6502
rect 24932 6500 24988 6502
rect 24692 5466 24748 5468
rect 24772 5466 24828 5468
rect 24852 5466 24908 5468
rect 24932 5466 24988 5468
rect 24692 5414 24738 5466
rect 24738 5414 24748 5466
rect 24772 5414 24802 5466
rect 24802 5414 24814 5466
rect 24814 5414 24828 5466
rect 24852 5414 24866 5466
rect 24866 5414 24878 5466
rect 24878 5414 24908 5466
rect 24932 5414 24942 5466
rect 24942 5414 24988 5466
rect 24692 5412 24748 5414
rect 24772 5412 24828 5414
rect 24852 5412 24908 5414
rect 24932 5412 24988 5414
rect 24692 4378 24748 4380
rect 24772 4378 24828 4380
rect 24852 4378 24908 4380
rect 24932 4378 24988 4380
rect 24692 4326 24738 4378
rect 24738 4326 24748 4378
rect 24772 4326 24802 4378
rect 24802 4326 24814 4378
rect 24814 4326 24828 4378
rect 24852 4326 24866 4378
rect 24866 4326 24878 4378
rect 24878 4326 24908 4378
rect 24932 4326 24942 4378
rect 24942 4326 24988 4378
rect 24692 4324 24748 4326
rect 24772 4324 24828 4326
rect 24852 4324 24908 4326
rect 24932 4324 24988 4326
rect 24692 3290 24748 3292
rect 24772 3290 24828 3292
rect 24852 3290 24908 3292
rect 24932 3290 24988 3292
rect 24692 3238 24738 3290
rect 24738 3238 24748 3290
rect 24772 3238 24802 3290
rect 24802 3238 24814 3290
rect 24814 3238 24828 3290
rect 24852 3238 24866 3290
rect 24866 3238 24878 3290
rect 24878 3238 24908 3290
rect 24932 3238 24942 3290
rect 24942 3238 24988 3290
rect 24692 3236 24748 3238
rect 24772 3236 24828 3238
rect 24852 3236 24908 3238
rect 24932 3236 24988 3238
rect 24692 2202 24748 2204
rect 24772 2202 24828 2204
rect 24852 2202 24908 2204
rect 24932 2202 24988 2204
rect 24692 2150 24738 2202
rect 24738 2150 24748 2202
rect 24772 2150 24802 2202
rect 24802 2150 24814 2202
rect 24814 2150 24828 2202
rect 24852 2150 24866 2202
rect 24866 2150 24878 2202
rect 24878 2150 24908 2202
rect 24932 2150 24942 2202
rect 24942 2150 24988 2202
rect 24692 2148 24748 2150
rect 24772 2148 24828 2150
rect 24852 2148 24908 2150
rect 24932 2148 24988 2150
rect 24692 1114 24748 1116
rect 24772 1114 24828 1116
rect 24852 1114 24908 1116
rect 24932 1114 24988 1116
rect 24692 1062 24738 1114
rect 24738 1062 24748 1114
rect 24772 1062 24802 1114
rect 24802 1062 24814 1114
rect 24814 1062 24828 1114
rect 24852 1062 24866 1114
rect 24866 1062 24878 1114
rect 24878 1062 24908 1114
rect 24932 1062 24942 1114
rect 24942 1062 24988 1114
rect 24692 1060 24748 1062
rect 24772 1060 24828 1062
rect 24852 1060 24908 1062
rect 24932 1060 24988 1062
rect 25318 3984 25374 4040
rect 25410 1808 25466 1864
<< metal3 >>
rect 23013 43890 23079 43893
rect 25840 43890 26000 43920
rect 23013 43888 26000 43890
rect 23013 43832 23018 43888
rect 23074 43832 26000 43888
rect 23013 43830 26000 43832
rect 23013 43827 23079 43830
rect 25840 43800 26000 43830
rect 6880 43552 7196 43553
rect 6880 43488 6886 43552
rect 6950 43488 6966 43552
rect 7030 43488 7046 43552
rect 7110 43488 7126 43552
rect 7190 43488 7196 43552
rect 6880 43487 7196 43488
rect 12814 43552 13130 43553
rect 12814 43488 12820 43552
rect 12884 43488 12900 43552
rect 12964 43488 12980 43552
rect 13044 43488 13060 43552
rect 13124 43488 13130 43552
rect 12814 43487 13130 43488
rect 18748 43552 19064 43553
rect 18748 43488 18754 43552
rect 18818 43488 18834 43552
rect 18898 43488 18914 43552
rect 18978 43488 18994 43552
rect 19058 43488 19064 43552
rect 18748 43487 19064 43488
rect 24682 43552 24998 43553
rect 24682 43488 24688 43552
rect 24752 43488 24768 43552
rect 24832 43488 24848 43552
rect 24912 43488 24928 43552
rect 24992 43488 24998 43552
rect 24682 43487 24998 43488
rect 23657 43346 23723 43349
rect 25840 43346 26000 43376
rect 23657 43344 26000 43346
rect 23657 43288 23662 43344
rect 23718 43288 26000 43344
rect 23657 43286 26000 43288
rect 23657 43283 23723 43286
rect 25840 43256 26000 43286
rect 20662 43148 20668 43212
rect 20732 43210 20738 43212
rect 22093 43210 22159 43213
rect 20732 43208 22159 43210
rect 20732 43152 22098 43208
rect 22154 43152 22159 43208
rect 20732 43150 22159 43152
rect 20732 43148 20738 43150
rect 22093 43147 22159 43150
rect 11462 43012 11468 43076
rect 11532 43074 11538 43076
rect 12893 43074 12959 43077
rect 11532 43072 12959 43074
rect 11532 43016 12898 43072
rect 12954 43016 12959 43072
rect 11532 43014 12959 43016
rect 11532 43012 11538 43014
rect 12893 43011 12959 43014
rect 13077 43074 13143 43077
rect 13670 43074 13676 43076
rect 13077 43072 13676 43074
rect 13077 43016 13082 43072
rect 13138 43016 13676 43072
rect 13077 43014 13676 43016
rect 13077 43011 13143 43014
rect 13670 43012 13676 43014
rect 13740 43012 13746 43076
rect 3913 43008 4229 43009
rect 3913 42944 3919 43008
rect 3983 42944 3999 43008
rect 4063 42944 4079 43008
rect 4143 42944 4159 43008
rect 4223 42944 4229 43008
rect 3913 42943 4229 42944
rect 9847 43008 10163 43009
rect 9847 42944 9853 43008
rect 9917 42944 9933 43008
rect 9997 42944 10013 43008
rect 10077 42944 10093 43008
rect 10157 42944 10163 43008
rect 9847 42943 10163 42944
rect 15781 43008 16097 43009
rect 15781 42944 15787 43008
rect 15851 42944 15867 43008
rect 15931 42944 15947 43008
rect 16011 42944 16027 43008
rect 16091 42944 16097 43008
rect 15781 42943 16097 42944
rect 21715 43008 22031 43009
rect 21715 42944 21721 43008
rect 21785 42944 21801 43008
rect 21865 42944 21881 43008
rect 21945 42944 21961 43008
rect 22025 42944 22031 43008
rect 21715 42943 22031 42944
rect 10409 42938 10475 42941
rect 12249 42940 12315 42941
rect 11646 42938 11652 42940
rect 10409 42936 11652 42938
rect 10409 42880 10414 42936
rect 10470 42880 11652 42936
rect 10409 42878 11652 42880
rect 10409 42875 10475 42878
rect 11646 42876 11652 42878
rect 11716 42876 11722 42940
rect 12198 42938 12204 42940
rect 12158 42878 12204 42938
rect 12268 42936 12315 42940
rect 12310 42880 12315 42936
rect 12198 42876 12204 42878
rect 12268 42876 12315 42880
rect 13302 42876 13308 42940
rect 13372 42938 13378 42940
rect 13813 42938 13879 42941
rect 13372 42936 13879 42938
rect 13372 42880 13818 42936
rect 13874 42880 13879 42936
rect 13372 42878 13879 42880
rect 13372 42876 13378 42878
rect 12249 42875 12315 42876
rect 13813 42875 13879 42878
rect 14273 42938 14339 42941
rect 14917 42940 14983 42941
rect 15285 42940 15351 42941
rect 14406 42938 14412 42940
rect 14273 42936 14412 42938
rect 14273 42880 14278 42936
rect 14334 42880 14412 42936
rect 14273 42878 14412 42880
rect 14273 42875 14339 42878
rect 14406 42876 14412 42878
rect 14476 42876 14482 42940
rect 14917 42936 14964 42940
rect 15028 42938 15034 42940
rect 14917 42880 14922 42936
rect 14917 42876 14964 42880
rect 15028 42878 15074 42938
rect 15285 42936 15332 42940
rect 15396 42938 15402 42940
rect 15285 42880 15290 42936
rect 15028 42876 15034 42878
rect 15285 42876 15332 42880
rect 15396 42878 15442 42938
rect 15396 42876 15402 42878
rect 14917 42875 14983 42876
rect 15285 42875 15351 42876
rect 18413 42802 18479 42805
rect 23105 42802 23171 42805
rect 18413 42800 23171 42802
rect 18413 42744 18418 42800
rect 18474 42744 23110 42800
rect 23166 42744 23171 42800
rect 18413 42742 23171 42744
rect 18413 42739 18479 42742
rect 23105 42739 23171 42742
rect 24117 42802 24183 42805
rect 25840 42802 26000 42832
rect 24117 42800 26000 42802
rect 24117 42744 24122 42800
rect 24178 42744 26000 42800
rect 24117 42742 26000 42744
rect 24117 42739 24183 42742
rect 25840 42712 26000 42742
rect 6880 42464 7196 42465
rect 6880 42400 6886 42464
rect 6950 42400 6966 42464
rect 7030 42400 7046 42464
rect 7110 42400 7126 42464
rect 7190 42400 7196 42464
rect 6880 42399 7196 42400
rect 12814 42464 13130 42465
rect 12814 42400 12820 42464
rect 12884 42400 12900 42464
rect 12964 42400 12980 42464
rect 13044 42400 13060 42464
rect 13124 42400 13130 42464
rect 12814 42399 13130 42400
rect 18748 42464 19064 42465
rect 18748 42400 18754 42464
rect 18818 42400 18834 42464
rect 18898 42400 18914 42464
rect 18978 42400 18994 42464
rect 19058 42400 19064 42464
rect 18748 42399 19064 42400
rect 24682 42464 24998 42465
rect 24682 42400 24688 42464
rect 24752 42400 24768 42464
rect 24832 42400 24848 42464
rect 24912 42400 24928 42464
rect 24992 42400 24998 42464
rect 24682 42399 24998 42400
rect 2497 42258 2563 42261
rect 15285 42258 15351 42261
rect 2497 42256 15351 42258
rect 2497 42200 2502 42256
rect 2558 42200 15290 42256
rect 15346 42200 15351 42256
rect 2497 42198 15351 42200
rect 2497 42195 2563 42198
rect 15285 42195 15351 42198
rect 16297 42258 16363 42261
rect 17585 42258 17651 42261
rect 16297 42256 17651 42258
rect 16297 42200 16302 42256
rect 16358 42200 17590 42256
rect 17646 42200 17651 42256
rect 16297 42198 17651 42200
rect 16297 42195 16363 42198
rect 17585 42195 17651 42198
rect 24025 42258 24091 42261
rect 25840 42258 26000 42288
rect 24025 42256 26000 42258
rect 24025 42200 24030 42256
rect 24086 42200 26000 42256
rect 24025 42198 26000 42200
rect 24025 42195 24091 42198
rect 25840 42168 26000 42198
rect 2221 42122 2287 42125
rect 8109 42124 8175 42125
rect 2221 42120 7298 42122
rect 2221 42064 2226 42120
rect 2282 42064 7298 42120
rect 2221 42062 7298 42064
rect 2221 42059 2287 42062
rect 3913 41920 4229 41921
rect 3913 41856 3919 41920
rect 3983 41856 3999 41920
rect 4063 41856 4079 41920
rect 4143 41856 4159 41920
rect 4223 41856 4229 41920
rect 3913 41855 4229 41856
rect 6177 41850 6243 41853
rect 6310 41850 6316 41852
rect 6177 41848 6316 41850
rect 6177 41792 6182 41848
rect 6238 41792 6316 41848
rect 6177 41790 6316 41792
rect 6177 41787 6243 41790
rect 6310 41788 6316 41790
rect 6380 41788 6386 41852
rect 6494 41788 6500 41852
rect 6564 41850 6570 41852
rect 6637 41850 6703 41853
rect 6564 41848 6703 41850
rect 6564 41792 6642 41848
rect 6698 41792 6703 41848
rect 6564 41790 6703 41792
rect 6564 41788 6570 41790
rect 6637 41787 6703 41790
rect 1025 41714 1091 41717
rect 4705 41714 4771 41717
rect 1025 41712 4771 41714
rect 1025 41656 1030 41712
rect 1086 41656 4710 41712
rect 4766 41656 4771 41712
rect 1025 41654 4771 41656
rect 7238 41714 7298 42062
rect 8109 42120 8156 42124
rect 8220 42122 8226 42124
rect 8109 42064 8114 42120
rect 8109 42060 8156 42064
rect 8220 42062 8266 42122
rect 8220 42060 8226 42062
rect 21030 42060 21036 42124
rect 21100 42122 21106 42124
rect 21357 42122 21423 42125
rect 21100 42120 21423 42122
rect 21100 42064 21362 42120
rect 21418 42064 21423 42120
rect 21100 42062 21423 42064
rect 21100 42060 21106 42062
rect 8109 42059 8175 42060
rect 21357 42059 21423 42062
rect 19333 41986 19399 41989
rect 16622 41984 19399 41986
rect 16622 41928 19338 41984
rect 19394 41928 19399 41984
rect 16622 41926 19399 41928
rect 9847 41920 10163 41921
rect 9847 41856 9853 41920
rect 9917 41856 9933 41920
rect 9997 41856 10013 41920
rect 10077 41856 10093 41920
rect 10157 41856 10163 41920
rect 9847 41855 10163 41856
rect 15781 41920 16097 41921
rect 15781 41856 15787 41920
rect 15851 41856 15867 41920
rect 15931 41856 15947 41920
rect 16011 41856 16027 41920
rect 16091 41856 16097 41920
rect 15781 41855 16097 41856
rect 7373 41850 7439 41853
rect 7966 41850 7972 41852
rect 7373 41848 7972 41850
rect 7373 41792 7378 41848
rect 7434 41792 7972 41848
rect 7373 41790 7972 41792
rect 7373 41787 7439 41790
rect 7966 41788 7972 41790
rect 8036 41788 8042 41852
rect 12525 41714 12591 41717
rect 7238 41712 12591 41714
rect 7238 41656 12530 41712
rect 12586 41656 12591 41712
rect 7238 41654 12591 41656
rect 1025 41651 1091 41654
rect 4705 41651 4771 41654
rect 12525 41651 12591 41654
rect 14590 41652 14596 41716
rect 14660 41714 14666 41716
rect 16622 41714 16682 41926
rect 19333 41923 19399 41926
rect 21715 41920 22031 41921
rect 21715 41856 21721 41920
rect 21785 41856 21801 41920
rect 21865 41856 21881 41920
rect 21945 41856 21961 41920
rect 22025 41856 22031 41920
rect 21715 41855 22031 41856
rect 17309 41850 17375 41853
rect 17718 41850 17724 41852
rect 17309 41848 17724 41850
rect 17309 41792 17314 41848
rect 17370 41792 17724 41848
rect 17309 41790 17724 41792
rect 17309 41787 17375 41790
rect 17718 41788 17724 41790
rect 17788 41788 17794 41852
rect 18270 41788 18276 41852
rect 18340 41850 18346 41852
rect 19057 41850 19123 41853
rect 18340 41848 19123 41850
rect 18340 41792 19062 41848
rect 19118 41792 19123 41848
rect 18340 41790 19123 41792
rect 18340 41788 18346 41790
rect 19057 41787 19123 41790
rect 17585 41716 17651 41717
rect 17534 41714 17540 41716
rect 14660 41654 16682 41714
rect 17494 41654 17540 41714
rect 17604 41712 17651 41716
rect 17953 41714 18019 41717
rect 22185 41714 22251 41717
rect 17646 41656 17651 41712
rect 14660 41652 14666 41654
rect 17534 41652 17540 41654
rect 17604 41652 17651 41656
rect 17585 41651 17651 41652
rect 17726 41712 18019 41714
rect 17726 41656 17958 41712
rect 18014 41656 18019 41712
rect 17726 41654 18019 41656
rect 1158 41516 1164 41580
rect 1228 41578 1234 41580
rect 1228 41518 2790 41578
rect 1228 41516 1234 41518
rect 2730 41442 2790 41518
rect 4838 41516 4844 41580
rect 4908 41578 4914 41580
rect 5165 41578 5231 41581
rect 6729 41578 6795 41581
rect 4908 41576 5231 41578
rect 4908 41520 5170 41576
rect 5226 41520 5231 41576
rect 4908 41518 5231 41520
rect 4908 41516 4914 41518
rect 5165 41515 5231 41518
rect 5398 41576 6795 41578
rect 5398 41520 6734 41576
rect 6790 41520 6795 41576
rect 5398 41518 6795 41520
rect 5398 41442 5458 41518
rect 6729 41515 6795 41518
rect 14774 41516 14780 41580
rect 14844 41578 14850 41580
rect 17726 41578 17786 41654
rect 17953 41651 18019 41654
rect 19014 41712 22251 41714
rect 19014 41656 22190 41712
rect 22246 41656 22251 41712
rect 19014 41654 22251 41656
rect 14844 41518 17786 41578
rect 18689 41578 18755 41581
rect 19014 41578 19074 41654
rect 22185 41651 22251 41654
rect 23197 41714 23263 41717
rect 25840 41714 26000 41744
rect 23197 41712 26000 41714
rect 23197 41656 23202 41712
rect 23258 41656 26000 41712
rect 23197 41654 26000 41656
rect 23197 41651 23263 41654
rect 25840 41624 26000 41654
rect 18689 41576 19074 41578
rect 18689 41520 18694 41576
rect 18750 41520 19074 41576
rect 18689 41518 19074 41520
rect 14844 41516 14850 41518
rect 18689 41515 18755 41518
rect 19190 41516 19196 41580
rect 19260 41578 19266 41580
rect 22001 41578 22067 41581
rect 19260 41576 22067 41578
rect 19260 41520 22006 41576
rect 22062 41520 22067 41576
rect 19260 41518 22067 41520
rect 19260 41516 19266 41518
rect 22001 41515 22067 41518
rect 2730 41382 5458 41442
rect 9254 41380 9260 41444
rect 9324 41442 9330 41444
rect 9397 41442 9463 41445
rect 9324 41440 9463 41442
rect 9324 41384 9402 41440
rect 9458 41384 9463 41440
rect 9324 41382 9463 41384
rect 9324 41380 9330 41382
rect 9397 41379 9463 41382
rect 16205 41444 16271 41445
rect 16205 41440 16252 41444
rect 16316 41442 16322 41444
rect 20989 41442 21055 41445
rect 22461 41442 22527 41445
rect 16205 41384 16210 41440
rect 16205 41380 16252 41384
rect 16316 41382 16362 41442
rect 20989 41440 22527 41442
rect 20989 41384 20994 41440
rect 21050 41384 22466 41440
rect 22522 41384 22527 41440
rect 20989 41382 22527 41384
rect 16316 41380 16322 41382
rect 16205 41379 16271 41380
rect 20989 41379 21055 41382
rect 22461 41379 22527 41382
rect 6880 41376 7196 41377
rect 6880 41312 6886 41376
rect 6950 41312 6966 41376
rect 7030 41312 7046 41376
rect 7110 41312 7126 41376
rect 7190 41312 7196 41376
rect 6880 41311 7196 41312
rect 12814 41376 13130 41377
rect 12814 41312 12820 41376
rect 12884 41312 12900 41376
rect 12964 41312 12980 41376
rect 13044 41312 13060 41376
rect 13124 41312 13130 41376
rect 12814 41311 13130 41312
rect 18748 41376 19064 41377
rect 18748 41312 18754 41376
rect 18818 41312 18834 41376
rect 18898 41312 18914 41376
rect 18978 41312 18994 41376
rect 19058 41312 19064 41376
rect 18748 41311 19064 41312
rect 24682 41376 24998 41377
rect 24682 41312 24688 41376
rect 24752 41312 24768 41376
rect 24832 41312 24848 41376
rect 24912 41312 24928 41376
rect 24992 41312 24998 41376
rect 24682 41311 24998 41312
rect 20529 41306 20595 41309
rect 23841 41306 23907 41309
rect 20529 41304 23907 41306
rect 20529 41248 20534 41304
rect 20590 41248 23846 41304
rect 23902 41248 23907 41304
rect 20529 41246 23907 41248
rect 20529 41243 20595 41246
rect 23841 41243 23907 41246
rect 3877 41170 3943 41173
rect 9121 41170 9187 41173
rect 3877 41168 9187 41170
rect 3877 41112 3882 41168
rect 3938 41112 9126 41168
rect 9182 41112 9187 41168
rect 3877 41110 9187 41112
rect 3877 41107 3943 41110
rect 9121 41107 9187 41110
rect 10225 41170 10291 41173
rect 22277 41170 22343 41173
rect 10225 41168 22343 41170
rect 10225 41112 10230 41168
rect 10286 41112 22282 41168
rect 22338 41112 22343 41168
rect 10225 41110 22343 41112
rect 10225 41107 10291 41110
rect 22277 41107 22343 41110
rect 25037 41170 25103 41173
rect 25840 41170 26000 41200
rect 25037 41168 26000 41170
rect 25037 41112 25042 41168
rect 25098 41112 26000 41168
rect 25037 41110 26000 41112
rect 25037 41107 25103 41110
rect 25840 41080 26000 41110
rect 1669 41034 1735 41037
rect 13486 41034 13492 41036
rect 1669 41032 13492 41034
rect 1669 40976 1674 41032
rect 1730 40976 13492 41032
rect 1669 40974 13492 40976
rect 1669 40971 1735 40974
rect 13486 40972 13492 40974
rect 13556 40972 13562 41036
rect 20897 41034 20963 41037
rect 22645 41034 22711 41037
rect 20897 41032 22711 41034
rect 20897 40976 20902 41032
rect 20958 40976 22650 41032
rect 22706 40976 22711 41032
rect 20897 40974 22711 40976
rect 20897 40971 20963 40974
rect 22645 40971 22711 40974
rect 3913 40832 4229 40833
rect 3913 40768 3919 40832
rect 3983 40768 3999 40832
rect 4063 40768 4079 40832
rect 4143 40768 4159 40832
rect 4223 40768 4229 40832
rect 3913 40767 4229 40768
rect 9847 40832 10163 40833
rect 9847 40768 9853 40832
rect 9917 40768 9933 40832
rect 9997 40768 10013 40832
rect 10077 40768 10093 40832
rect 10157 40768 10163 40832
rect 9847 40767 10163 40768
rect 15781 40832 16097 40833
rect 15781 40768 15787 40832
rect 15851 40768 15867 40832
rect 15931 40768 15947 40832
rect 16011 40768 16027 40832
rect 16091 40768 16097 40832
rect 15781 40767 16097 40768
rect 21715 40832 22031 40833
rect 21715 40768 21721 40832
rect 21785 40768 21801 40832
rect 21865 40768 21881 40832
rect 21945 40768 21961 40832
rect 22025 40768 22031 40832
rect 21715 40767 22031 40768
rect 20529 40762 20595 40765
rect 21449 40762 21515 40765
rect 20529 40760 21515 40762
rect 20529 40704 20534 40760
rect 20590 40704 21454 40760
rect 21510 40704 21515 40760
rect 20529 40702 21515 40704
rect 20529 40699 20595 40702
rect 21449 40699 21515 40702
rect 2221 40626 2287 40629
rect 2589 40626 2655 40629
rect 6821 40626 6887 40629
rect 17953 40626 18019 40629
rect 2221 40624 18019 40626
rect 2221 40568 2226 40624
rect 2282 40568 2594 40624
rect 2650 40568 6826 40624
rect 6882 40568 17958 40624
rect 18014 40568 18019 40624
rect 2221 40566 18019 40568
rect 2221 40563 2287 40566
rect 2589 40563 2655 40566
rect 6821 40563 6887 40566
rect 17953 40563 18019 40566
rect 20253 40626 20319 40629
rect 20662 40626 20668 40628
rect 20253 40624 20668 40626
rect 20253 40568 20258 40624
rect 20314 40568 20668 40624
rect 20253 40566 20668 40568
rect 20253 40563 20319 40566
rect 20662 40564 20668 40566
rect 20732 40564 20738 40628
rect 21265 40626 21331 40629
rect 23473 40626 23539 40629
rect 21265 40624 23539 40626
rect 21265 40568 21270 40624
rect 21326 40568 23478 40624
rect 23534 40568 23539 40624
rect 21265 40566 23539 40568
rect 21265 40563 21331 40566
rect 23473 40563 23539 40566
rect 23657 40626 23723 40629
rect 25840 40626 26000 40656
rect 23657 40624 26000 40626
rect 23657 40568 23662 40624
rect 23718 40568 26000 40624
rect 23657 40566 26000 40568
rect 23657 40563 23723 40566
rect 25840 40536 26000 40566
rect 2078 40428 2084 40492
rect 2148 40490 2154 40492
rect 2681 40490 2747 40493
rect 3877 40490 3943 40493
rect 2148 40488 3943 40490
rect 2148 40432 2686 40488
rect 2742 40432 3882 40488
rect 3938 40432 3943 40488
rect 2148 40430 3943 40432
rect 2148 40428 2154 40430
rect 2681 40427 2747 40430
rect 3877 40427 3943 40430
rect 4153 40490 4219 40493
rect 6913 40490 6979 40493
rect 4153 40488 6979 40490
rect 4153 40432 4158 40488
rect 4214 40432 6918 40488
rect 6974 40432 6979 40488
rect 4153 40430 6979 40432
rect 4153 40427 4219 40430
rect 6913 40427 6979 40430
rect 8293 40490 8359 40493
rect 10225 40490 10291 40493
rect 21081 40490 21147 40493
rect 8293 40488 10291 40490
rect 8293 40432 8298 40488
rect 8354 40432 10230 40488
rect 10286 40432 10291 40488
rect 8293 40430 10291 40432
rect 8293 40427 8359 40430
rect 10225 40427 10291 40430
rect 12390 40488 21147 40490
rect 12390 40432 21086 40488
rect 21142 40432 21147 40488
rect 12390 40430 21147 40432
rect 1710 40292 1716 40356
rect 1780 40354 1786 40356
rect 2037 40354 2103 40357
rect 5257 40354 5323 40357
rect 1780 40352 5323 40354
rect 1780 40296 2042 40352
rect 2098 40296 5262 40352
rect 5318 40296 5323 40352
rect 1780 40294 5323 40296
rect 1780 40292 1786 40294
rect 2037 40291 2103 40294
rect 5257 40291 5323 40294
rect 10317 40354 10383 40357
rect 12390 40354 12450 40430
rect 21081 40427 21147 40430
rect 21265 40490 21331 40493
rect 22277 40490 22343 40493
rect 21265 40488 22343 40490
rect 21265 40432 21270 40488
rect 21326 40432 22282 40488
rect 22338 40432 22343 40488
rect 21265 40430 22343 40432
rect 21265 40427 21331 40430
rect 22277 40427 22343 40430
rect 22093 40354 22159 40357
rect 10317 40352 12450 40354
rect 10317 40296 10322 40352
rect 10378 40296 12450 40352
rect 10317 40294 12450 40296
rect 19198 40352 22159 40354
rect 19198 40296 22098 40352
rect 22154 40296 22159 40352
rect 19198 40294 22159 40296
rect 10317 40291 10383 40294
rect 6880 40288 7196 40289
rect 6880 40224 6886 40288
rect 6950 40224 6966 40288
rect 7030 40224 7046 40288
rect 7110 40224 7126 40288
rect 7190 40224 7196 40288
rect 6880 40223 7196 40224
rect 12814 40288 13130 40289
rect 12814 40224 12820 40288
rect 12884 40224 12900 40288
rect 12964 40224 12980 40288
rect 13044 40224 13060 40288
rect 13124 40224 13130 40288
rect 12814 40223 13130 40224
rect 18748 40288 19064 40289
rect 18748 40224 18754 40288
rect 18818 40224 18834 40288
rect 18898 40224 18914 40288
rect 18978 40224 18994 40288
rect 19058 40224 19064 40288
rect 18748 40223 19064 40224
rect 657 40218 723 40221
rect 5441 40218 5507 40221
rect 657 40216 5507 40218
rect 657 40160 662 40216
rect 718 40160 5446 40216
rect 5502 40160 5507 40216
rect 657 40158 5507 40160
rect 657 40155 723 40158
rect 5441 40155 5507 40158
rect 933 40082 999 40085
rect 4245 40082 4311 40085
rect 933 40080 4311 40082
rect 933 40024 938 40080
rect 994 40024 4250 40080
rect 4306 40024 4311 40080
rect 933 40022 4311 40024
rect 933 40019 999 40022
rect 4245 40019 4311 40022
rect 7782 40020 7788 40084
rect 7852 40082 7858 40084
rect 8201 40082 8267 40085
rect 9673 40084 9739 40085
rect 9622 40082 9628 40084
rect 7852 40080 8267 40082
rect 7852 40024 8206 40080
rect 8262 40024 8267 40080
rect 7852 40022 8267 40024
rect 9582 40022 9628 40082
rect 9692 40080 9739 40084
rect 9734 40024 9739 40080
rect 7852 40020 7858 40022
rect 8201 40019 8267 40022
rect 9622 40020 9628 40022
rect 9692 40020 9739 40024
rect 9673 40019 9739 40020
rect 10225 40082 10291 40085
rect 10685 40082 10751 40085
rect 10225 40080 10751 40082
rect 10225 40024 10230 40080
rect 10286 40024 10690 40080
rect 10746 40024 10751 40080
rect 10225 40022 10751 40024
rect 10225 40019 10291 40022
rect 10685 40019 10751 40022
rect 16849 40082 16915 40085
rect 19198 40082 19258 40294
rect 22093 40291 22159 40294
rect 24682 40288 24998 40289
rect 24682 40224 24688 40288
rect 24752 40224 24768 40288
rect 24832 40224 24848 40288
rect 24912 40224 24928 40288
rect 24992 40224 24998 40288
rect 24682 40223 24998 40224
rect 19885 40218 19951 40221
rect 23473 40218 23539 40221
rect 19885 40216 23539 40218
rect 19885 40160 19890 40216
rect 19946 40160 23478 40216
rect 23534 40160 23539 40216
rect 19885 40158 23539 40160
rect 19885 40155 19951 40158
rect 23473 40155 23539 40158
rect 16849 40080 19258 40082
rect 16849 40024 16854 40080
rect 16910 40024 19258 40080
rect 16849 40022 19258 40024
rect 19425 40082 19491 40085
rect 19558 40082 19564 40084
rect 19425 40080 19564 40082
rect 19425 40024 19430 40080
rect 19486 40024 19564 40080
rect 19425 40022 19564 40024
rect 16849 40019 16915 40022
rect 19425 40019 19491 40022
rect 19558 40020 19564 40022
rect 19628 40020 19634 40084
rect 20897 40082 20963 40085
rect 21725 40082 21791 40085
rect 20897 40080 21791 40082
rect 20897 40024 20902 40080
rect 20958 40024 21730 40080
rect 21786 40024 21791 40080
rect 20897 40022 21791 40024
rect 20897 40019 20963 40022
rect 21725 40019 21791 40022
rect 24209 40082 24275 40085
rect 25840 40082 26000 40112
rect 24209 40080 26000 40082
rect 24209 40024 24214 40080
rect 24270 40024 26000 40080
rect 24209 40022 26000 40024
rect 24209 40019 24275 40022
rect 25840 39992 26000 40022
rect 3969 39946 4035 39949
rect 10542 39946 10548 39948
rect 3969 39944 10548 39946
rect 3969 39888 3974 39944
rect 4030 39888 10548 39944
rect 3969 39886 10548 39888
rect 3969 39883 4035 39886
rect 10542 39884 10548 39886
rect 10612 39884 10618 39948
rect 20161 39946 20227 39949
rect 23749 39946 23815 39949
rect 20161 39944 23815 39946
rect 20161 39888 20166 39944
rect 20222 39888 23754 39944
rect 23810 39888 23815 39944
rect 20161 39886 23815 39888
rect 20161 39883 20227 39886
rect 23749 39883 23815 39886
rect 0 39810 160 39840
rect 2405 39810 2471 39813
rect 0 39808 2471 39810
rect 0 39752 2410 39808
rect 2466 39752 2471 39808
rect 0 39750 2471 39752
rect 0 39720 160 39750
rect 2405 39747 2471 39750
rect 3913 39744 4229 39745
rect 3913 39680 3919 39744
rect 3983 39680 3999 39744
rect 4063 39680 4079 39744
rect 4143 39680 4159 39744
rect 4223 39680 4229 39744
rect 3913 39679 4229 39680
rect 9847 39744 10163 39745
rect 9847 39680 9853 39744
rect 9917 39680 9933 39744
rect 9997 39680 10013 39744
rect 10077 39680 10093 39744
rect 10157 39680 10163 39744
rect 9847 39679 10163 39680
rect 15781 39744 16097 39745
rect 15781 39680 15787 39744
rect 15851 39680 15867 39744
rect 15931 39680 15947 39744
rect 16011 39680 16027 39744
rect 16091 39680 16097 39744
rect 15781 39679 16097 39680
rect 21715 39744 22031 39745
rect 21715 39680 21721 39744
rect 21785 39680 21801 39744
rect 21865 39680 21881 39744
rect 21945 39680 21961 39744
rect 22025 39680 22031 39744
rect 21715 39679 22031 39680
rect 0 39538 160 39568
rect 1393 39538 1459 39541
rect 0 39536 1459 39538
rect 0 39480 1398 39536
rect 1454 39480 1459 39536
rect 0 39478 1459 39480
rect 0 39448 160 39478
rect 1393 39475 1459 39478
rect 2497 39538 2563 39541
rect 3601 39538 3667 39541
rect 6821 39538 6887 39541
rect 2497 39536 6887 39538
rect 2497 39480 2502 39536
rect 2558 39480 3606 39536
rect 3662 39480 6826 39536
rect 6882 39480 6887 39536
rect 2497 39478 6887 39480
rect 2497 39475 2563 39478
rect 3601 39475 3667 39478
rect 6821 39475 6887 39478
rect 7005 39538 7071 39541
rect 9397 39538 9463 39541
rect 7005 39536 9463 39538
rect 7005 39480 7010 39536
rect 7066 39480 9402 39536
rect 9458 39480 9463 39536
rect 7005 39478 9463 39480
rect 7005 39475 7071 39478
rect 9397 39475 9463 39478
rect 20069 39538 20135 39541
rect 23473 39538 23539 39541
rect 20069 39536 23539 39538
rect 20069 39480 20074 39536
rect 20130 39480 23478 39536
rect 23534 39480 23539 39536
rect 20069 39478 23539 39480
rect 20069 39475 20135 39478
rect 23473 39475 23539 39478
rect 24393 39538 24459 39541
rect 25840 39538 26000 39568
rect 24393 39536 26000 39538
rect 24393 39480 24398 39536
rect 24454 39480 26000 39536
rect 24393 39478 26000 39480
rect 24393 39475 24459 39478
rect 25840 39448 26000 39478
rect 7966 39340 7972 39404
rect 8036 39402 8042 39404
rect 19742 39402 19748 39404
rect 8036 39342 19748 39402
rect 8036 39340 8042 39342
rect 19742 39340 19748 39342
rect 19812 39340 19818 39404
rect 21357 39402 21423 39405
rect 22277 39402 22343 39405
rect 21357 39400 22343 39402
rect 21357 39344 21362 39400
rect 21418 39344 22282 39400
rect 22338 39344 22343 39400
rect 21357 39342 22343 39344
rect 21357 39339 21423 39342
rect 22277 39339 22343 39342
rect 22461 39402 22527 39405
rect 24577 39402 24643 39405
rect 22461 39400 24643 39402
rect 22461 39344 22466 39400
rect 22522 39344 24582 39400
rect 24638 39344 24643 39400
rect 22461 39342 24643 39344
rect 22461 39339 22527 39342
rect 24577 39339 24643 39342
rect 0 39266 160 39296
rect 2313 39266 2379 39269
rect 0 39264 2379 39266
rect 0 39208 2318 39264
rect 2374 39208 2379 39264
rect 0 39206 2379 39208
rect 0 39176 160 39206
rect 2313 39203 2379 39206
rect 20805 39266 20871 39269
rect 23841 39266 23907 39269
rect 20805 39264 23907 39266
rect 20805 39208 20810 39264
rect 20866 39208 23846 39264
rect 23902 39208 23907 39264
rect 20805 39206 23907 39208
rect 20805 39203 20871 39206
rect 23841 39203 23907 39206
rect 6880 39200 7196 39201
rect 6880 39136 6886 39200
rect 6950 39136 6966 39200
rect 7030 39136 7046 39200
rect 7110 39136 7126 39200
rect 7190 39136 7196 39200
rect 6880 39135 7196 39136
rect 12814 39200 13130 39201
rect 12814 39136 12820 39200
rect 12884 39136 12900 39200
rect 12964 39136 12980 39200
rect 13044 39136 13060 39200
rect 13124 39136 13130 39200
rect 12814 39135 13130 39136
rect 18748 39200 19064 39201
rect 18748 39136 18754 39200
rect 18818 39136 18834 39200
rect 18898 39136 18914 39200
rect 18978 39136 18994 39200
rect 19058 39136 19064 39200
rect 18748 39135 19064 39136
rect 24682 39200 24998 39201
rect 24682 39136 24688 39200
rect 24752 39136 24768 39200
rect 24832 39136 24848 39200
rect 24912 39136 24928 39200
rect 24992 39136 24998 39200
rect 24682 39135 24998 39136
rect 1485 39130 1551 39133
rect 798 39128 1551 39130
rect 798 39072 1490 39128
rect 1546 39072 1551 39128
rect 798 39070 1551 39072
rect 0 38994 160 39024
rect 798 38994 858 39070
rect 1485 39067 1551 39070
rect 0 38934 858 38994
rect 3417 38994 3483 38997
rect 6637 38994 6703 38997
rect 3417 38992 6703 38994
rect 3417 38936 3422 38992
rect 3478 38936 6642 38992
rect 6698 38936 6703 38992
rect 3417 38934 6703 38936
rect 0 38904 160 38934
rect 3417 38931 3483 38934
rect 6637 38931 6703 38934
rect 7281 38994 7347 38997
rect 8201 38994 8267 38997
rect 7281 38992 8267 38994
rect 7281 38936 7286 38992
rect 7342 38936 8206 38992
rect 8262 38936 8267 38992
rect 7281 38934 8267 38936
rect 7281 38931 7347 38934
rect 8201 38931 8267 38934
rect 13670 38932 13676 38996
rect 13740 38994 13746 38996
rect 22502 38994 22508 38996
rect 13740 38934 22508 38994
rect 13740 38932 13746 38934
rect 22502 38932 22508 38934
rect 22572 38932 22578 38996
rect 24117 38994 24183 38997
rect 25840 38994 26000 39024
rect 24117 38992 26000 38994
rect 24117 38936 24122 38992
rect 24178 38936 26000 38992
rect 24117 38934 26000 38936
rect 24117 38931 24183 38934
rect 25840 38904 26000 38934
rect 11789 38858 11855 38861
rect 22318 38858 22324 38860
rect 3742 38798 4354 38858
rect 0 38722 160 38752
rect 1393 38722 1459 38725
rect 1945 38724 2011 38725
rect 1894 38722 1900 38724
rect 0 38720 1459 38722
rect 0 38664 1398 38720
rect 1454 38664 1459 38720
rect 0 38662 1459 38664
rect 1854 38662 1900 38722
rect 1964 38720 2011 38724
rect 2006 38664 2011 38720
rect 0 38632 160 38662
rect 1393 38659 1459 38662
rect 1894 38660 1900 38662
rect 1964 38660 2011 38664
rect 1945 38659 2011 38660
rect 606 38524 612 38588
rect 676 38586 682 38588
rect 3742 38586 3802 38798
rect 3913 38656 4229 38657
rect 3913 38592 3919 38656
rect 3983 38592 3999 38656
rect 4063 38592 4079 38656
rect 4143 38592 4159 38656
rect 4223 38592 4229 38656
rect 3913 38591 4229 38592
rect 676 38526 3802 38586
rect 4294 38586 4354 38798
rect 11789 38856 22324 38858
rect 11789 38800 11794 38856
rect 11850 38800 22324 38856
rect 11789 38798 22324 38800
rect 11789 38795 11855 38798
rect 22318 38796 22324 38798
rect 22388 38796 22394 38860
rect 11329 38722 11395 38725
rect 14089 38722 14155 38725
rect 11329 38720 14155 38722
rect 11329 38664 11334 38720
rect 11390 38664 14094 38720
rect 14150 38664 14155 38720
rect 11329 38662 14155 38664
rect 11329 38659 11395 38662
rect 14089 38659 14155 38662
rect 16665 38722 16731 38725
rect 19190 38722 19196 38724
rect 16665 38720 19196 38722
rect 16665 38664 16670 38720
rect 16726 38664 19196 38720
rect 16665 38662 19196 38664
rect 16665 38659 16731 38662
rect 19190 38660 19196 38662
rect 19260 38660 19266 38724
rect 21265 38722 21331 38725
rect 21398 38722 21404 38724
rect 21265 38720 21404 38722
rect 21265 38664 21270 38720
rect 21326 38664 21404 38720
rect 21265 38662 21404 38664
rect 21265 38659 21331 38662
rect 21398 38660 21404 38662
rect 21468 38660 21474 38724
rect 9847 38656 10163 38657
rect 9847 38592 9853 38656
rect 9917 38592 9933 38656
rect 9997 38592 10013 38656
rect 10077 38592 10093 38656
rect 10157 38592 10163 38656
rect 9847 38591 10163 38592
rect 15781 38656 16097 38657
rect 15781 38592 15787 38656
rect 15851 38592 15867 38656
rect 15931 38592 15947 38656
rect 16011 38592 16027 38656
rect 16091 38592 16097 38656
rect 15781 38591 16097 38592
rect 21715 38656 22031 38657
rect 21715 38592 21721 38656
rect 21785 38592 21801 38656
rect 21865 38592 21881 38656
rect 21945 38592 21961 38656
rect 22025 38592 22031 38656
rect 21715 38591 22031 38592
rect 7373 38586 7439 38589
rect 4294 38584 7439 38586
rect 4294 38528 7378 38584
rect 7434 38528 7439 38584
rect 4294 38526 7439 38528
rect 676 38524 682 38526
rect 7373 38523 7439 38526
rect 24393 38586 24459 38589
rect 24393 38584 25146 38586
rect 24393 38528 24398 38584
rect 24454 38528 25146 38584
rect 24393 38526 25146 38528
rect 24393 38523 24459 38526
rect 0 38450 160 38480
rect 1485 38450 1551 38453
rect 12566 38450 12572 38452
rect 0 38448 1551 38450
rect 0 38392 1490 38448
rect 1546 38392 1551 38448
rect 0 38390 1551 38392
rect 0 38360 160 38390
rect 1485 38387 1551 38390
rect 2730 38390 12572 38450
rect 1669 38314 1735 38317
rect 2730 38314 2790 38390
rect 12566 38388 12572 38390
rect 12636 38388 12642 38452
rect 25086 38450 25146 38526
rect 25840 38450 26000 38480
rect 25086 38390 26000 38450
rect 25840 38360 26000 38390
rect 1669 38312 2790 38314
rect 1669 38256 1674 38312
rect 1730 38256 2790 38312
rect 1669 38254 2790 38256
rect 1669 38251 1735 38254
rect 2998 38252 3004 38316
rect 3068 38314 3074 38316
rect 3233 38314 3299 38317
rect 8201 38314 8267 38317
rect 3068 38312 8267 38314
rect 3068 38256 3238 38312
rect 3294 38256 8206 38312
rect 8262 38256 8267 38312
rect 3068 38254 8267 38256
rect 3068 38252 3074 38254
rect 3233 38251 3299 38254
rect 8201 38251 8267 38254
rect 0 38178 160 38208
rect 1301 38178 1367 38181
rect 0 38176 1367 38178
rect 0 38120 1306 38176
rect 1362 38120 1367 38176
rect 0 38118 1367 38120
rect 0 38088 160 38118
rect 1301 38115 1367 38118
rect 6880 38112 7196 38113
rect 6880 38048 6886 38112
rect 6950 38048 6966 38112
rect 7030 38048 7046 38112
rect 7110 38048 7126 38112
rect 7190 38048 7196 38112
rect 6880 38047 7196 38048
rect 12814 38112 13130 38113
rect 12814 38048 12820 38112
rect 12884 38048 12900 38112
rect 12964 38048 12980 38112
rect 13044 38048 13060 38112
rect 13124 38048 13130 38112
rect 12814 38047 13130 38048
rect 18748 38112 19064 38113
rect 18748 38048 18754 38112
rect 18818 38048 18834 38112
rect 18898 38048 18914 38112
rect 18978 38048 18994 38112
rect 19058 38048 19064 38112
rect 18748 38047 19064 38048
rect 24682 38112 24998 38113
rect 24682 38048 24688 38112
rect 24752 38048 24768 38112
rect 24832 38048 24848 38112
rect 24912 38048 24928 38112
rect 24992 38048 24998 38112
rect 24682 38047 24998 38048
rect 974 37980 980 38044
rect 1044 38042 1050 38044
rect 4613 38042 4679 38045
rect 1044 38040 4679 38042
rect 1044 37984 4618 38040
rect 4674 37984 4679 38040
rect 1044 37982 4679 37984
rect 1044 37980 1050 37982
rect 4613 37979 4679 37982
rect 0 37906 160 37936
rect 2865 37906 2931 37909
rect 0 37904 2931 37906
rect 0 37848 2870 37904
rect 2926 37848 2931 37904
rect 0 37846 2931 37848
rect 0 37816 160 37846
rect 2865 37843 2931 37846
rect 3550 37844 3556 37908
rect 3620 37906 3626 37908
rect 4061 37906 4127 37909
rect 3620 37904 4127 37906
rect 3620 37848 4066 37904
rect 4122 37848 4127 37904
rect 3620 37846 4127 37848
rect 3620 37844 3626 37846
rect 4061 37843 4127 37846
rect 6085 37906 6151 37909
rect 16614 37906 16620 37908
rect 6085 37904 16620 37906
rect 6085 37848 6090 37904
rect 6146 37848 16620 37904
rect 6085 37846 16620 37848
rect 6085 37843 6151 37846
rect 16614 37844 16620 37846
rect 16684 37844 16690 37908
rect 24117 37906 24183 37909
rect 25840 37906 26000 37936
rect 24117 37904 26000 37906
rect 24117 37848 24122 37904
rect 24178 37848 26000 37904
rect 24117 37846 26000 37848
rect 24117 37843 24183 37846
rect 25840 37816 26000 37846
rect 4153 37770 4219 37773
rect 4654 37770 4660 37772
rect 4153 37768 4660 37770
rect 4153 37712 4158 37768
rect 4214 37712 4660 37768
rect 4153 37710 4660 37712
rect 4153 37707 4219 37710
rect 4654 37708 4660 37710
rect 4724 37708 4730 37772
rect 8017 37770 8083 37773
rect 8886 37770 8892 37772
rect 8017 37768 8892 37770
rect 8017 37712 8022 37768
rect 8078 37712 8892 37768
rect 8017 37710 8892 37712
rect 8017 37707 8083 37710
rect 8886 37708 8892 37710
rect 8956 37708 8962 37772
rect 0 37634 160 37664
rect 1209 37634 1275 37637
rect 0 37632 1275 37634
rect 0 37576 1214 37632
rect 1270 37576 1275 37632
rect 0 37574 1275 37576
rect 0 37544 160 37574
rect 1209 37571 1275 37574
rect 3913 37568 4229 37569
rect 3913 37504 3919 37568
rect 3983 37504 3999 37568
rect 4063 37504 4079 37568
rect 4143 37504 4159 37568
rect 4223 37504 4229 37568
rect 3913 37503 4229 37504
rect 9847 37568 10163 37569
rect 9847 37504 9853 37568
rect 9917 37504 9933 37568
rect 9997 37504 10013 37568
rect 10077 37504 10093 37568
rect 10157 37504 10163 37568
rect 9847 37503 10163 37504
rect 15781 37568 16097 37569
rect 15781 37504 15787 37568
rect 15851 37504 15867 37568
rect 15931 37504 15947 37568
rect 16011 37504 16027 37568
rect 16091 37504 16097 37568
rect 15781 37503 16097 37504
rect 21715 37568 22031 37569
rect 21715 37504 21721 37568
rect 21785 37504 21801 37568
rect 21865 37504 21881 37568
rect 21945 37504 21961 37568
rect 22025 37504 22031 37568
rect 21715 37503 22031 37504
rect 0 37362 160 37392
rect 2773 37362 2839 37365
rect 0 37360 2839 37362
rect 0 37304 2778 37360
rect 2834 37304 2839 37360
rect 0 37302 2839 37304
rect 0 37272 160 37302
rect 2773 37299 2839 37302
rect 7741 37362 7807 37365
rect 8518 37362 8524 37364
rect 7741 37360 8524 37362
rect 7741 37304 7746 37360
rect 7802 37304 8524 37360
rect 7741 37302 8524 37304
rect 7741 37299 7807 37302
rect 8518 37300 8524 37302
rect 8588 37300 8594 37364
rect 24393 37362 24459 37365
rect 25840 37362 26000 37392
rect 24393 37360 26000 37362
rect 24393 37304 24398 37360
rect 24454 37304 26000 37360
rect 24393 37302 26000 37304
rect 24393 37299 24459 37302
rect 25840 37272 26000 37302
rect 0 37090 160 37120
rect 1577 37090 1643 37093
rect 0 37088 1643 37090
rect 0 37032 1582 37088
rect 1638 37032 1643 37088
rect 0 37030 1643 37032
rect 0 37000 160 37030
rect 1577 37027 1643 37030
rect 6880 37024 7196 37025
rect 6880 36960 6886 37024
rect 6950 36960 6966 37024
rect 7030 36960 7046 37024
rect 7110 36960 7126 37024
rect 7190 36960 7196 37024
rect 6880 36959 7196 36960
rect 12814 37024 13130 37025
rect 12814 36960 12820 37024
rect 12884 36960 12900 37024
rect 12964 36960 12980 37024
rect 13044 36960 13060 37024
rect 13124 36960 13130 37024
rect 12814 36959 13130 36960
rect 18748 37024 19064 37025
rect 18748 36960 18754 37024
rect 18818 36960 18834 37024
rect 18898 36960 18914 37024
rect 18978 36960 18994 37024
rect 19058 36960 19064 37024
rect 18748 36959 19064 36960
rect 24682 37024 24998 37025
rect 24682 36960 24688 37024
rect 24752 36960 24768 37024
rect 24832 36960 24848 37024
rect 24912 36960 24928 37024
rect 24992 36960 24998 37024
rect 24682 36959 24998 36960
rect 0 36818 160 36848
rect 3877 36818 3943 36821
rect 0 36816 3943 36818
rect 0 36760 3882 36816
rect 3938 36760 3943 36816
rect 0 36758 3943 36760
rect 0 36728 160 36758
rect 3877 36755 3943 36758
rect 24117 36818 24183 36821
rect 25840 36818 26000 36848
rect 24117 36816 26000 36818
rect 24117 36760 24122 36816
rect 24178 36760 26000 36816
rect 24117 36758 26000 36760
rect 24117 36755 24183 36758
rect 25840 36728 26000 36758
rect 790 36620 796 36684
rect 860 36682 866 36684
rect 1669 36682 1735 36685
rect 860 36680 1735 36682
rect 860 36624 1674 36680
rect 1730 36624 1735 36680
rect 860 36622 1735 36624
rect 860 36620 866 36622
rect 1669 36619 1735 36622
rect 0 36546 160 36576
rect 3233 36546 3299 36549
rect 0 36544 3299 36546
rect 0 36488 3238 36544
rect 3294 36488 3299 36544
rect 0 36486 3299 36488
rect 0 36456 160 36486
rect 3233 36483 3299 36486
rect 3913 36480 4229 36481
rect 3913 36416 3919 36480
rect 3983 36416 3999 36480
rect 4063 36416 4079 36480
rect 4143 36416 4159 36480
rect 4223 36416 4229 36480
rect 3913 36415 4229 36416
rect 9847 36480 10163 36481
rect 9847 36416 9853 36480
rect 9917 36416 9933 36480
rect 9997 36416 10013 36480
rect 10077 36416 10093 36480
rect 10157 36416 10163 36480
rect 9847 36415 10163 36416
rect 15781 36480 16097 36481
rect 15781 36416 15787 36480
rect 15851 36416 15867 36480
rect 15931 36416 15947 36480
rect 16011 36416 16027 36480
rect 16091 36416 16097 36480
rect 15781 36415 16097 36416
rect 21715 36480 22031 36481
rect 21715 36416 21721 36480
rect 21785 36416 21801 36480
rect 21865 36416 21881 36480
rect 21945 36416 21961 36480
rect 22025 36416 22031 36480
rect 21715 36415 22031 36416
rect 0 36274 160 36304
rect 3049 36274 3115 36277
rect 0 36272 3115 36274
rect 0 36216 3054 36272
rect 3110 36216 3115 36272
rect 0 36214 3115 36216
rect 0 36184 160 36214
rect 3049 36211 3115 36214
rect 4337 36272 4403 36277
rect 4337 36216 4342 36272
rect 4398 36216 4403 36272
rect 4337 36211 4403 36216
rect 4521 36274 4587 36277
rect 12433 36274 12499 36277
rect 4521 36272 12499 36274
rect 4521 36216 4526 36272
rect 4582 36216 12438 36272
rect 12494 36216 12499 36272
rect 4521 36214 12499 36216
rect 4521 36211 4587 36214
rect 12433 36211 12499 36214
rect 24393 36274 24459 36277
rect 25840 36274 26000 36304
rect 24393 36272 26000 36274
rect 24393 36216 24398 36272
rect 24454 36216 26000 36272
rect 24393 36214 26000 36216
rect 24393 36211 24459 36214
rect 473 36138 539 36141
rect 4340 36138 4400 36211
rect 25840 36184 26000 36214
rect 473 36136 4400 36138
rect 473 36080 478 36136
rect 534 36080 4400 36136
rect 473 36078 4400 36080
rect 5165 36138 5231 36141
rect 8017 36138 8083 36141
rect 5165 36136 8083 36138
rect 5165 36080 5170 36136
rect 5226 36080 8022 36136
rect 8078 36080 8083 36136
rect 5165 36078 8083 36080
rect 473 36075 539 36078
rect 5165 36075 5231 36078
rect 8017 36075 8083 36078
rect 21214 36076 21220 36140
rect 21284 36138 21290 36140
rect 23013 36138 23079 36141
rect 21284 36136 23079 36138
rect 21284 36080 23018 36136
rect 23074 36080 23079 36136
rect 21284 36078 23079 36080
rect 21284 36076 21290 36078
rect 23013 36075 23079 36078
rect 0 36002 160 36032
rect 1301 36002 1367 36005
rect 0 36000 1367 36002
rect 0 35944 1306 36000
rect 1362 35944 1367 36000
rect 0 35942 1367 35944
rect 0 35912 160 35942
rect 1301 35939 1367 35942
rect 3969 36002 4035 36005
rect 4797 36002 4863 36005
rect 3969 36000 4863 36002
rect 3969 35944 3974 36000
rect 4030 35944 4802 36000
rect 4858 35944 4863 36000
rect 3969 35942 4863 35944
rect 3969 35939 4035 35942
rect 4797 35939 4863 35942
rect 7925 36002 7991 36005
rect 10041 36002 10107 36005
rect 10358 36002 10364 36004
rect 7925 36000 10364 36002
rect 7925 35944 7930 36000
rect 7986 35944 10046 36000
rect 10102 35944 10364 36000
rect 7925 35942 10364 35944
rect 7925 35939 7991 35942
rect 10041 35939 10107 35942
rect 10358 35940 10364 35942
rect 10428 35940 10434 36004
rect 6880 35936 7196 35937
rect 6880 35872 6886 35936
rect 6950 35872 6966 35936
rect 7030 35872 7046 35936
rect 7110 35872 7126 35936
rect 7190 35872 7196 35936
rect 6880 35871 7196 35872
rect 12814 35936 13130 35937
rect 12814 35872 12820 35936
rect 12884 35872 12900 35936
rect 12964 35872 12980 35936
rect 13044 35872 13060 35936
rect 13124 35872 13130 35936
rect 12814 35871 13130 35872
rect 18748 35936 19064 35937
rect 18748 35872 18754 35936
rect 18818 35872 18834 35936
rect 18898 35872 18914 35936
rect 18978 35872 18994 35936
rect 19058 35872 19064 35936
rect 18748 35871 19064 35872
rect 24682 35936 24998 35937
rect 24682 35872 24688 35936
rect 24752 35872 24768 35936
rect 24832 35872 24848 35936
rect 24912 35872 24928 35936
rect 24992 35872 24998 35936
rect 24682 35871 24998 35872
rect 3182 35804 3188 35868
rect 3252 35866 3258 35868
rect 3785 35866 3851 35869
rect 3252 35864 3851 35866
rect 3252 35808 3790 35864
rect 3846 35808 3851 35864
rect 3252 35806 3851 35808
rect 3252 35804 3258 35806
rect 3785 35803 3851 35806
rect 24117 35866 24183 35869
rect 24117 35864 24594 35866
rect 24117 35808 24122 35864
rect 24178 35808 24594 35864
rect 24117 35806 24594 35808
rect 24117 35803 24183 35806
rect 0 35730 160 35760
rect 4337 35730 4403 35733
rect 0 35728 4403 35730
rect 0 35672 4342 35728
rect 4398 35672 4403 35728
rect 0 35670 4403 35672
rect 24534 35730 24594 35806
rect 25840 35730 26000 35760
rect 24534 35670 26000 35730
rect 0 35640 160 35670
rect 4337 35667 4403 35670
rect 25840 35640 26000 35670
rect 1669 35594 1735 35597
rect 4061 35594 4127 35597
rect 6637 35594 6703 35597
rect 8753 35596 8819 35597
rect 1669 35592 3802 35594
rect 1669 35536 1674 35592
rect 1730 35536 3802 35592
rect 1669 35534 3802 35536
rect 1669 35531 1735 35534
rect 0 35458 160 35488
rect 2773 35458 2839 35461
rect 0 35456 2839 35458
rect 0 35400 2778 35456
rect 2834 35400 2839 35456
rect 0 35398 2839 35400
rect 0 35368 160 35398
rect 2773 35395 2839 35398
rect 0 35186 160 35216
rect 3182 35186 3188 35188
rect 0 35126 3188 35186
rect 0 35096 160 35126
rect 3182 35124 3188 35126
rect 3252 35124 3258 35188
rect 3742 35186 3802 35534
rect 4061 35592 6703 35594
rect 4061 35536 4066 35592
rect 4122 35536 6642 35592
rect 6698 35536 6703 35592
rect 4061 35534 6703 35536
rect 4061 35531 4127 35534
rect 6637 35531 6703 35534
rect 8702 35532 8708 35596
rect 8772 35594 8819 35596
rect 11973 35594 12039 35597
rect 15285 35594 15351 35597
rect 8772 35592 8864 35594
rect 8814 35536 8864 35592
rect 8772 35534 8864 35536
rect 11973 35592 15351 35594
rect 11973 35536 11978 35592
rect 12034 35536 15290 35592
rect 15346 35536 15351 35592
rect 11973 35534 15351 35536
rect 8772 35532 8819 35534
rect 8753 35531 8819 35532
rect 11973 35531 12039 35534
rect 15285 35531 15351 35534
rect 3913 35392 4229 35393
rect 3913 35328 3919 35392
rect 3983 35328 3999 35392
rect 4063 35328 4079 35392
rect 4143 35328 4159 35392
rect 4223 35328 4229 35392
rect 3913 35327 4229 35328
rect 9847 35392 10163 35393
rect 9847 35328 9853 35392
rect 9917 35328 9933 35392
rect 9997 35328 10013 35392
rect 10077 35328 10093 35392
rect 10157 35328 10163 35392
rect 9847 35327 10163 35328
rect 15781 35392 16097 35393
rect 15781 35328 15787 35392
rect 15851 35328 15867 35392
rect 15931 35328 15947 35392
rect 16011 35328 16027 35392
rect 16091 35328 16097 35392
rect 15781 35327 16097 35328
rect 21715 35392 22031 35393
rect 21715 35328 21721 35392
rect 21785 35328 21801 35392
rect 21865 35328 21881 35392
rect 21945 35328 21961 35392
rect 22025 35328 22031 35392
rect 21715 35327 22031 35328
rect 10317 35186 10383 35189
rect 3742 35184 10383 35186
rect 3742 35128 10322 35184
rect 10378 35128 10383 35184
rect 3742 35126 10383 35128
rect 10317 35123 10383 35126
rect 24393 35186 24459 35189
rect 25840 35186 26000 35216
rect 24393 35184 26000 35186
rect 24393 35128 24398 35184
rect 24454 35128 26000 35184
rect 24393 35126 26000 35128
rect 24393 35123 24459 35126
rect 25840 35096 26000 35126
rect 3141 35050 3207 35053
rect 3785 35050 3851 35053
rect 4613 35050 4679 35053
rect 3141 35048 4679 35050
rect 3141 34992 3146 35048
rect 3202 34992 3790 35048
rect 3846 34992 4618 35048
rect 4674 34992 4679 35048
rect 3141 34990 4679 34992
rect 3141 34987 3207 34990
rect 3785 34987 3851 34990
rect 4613 34987 4679 34990
rect 13997 35050 14063 35053
rect 20621 35050 20687 35053
rect 13997 35048 20687 35050
rect 13997 34992 14002 35048
rect 14058 34992 20626 35048
rect 20682 34992 20687 35048
rect 13997 34990 20687 34992
rect 13997 34987 14063 34990
rect 20621 34987 20687 34990
rect 0 34914 160 34944
rect 1301 34914 1367 34917
rect 0 34912 1367 34914
rect 0 34856 1306 34912
rect 1362 34856 1367 34912
rect 0 34854 1367 34856
rect 0 34824 160 34854
rect 1301 34851 1367 34854
rect 4797 34914 4863 34917
rect 5574 34914 5580 34916
rect 4797 34912 5580 34914
rect 4797 34856 4802 34912
rect 4858 34856 5580 34912
rect 4797 34854 5580 34856
rect 4797 34851 4863 34854
rect 5574 34852 5580 34854
rect 5644 34852 5650 34916
rect 13445 34914 13511 34917
rect 18229 34914 18295 34917
rect 13445 34912 18295 34914
rect 13445 34856 13450 34912
rect 13506 34856 18234 34912
rect 18290 34856 18295 34912
rect 13445 34854 18295 34856
rect 13445 34851 13511 34854
rect 18229 34851 18295 34854
rect 6880 34848 7196 34849
rect 6880 34784 6886 34848
rect 6950 34784 6966 34848
rect 7030 34784 7046 34848
rect 7110 34784 7126 34848
rect 7190 34784 7196 34848
rect 6880 34783 7196 34784
rect 12814 34848 13130 34849
rect 12814 34784 12820 34848
rect 12884 34784 12900 34848
rect 12964 34784 12980 34848
rect 13044 34784 13060 34848
rect 13124 34784 13130 34848
rect 12814 34783 13130 34784
rect 18748 34848 19064 34849
rect 18748 34784 18754 34848
rect 18818 34784 18834 34848
rect 18898 34784 18914 34848
rect 18978 34784 18994 34848
rect 19058 34784 19064 34848
rect 18748 34783 19064 34784
rect 24682 34848 24998 34849
rect 24682 34784 24688 34848
rect 24752 34784 24768 34848
rect 24832 34784 24848 34848
rect 24912 34784 24928 34848
rect 24992 34784 24998 34848
rect 24682 34783 24998 34784
rect 0 34642 160 34672
rect 2865 34642 2931 34645
rect 0 34640 2931 34642
rect 0 34584 2870 34640
rect 2926 34584 2931 34640
rect 0 34582 2931 34584
rect 0 34552 160 34582
rect 2865 34579 2931 34582
rect 6637 34642 6703 34645
rect 11329 34642 11395 34645
rect 6637 34640 11395 34642
rect 6637 34584 6642 34640
rect 6698 34584 11334 34640
rect 11390 34584 11395 34640
rect 6637 34582 11395 34584
rect 6637 34579 6703 34582
rect 11329 34579 11395 34582
rect 16113 34642 16179 34645
rect 17861 34642 17927 34645
rect 16113 34640 17927 34642
rect 16113 34584 16118 34640
rect 16174 34584 17866 34640
rect 17922 34584 17927 34640
rect 16113 34582 17927 34584
rect 16113 34579 16179 34582
rect 17861 34579 17927 34582
rect 24209 34642 24275 34645
rect 25840 34642 26000 34672
rect 24209 34640 26000 34642
rect 24209 34584 24214 34640
rect 24270 34584 26000 34640
rect 24209 34582 26000 34584
rect 24209 34579 24275 34582
rect 25840 34552 26000 34582
rect 1209 34506 1275 34509
rect 798 34504 1275 34506
rect 798 34448 1214 34504
rect 1270 34448 1275 34504
rect 798 34446 1275 34448
rect 0 34370 160 34400
rect 798 34370 858 34446
rect 1209 34443 1275 34446
rect 6637 34506 6703 34509
rect 8845 34506 8911 34509
rect 6637 34504 8911 34506
rect 6637 34448 6642 34504
rect 6698 34448 8850 34504
rect 8906 34448 8911 34504
rect 6637 34446 8911 34448
rect 6637 34443 6703 34446
rect 8845 34443 8911 34446
rect 9489 34506 9555 34509
rect 12065 34506 12131 34509
rect 9489 34504 12131 34506
rect 9489 34448 9494 34504
rect 9550 34448 12070 34504
rect 12126 34448 12131 34504
rect 9489 34446 12131 34448
rect 9489 34443 9555 34446
rect 12065 34443 12131 34446
rect 24393 34506 24459 34509
rect 24393 34504 25146 34506
rect 24393 34448 24398 34504
rect 24454 34448 25146 34504
rect 24393 34446 25146 34448
rect 24393 34443 24459 34446
rect 0 34310 858 34370
rect 0 34280 160 34310
rect 3913 34304 4229 34305
rect 3913 34240 3919 34304
rect 3983 34240 3999 34304
rect 4063 34240 4079 34304
rect 4143 34240 4159 34304
rect 4223 34240 4229 34304
rect 3913 34239 4229 34240
rect 9847 34304 10163 34305
rect 9847 34240 9853 34304
rect 9917 34240 9933 34304
rect 9997 34240 10013 34304
rect 10077 34240 10093 34304
rect 10157 34240 10163 34304
rect 9847 34239 10163 34240
rect 15781 34304 16097 34305
rect 15781 34240 15787 34304
rect 15851 34240 15867 34304
rect 15931 34240 15947 34304
rect 16011 34240 16027 34304
rect 16091 34240 16097 34304
rect 15781 34239 16097 34240
rect 21715 34304 22031 34305
rect 21715 34240 21721 34304
rect 21785 34240 21801 34304
rect 21865 34240 21881 34304
rect 21945 34240 21961 34304
rect 22025 34240 22031 34304
rect 21715 34239 22031 34240
rect 0 34098 160 34128
rect 1393 34098 1459 34101
rect 0 34096 1459 34098
rect 0 34040 1398 34096
rect 1454 34040 1459 34096
rect 0 34038 1459 34040
rect 0 34008 160 34038
rect 1393 34035 1459 34038
rect 3233 34098 3299 34101
rect 6545 34098 6611 34101
rect 3233 34096 6611 34098
rect 3233 34040 3238 34096
rect 3294 34040 6550 34096
rect 6606 34040 6611 34096
rect 3233 34038 6611 34040
rect 25086 34098 25146 34446
rect 25840 34098 26000 34128
rect 25086 34038 26000 34098
rect 3233 34035 3299 34038
rect 6545 34035 6611 34038
rect 25840 34008 26000 34038
rect 2221 33962 2287 33965
rect 7598 33962 7604 33964
rect 2221 33960 7604 33962
rect 2221 33904 2226 33960
rect 2282 33904 7604 33960
rect 2221 33902 7604 33904
rect 2221 33899 2287 33902
rect 7598 33900 7604 33902
rect 7668 33900 7674 33964
rect 9121 33962 9187 33965
rect 10501 33962 10567 33965
rect 9121 33960 10567 33962
rect 9121 33904 9126 33960
rect 9182 33904 10506 33960
rect 10562 33904 10567 33960
rect 9121 33902 10567 33904
rect 9121 33899 9187 33902
rect 10501 33899 10567 33902
rect 14590 33900 14596 33964
rect 14660 33962 14666 33964
rect 22870 33962 22876 33964
rect 14660 33902 22876 33962
rect 14660 33900 14666 33902
rect 22870 33900 22876 33902
rect 22940 33900 22946 33964
rect 0 33826 160 33856
rect 3877 33826 3943 33829
rect 0 33824 3943 33826
rect 0 33768 3882 33824
rect 3938 33768 3943 33824
rect 0 33766 3943 33768
rect 0 33736 160 33766
rect 3877 33763 3943 33766
rect 9397 33826 9463 33829
rect 9765 33826 9831 33829
rect 9397 33824 9831 33826
rect 9397 33768 9402 33824
rect 9458 33768 9770 33824
rect 9826 33768 9831 33824
rect 9397 33766 9831 33768
rect 9397 33763 9463 33766
rect 9765 33763 9831 33766
rect 9949 33826 10015 33829
rect 10593 33826 10659 33829
rect 9949 33824 10659 33826
rect 9949 33768 9954 33824
rect 10010 33768 10598 33824
rect 10654 33768 10659 33824
rect 9949 33766 10659 33768
rect 9949 33763 10015 33766
rect 10593 33763 10659 33766
rect 6880 33760 7196 33761
rect 6880 33696 6886 33760
rect 6950 33696 6966 33760
rect 7030 33696 7046 33760
rect 7110 33696 7126 33760
rect 7190 33696 7196 33760
rect 6880 33695 7196 33696
rect 12814 33760 13130 33761
rect 12814 33696 12820 33760
rect 12884 33696 12900 33760
rect 12964 33696 12980 33760
rect 13044 33696 13060 33760
rect 13124 33696 13130 33760
rect 12814 33695 13130 33696
rect 18748 33760 19064 33761
rect 18748 33696 18754 33760
rect 18818 33696 18834 33760
rect 18898 33696 18914 33760
rect 18978 33696 18994 33760
rect 19058 33696 19064 33760
rect 18748 33695 19064 33696
rect 24682 33760 24998 33761
rect 24682 33696 24688 33760
rect 24752 33696 24768 33760
rect 24832 33696 24848 33760
rect 24912 33696 24928 33760
rect 24992 33696 24998 33760
rect 24682 33695 24998 33696
rect 1669 33690 1735 33693
rect 1894 33690 1900 33692
rect 1669 33688 1900 33690
rect 1669 33632 1674 33688
rect 1730 33632 1900 33688
rect 1669 33630 1900 33632
rect 1669 33627 1735 33630
rect 1894 33628 1900 33630
rect 1964 33628 1970 33692
rect 9765 33690 9831 33693
rect 10777 33690 10843 33693
rect 9765 33688 10843 33690
rect 9765 33632 9770 33688
rect 9826 33632 10782 33688
rect 10838 33632 10843 33688
rect 9765 33630 10843 33632
rect 9765 33627 9831 33630
rect 10777 33627 10843 33630
rect 0 33554 160 33584
rect 1577 33554 1643 33557
rect 0 33552 1643 33554
rect 0 33496 1582 33552
rect 1638 33496 1643 33552
rect 0 33494 1643 33496
rect 0 33464 160 33494
rect 1577 33491 1643 33494
rect 9213 33554 9279 33557
rect 14917 33554 14983 33557
rect 9213 33552 14983 33554
rect 9213 33496 9218 33552
rect 9274 33496 14922 33552
rect 14978 33496 14983 33552
rect 9213 33494 14983 33496
rect 9213 33491 9279 33494
rect 14917 33491 14983 33494
rect 24117 33554 24183 33557
rect 25840 33554 26000 33584
rect 24117 33552 26000 33554
rect 24117 33496 24122 33552
rect 24178 33496 26000 33552
rect 24117 33494 26000 33496
rect 24117 33491 24183 33494
rect 25840 33464 26000 33494
rect 3785 33418 3851 33421
rect 7925 33420 7991 33421
rect 7925 33418 7972 33420
rect 1902 33416 3851 33418
rect 1902 33360 3790 33416
rect 3846 33360 3851 33416
rect 1902 33358 3851 33360
rect 7880 33416 7972 33418
rect 7880 33360 7930 33416
rect 7880 33358 7972 33360
rect 0 33282 160 33312
rect 1902 33282 1962 33358
rect 3785 33355 3851 33358
rect 7925 33356 7972 33358
rect 8036 33356 8042 33420
rect 8293 33418 8359 33421
rect 9949 33418 10015 33421
rect 8293 33416 10015 33418
rect 8293 33360 8298 33416
rect 8354 33360 9954 33416
rect 10010 33360 10015 33416
rect 8293 33358 10015 33360
rect 7925 33355 7991 33356
rect 8293 33355 8359 33358
rect 9949 33355 10015 33358
rect 0 33222 1962 33282
rect 5073 33282 5139 33285
rect 9581 33282 9647 33285
rect 5073 33280 9647 33282
rect 5073 33224 5078 33280
rect 5134 33224 9586 33280
rect 9642 33224 9647 33280
rect 5073 33222 9647 33224
rect 0 33192 160 33222
rect 5073 33219 5139 33222
rect 9581 33219 9647 33222
rect 3913 33216 4229 33217
rect 3913 33152 3919 33216
rect 3983 33152 3999 33216
rect 4063 33152 4079 33216
rect 4143 33152 4159 33216
rect 4223 33152 4229 33216
rect 3913 33151 4229 33152
rect 9847 33216 10163 33217
rect 9847 33152 9853 33216
rect 9917 33152 9933 33216
rect 9997 33152 10013 33216
rect 10077 33152 10093 33216
rect 10157 33152 10163 33216
rect 9847 33151 10163 33152
rect 15781 33216 16097 33217
rect 15781 33152 15787 33216
rect 15851 33152 15867 33216
rect 15931 33152 15947 33216
rect 16011 33152 16027 33216
rect 16091 33152 16097 33216
rect 15781 33151 16097 33152
rect 21715 33216 22031 33217
rect 21715 33152 21721 33216
rect 21785 33152 21801 33216
rect 21865 33152 21881 33216
rect 21945 33152 21961 33216
rect 22025 33152 22031 33216
rect 21715 33151 22031 33152
rect 4337 33146 4403 33149
rect 4470 33146 4476 33148
rect 4337 33144 4476 33146
rect 4337 33088 4342 33144
rect 4398 33088 4476 33144
rect 4337 33086 4476 33088
rect 4337 33083 4403 33086
rect 4470 33084 4476 33086
rect 4540 33084 4546 33148
rect 21030 33084 21036 33148
rect 21100 33146 21106 33148
rect 21541 33146 21607 33149
rect 21100 33144 21607 33146
rect 21100 33088 21546 33144
rect 21602 33088 21607 33144
rect 21100 33086 21607 33088
rect 21100 33084 21106 33086
rect 21541 33083 21607 33086
rect 24393 33146 24459 33149
rect 24393 33144 25146 33146
rect 24393 33088 24398 33144
rect 24454 33088 25146 33144
rect 24393 33086 25146 33088
rect 24393 33083 24459 33086
rect 0 33010 160 33040
rect 2773 33010 2839 33013
rect 0 33008 2839 33010
rect 0 32952 2778 33008
rect 2834 32952 2839 33008
rect 0 32950 2839 32952
rect 0 32920 160 32950
rect 2773 32947 2839 32950
rect 3601 33010 3667 33013
rect 7097 33010 7163 33013
rect 7414 33010 7420 33012
rect 3601 33008 7420 33010
rect 3601 32952 3606 33008
rect 3662 32952 7102 33008
rect 7158 32952 7420 33008
rect 3601 32950 7420 32952
rect 3601 32947 3667 32950
rect 7097 32947 7163 32950
rect 7414 32948 7420 32950
rect 7484 32948 7490 33012
rect 10041 33010 10107 33013
rect 10501 33010 10567 33013
rect 10041 33008 10567 33010
rect 10041 32952 10046 33008
rect 10102 32952 10506 33008
rect 10562 32952 10567 33008
rect 10041 32950 10567 32952
rect 10041 32947 10107 32950
rect 10501 32947 10567 32950
rect 11697 33010 11763 33013
rect 17217 33010 17283 33013
rect 11697 33008 17283 33010
rect 11697 32952 11702 33008
rect 11758 32952 17222 33008
rect 17278 32952 17283 33008
rect 11697 32950 17283 32952
rect 25086 33010 25146 33086
rect 25840 33010 26000 33040
rect 25086 32950 26000 33010
rect 11697 32947 11763 32950
rect 17217 32947 17283 32950
rect 25840 32920 26000 32950
rect 2497 32874 2563 32877
rect 1304 32872 2563 32874
rect 1304 32816 2502 32872
rect 2558 32816 2563 32872
rect 1304 32814 2563 32816
rect 0 32738 160 32768
rect 1304 32738 1364 32814
rect 2497 32811 2563 32814
rect 2773 32874 2839 32877
rect 2998 32874 3004 32876
rect 2773 32872 3004 32874
rect 2773 32816 2778 32872
rect 2834 32816 3004 32872
rect 2773 32814 3004 32816
rect 2773 32811 2839 32814
rect 2998 32812 3004 32814
rect 3068 32812 3074 32876
rect 3550 32812 3556 32876
rect 3620 32874 3626 32876
rect 3969 32874 4035 32877
rect 4286 32874 4292 32876
rect 3620 32872 4292 32874
rect 3620 32816 3974 32872
rect 4030 32816 4292 32872
rect 3620 32814 4292 32816
rect 3620 32812 3626 32814
rect 0 32678 1364 32738
rect 2681 32738 2747 32741
rect 3558 32738 3618 32812
rect 3969 32811 4035 32814
rect 4286 32812 4292 32814
rect 4356 32812 4362 32876
rect 5717 32874 5783 32877
rect 6913 32874 6979 32877
rect 8661 32874 8727 32877
rect 5717 32872 8727 32874
rect 5717 32816 5722 32872
rect 5778 32816 6918 32872
rect 6974 32816 8666 32872
rect 8722 32816 8727 32872
rect 5717 32814 8727 32816
rect 5717 32811 5783 32814
rect 6913 32811 6979 32814
rect 8661 32811 8727 32814
rect 13077 32874 13143 32877
rect 18137 32874 18203 32877
rect 13077 32872 18203 32874
rect 13077 32816 13082 32872
rect 13138 32816 18142 32872
rect 18198 32816 18203 32872
rect 13077 32814 18203 32816
rect 13077 32811 13143 32814
rect 18137 32811 18203 32814
rect 2681 32736 3618 32738
rect 2681 32680 2686 32736
rect 2742 32680 3618 32736
rect 2681 32678 3618 32680
rect 0 32648 160 32678
rect 2681 32675 2747 32678
rect 6880 32672 7196 32673
rect 6880 32608 6886 32672
rect 6950 32608 6966 32672
rect 7030 32608 7046 32672
rect 7110 32608 7126 32672
rect 7190 32608 7196 32672
rect 6880 32607 7196 32608
rect 12814 32672 13130 32673
rect 12814 32608 12820 32672
rect 12884 32608 12900 32672
rect 12964 32608 12980 32672
rect 13044 32608 13060 32672
rect 13124 32608 13130 32672
rect 12814 32607 13130 32608
rect 18748 32672 19064 32673
rect 18748 32608 18754 32672
rect 18818 32608 18834 32672
rect 18898 32608 18914 32672
rect 18978 32608 18994 32672
rect 19058 32608 19064 32672
rect 18748 32607 19064 32608
rect 24682 32672 24998 32673
rect 24682 32608 24688 32672
rect 24752 32608 24768 32672
rect 24832 32608 24848 32672
rect 24912 32608 24928 32672
rect 24992 32608 24998 32672
rect 24682 32607 24998 32608
rect 2129 32602 2195 32605
rect 6729 32602 6795 32605
rect 16757 32602 16823 32605
rect 2129 32600 6795 32602
rect 2129 32544 2134 32600
rect 2190 32544 6734 32600
rect 6790 32544 6795 32600
rect 2129 32542 6795 32544
rect 2129 32539 2195 32542
rect 6729 32539 6795 32542
rect 15150 32600 16823 32602
rect 15150 32544 16762 32600
rect 16818 32544 16823 32600
rect 15150 32542 16823 32544
rect 0 32466 160 32496
rect 1301 32466 1367 32469
rect 0 32464 1367 32466
rect 0 32408 1306 32464
rect 1362 32408 1367 32464
rect 0 32406 1367 32408
rect 0 32376 160 32406
rect 1301 32403 1367 32406
rect 1669 32464 1735 32469
rect 1669 32408 1674 32464
rect 1730 32408 1735 32464
rect 1669 32403 1735 32408
rect 2865 32466 2931 32469
rect 7557 32466 7623 32469
rect 2865 32464 7623 32466
rect 2865 32408 2870 32464
rect 2926 32408 7562 32464
rect 7618 32408 7623 32464
rect 2865 32406 7623 32408
rect 2865 32403 2931 32406
rect 7557 32403 7623 32406
rect 9489 32466 9555 32469
rect 11237 32466 11303 32469
rect 9489 32464 11303 32466
rect 9489 32408 9494 32464
rect 9550 32408 11242 32464
rect 11298 32408 11303 32464
rect 9489 32406 11303 32408
rect 9489 32403 9555 32406
rect 11237 32403 11303 32406
rect 11789 32466 11855 32469
rect 15150 32466 15210 32542
rect 16757 32539 16823 32542
rect 11789 32464 15210 32466
rect 11789 32408 11794 32464
rect 11850 32408 15210 32464
rect 11789 32406 15210 32408
rect 15377 32466 15443 32469
rect 15653 32466 15719 32469
rect 17033 32466 17099 32469
rect 15377 32464 17099 32466
rect 15377 32408 15382 32464
rect 15438 32408 15658 32464
rect 15714 32408 17038 32464
rect 17094 32408 17099 32464
rect 15377 32406 17099 32408
rect 11789 32403 11855 32406
rect 15377 32403 15443 32406
rect 15653 32403 15719 32406
rect 17033 32403 17099 32406
rect 24117 32466 24183 32469
rect 25840 32466 26000 32496
rect 24117 32464 26000 32466
rect 24117 32408 24122 32464
rect 24178 32408 26000 32464
rect 24117 32406 26000 32408
rect 24117 32403 24183 32406
rect 1672 32330 1732 32403
rect 25840 32376 26000 32406
rect 4245 32330 4311 32333
rect 1672 32328 4311 32330
rect 1672 32272 4250 32328
rect 4306 32272 4311 32328
rect 1672 32270 4311 32272
rect 4245 32267 4311 32270
rect 5717 32330 5783 32333
rect 7925 32330 7991 32333
rect 5717 32328 7991 32330
rect 5717 32272 5722 32328
rect 5778 32272 7930 32328
rect 7986 32272 7991 32328
rect 5717 32270 7991 32272
rect 5717 32267 5783 32270
rect 7925 32267 7991 32270
rect 11881 32330 11947 32333
rect 19374 32330 19380 32332
rect 11881 32328 19380 32330
rect 11881 32272 11886 32328
rect 11942 32272 19380 32328
rect 11881 32270 19380 32272
rect 11881 32267 11947 32270
rect 19374 32268 19380 32270
rect 19444 32268 19450 32332
rect 0 32194 160 32224
rect 1945 32194 2011 32197
rect 0 32192 2011 32194
rect 0 32136 1950 32192
rect 2006 32136 2011 32192
rect 0 32134 2011 32136
rect 0 32104 160 32134
rect 1945 32131 2011 32134
rect 3913 32128 4229 32129
rect 3913 32064 3919 32128
rect 3983 32064 3999 32128
rect 4063 32064 4079 32128
rect 4143 32064 4159 32128
rect 4223 32064 4229 32128
rect 3913 32063 4229 32064
rect 9847 32128 10163 32129
rect 9847 32064 9853 32128
rect 9917 32064 9933 32128
rect 9997 32064 10013 32128
rect 10077 32064 10093 32128
rect 10157 32064 10163 32128
rect 9847 32063 10163 32064
rect 15781 32128 16097 32129
rect 15781 32064 15787 32128
rect 15851 32064 15867 32128
rect 15931 32064 15947 32128
rect 16011 32064 16027 32128
rect 16091 32064 16097 32128
rect 15781 32063 16097 32064
rect 21715 32128 22031 32129
rect 21715 32064 21721 32128
rect 21785 32064 21801 32128
rect 21865 32064 21881 32128
rect 21945 32064 21961 32128
rect 22025 32064 22031 32128
rect 21715 32063 22031 32064
rect 1393 32058 1459 32061
rect 798 32056 1459 32058
rect 798 32000 1398 32056
rect 1454 32000 1459 32056
rect 798 31998 1459 32000
rect 0 31922 160 31952
rect 798 31922 858 31998
rect 1393 31995 1459 31998
rect 4613 32058 4679 32061
rect 9581 32058 9647 32061
rect 15561 32060 15627 32061
rect 4613 32056 9647 32058
rect 4613 32000 4618 32056
rect 4674 32000 9586 32056
rect 9642 32000 9647 32056
rect 4613 31998 9647 32000
rect 4613 31995 4679 31998
rect 9581 31995 9647 31998
rect 12382 31996 12388 32060
rect 12452 32058 12458 32060
rect 13486 32058 13492 32060
rect 12452 31998 13492 32058
rect 12452 31996 12458 31998
rect 13486 31996 13492 31998
rect 13556 31996 13562 32060
rect 15510 32058 15516 32060
rect 15470 31998 15516 32058
rect 15580 32056 15627 32060
rect 15622 32000 15627 32056
rect 15510 31996 15516 31998
rect 15580 31996 15627 32000
rect 15561 31995 15627 31996
rect 0 31862 858 31922
rect 0 31832 160 31862
rect 4470 31860 4476 31924
rect 4540 31922 4546 31924
rect 7557 31922 7623 31925
rect 16021 31922 16087 31925
rect 23657 31922 23723 31925
rect 4540 31920 23723 31922
rect 4540 31864 7562 31920
rect 7618 31864 16026 31920
rect 16082 31864 23662 31920
rect 23718 31864 23723 31920
rect 4540 31862 23723 31864
rect 4540 31860 4546 31862
rect 7557 31859 7623 31862
rect 16021 31859 16087 31862
rect 23657 31859 23723 31862
rect 24393 31922 24459 31925
rect 25840 31922 26000 31952
rect 24393 31920 26000 31922
rect 24393 31864 24398 31920
rect 24454 31864 26000 31920
rect 24393 31862 26000 31864
rect 24393 31859 24459 31862
rect 25840 31832 26000 31862
rect 3325 31786 3391 31789
rect 3550 31786 3556 31788
rect 3325 31784 3556 31786
rect 3325 31728 3330 31784
rect 3386 31728 3556 31784
rect 3325 31726 3556 31728
rect 3325 31723 3391 31726
rect 3550 31724 3556 31726
rect 3620 31786 3626 31788
rect 6177 31786 6243 31789
rect 3620 31784 6243 31786
rect 3620 31728 6182 31784
rect 6238 31728 6243 31784
rect 3620 31726 6243 31728
rect 3620 31724 3626 31726
rect 6177 31723 6243 31726
rect 7598 31724 7604 31788
rect 7668 31786 7674 31788
rect 11237 31786 11303 31789
rect 7668 31784 11303 31786
rect 7668 31728 11242 31784
rect 11298 31728 11303 31784
rect 7668 31726 11303 31728
rect 7668 31724 7674 31726
rect 11237 31723 11303 31726
rect 11881 31786 11947 31789
rect 14181 31786 14247 31789
rect 11881 31784 14247 31786
rect 11881 31728 11886 31784
rect 11942 31728 14186 31784
rect 14242 31728 14247 31784
rect 11881 31726 14247 31728
rect 11881 31723 11947 31726
rect 14181 31723 14247 31726
rect 0 31650 160 31680
rect 2221 31650 2287 31653
rect 5717 31650 5783 31653
rect 0 31590 858 31650
rect 0 31560 160 31590
rect 798 31514 858 31590
rect 2221 31648 5783 31650
rect 2221 31592 2226 31648
rect 2282 31592 5722 31648
rect 5778 31592 5783 31648
rect 2221 31590 5783 31592
rect 2221 31587 2287 31590
rect 5717 31587 5783 31590
rect 12382 31588 12388 31652
rect 12452 31588 12458 31652
rect 13905 31650 13971 31653
rect 18321 31650 18387 31653
rect 13905 31648 18387 31650
rect 13905 31592 13910 31648
rect 13966 31592 18326 31648
rect 18382 31592 18387 31648
rect 13905 31590 18387 31592
rect 6880 31584 7196 31585
rect 6880 31520 6886 31584
rect 6950 31520 6966 31584
rect 7030 31520 7046 31584
rect 7110 31520 7126 31584
rect 7190 31520 7196 31584
rect 6880 31519 7196 31520
rect 1485 31514 1551 31517
rect 798 31512 1551 31514
rect 798 31456 1490 31512
rect 1546 31456 1551 31512
rect 798 31454 1551 31456
rect 1485 31451 1551 31454
rect 4613 31514 4679 31517
rect 5533 31514 5599 31517
rect 4613 31512 5599 31514
rect 4613 31456 4618 31512
rect 4674 31456 5538 31512
rect 5594 31456 5599 31512
rect 4613 31454 5599 31456
rect 4613 31451 4679 31454
rect 5533 31451 5599 31454
rect 7741 31514 7807 31517
rect 8845 31514 8911 31517
rect 7741 31512 8911 31514
rect 7741 31456 7746 31512
rect 7802 31456 8850 31512
rect 8906 31456 8911 31512
rect 7741 31454 8911 31456
rect 7741 31451 7807 31454
rect 8845 31451 8911 31454
rect 0 31378 160 31408
rect 2773 31378 2839 31381
rect 3877 31378 3943 31381
rect 0 31376 2839 31378
rect 0 31320 2778 31376
rect 2834 31320 2839 31376
rect 0 31318 2839 31320
rect 0 31288 160 31318
rect 2773 31315 2839 31318
rect 3374 31376 3943 31378
rect 3374 31320 3882 31376
rect 3938 31320 3943 31376
rect 3374 31318 3943 31320
rect 3049 31242 3115 31245
rect 3182 31242 3188 31244
rect 3049 31240 3188 31242
rect 3049 31184 3054 31240
rect 3110 31184 3188 31240
rect 3049 31182 3188 31184
rect 3049 31179 3115 31182
rect 3182 31180 3188 31182
rect 3252 31180 3258 31244
rect 0 31106 160 31136
rect 3374 31106 3434 31318
rect 3877 31315 3943 31318
rect 4654 31316 4660 31380
rect 4724 31378 4730 31380
rect 9029 31378 9095 31381
rect 4724 31376 9095 31378
rect 4724 31320 9034 31376
rect 9090 31320 9095 31376
rect 4724 31318 9095 31320
rect 12390 31378 12450 31588
rect 13905 31587 13971 31590
rect 18321 31587 18387 31590
rect 24209 31650 24275 31653
rect 24209 31648 24594 31650
rect 24209 31592 24214 31648
rect 24270 31592 24594 31648
rect 24209 31590 24594 31592
rect 24209 31587 24275 31590
rect 12814 31584 13130 31585
rect 12814 31520 12820 31584
rect 12884 31520 12900 31584
rect 12964 31520 12980 31584
rect 13044 31520 13060 31584
rect 13124 31520 13130 31584
rect 12814 31519 13130 31520
rect 18748 31584 19064 31585
rect 18748 31520 18754 31584
rect 18818 31520 18834 31584
rect 18898 31520 18914 31584
rect 18978 31520 18994 31584
rect 19058 31520 19064 31584
rect 18748 31519 19064 31520
rect 13486 31378 13492 31380
rect 12390 31318 13492 31378
rect 4724 31316 4730 31318
rect 9029 31315 9095 31318
rect 13486 31316 13492 31318
rect 13556 31316 13562 31380
rect 24534 31378 24594 31590
rect 24682 31584 24998 31585
rect 24682 31520 24688 31584
rect 24752 31520 24768 31584
rect 24832 31520 24848 31584
rect 24912 31520 24928 31584
rect 24992 31520 24998 31584
rect 24682 31519 24998 31520
rect 25840 31378 26000 31408
rect 24534 31318 26000 31378
rect 25840 31288 26000 31318
rect 5257 31242 5323 31245
rect 5441 31242 5507 31245
rect 8661 31242 8727 31245
rect 5257 31240 8727 31242
rect 5257 31184 5262 31240
rect 5318 31184 5446 31240
rect 5502 31184 8666 31240
rect 8722 31184 8727 31240
rect 5257 31182 8727 31184
rect 5257 31179 5323 31182
rect 5441 31179 5507 31182
rect 8661 31179 8727 31182
rect 11881 31242 11947 31245
rect 13077 31242 13143 31245
rect 11881 31240 13143 31242
rect 11881 31184 11886 31240
rect 11942 31184 13082 31240
rect 13138 31184 13143 31240
rect 11881 31182 13143 31184
rect 11881 31179 11947 31182
rect 13077 31179 13143 31182
rect 0 31046 3434 31106
rect 4613 31106 4679 31109
rect 6177 31106 6243 31109
rect 4613 31104 6243 31106
rect 4613 31048 4618 31104
rect 4674 31048 6182 31104
rect 6238 31048 6243 31104
rect 4613 31046 6243 31048
rect 0 31016 160 31046
rect 4613 31043 4679 31046
rect 6177 31043 6243 31046
rect 3913 31040 4229 31041
rect 3913 30976 3919 31040
rect 3983 30976 3999 31040
rect 4063 30976 4079 31040
rect 4143 30976 4159 31040
rect 4223 30976 4229 31040
rect 3913 30975 4229 30976
rect 9847 31040 10163 31041
rect 9847 30976 9853 31040
rect 9917 30976 9933 31040
rect 9997 30976 10013 31040
rect 10077 30976 10093 31040
rect 10157 30976 10163 31040
rect 9847 30975 10163 30976
rect 15781 31040 16097 31041
rect 15781 30976 15787 31040
rect 15851 30976 15867 31040
rect 15931 30976 15947 31040
rect 16011 30976 16027 31040
rect 16091 30976 16097 31040
rect 15781 30975 16097 30976
rect 21715 31040 22031 31041
rect 21715 30976 21721 31040
rect 21785 30976 21801 31040
rect 21865 30976 21881 31040
rect 21945 30976 21961 31040
rect 22025 30976 22031 31040
rect 21715 30975 22031 30976
rect 6085 30970 6151 30973
rect 4294 30968 6151 30970
rect 4294 30912 6090 30968
rect 6146 30912 6151 30968
rect 4294 30910 6151 30912
rect 0 30834 160 30864
rect 1117 30834 1183 30837
rect 0 30832 1183 30834
rect 0 30776 1122 30832
rect 1178 30776 1183 30832
rect 0 30774 1183 30776
rect 0 30744 160 30774
rect 1117 30771 1183 30774
rect 2221 30834 2287 30837
rect 4294 30834 4354 30910
rect 6085 30907 6151 30910
rect 2221 30832 4354 30834
rect 2221 30776 2226 30832
rect 2282 30776 4354 30832
rect 2221 30774 4354 30776
rect 4797 30834 4863 30837
rect 9029 30834 9095 30837
rect 4797 30832 9095 30834
rect 4797 30776 4802 30832
rect 4858 30776 9034 30832
rect 9090 30776 9095 30832
rect 4797 30774 9095 30776
rect 2221 30771 2287 30774
rect 4797 30771 4863 30774
rect 9029 30771 9095 30774
rect 24393 30834 24459 30837
rect 25840 30834 26000 30864
rect 24393 30832 26000 30834
rect 24393 30776 24398 30832
rect 24454 30776 26000 30832
rect 24393 30774 26000 30776
rect 24393 30771 24459 30774
rect 25840 30744 26000 30774
rect 5073 30698 5139 30701
rect 7833 30698 7899 30701
rect 5073 30696 7899 30698
rect 5073 30640 5078 30696
rect 5134 30640 7838 30696
rect 7894 30640 7899 30696
rect 5073 30638 7899 30640
rect 5073 30635 5139 30638
rect 7833 30635 7899 30638
rect 0 30562 160 30592
rect 1301 30562 1367 30565
rect 0 30560 1367 30562
rect 0 30504 1306 30560
rect 1362 30504 1367 30560
rect 0 30502 1367 30504
rect 0 30472 160 30502
rect 1301 30499 1367 30502
rect 3601 30562 3667 30565
rect 5901 30562 5967 30565
rect 3601 30560 5967 30562
rect 3601 30504 3606 30560
rect 3662 30504 5906 30560
rect 5962 30504 5967 30560
rect 3601 30502 5967 30504
rect 3601 30499 3667 30502
rect 5901 30499 5967 30502
rect 13905 30562 13971 30565
rect 14038 30562 14044 30564
rect 13905 30560 14044 30562
rect 13905 30504 13910 30560
rect 13966 30504 14044 30560
rect 13905 30502 14044 30504
rect 13905 30499 13971 30502
rect 14038 30500 14044 30502
rect 14108 30500 14114 30564
rect 6880 30496 7196 30497
rect 6880 30432 6886 30496
rect 6950 30432 6966 30496
rect 7030 30432 7046 30496
rect 7110 30432 7126 30496
rect 7190 30432 7196 30496
rect 6880 30431 7196 30432
rect 12814 30496 13130 30497
rect 12814 30432 12820 30496
rect 12884 30432 12900 30496
rect 12964 30432 12980 30496
rect 13044 30432 13060 30496
rect 13124 30432 13130 30496
rect 12814 30431 13130 30432
rect 18748 30496 19064 30497
rect 18748 30432 18754 30496
rect 18818 30432 18834 30496
rect 18898 30432 18914 30496
rect 18978 30432 18994 30496
rect 19058 30432 19064 30496
rect 18748 30431 19064 30432
rect 24682 30496 24998 30497
rect 24682 30432 24688 30496
rect 24752 30432 24768 30496
rect 24832 30432 24848 30496
rect 24912 30432 24928 30496
rect 24992 30432 24998 30496
rect 24682 30431 24998 30432
rect 2129 30426 2195 30429
rect 3233 30426 3299 30429
rect 9949 30426 10015 30429
rect 11605 30426 11671 30429
rect 12014 30426 12020 30428
rect 2129 30424 5090 30426
rect 2129 30368 2134 30424
rect 2190 30368 3238 30424
rect 3294 30368 5090 30424
rect 2129 30366 5090 30368
rect 2129 30363 2195 30366
rect 3233 30363 3299 30366
rect 0 30290 160 30320
rect 1393 30290 1459 30293
rect 1577 30290 1643 30293
rect 4797 30292 4863 30293
rect 4797 30290 4844 30292
rect 0 30288 1459 30290
rect 0 30232 1398 30288
rect 1454 30232 1459 30288
rect 0 30230 1459 30232
rect 0 30200 160 30230
rect 1393 30227 1459 30230
rect 1534 30288 1643 30290
rect 1534 30232 1582 30288
rect 1638 30232 1643 30288
rect 1534 30227 1643 30232
rect 4752 30288 4844 30290
rect 4752 30232 4802 30288
rect 4752 30230 4844 30232
rect 4797 30228 4844 30230
rect 4908 30228 4914 30292
rect 5030 30290 5090 30366
rect 9949 30424 10978 30426
rect 9949 30368 9954 30424
rect 10010 30368 10978 30424
rect 9949 30366 10978 30368
rect 9949 30363 10015 30366
rect 9029 30290 9095 30293
rect 5030 30288 9095 30290
rect 5030 30232 9034 30288
rect 9090 30232 9095 30288
rect 5030 30230 9095 30232
rect 4797 30227 4863 30228
rect 9029 30227 9095 30230
rect 9489 30290 9555 30293
rect 10041 30290 10107 30293
rect 9489 30288 10107 30290
rect 9489 30232 9494 30288
rect 9550 30232 10046 30288
rect 10102 30232 10107 30288
rect 9489 30230 10107 30232
rect 10918 30290 10978 30366
rect 11605 30424 12020 30426
rect 11605 30368 11610 30424
rect 11666 30368 12020 30424
rect 11605 30366 12020 30368
rect 11605 30363 11671 30366
rect 12014 30364 12020 30366
rect 12084 30364 12090 30428
rect 14089 30426 14155 30429
rect 14406 30426 14412 30428
rect 14089 30424 14412 30426
rect 14089 30368 14094 30424
rect 14150 30368 14412 30424
rect 14089 30366 14412 30368
rect 14089 30363 14155 30366
rect 14406 30364 14412 30366
rect 14476 30364 14482 30428
rect 20437 30426 20503 30429
rect 23013 30426 23079 30429
rect 20437 30424 23079 30426
rect 20437 30368 20442 30424
rect 20498 30368 23018 30424
rect 23074 30368 23079 30424
rect 20437 30366 23079 30368
rect 20437 30363 20503 30366
rect 23013 30363 23079 30366
rect 11605 30290 11671 30293
rect 10918 30288 11671 30290
rect 10918 30232 11610 30288
rect 11666 30232 11671 30288
rect 10918 30230 11671 30232
rect 9489 30227 9555 30230
rect 10041 30227 10107 30230
rect 11605 30227 11671 30230
rect 20989 30290 21055 30293
rect 23197 30290 23263 30293
rect 20989 30288 23263 30290
rect 20989 30232 20994 30288
rect 21050 30232 23202 30288
rect 23258 30232 23263 30288
rect 20989 30230 23263 30232
rect 20989 30227 21055 30230
rect 23197 30227 23263 30230
rect 24209 30290 24275 30293
rect 25840 30290 26000 30320
rect 24209 30288 26000 30290
rect 24209 30232 24214 30288
rect 24270 30232 26000 30288
rect 24209 30230 26000 30232
rect 24209 30227 24275 30230
rect 0 30018 160 30048
rect 1534 30018 1594 30227
rect 25840 30200 26000 30230
rect 3190 30094 5458 30154
rect 3190 30020 3250 30094
rect 5165 30020 5231 30021
rect 0 29958 1594 30018
rect 0 29928 160 29958
rect 3182 29956 3188 30020
rect 3252 29956 3258 30020
rect 5165 30016 5212 30020
rect 5276 30018 5282 30020
rect 5398 30018 5458 30094
rect 6126 30092 6132 30156
rect 6196 30154 6202 30156
rect 6269 30154 6335 30157
rect 10358 30154 10364 30156
rect 6196 30152 6335 30154
rect 6196 30096 6274 30152
rect 6330 30096 6335 30152
rect 6196 30094 6335 30096
rect 6196 30092 6202 30094
rect 6269 30091 6335 30094
rect 9630 30094 10364 30154
rect 9630 30018 9690 30094
rect 10358 30092 10364 30094
rect 10428 30154 10434 30156
rect 10428 30094 14428 30154
rect 10428 30092 10434 30094
rect 14368 30021 14428 30094
rect 10409 30020 10475 30021
rect 5165 29960 5170 30016
rect 5165 29956 5212 29960
rect 5276 29958 5322 30018
rect 5398 29958 9690 30018
rect 5276 29956 5282 29958
rect 10358 29956 10364 30020
rect 10428 30018 10475 30020
rect 10428 30016 10520 30018
rect 10470 29960 10520 30016
rect 10428 29958 10520 29960
rect 14365 30016 14431 30021
rect 14365 29960 14370 30016
rect 14426 29960 14431 30016
rect 10428 29956 10475 29958
rect 5165 29955 5231 29956
rect 10409 29955 10475 29956
rect 14365 29955 14431 29960
rect 3913 29952 4229 29953
rect 3913 29888 3919 29952
rect 3983 29888 3999 29952
rect 4063 29888 4079 29952
rect 4143 29888 4159 29952
rect 4223 29888 4229 29952
rect 3913 29887 4229 29888
rect 9847 29952 10163 29953
rect 9847 29888 9853 29952
rect 9917 29888 9933 29952
rect 9997 29888 10013 29952
rect 10077 29888 10093 29952
rect 10157 29888 10163 29952
rect 9847 29887 10163 29888
rect 15781 29952 16097 29953
rect 15781 29888 15787 29952
rect 15851 29888 15867 29952
rect 15931 29888 15947 29952
rect 16011 29888 16027 29952
rect 16091 29888 16097 29952
rect 15781 29887 16097 29888
rect 21715 29952 22031 29953
rect 21715 29888 21721 29952
rect 21785 29888 21801 29952
rect 21865 29888 21881 29952
rect 21945 29888 21961 29952
rect 22025 29888 22031 29952
rect 21715 29887 22031 29888
rect 7189 29882 7255 29885
rect 7833 29882 7899 29885
rect 7189 29880 7899 29882
rect 7189 29824 7194 29880
rect 7250 29824 7838 29880
rect 7894 29824 7899 29880
rect 7189 29822 7899 29824
rect 7189 29819 7255 29822
rect 7833 29819 7899 29822
rect 7966 29820 7972 29884
rect 8036 29882 8042 29884
rect 8109 29882 8175 29885
rect 8036 29880 8175 29882
rect 8036 29824 8114 29880
rect 8170 29824 8175 29880
rect 8036 29822 8175 29824
rect 8036 29820 8042 29822
rect 8109 29819 8175 29822
rect 0 29746 160 29776
rect 1117 29746 1183 29749
rect 0 29744 1183 29746
rect 0 29688 1122 29744
rect 1178 29688 1183 29744
rect 0 29686 1183 29688
rect 0 29656 160 29686
rect 1117 29683 1183 29686
rect 2773 29746 2839 29749
rect 11881 29746 11947 29749
rect 2773 29744 11947 29746
rect 2773 29688 2778 29744
rect 2834 29688 11886 29744
rect 11942 29688 11947 29744
rect 2773 29686 11947 29688
rect 2773 29683 2839 29686
rect 11881 29683 11947 29686
rect 24393 29746 24459 29749
rect 25840 29746 26000 29776
rect 24393 29744 26000 29746
rect 24393 29688 24398 29744
rect 24454 29688 26000 29744
rect 24393 29686 26000 29688
rect 24393 29683 24459 29686
rect 25840 29656 26000 29686
rect 2446 29548 2452 29612
rect 2516 29610 2522 29612
rect 8845 29610 8911 29613
rect 2516 29608 8911 29610
rect 2516 29552 8850 29608
rect 8906 29552 8911 29608
rect 2516 29550 8911 29552
rect 2516 29548 2522 29550
rect 8845 29547 8911 29550
rect 9213 29610 9279 29613
rect 13169 29610 13235 29613
rect 9213 29608 13235 29610
rect 9213 29552 9218 29608
rect 9274 29552 13174 29608
rect 13230 29552 13235 29608
rect 9213 29550 13235 29552
rect 9213 29547 9279 29550
rect 13169 29547 13235 29550
rect 0 29474 160 29504
rect 1301 29474 1367 29477
rect 2129 29476 2195 29477
rect 0 29472 1367 29474
rect 0 29416 1306 29472
rect 1362 29416 1367 29472
rect 0 29414 1367 29416
rect 0 29384 160 29414
rect 1301 29411 1367 29414
rect 2078 29412 2084 29476
rect 2148 29474 2195 29476
rect 4889 29474 4955 29477
rect 2148 29472 2240 29474
rect 2190 29416 2240 29472
rect 2148 29414 2240 29416
rect 3880 29472 4955 29474
rect 3880 29416 4894 29472
rect 4950 29416 4955 29472
rect 3880 29414 4955 29416
rect 2148 29412 2195 29414
rect 2129 29411 2195 29412
rect 0 29202 160 29232
rect 3880 29202 3940 29414
rect 4889 29411 4955 29414
rect 6880 29408 7196 29409
rect 6880 29344 6886 29408
rect 6950 29344 6966 29408
rect 7030 29344 7046 29408
rect 7110 29344 7126 29408
rect 7190 29344 7196 29408
rect 6880 29343 7196 29344
rect 12814 29408 13130 29409
rect 12814 29344 12820 29408
rect 12884 29344 12900 29408
rect 12964 29344 12980 29408
rect 13044 29344 13060 29408
rect 13124 29344 13130 29408
rect 12814 29343 13130 29344
rect 18748 29408 19064 29409
rect 18748 29344 18754 29408
rect 18818 29344 18834 29408
rect 18898 29344 18914 29408
rect 18978 29344 18994 29408
rect 19058 29344 19064 29408
rect 18748 29343 19064 29344
rect 24682 29408 24998 29409
rect 24682 29344 24688 29408
rect 24752 29344 24768 29408
rect 24832 29344 24848 29408
rect 24912 29344 24928 29408
rect 24992 29344 24998 29408
rect 24682 29343 24998 29344
rect 4286 29276 4292 29340
rect 4356 29338 4362 29340
rect 4889 29338 4955 29341
rect 4356 29336 4955 29338
rect 4356 29280 4894 29336
rect 4950 29280 4955 29336
rect 4356 29278 4955 29280
rect 4356 29276 4362 29278
rect 4889 29275 4955 29278
rect 0 29142 3940 29202
rect 5901 29202 5967 29205
rect 9581 29202 9647 29205
rect 5901 29200 9647 29202
rect 5901 29144 5906 29200
rect 5962 29144 9586 29200
rect 9642 29144 9647 29200
rect 5901 29142 9647 29144
rect 0 29112 160 29142
rect 5901 29139 5967 29142
rect 9581 29139 9647 29142
rect 12985 29202 13051 29205
rect 13445 29202 13511 29205
rect 12985 29200 13511 29202
rect 12985 29144 12990 29200
rect 13046 29144 13450 29200
rect 13506 29144 13511 29200
rect 12985 29142 13511 29144
rect 12985 29139 13051 29142
rect 13445 29139 13511 29142
rect 13997 29202 14063 29205
rect 14917 29202 14983 29205
rect 17861 29202 17927 29205
rect 13997 29200 17927 29202
rect 13997 29144 14002 29200
rect 14058 29144 14922 29200
rect 14978 29144 17866 29200
rect 17922 29144 17927 29200
rect 13997 29142 17927 29144
rect 13997 29139 14063 29142
rect 14917 29139 14983 29142
rect 17861 29139 17927 29142
rect 18413 29202 18479 29205
rect 21725 29202 21791 29205
rect 22461 29202 22527 29205
rect 23289 29202 23355 29205
rect 18413 29200 18706 29202
rect 18413 29144 18418 29200
rect 18474 29144 18706 29200
rect 18413 29142 18706 29144
rect 18413 29139 18479 29142
rect 18646 29069 18706 29142
rect 21725 29200 23355 29202
rect 21725 29144 21730 29200
rect 21786 29144 22466 29200
rect 22522 29144 23294 29200
rect 23350 29144 23355 29200
rect 21725 29142 23355 29144
rect 21725 29139 21791 29142
rect 22461 29139 22527 29142
rect 23289 29139 23355 29142
rect 24209 29202 24275 29205
rect 25840 29202 26000 29232
rect 24209 29200 26000 29202
rect 24209 29144 24214 29200
rect 24270 29144 26000 29200
rect 24209 29142 26000 29144
rect 24209 29139 24275 29142
rect 25840 29112 26000 29142
rect 12157 29066 12223 29069
rect 14181 29066 14247 29069
rect 12157 29064 14247 29066
rect 0 28930 160 28960
rect 3788 28950 4354 29010
rect 12157 29008 12162 29064
rect 12218 29008 14186 29064
rect 14242 29008 14247 29064
rect 12157 29006 14247 29008
rect 12157 29003 12223 29006
rect 14181 29003 14247 29006
rect 14774 29004 14780 29068
rect 14844 29066 14850 29068
rect 18454 29066 18460 29068
rect 14844 29006 18460 29066
rect 14844 29004 14850 29006
rect 18454 29004 18460 29006
rect 18524 29004 18530 29068
rect 18646 29064 18755 29069
rect 18646 29008 18694 29064
rect 18750 29008 18755 29064
rect 18646 29006 18755 29008
rect 18689 29003 18755 29006
rect 21633 29066 21699 29069
rect 24117 29066 24183 29069
rect 21633 29064 24183 29066
rect 21633 29008 21638 29064
rect 21694 29008 24122 29064
rect 24178 29008 24183 29064
rect 21633 29006 24183 29008
rect 21633 29003 21699 29006
rect 24117 29003 24183 29006
rect 1669 28930 1735 28933
rect 0 28928 1735 28930
rect 0 28872 1674 28928
rect 1730 28872 1735 28928
rect 0 28870 1735 28872
rect 0 28840 160 28870
rect 1669 28867 1735 28870
rect 2129 28930 2195 28933
rect 3788 28930 3848 28950
rect 2129 28928 3848 28930
rect 2129 28872 2134 28928
rect 2190 28872 3848 28928
rect 2129 28870 3848 28872
rect 4294 28930 4354 28950
rect 8661 28930 8727 28933
rect 4294 28928 8727 28930
rect 4294 28872 8666 28928
rect 8722 28872 8727 28928
rect 4294 28870 8727 28872
rect 2129 28867 2195 28870
rect 8661 28867 8727 28870
rect 18229 28930 18295 28933
rect 18229 28928 19258 28930
rect 18229 28872 18234 28928
rect 18290 28872 19258 28928
rect 18229 28870 19258 28872
rect 18229 28867 18295 28870
rect 3913 28864 4229 28865
rect 3913 28800 3919 28864
rect 3983 28800 3999 28864
rect 4063 28800 4079 28864
rect 4143 28800 4159 28864
rect 4223 28800 4229 28864
rect 3913 28799 4229 28800
rect 9847 28864 10163 28865
rect 9847 28800 9853 28864
rect 9917 28800 9933 28864
rect 9997 28800 10013 28864
rect 10077 28800 10093 28864
rect 10157 28800 10163 28864
rect 9847 28799 10163 28800
rect 15781 28864 16097 28865
rect 15781 28800 15787 28864
rect 15851 28800 15867 28864
rect 15931 28800 15947 28864
rect 16011 28800 16027 28864
rect 16091 28800 16097 28864
rect 15781 28799 16097 28800
rect 4889 28794 4955 28797
rect 5901 28794 5967 28797
rect 4889 28792 5967 28794
rect 4889 28736 4894 28792
rect 4950 28736 5906 28792
rect 5962 28736 5967 28792
rect 4889 28734 5967 28736
rect 4889 28731 4955 28734
rect 5901 28731 5967 28734
rect 6269 28794 6335 28797
rect 7465 28794 7531 28797
rect 9673 28796 9739 28797
rect 9622 28794 9628 28796
rect 6269 28792 7531 28794
rect 6269 28736 6274 28792
rect 6330 28736 7470 28792
rect 7526 28736 7531 28792
rect 6269 28734 7531 28736
rect 9582 28734 9628 28794
rect 9692 28792 9739 28796
rect 9734 28736 9739 28792
rect 6269 28731 6335 28734
rect 7465 28731 7531 28734
rect 9622 28732 9628 28734
rect 9692 28732 9739 28736
rect 9673 28731 9739 28732
rect 16757 28794 16823 28797
rect 18137 28794 18203 28797
rect 16757 28792 18203 28794
rect 16757 28736 16762 28792
rect 16818 28736 18142 28792
rect 18198 28736 18203 28792
rect 16757 28734 18203 28736
rect 16757 28731 16823 28734
rect 18137 28731 18203 28734
rect 0 28658 160 28688
rect 1209 28658 1275 28661
rect 15469 28658 15535 28661
rect 18597 28658 18663 28661
rect 19198 28660 19258 28870
rect 24393 28928 24459 28933
rect 24393 28872 24398 28928
rect 24454 28872 24459 28928
rect 24393 28867 24459 28872
rect 21715 28864 22031 28865
rect 21715 28800 21721 28864
rect 21785 28800 21801 28864
rect 21865 28800 21881 28864
rect 21945 28800 21961 28864
rect 22025 28800 22031 28864
rect 21715 28799 22031 28800
rect 0 28656 1275 28658
rect 0 28600 1214 28656
rect 1270 28600 1275 28656
rect 0 28598 1275 28600
rect 0 28568 160 28598
rect 1209 28595 1275 28598
rect 2730 28656 15535 28658
rect 2730 28600 15474 28656
rect 15530 28600 15535 28656
rect 2730 28598 15535 28600
rect 2078 28460 2084 28524
rect 2148 28522 2154 28524
rect 2730 28522 2790 28598
rect 15469 28595 15535 28598
rect 18094 28656 18663 28658
rect 18094 28600 18602 28656
rect 18658 28600 18663 28656
rect 18094 28598 18663 28600
rect 2148 28462 2790 28522
rect 3877 28522 3943 28525
rect 4889 28522 4955 28525
rect 3877 28520 4955 28522
rect 3877 28464 3882 28520
rect 3938 28464 4894 28520
rect 4950 28464 4955 28520
rect 3877 28462 4955 28464
rect 2148 28460 2154 28462
rect 3877 28459 3943 28462
rect 4889 28459 4955 28462
rect 5349 28522 5415 28525
rect 10593 28522 10659 28525
rect 5349 28520 10659 28522
rect 5349 28464 5354 28520
rect 5410 28464 10598 28520
rect 10654 28464 10659 28520
rect 5349 28462 10659 28464
rect 5349 28459 5415 28462
rect 10593 28459 10659 28462
rect 12525 28522 12591 28525
rect 18094 28522 18154 28598
rect 18597 28595 18663 28598
rect 19190 28596 19196 28660
rect 19260 28596 19266 28660
rect 24396 28658 24456 28867
rect 25840 28658 26000 28688
rect 24396 28598 26000 28658
rect 25840 28568 26000 28598
rect 12525 28520 18154 28522
rect 12525 28464 12530 28520
rect 12586 28464 18154 28520
rect 12525 28462 18154 28464
rect 12525 28459 12591 28462
rect 0 28386 160 28416
rect 3049 28386 3115 28389
rect 6545 28386 6611 28389
rect 0 28384 3115 28386
rect 0 28328 3054 28384
rect 3110 28328 3115 28384
rect 0 28326 3115 28328
rect 0 28296 160 28326
rect 3049 28323 3115 28326
rect 3190 28384 6611 28386
rect 3190 28328 6550 28384
rect 6606 28328 6611 28384
rect 3190 28326 6611 28328
rect 2405 28250 2471 28253
rect 3190 28250 3250 28326
rect 6545 28323 6611 28326
rect 15009 28386 15075 28389
rect 17493 28386 17559 28389
rect 18229 28386 18295 28389
rect 15009 28384 18295 28386
rect 15009 28328 15014 28384
rect 15070 28328 17498 28384
rect 17554 28328 18234 28384
rect 18290 28328 18295 28384
rect 15009 28326 18295 28328
rect 15009 28323 15075 28326
rect 17493 28323 17559 28326
rect 18229 28323 18295 28326
rect 6880 28320 7196 28321
rect 6880 28256 6886 28320
rect 6950 28256 6966 28320
rect 7030 28256 7046 28320
rect 7110 28256 7126 28320
rect 7190 28256 7196 28320
rect 6880 28255 7196 28256
rect 12814 28320 13130 28321
rect 12814 28256 12820 28320
rect 12884 28256 12900 28320
rect 12964 28256 12980 28320
rect 13044 28256 13060 28320
rect 13124 28256 13130 28320
rect 12814 28255 13130 28256
rect 18748 28320 19064 28321
rect 18748 28256 18754 28320
rect 18818 28256 18834 28320
rect 18898 28256 18914 28320
rect 18978 28256 18994 28320
rect 19058 28256 19064 28320
rect 18748 28255 19064 28256
rect 24682 28320 24998 28321
rect 24682 28256 24688 28320
rect 24752 28256 24768 28320
rect 24832 28256 24848 28320
rect 24912 28256 24928 28320
rect 24992 28256 24998 28320
rect 24682 28255 24998 28256
rect 2405 28248 3250 28250
rect 2405 28192 2410 28248
rect 2466 28192 3250 28248
rect 2405 28190 3250 28192
rect 4889 28250 4955 28253
rect 6545 28250 6611 28253
rect 4889 28248 6611 28250
rect 4889 28192 4894 28248
rect 4950 28192 6550 28248
rect 6606 28192 6611 28248
rect 4889 28190 6611 28192
rect 2405 28187 2471 28190
rect 4889 28187 4955 28190
rect 6545 28187 6611 28190
rect 19609 28250 19675 28253
rect 20529 28250 20595 28253
rect 19609 28248 20595 28250
rect 19609 28192 19614 28248
rect 19670 28192 20534 28248
rect 20590 28192 20595 28248
rect 19609 28190 20595 28192
rect 19609 28187 19675 28190
rect 20529 28187 20595 28190
rect 0 28114 160 28144
rect 749 28114 815 28117
rect 0 28112 815 28114
rect 0 28056 754 28112
rect 810 28056 815 28112
rect 0 28054 815 28056
rect 0 28024 160 28054
rect 749 28051 815 28054
rect 1393 28114 1459 28117
rect 3601 28114 3667 28117
rect 6913 28114 6979 28117
rect 1393 28112 6979 28114
rect 1393 28056 1398 28112
rect 1454 28056 3606 28112
rect 3662 28056 6918 28112
rect 6974 28056 6979 28112
rect 1393 28054 6979 28056
rect 1393 28051 1459 28054
rect 3601 28051 3667 28054
rect 6913 28051 6979 28054
rect 11053 28114 11119 28117
rect 15285 28114 15351 28117
rect 11053 28112 15351 28114
rect 11053 28056 11058 28112
rect 11114 28056 15290 28112
rect 15346 28056 15351 28112
rect 11053 28054 15351 28056
rect 11053 28051 11119 28054
rect 15285 28051 15351 28054
rect 15745 28114 15811 28117
rect 18781 28114 18847 28117
rect 15745 28112 18847 28114
rect 15745 28056 15750 28112
rect 15806 28056 18786 28112
rect 18842 28056 18847 28112
rect 15745 28054 18847 28056
rect 15745 28051 15811 28054
rect 18781 28051 18847 28054
rect 24117 28114 24183 28117
rect 25840 28114 26000 28144
rect 24117 28112 26000 28114
rect 24117 28056 24122 28112
rect 24178 28056 26000 28112
rect 24117 28054 26000 28056
rect 24117 28051 24183 28054
rect 25840 28024 26000 28054
rect 1577 27978 1643 27981
rect 1710 27978 1716 27980
rect 1577 27976 1716 27978
rect 1577 27920 1582 27976
rect 1638 27920 1716 27976
rect 1577 27918 1716 27920
rect 1577 27915 1643 27918
rect 1710 27916 1716 27918
rect 1780 27916 1786 27980
rect 4613 27978 4679 27981
rect 5165 27978 5231 27981
rect 4613 27976 5231 27978
rect 4613 27920 4618 27976
rect 4674 27920 5170 27976
rect 5226 27920 5231 27976
rect 4613 27918 5231 27920
rect 4613 27915 4679 27918
rect 5165 27915 5231 27918
rect 5901 27978 5967 27981
rect 18229 27978 18295 27981
rect 5901 27976 18295 27978
rect 5901 27920 5906 27976
rect 5962 27920 18234 27976
rect 18290 27920 18295 27976
rect 5901 27918 18295 27920
rect 5901 27915 5967 27918
rect 18229 27915 18295 27918
rect 0 27842 160 27872
rect 3785 27842 3851 27845
rect 0 27840 3851 27842
rect 0 27784 3790 27840
rect 3846 27784 3851 27840
rect 0 27782 3851 27784
rect 0 27752 160 27782
rect 3785 27779 3851 27782
rect 4613 27842 4679 27845
rect 8569 27842 8635 27845
rect 4613 27840 8635 27842
rect 4613 27784 4618 27840
rect 4674 27784 8574 27840
rect 8630 27784 8635 27840
rect 4613 27782 8635 27784
rect 4613 27779 4679 27782
rect 8569 27779 8635 27782
rect 10593 27842 10659 27845
rect 10726 27842 10732 27844
rect 10593 27840 10732 27842
rect 10593 27784 10598 27840
rect 10654 27784 10732 27840
rect 10593 27782 10732 27784
rect 10593 27779 10659 27782
rect 10726 27780 10732 27782
rect 10796 27780 10802 27844
rect 3913 27776 4229 27777
rect 3913 27712 3919 27776
rect 3983 27712 3999 27776
rect 4063 27712 4079 27776
rect 4143 27712 4159 27776
rect 4223 27712 4229 27776
rect 3913 27711 4229 27712
rect 9847 27776 10163 27777
rect 9847 27712 9853 27776
rect 9917 27712 9933 27776
rect 9997 27712 10013 27776
rect 10077 27712 10093 27776
rect 10157 27712 10163 27776
rect 9847 27711 10163 27712
rect 15781 27776 16097 27777
rect 15781 27712 15787 27776
rect 15851 27712 15867 27776
rect 15931 27712 15947 27776
rect 16011 27712 16027 27776
rect 16091 27712 16097 27776
rect 15781 27711 16097 27712
rect 21715 27776 22031 27777
rect 21715 27712 21721 27776
rect 21785 27712 21801 27776
rect 21865 27712 21881 27776
rect 21945 27712 21961 27776
rect 22025 27712 22031 27776
rect 21715 27711 22031 27712
rect 3049 27706 3115 27709
rect 1350 27646 2652 27706
rect 0 27570 160 27600
rect 1350 27570 1410 27646
rect 2592 27573 2652 27646
rect 3049 27704 3250 27706
rect 3049 27648 3054 27704
rect 3110 27648 3250 27704
rect 3049 27646 3250 27648
rect 3049 27643 3115 27646
rect 0 27510 1410 27570
rect 1488 27510 1916 27570
rect 0 27480 160 27510
rect 1209 27434 1275 27437
rect 1488 27434 1548 27510
rect 1209 27432 1548 27434
rect 1209 27376 1214 27432
rect 1270 27376 1548 27432
rect 1209 27374 1548 27376
rect 1856 27434 1916 27510
rect 2589 27568 2655 27573
rect 2589 27512 2594 27568
rect 2650 27512 2655 27568
rect 2589 27507 2655 27512
rect 2957 27434 3023 27437
rect 1856 27432 3023 27434
rect 1856 27376 2962 27432
rect 3018 27376 3023 27432
rect 1856 27374 3023 27376
rect 1209 27371 1275 27374
rect 2957 27371 3023 27374
rect 0 27298 160 27328
rect 2773 27298 2839 27301
rect 0 27296 2839 27298
rect 0 27240 2778 27296
rect 2834 27240 2839 27296
rect 0 27238 2839 27240
rect 0 27208 160 27238
rect 2773 27235 2839 27238
rect 2957 27298 3023 27301
rect 3190 27298 3250 27646
rect 5390 27644 5396 27708
rect 5460 27706 5466 27708
rect 8201 27706 8267 27709
rect 13813 27706 13879 27709
rect 14733 27706 14799 27709
rect 5460 27704 8267 27706
rect 5460 27648 8206 27704
rect 8262 27648 8267 27704
rect 5460 27646 8267 27648
rect 5460 27644 5466 27646
rect 8201 27643 8267 27646
rect 10320 27704 14799 27706
rect 10320 27648 13818 27704
rect 13874 27648 14738 27704
rect 14794 27648 14799 27704
rect 10320 27646 14799 27648
rect 3601 27570 3667 27573
rect 7373 27570 7439 27573
rect 10320 27570 10380 27646
rect 13813 27643 13879 27646
rect 14733 27643 14799 27646
rect 17769 27706 17835 27709
rect 20713 27706 20779 27709
rect 17769 27704 20779 27706
rect 17769 27648 17774 27704
rect 17830 27648 20718 27704
rect 20774 27648 20779 27704
rect 17769 27646 20779 27648
rect 17769 27643 17835 27646
rect 20713 27643 20779 27646
rect 10501 27572 10567 27573
rect 10501 27570 10548 27572
rect 3601 27568 7439 27570
rect 3601 27512 3606 27568
rect 3662 27512 7378 27568
rect 7434 27512 7439 27568
rect 3601 27510 7439 27512
rect 3601 27507 3667 27510
rect 7373 27507 7439 27510
rect 9630 27510 10380 27570
rect 10456 27568 10548 27570
rect 10456 27512 10506 27568
rect 10456 27510 10548 27512
rect 5165 27434 5231 27437
rect 5441 27434 5507 27437
rect 5165 27432 5507 27434
rect 5165 27376 5170 27432
rect 5226 27376 5446 27432
rect 5502 27376 5507 27432
rect 5165 27374 5507 27376
rect 5165 27371 5231 27374
rect 5441 27371 5507 27374
rect 5901 27434 5967 27437
rect 9630 27434 9690 27510
rect 10501 27508 10548 27510
rect 10612 27508 10618 27572
rect 24393 27570 24459 27573
rect 25840 27570 26000 27600
rect 24393 27568 26000 27570
rect 24393 27512 24398 27568
rect 24454 27512 26000 27568
rect 24393 27510 26000 27512
rect 10501 27507 10567 27508
rect 24393 27507 24459 27510
rect 25840 27480 26000 27510
rect 5901 27432 9690 27434
rect 5901 27376 5906 27432
rect 5962 27376 9690 27432
rect 5901 27374 9690 27376
rect 5901 27371 5967 27374
rect 2957 27296 3250 27298
rect 2957 27240 2962 27296
rect 3018 27240 3250 27296
rect 2957 27238 3250 27240
rect 2957 27235 3023 27238
rect 6880 27232 7196 27233
rect 6880 27168 6886 27232
rect 6950 27168 6966 27232
rect 7030 27168 7046 27232
rect 7110 27168 7126 27232
rect 7190 27168 7196 27232
rect 6880 27167 7196 27168
rect 12814 27232 13130 27233
rect 12814 27168 12820 27232
rect 12884 27168 12900 27232
rect 12964 27168 12980 27232
rect 13044 27168 13060 27232
rect 13124 27168 13130 27232
rect 12814 27167 13130 27168
rect 18748 27232 19064 27233
rect 18748 27168 18754 27232
rect 18818 27168 18834 27232
rect 18898 27168 18914 27232
rect 18978 27168 18994 27232
rect 19058 27168 19064 27232
rect 18748 27167 19064 27168
rect 24682 27232 24998 27233
rect 24682 27168 24688 27232
rect 24752 27168 24768 27232
rect 24832 27168 24848 27232
rect 24912 27168 24928 27232
rect 24992 27168 24998 27232
rect 24682 27167 24998 27168
rect 1669 27162 1735 27165
rect 2262 27162 2268 27164
rect 1669 27160 2268 27162
rect 1669 27104 1674 27160
rect 1730 27104 2268 27160
rect 1669 27102 2268 27104
rect 1669 27099 1735 27102
rect 2262 27100 2268 27102
rect 2332 27162 2338 27164
rect 5901 27162 5967 27165
rect 2332 27160 5967 27162
rect 2332 27104 5906 27160
rect 5962 27104 5967 27160
rect 2332 27102 5967 27104
rect 2332 27100 2338 27102
rect 5901 27099 5967 27102
rect 0 27026 160 27056
rect 1209 27026 1275 27029
rect 7465 27026 7531 27029
rect 12341 27026 12407 27029
rect 0 27024 1275 27026
rect 0 26968 1214 27024
rect 1270 26968 1275 27024
rect 0 26966 1275 26968
rect 0 26936 160 26966
rect 1209 26963 1275 26966
rect 1350 27024 7531 27026
rect 1350 26968 7470 27024
rect 7526 26968 7531 27024
rect 1350 26966 7531 26968
rect 473 26890 539 26893
rect 1350 26890 1410 26966
rect 7465 26963 7531 26966
rect 7744 27024 12407 27026
rect 7744 26968 12346 27024
rect 12402 26968 12407 27024
rect 7744 26966 12407 26968
rect 473 26888 1410 26890
rect 473 26832 478 26888
rect 534 26832 1410 26888
rect 473 26830 1410 26832
rect 2497 26890 2563 26893
rect 7557 26890 7623 26893
rect 2497 26888 7623 26890
rect 2497 26832 2502 26888
rect 2558 26832 7562 26888
rect 7618 26832 7623 26888
rect 2497 26830 7623 26832
rect 473 26827 539 26830
rect 2497 26827 2563 26830
rect 7557 26827 7623 26830
rect 0 26754 160 26784
rect 7744 26757 7804 26966
rect 12341 26963 12407 26966
rect 23565 27026 23631 27029
rect 25840 27026 26000 27056
rect 23565 27024 26000 27026
rect 23565 26968 23570 27024
rect 23626 26968 26000 27024
rect 23565 26966 26000 26968
rect 23565 26963 23631 26966
rect 25840 26936 26000 26966
rect 16849 26890 16915 26893
rect 17217 26890 17283 26893
rect 17401 26892 17467 26893
rect 16849 26888 17283 26890
rect 16849 26832 16854 26888
rect 16910 26832 17222 26888
rect 17278 26832 17283 26888
rect 16849 26830 17283 26832
rect 16849 26827 16915 26830
rect 17217 26827 17283 26830
rect 17350 26828 17356 26892
rect 17420 26890 17467 26892
rect 17420 26888 17512 26890
rect 17462 26832 17512 26888
rect 17420 26830 17512 26832
rect 17420 26828 17467 26830
rect 17401 26827 17467 26828
rect 1301 26754 1367 26757
rect 0 26752 1367 26754
rect 0 26696 1306 26752
rect 1362 26696 1367 26752
rect 0 26694 1367 26696
rect 0 26664 160 26694
rect 1301 26691 1367 26694
rect 2037 26754 2103 26757
rect 2865 26754 2931 26757
rect 2037 26752 2931 26754
rect 2037 26696 2042 26752
rect 2098 26696 2870 26752
rect 2926 26696 2931 26752
rect 2037 26694 2931 26696
rect 2037 26691 2103 26694
rect 2865 26691 2931 26694
rect 6913 26754 6979 26757
rect 7741 26754 7807 26757
rect 6913 26752 7807 26754
rect 6913 26696 6918 26752
rect 6974 26696 7746 26752
rect 7802 26696 7807 26752
rect 6913 26694 7807 26696
rect 6913 26691 6979 26694
rect 7741 26691 7807 26694
rect 3913 26688 4229 26689
rect 3913 26624 3919 26688
rect 3983 26624 3999 26688
rect 4063 26624 4079 26688
rect 4143 26624 4159 26688
rect 4223 26624 4229 26688
rect 3913 26623 4229 26624
rect 9847 26688 10163 26689
rect 9847 26624 9853 26688
rect 9917 26624 9933 26688
rect 9997 26624 10013 26688
rect 10077 26624 10093 26688
rect 10157 26624 10163 26688
rect 9847 26623 10163 26624
rect 15781 26688 16097 26689
rect 15781 26624 15787 26688
rect 15851 26624 15867 26688
rect 15931 26624 15947 26688
rect 16011 26624 16027 26688
rect 16091 26624 16097 26688
rect 15781 26623 16097 26624
rect 21715 26688 22031 26689
rect 21715 26624 21721 26688
rect 21785 26624 21801 26688
rect 21865 26624 21881 26688
rect 21945 26624 21961 26688
rect 22025 26624 22031 26688
rect 21715 26623 22031 26624
rect 2221 26618 2287 26621
rect 1396 26616 2287 26618
rect 1396 26560 2226 26616
rect 2282 26560 2287 26616
rect 1396 26558 2287 26560
rect 0 26482 160 26512
rect 1396 26482 1456 26558
rect 2221 26555 2287 26558
rect 6453 26618 6519 26621
rect 6678 26618 6684 26620
rect 6453 26616 6684 26618
rect 6453 26560 6458 26616
rect 6514 26560 6684 26616
rect 6453 26558 6684 26560
rect 6453 26555 6519 26558
rect 6678 26556 6684 26558
rect 6748 26556 6754 26620
rect 0 26422 1456 26482
rect 2129 26482 2195 26485
rect 6729 26482 6795 26485
rect 2129 26480 6795 26482
rect 2129 26424 2134 26480
rect 2190 26424 6734 26480
rect 6790 26424 6795 26480
rect 2129 26422 6795 26424
rect 0 26392 160 26422
rect 2129 26419 2195 26422
rect 6729 26419 6795 26422
rect 11973 26482 12039 26485
rect 12525 26482 12591 26485
rect 13670 26482 13676 26484
rect 11973 26480 13676 26482
rect 11973 26424 11978 26480
rect 12034 26424 12530 26480
rect 12586 26424 13676 26480
rect 11973 26422 13676 26424
rect 11973 26419 12039 26422
rect 12525 26419 12591 26422
rect 13670 26420 13676 26422
rect 13740 26420 13746 26484
rect 24209 26482 24275 26485
rect 25840 26482 26000 26512
rect 24209 26480 26000 26482
rect 24209 26424 24214 26480
rect 24270 26424 26000 26480
rect 24209 26422 26000 26424
rect 24209 26419 24275 26422
rect 25840 26392 26000 26422
rect 1577 26346 1643 26349
rect 15469 26346 15535 26349
rect 1577 26344 15535 26346
rect 1577 26288 1582 26344
rect 1638 26288 15474 26344
rect 15530 26288 15535 26344
rect 1577 26286 15535 26288
rect 1577 26283 1643 26286
rect 15469 26283 15535 26286
rect 0 26210 160 26240
rect 2497 26210 2563 26213
rect 0 26208 2563 26210
rect 0 26152 2502 26208
rect 2558 26152 2563 26208
rect 0 26150 2563 26152
rect 0 26120 160 26150
rect 2497 26147 2563 26150
rect 8109 26208 8175 26213
rect 8109 26152 8114 26208
rect 8170 26152 8175 26208
rect 8109 26147 8175 26152
rect 9765 26210 9831 26213
rect 10726 26210 10732 26212
rect 9765 26208 10732 26210
rect 9765 26152 9770 26208
rect 9826 26152 10732 26208
rect 9765 26150 10732 26152
rect 9765 26147 9831 26150
rect 10726 26148 10732 26150
rect 10796 26148 10802 26212
rect 14549 26210 14615 26213
rect 16389 26212 16455 26213
rect 15326 26210 15332 26212
rect 14549 26208 15332 26210
rect 14549 26152 14554 26208
rect 14610 26152 15332 26208
rect 14549 26150 15332 26152
rect 14549 26147 14615 26150
rect 15326 26148 15332 26150
rect 15396 26148 15402 26212
rect 16389 26208 16436 26212
rect 16500 26210 16506 26212
rect 16389 26152 16394 26208
rect 16389 26148 16436 26152
rect 16500 26150 16546 26210
rect 16500 26148 16506 26150
rect 19190 26148 19196 26212
rect 19260 26210 19266 26212
rect 20110 26210 20116 26212
rect 19260 26150 20116 26210
rect 19260 26148 19266 26150
rect 20110 26148 20116 26150
rect 20180 26148 20186 26212
rect 16389 26147 16455 26148
rect 6880 26144 7196 26145
rect 6880 26080 6886 26144
rect 6950 26080 6966 26144
rect 7030 26080 7046 26144
rect 7110 26080 7126 26144
rect 7190 26080 7196 26144
rect 6880 26079 7196 26080
rect 657 26074 723 26077
rect 3601 26074 3667 26077
rect 657 26072 3667 26074
rect 657 26016 662 26072
rect 718 26016 3606 26072
rect 3662 26016 3667 26072
rect 657 26014 3667 26016
rect 657 26011 723 26014
rect 3601 26011 3667 26014
rect 4153 26074 4219 26077
rect 5625 26074 5691 26077
rect 4153 26072 5691 26074
rect 4153 26016 4158 26072
rect 4214 26016 5630 26072
rect 5686 26016 5691 26072
rect 4153 26014 5691 26016
rect 4153 26011 4219 26014
rect 5625 26011 5691 26014
rect 0 25938 160 25968
rect 2129 25938 2195 25941
rect 8112 25938 8172 26147
rect 12814 26144 13130 26145
rect 12814 26080 12820 26144
rect 12884 26080 12900 26144
rect 12964 26080 12980 26144
rect 13044 26080 13060 26144
rect 13124 26080 13130 26144
rect 12814 26079 13130 26080
rect 18748 26144 19064 26145
rect 18748 26080 18754 26144
rect 18818 26080 18834 26144
rect 18898 26080 18914 26144
rect 18978 26080 18994 26144
rect 19058 26080 19064 26144
rect 18748 26079 19064 26080
rect 24682 26144 24998 26145
rect 24682 26080 24688 26144
rect 24752 26080 24768 26144
rect 24832 26080 24848 26144
rect 24912 26080 24928 26144
rect 24992 26080 24998 26144
rect 24682 26079 24998 26080
rect 0 25878 1226 25938
rect 0 25848 160 25878
rect 1166 25802 1226 25878
rect 2129 25936 8172 25938
rect 2129 25880 2134 25936
rect 2190 25880 8172 25936
rect 2129 25878 8172 25880
rect 25129 25938 25195 25941
rect 25840 25938 26000 25968
rect 25129 25936 26000 25938
rect 25129 25880 25134 25936
rect 25190 25880 26000 25936
rect 25129 25878 26000 25880
rect 2129 25875 2195 25878
rect 25129 25875 25195 25878
rect 25840 25848 26000 25878
rect 2221 25802 2287 25805
rect 1166 25800 2287 25802
rect 1166 25744 2226 25800
rect 2282 25744 2287 25800
rect 1166 25742 2287 25744
rect 2221 25739 2287 25742
rect 2405 25802 2471 25805
rect 5441 25802 5507 25805
rect 15653 25802 15719 25805
rect 2405 25800 5274 25802
rect 2405 25744 2410 25800
rect 2466 25744 5274 25800
rect 2405 25742 5274 25744
rect 2405 25739 2471 25742
rect 0 25666 160 25696
rect 1393 25666 1459 25669
rect 0 25664 1459 25666
rect 0 25608 1398 25664
rect 1454 25608 1459 25664
rect 0 25606 1459 25608
rect 5214 25666 5274 25742
rect 5441 25800 15719 25802
rect 5441 25744 5446 25800
rect 5502 25744 15658 25800
rect 15714 25744 15719 25800
rect 5441 25742 15719 25744
rect 5441 25739 5507 25742
rect 15653 25739 15719 25742
rect 7465 25666 7531 25669
rect 5214 25664 7531 25666
rect 5214 25608 7470 25664
rect 7526 25608 7531 25664
rect 5214 25606 7531 25608
rect 0 25576 160 25606
rect 1393 25603 1459 25606
rect 7465 25603 7531 25606
rect 3913 25600 4229 25601
rect 3913 25536 3919 25600
rect 3983 25536 3999 25600
rect 4063 25536 4079 25600
rect 4143 25536 4159 25600
rect 4223 25536 4229 25600
rect 3913 25535 4229 25536
rect 9847 25600 10163 25601
rect 9847 25536 9853 25600
rect 9917 25536 9933 25600
rect 9997 25536 10013 25600
rect 10077 25536 10093 25600
rect 10157 25536 10163 25600
rect 9847 25535 10163 25536
rect 15781 25600 16097 25601
rect 15781 25536 15787 25600
rect 15851 25536 15867 25600
rect 15931 25536 15947 25600
rect 16011 25536 16027 25600
rect 16091 25536 16097 25600
rect 15781 25535 16097 25536
rect 21715 25600 22031 25601
rect 21715 25536 21721 25600
rect 21785 25536 21801 25600
rect 21865 25536 21881 25600
rect 21945 25536 21961 25600
rect 22025 25536 22031 25600
rect 21715 25535 22031 25536
rect 0 25394 160 25424
rect 933 25394 999 25397
rect 0 25392 999 25394
rect 0 25336 938 25392
rect 994 25336 999 25392
rect 0 25334 999 25336
rect 0 25304 160 25334
rect 933 25331 999 25334
rect 6269 25394 6335 25397
rect 8293 25394 8359 25397
rect 6269 25392 8359 25394
rect 6269 25336 6274 25392
rect 6330 25336 8298 25392
rect 8354 25336 8359 25392
rect 6269 25334 8359 25336
rect 6269 25331 6335 25334
rect 8293 25331 8359 25334
rect 11053 25394 11119 25397
rect 14774 25394 14780 25396
rect 11053 25392 14780 25394
rect 11053 25336 11058 25392
rect 11114 25336 14780 25392
rect 11053 25334 14780 25336
rect 11053 25331 11119 25334
rect 14774 25332 14780 25334
rect 14844 25332 14850 25396
rect 24393 25394 24459 25397
rect 25840 25394 26000 25424
rect 24393 25392 26000 25394
rect 24393 25336 24398 25392
rect 24454 25336 26000 25392
rect 24393 25334 26000 25336
rect 24393 25331 24459 25334
rect 25840 25304 26000 25334
rect 2681 25258 2747 25261
rect 4838 25258 4844 25260
rect 2681 25256 4844 25258
rect 2681 25200 2686 25256
rect 2742 25200 4844 25256
rect 2681 25198 4844 25200
rect 2681 25195 2747 25198
rect 4838 25196 4844 25198
rect 4908 25258 4914 25260
rect 7557 25258 7623 25261
rect 19333 25258 19399 25261
rect 4908 25198 7436 25258
rect 4908 25196 4914 25198
rect 0 25122 160 25152
rect 841 25122 907 25125
rect 0 25120 907 25122
rect 0 25064 846 25120
rect 902 25064 907 25120
rect 0 25062 907 25064
rect 0 25032 160 25062
rect 841 25059 907 25062
rect 1577 25122 1643 25125
rect 5625 25122 5691 25125
rect 1577 25120 5691 25122
rect 1577 25064 1582 25120
rect 1638 25064 5630 25120
rect 5686 25064 5691 25120
rect 1577 25062 5691 25064
rect 7376 25122 7436 25198
rect 7557 25256 19399 25258
rect 7557 25200 7562 25256
rect 7618 25200 19338 25256
rect 19394 25200 19399 25256
rect 7557 25198 19399 25200
rect 7557 25195 7623 25198
rect 19333 25195 19399 25198
rect 7598 25122 7604 25124
rect 7376 25062 7604 25122
rect 1577 25059 1643 25062
rect 5625 25059 5691 25062
rect 7598 25060 7604 25062
rect 7668 25060 7674 25124
rect 6880 25056 7196 25057
rect 6880 24992 6886 25056
rect 6950 24992 6966 25056
rect 7030 24992 7046 25056
rect 7110 24992 7126 25056
rect 7190 24992 7196 25056
rect 6880 24991 7196 24992
rect 12814 25056 13130 25057
rect 12814 24992 12820 25056
rect 12884 24992 12900 25056
rect 12964 24992 12980 25056
rect 13044 24992 13060 25056
rect 13124 24992 13130 25056
rect 12814 24991 13130 24992
rect 18748 25056 19064 25057
rect 18748 24992 18754 25056
rect 18818 24992 18834 25056
rect 18898 24992 18914 25056
rect 18978 24992 18994 25056
rect 19058 24992 19064 25056
rect 18748 24991 19064 24992
rect 24682 25056 24998 25057
rect 24682 24992 24688 25056
rect 24752 24992 24768 25056
rect 24832 24992 24848 25056
rect 24912 24992 24928 25056
rect 24992 24992 24998 25056
rect 24682 24991 24998 24992
rect 8937 24986 9003 24989
rect 9070 24986 9076 24988
rect 8937 24984 9076 24986
rect 8937 24928 8942 24984
rect 8998 24928 9076 24984
rect 8937 24926 9076 24928
rect 8937 24923 9003 24926
rect 9070 24924 9076 24926
rect 9140 24924 9146 24988
rect 9397 24986 9463 24989
rect 10358 24986 10364 24988
rect 9397 24984 10364 24986
rect 9397 24928 9402 24984
rect 9458 24928 10364 24984
rect 9397 24926 10364 24928
rect 9397 24923 9463 24926
rect 10358 24924 10364 24926
rect 10428 24924 10434 24988
rect 0 24850 160 24880
rect 1301 24850 1367 24853
rect 0 24848 1367 24850
rect 0 24792 1306 24848
rect 1362 24792 1367 24848
rect 0 24790 1367 24792
rect 0 24760 160 24790
rect 1301 24787 1367 24790
rect 1853 24850 1919 24853
rect 2078 24850 2084 24852
rect 1853 24848 2084 24850
rect 1853 24792 1858 24848
rect 1914 24792 2084 24848
rect 1853 24790 2084 24792
rect 1853 24787 1919 24790
rect 2078 24788 2084 24790
rect 2148 24788 2154 24852
rect 2589 24850 2655 24853
rect 4654 24850 4660 24852
rect 2589 24848 4660 24850
rect 2589 24792 2594 24848
rect 2650 24792 4660 24848
rect 2589 24790 4660 24792
rect 2589 24787 2655 24790
rect 4654 24788 4660 24790
rect 4724 24788 4730 24852
rect 5901 24850 5967 24853
rect 11329 24850 11395 24853
rect 5901 24848 11395 24850
rect 5901 24792 5906 24848
rect 5962 24792 11334 24848
rect 11390 24792 11395 24848
rect 5901 24790 11395 24792
rect 5901 24787 5967 24790
rect 11329 24787 11395 24790
rect 24117 24850 24183 24853
rect 25840 24850 26000 24880
rect 24117 24848 26000 24850
rect 24117 24792 24122 24848
rect 24178 24792 26000 24848
rect 24117 24790 26000 24792
rect 24117 24787 24183 24790
rect 25840 24760 26000 24790
rect 841 24714 907 24717
rect 3049 24714 3115 24717
rect 841 24712 3115 24714
rect 841 24656 846 24712
rect 902 24656 3054 24712
rect 3110 24656 3115 24712
rect 841 24654 3115 24656
rect 841 24651 907 24654
rect 3049 24651 3115 24654
rect 4705 24714 4771 24717
rect 21357 24714 21423 24717
rect 4705 24712 21423 24714
rect 4705 24656 4710 24712
rect 4766 24656 21362 24712
rect 21418 24656 21423 24712
rect 4705 24654 21423 24656
rect 4705 24651 4771 24654
rect 21357 24651 21423 24654
rect 0 24578 160 24608
rect 1301 24578 1367 24581
rect 0 24576 1367 24578
rect 0 24520 1306 24576
rect 1362 24520 1367 24576
rect 0 24518 1367 24520
rect 0 24488 160 24518
rect 1301 24515 1367 24518
rect 10501 24578 10567 24581
rect 14181 24578 14247 24581
rect 10501 24576 14247 24578
rect 10501 24520 10506 24576
rect 10562 24520 14186 24576
rect 14242 24520 14247 24576
rect 10501 24518 14247 24520
rect 10501 24515 10567 24518
rect 14181 24515 14247 24518
rect 3913 24512 4229 24513
rect 3913 24448 3919 24512
rect 3983 24448 3999 24512
rect 4063 24448 4079 24512
rect 4143 24448 4159 24512
rect 4223 24448 4229 24512
rect 3913 24447 4229 24448
rect 9847 24512 10163 24513
rect 9847 24448 9853 24512
rect 9917 24448 9933 24512
rect 9997 24448 10013 24512
rect 10077 24448 10093 24512
rect 10157 24448 10163 24512
rect 9847 24447 10163 24448
rect 15781 24512 16097 24513
rect 15781 24448 15787 24512
rect 15851 24448 15867 24512
rect 15931 24448 15947 24512
rect 16011 24448 16027 24512
rect 16091 24448 16097 24512
rect 15781 24447 16097 24448
rect 21715 24512 22031 24513
rect 21715 24448 21721 24512
rect 21785 24448 21801 24512
rect 21865 24448 21881 24512
rect 21945 24448 21961 24512
rect 22025 24448 22031 24512
rect 21715 24447 22031 24448
rect 10501 24442 10567 24445
rect 10910 24442 10916 24444
rect 10501 24440 10916 24442
rect 10501 24384 10506 24440
rect 10562 24384 10916 24440
rect 10501 24382 10916 24384
rect 10501 24379 10567 24382
rect 10910 24380 10916 24382
rect 10980 24380 10986 24444
rect 0 24306 160 24336
rect 1945 24306 2011 24309
rect 0 24304 2011 24306
rect 0 24248 1950 24304
rect 2006 24248 2011 24304
rect 0 24246 2011 24248
rect 0 24216 160 24246
rect 1945 24243 2011 24246
rect 24393 24306 24459 24309
rect 25840 24306 26000 24336
rect 24393 24304 26000 24306
rect 24393 24248 24398 24304
rect 24454 24248 26000 24304
rect 24393 24246 26000 24248
rect 24393 24243 24459 24246
rect 25840 24216 26000 24246
rect 2773 24170 2839 24173
rect 13905 24170 13971 24173
rect 2773 24168 13971 24170
rect 2773 24112 2778 24168
rect 2834 24112 13910 24168
rect 13966 24112 13971 24168
rect 2773 24110 13971 24112
rect 2773 24107 2839 24110
rect 13905 24107 13971 24110
rect 24025 24170 24091 24173
rect 24158 24170 24164 24172
rect 24025 24168 24164 24170
rect 24025 24112 24030 24168
rect 24086 24112 24164 24168
rect 24025 24110 24164 24112
rect 24025 24107 24091 24110
rect 24158 24108 24164 24110
rect 24228 24108 24234 24172
rect 0 24034 160 24064
rect 1669 24034 1735 24037
rect 0 24032 1735 24034
rect 0 23976 1674 24032
rect 1730 23976 1735 24032
rect 0 23974 1735 23976
rect 0 23944 160 23974
rect 1669 23971 1735 23974
rect 6880 23968 7196 23969
rect 6880 23904 6886 23968
rect 6950 23904 6966 23968
rect 7030 23904 7046 23968
rect 7110 23904 7126 23968
rect 7190 23904 7196 23968
rect 6880 23903 7196 23904
rect 12814 23968 13130 23969
rect 12814 23904 12820 23968
rect 12884 23904 12900 23968
rect 12964 23904 12980 23968
rect 13044 23904 13060 23968
rect 13124 23904 13130 23968
rect 12814 23903 13130 23904
rect 18748 23968 19064 23969
rect 18748 23904 18754 23968
rect 18818 23904 18834 23968
rect 18898 23904 18914 23968
rect 18978 23904 18994 23968
rect 19058 23904 19064 23968
rect 18748 23903 19064 23904
rect 24682 23968 24998 23969
rect 24682 23904 24688 23968
rect 24752 23904 24768 23968
rect 24832 23904 24848 23968
rect 24912 23904 24928 23968
rect 24992 23904 24998 23968
rect 24682 23903 24998 23904
rect 933 23898 999 23901
rect 7557 23900 7623 23901
rect 7557 23898 7604 23900
rect 798 23896 999 23898
rect 798 23840 938 23896
rect 994 23840 999 23896
rect 798 23838 999 23840
rect 7512 23896 7604 23898
rect 7512 23840 7562 23896
rect 7512 23838 7604 23840
rect 0 23762 160 23792
rect 798 23762 858 23838
rect 933 23835 999 23838
rect 7557 23836 7604 23838
rect 7668 23836 7674 23900
rect 7557 23835 7623 23836
rect 0 23702 858 23762
rect 1669 23762 1735 23765
rect 7833 23762 7899 23765
rect 1669 23760 7899 23762
rect 1669 23704 1674 23760
rect 1730 23704 7838 23760
rect 7894 23704 7899 23760
rect 1669 23702 7899 23704
rect 0 23672 160 23702
rect 1669 23699 1735 23702
rect 7833 23699 7899 23702
rect 24117 23762 24183 23765
rect 25840 23762 26000 23792
rect 24117 23760 26000 23762
rect 24117 23704 24122 23760
rect 24178 23704 26000 23760
rect 24117 23702 26000 23704
rect 24117 23699 24183 23702
rect 25840 23672 26000 23702
rect 15285 23626 15351 23629
rect 18781 23626 18847 23629
rect 15285 23624 18847 23626
rect 15285 23568 15290 23624
rect 15346 23568 18786 23624
rect 18842 23568 18847 23624
rect 15285 23566 18847 23568
rect 15285 23563 15351 23566
rect 18781 23563 18847 23566
rect 0 23490 160 23520
rect 1301 23490 1367 23493
rect 0 23488 1367 23490
rect 0 23432 1306 23488
rect 1362 23432 1367 23488
rect 0 23430 1367 23432
rect 0 23400 160 23430
rect 1301 23427 1367 23430
rect 4654 23428 4660 23492
rect 4724 23490 4730 23492
rect 6361 23490 6427 23493
rect 4724 23488 6427 23490
rect 4724 23432 6366 23488
rect 6422 23432 6427 23488
rect 4724 23430 6427 23432
rect 4724 23428 4730 23430
rect 6361 23427 6427 23430
rect 7414 23428 7420 23492
rect 7484 23490 7490 23492
rect 9305 23490 9371 23493
rect 7484 23488 9371 23490
rect 7484 23432 9310 23488
rect 9366 23432 9371 23488
rect 7484 23430 9371 23432
rect 7484 23428 7490 23430
rect 9305 23427 9371 23430
rect 10225 23490 10291 23493
rect 12198 23490 12204 23492
rect 10225 23488 12204 23490
rect 10225 23432 10230 23488
rect 10286 23432 12204 23488
rect 10225 23430 12204 23432
rect 10225 23427 10291 23430
rect 12198 23428 12204 23430
rect 12268 23428 12274 23492
rect 14038 23490 14044 23492
rect 12390 23430 14044 23490
rect 3913 23424 4229 23425
rect 3913 23360 3919 23424
rect 3983 23360 3999 23424
rect 4063 23360 4079 23424
rect 4143 23360 4159 23424
rect 4223 23360 4229 23424
rect 3913 23359 4229 23360
rect 9847 23424 10163 23425
rect 9847 23360 9853 23424
rect 9917 23360 9933 23424
rect 9997 23360 10013 23424
rect 10077 23360 10093 23424
rect 10157 23360 10163 23424
rect 9847 23359 10163 23360
rect 5441 23356 5507 23357
rect 5390 23354 5396 23356
rect 5350 23294 5396 23354
rect 5460 23352 5507 23356
rect 5502 23296 5507 23352
rect 5390 23292 5396 23294
rect 5460 23292 5507 23296
rect 5441 23291 5507 23292
rect 7833 23354 7899 23357
rect 8661 23354 8727 23357
rect 7833 23352 8727 23354
rect 7833 23296 7838 23352
rect 7894 23296 8666 23352
rect 8722 23296 8727 23352
rect 7833 23294 8727 23296
rect 7833 23291 7899 23294
rect 8661 23291 8727 23294
rect 0 23218 160 23248
rect 3417 23218 3483 23221
rect 12390 23218 12450 23430
rect 14038 23428 14044 23430
rect 14108 23490 14114 23492
rect 15193 23490 15259 23493
rect 16665 23492 16731 23493
rect 14108 23488 15259 23490
rect 14108 23432 15198 23488
rect 15254 23432 15259 23488
rect 14108 23430 15259 23432
rect 14108 23428 14114 23430
rect 15193 23427 15259 23430
rect 16614 23428 16620 23492
rect 16684 23490 16731 23492
rect 16684 23488 16776 23490
rect 16726 23432 16776 23488
rect 16684 23430 16776 23432
rect 16684 23428 16731 23430
rect 16982 23428 16988 23492
rect 17052 23490 17058 23492
rect 18689 23490 18755 23493
rect 17052 23488 18755 23490
rect 17052 23432 18694 23488
rect 18750 23432 18755 23488
rect 17052 23430 18755 23432
rect 17052 23428 17058 23430
rect 16665 23427 16731 23428
rect 18689 23427 18755 23430
rect 22502 23428 22508 23492
rect 22572 23490 22578 23492
rect 23105 23490 23171 23493
rect 22572 23488 23171 23490
rect 22572 23432 23110 23488
rect 23166 23432 23171 23488
rect 22572 23430 23171 23432
rect 22572 23428 22578 23430
rect 23105 23427 23171 23430
rect 24393 23488 24459 23493
rect 24393 23432 24398 23488
rect 24454 23432 24459 23488
rect 24393 23427 24459 23432
rect 15781 23424 16097 23425
rect 15781 23360 15787 23424
rect 15851 23360 15867 23424
rect 15931 23360 15947 23424
rect 16011 23360 16027 23424
rect 16091 23360 16097 23424
rect 15781 23359 16097 23360
rect 21715 23424 22031 23425
rect 21715 23360 21721 23424
rect 21785 23360 21801 23424
rect 21865 23360 21881 23424
rect 21945 23360 21961 23424
rect 22025 23360 22031 23424
rect 21715 23359 22031 23360
rect 0 23216 3483 23218
rect 0 23160 3422 23216
rect 3478 23160 3483 23216
rect 0 23158 3483 23160
rect 0 23128 160 23158
rect 3417 23155 3483 23158
rect 10182 23158 12450 23218
rect 24396 23218 24456 23427
rect 25840 23218 26000 23248
rect 24396 23158 26000 23218
rect 1117 23082 1183 23085
rect 3969 23082 4035 23085
rect 10182 23082 10242 23158
rect 25840 23128 26000 23158
rect 1117 23080 4035 23082
rect 1117 23024 1122 23080
rect 1178 23024 3974 23080
rect 4030 23024 4035 23080
rect 1117 23022 4035 23024
rect 1117 23019 1183 23022
rect 3969 23019 4035 23022
rect 6686 23022 10242 23082
rect 0 22946 160 22976
rect 1301 22946 1367 22949
rect 0 22944 1367 22946
rect 0 22888 1306 22944
rect 1362 22888 1367 22944
rect 0 22886 1367 22888
rect 0 22856 160 22886
rect 1301 22883 1367 22886
rect 3785 22946 3851 22949
rect 6686 22946 6746 23022
rect 3785 22944 6746 22946
rect 3785 22888 3790 22944
rect 3846 22888 6746 22944
rect 3785 22886 6746 22888
rect 3785 22883 3851 22886
rect 6880 22880 7196 22881
rect 6880 22816 6886 22880
rect 6950 22816 6966 22880
rect 7030 22816 7046 22880
rect 7110 22816 7126 22880
rect 7190 22816 7196 22880
rect 6880 22815 7196 22816
rect 12814 22880 13130 22881
rect 12814 22816 12820 22880
rect 12884 22816 12900 22880
rect 12964 22816 12980 22880
rect 13044 22816 13060 22880
rect 13124 22816 13130 22880
rect 12814 22815 13130 22816
rect 18748 22880 19064 22881
rect 18748 22816 18754 22880
rect 18818 22816 18834 22880
rect 18898 22816 18914 22880
rect 18978 22816 18994 22880
rect 19058 22816 19064 22880
rect 18748 22815 19064 22816
rect 24682 22880 24998 22881
rect 24682 22816 24688 22880
rect 24752 22816 24768 22880
rect 24832 22816 24848 22880
rect 24912 22816 24928 22880
rect 24992 22816 24998 22880
rect 24682 22815 24998 22816
rect 657 22810 723 22813
rect 5717 22810 5783 22813
rect 657 22808 5783 22810
rect 657 22752 662 22808
rect 718 22752 5722 22808
rect 5778 22752 5783 22808
rect 657 22750 5783 22752
rect 657 22747 723 22750
rect 5717 22747 5783 22750
rect 10133 22810 10199 22813
rect 10358 22810 10364 22812
rect 10133 22808 10364 22810
rect 10133 22752 10138 22808
rect 10194 22752 10364 22808
rect 10133 22750 10364 22752
rect 10133 22747 10199 22750
rect 10358 22748 10364 22750
rect 10428 22748 10434 22812
rect 0 22674 160 22704
rect 1485 22674 1551 22677
rect 4061 22674 4127 22677
rect 11145 22674 11211 22677
rect 0 22672 1551 22674
rect 0 22616 1490 22672
rect 1546 22616 1551 22672
rect 0 22614 1551 22616
rect 0 22584 160 22614
rect 1485 22611 1551 22614
rect 3788 22672 11211 22674
rect 3788 22616 4066 22672
rect 4122 22616 11150 22672
rect 11206 22616 11211 22672
rect 3788 22614 11211 22616
rect 2773 22538 2839 22541
rect 1396 22536 2839 22538
rect 1396 22480 2778 22536
rect 2834 22480 2839 22536
rect 1396 22478 2839 22480
rect 0 22402 160 22432
rect 1396 22402 1456 22478
rect 2773 22475 2839 22478
rect 0 22342 1456 22402
rect 0 22312 160 22342
rect 1301 22266 1367 22269
rect 2681 22266 2747 22269
rect 1301 22264 2747 22266
rect 1301 22208 1306 22264
rect 1362 22208 2686 22264
rect 2742 22208 2747 22264
rect 1301 22206 2747 22208
rect 1301 22203 1367 22206
rect 2681 22203 2747 22206
rect 0 22130 160 22160
rect 1301 22130 1367 22133
rect 0 22128 1367 22130
rect 0 22072 1306 22128
rect 1362 22072 1367 22128
rect 0 22070 1367 22072
rect 0 22040 160 22070
rect 1301 22067 1367 22070
rect 2630 22068 2636 22132
rect 2700 22130 2706 22132
rect 3788 22130 3848 22614
rect 4061 22611 4127 22614
rect 11145 22611 11211 22614
rect 22686 22612 22692 22676
rect 22756 22674 22762 22676
rect 23381 22674 23447 22677
rect 22756 22672 23447 22674
rect 22756 22616 23386 22672
rect 23442 22616 23447 22672
rect 22756 22614 23447 22616
rect 22756 22612 22762 22614
rect 23381 22611 23447 22614
rect 23657 22674 23723 22677
rect 25840 22674 26000 22704
rect 23657 22672 26000 22674
rect 23657 22616 23662 22672
rect 23718 22616 26000 22672
rect 23657 22614 26000 22616
rect 23657 22611 23723 22614
rect 25840 22584 26000 22614
rect 10409 22402 10475 22405
rect 15285 22402 15351 22405
rect 10409 22400 15351 22402
rect 10409 22344 10414 22400
rect 10470 22344 15290 22400
rect 15346 22344 15351 22400
rect 10409 22342 15351 22344
rect 10409 22339 10475 22342
rect 15285 22339 15351 22342
rect 3913 22336 4229 22337
rect 3913 22272 3919 22336
rect 3983 22272 3999 22336
rect 4063 22272 4079 22336
rect 4143 22272 4159 22336
rect 4223 22272 4229 22336
rect 3913 22271 4229 22272
rect 9847 22336 10163 22337
rect 9847 22272 9853 22336
rect 9917 22272 9933 22336
rect 9997 22272 10013 22336
rect 10077 22272 10093 22336
rect 10157 22272 10163 22336
rect 9847 22271 10163 22272
rect 15781 22336 16097 22337
rect 15781 22272 15787 22336
rect 15851 22272 15867 22336
rect 15931 22272 15947 22336
rect 16011 22272 16027 22336
rect 16091 22272 16097 22336
rect 15781 22271 16097 22272
rect 21715 22336 22031 22337
rect 21715 22272 21721 22336
rect 21785 22272 21801 22336
rect 21865 22272 21881 22336
rect 21945 22272 21961 22336
rect 22025 22272 22031 22336
rect 21715 22271 22031 22272
rect 11881 22268 11947 22269
rect 11830 22266 11836 22268
rect 11790 22206 11836 22266
rect 11900 22264 11947 22268
rect 11942 22208 11947 22264
rect 11830 22204 11836 22206
rect 11900 22204 11947 22208
rect 12382 22204 12388 22268
rect 12452 22266 12458 22268
rect 13486 22266 13492 22268
rect 12452 22206 13492 22266
rect 12452 22204 12458 22206
rect 13486 22204 13492 22206
rect 13556 22204 13562 22268
rect 11881 22203 11947 22204
rect 2700 22070 3848 22130
rect 4705 22130 4771 22133
rect 5390 22130 5396 22132
rect 4705 22128 5396 22130
rect 4705 22072 4710 22128
rect 4766 22072 5396 22128
rect 4705 22070 5396 22072
rect 2700 22068 2706 22070
rect 4705 22067 4771 22070
rect 5390 22068 5396 22070
rect 5460 22068 5466 22132
rect 7373 22130 7439 22133
rect 18086 22130 18092 22132
rect 7373 22128 18092 22130
rect 7373 22072 7378 22128
rect 7434 22072 18092 22128
rect 7373 22070 18092 22072
rect 7373 22067 7439 22070
rect 18086 22068 18092 22070
rect 18156 22068 18162 22132
rect 21398 22068 21404 22132
rect 21468 22130 21474 22132
rect 22502 22130 22508 22132
rect 21468 22070 22508 22130
rect 21468 22068 21474 22070
rect 22502 22068 22508 22070
rect 22572 22068 22578 22132
rect 24393 22130 24459 22133
rect 25840 22130 26000 22160
rect 24393 22128 26000 22130
rect 24393 22072 24398 22128
rect 24454 22072 26000 22128
rect 24393 22070 26000 22072
rect 24393 22067 24459 22070
rect 25840 22040 26000 22070
rect 1669 21994 1735 21997
rect 3785 21994 3851 21997
rect 4429 21996 4495 21997
rect 4429 21994 4476 21996
rect 1669 21992 3851 21994
rect 1669 21936 1674 21992
rect 1730 21936 3790 21992
rect 3846 21936 3851 21992
rect 1669 21934 3851 21936
rect 4384 21992 4476 21994
rect 4384 21936 4434 21992
rect 4384 21934 4476 21936
rect 1669 21931 1735 21934
rect 3785 21931 3851 21934
rect 4429 21932 4476 21934
rect 4540 21932 4546 21996
rect 8569 21994 8635 21997
rect 4616 21992 8635 21994
rect 4616 21936 8574 21992
rect 8630 21936 8635 21992
rect 4616 21934 8635 21936
rect 4429 21931 4495 21932
rect 0 21858 160 21888
rect 841 21858 907 21861
rect 0 21856 907 21858
rect 0 21800 846 21856
rect 902 21800 907 21856
rect 0 21798 907 21800
rect 0 21768 160 21798
rect 841 21795 907 21798
rect 2773 21858 2839 21861
rect 3233 21858 3299 21861
rect 4616 21858 4676 21934
rect 8569 21931 8635 21934
rect 12341 21994 12407 21997
rect 13486 21994 13492 21996
rect 12341 21992 13492 21994
rect 12341 21936 12346 21992
rect 12402 21936 13492 21992
rect 12341 21934 13492 21936
rect 12341 21931 12407 21934
rect 13486 21932 13492 21934
rect 13556 21994 13562 21996
rect 17217 21994 17283 21997
rect 20805 21994 20871 21997
rect 13556 21992 20871 21994
rect 13556 21936 17222 21992
rect 17278 21936 20810 21992
rect 20866 21936 20871 21992
rect 13556 21934 20871 21936
rect 13556 21932 13562 21934
rect 17217 21931 17283 21934
rect 20805 21931 20871 21934
rect 2773 21856 4676 21858
rect 2773 21800 2778 21856
rect 2834 21800 3238 21856
rect 3294 21800 4676 21856
rect 2773 21798 4676 21800
rect 2773 21795 2839 21798
rect 3233 21795 3299 21798
rect 6880 21792 7196 21793
rect 6880 21728 6886 21792
rect 6950 21728 6966 21792
rect 7030 21728 7046 21792
rect 7110 21728 7126 21792
rect 7190 21728 7196 21792
rect 6880 21727 7196 21728
rect 12814 21792 13130 21793
rect 12814 21728 12820 21792
rect 12884 21728 12900 21792
rect 12964 21728 12980 21792
rect 13044 21728 13060 21792
rect 13124 21728 13130 21792
rect 12814 21727 13130 21728
rect 18748 21792 19064 21793
rect 18748 21728 18754 21792
rect 18818 21728 18834 21792
rect 18898 21728 18914 21792
rect 18978 21728 18994 21792
rect 19058 21728 19064 21792
rect 18748 21727 19064 21728
rect 24682 21792 24998 21793
rect 24682 21728 24688 21792
rect 24752 21728 24768 21792
rect 24832 21728 24848 21792
rect 24912 21728 24928 21792
rect 24992 21728 24998 21792
rect 24682 21727 24998 21728
rect 13261 21722 13327 21725
rect 15101 21722 15167 21725
rect 15377 21722 15443 21725
rect 13261 21720 15443 21722
rect 13261 21664 13266 21720
rect 13322 21664 15106 21720
rect 15162 21664 15382 21720
rect 15438 21664 15443 21720
rect 13261 21662 15443 21664
rect 13261 21659 13327 21662
rect 15101 21659 15167 21662
rect 15377 21659 15443 21662
rect 0 21586 160 21616
rect 1025 21586 1091 21589
rect 0 21584 1091 21586
rect 0 21528 1030 21584
rect 1086 21528 1091 21584
rect 0 21526 1091 21528
rect 0 21496 160 21526
rect 1025 21523 1091 21526
rect 6453 21586 6519 21589
rect 8385 21586 8451 21589
rect 9070 21586 9076 21588
rect 6453 21584 9076 21586
rect 6453 21528 6458 21584
rect 6514 21528 8390 21584
rect 8446 21528 9076 21584
rect 6453 21526 9076 21528
rect 6453 21523 6519 21526
rect 8385 21523 8451 21526
rect 9070 21524 9076 21526
rect 9140 21586 9146 21588
rect 21030 21586 21036 21588
rect 9140 21526 21036 21586
rect 9140 21524 9146 21526
rect 21030 21524 21036 21526
rect 21100 21586 21106 21588
rect 23013 21586 23079 21589
rect 21100 21584 23079 21586
rect 21100 21528 23018 21584
rect 23074 21528 23079 21584
rect 21100 21526 23079 21528
rect 21100 21524 21106 21526
rect 23013 21523 23079 21526
rect 24117 21586 24183 21589
rect 25840 21586 26000 21616
rect 24117 21584 26000 21586
rect 24117 21528 24122 21584
rect 24178 21528 26000 21584
rect 24117 21526 26000 21528
rect 24117 21523 24183 21526
rect 25840 21496 26000 21526
rect 2129 21450 2195 21453
rect 2129 21448 5090 21450
rect 2129 21392 2134 21448
rect 2190 21392 5090 21448
rect 2129 21390 5090 21392
rect 2129 21387 2195 21390
rect 0 21314 160 21344
rect 933 21314 999 21317
rect 0 21312 999 21314
rect 0 21256 938 21312
rect 994 21256 999 21312
rect 0 21254 999 21256
rect 5030 21314 5090 21390
rect 6678 21388 6684 21452
rect 6748 21450 6754 21452
rect 7189 21450 7255 21453
rect 6748 21448 7255 21450
rect 6748 21392 7194 21448
rect 7250 21392 7255 21448
rect 6748 21390 7255 21392
rect 6748 21388 6754 21390
rect 7189 21387 7255 21390
rect 7373 21450 7439 21453
rect 9305 21450 9371 21453
rect 7373 21448 9371 21450
rect 7373 21392 7378 21448
rect 7434 21392 9310 21448
rect 9366 21392 9371 21448
rect 7373 21390 9371 21392
rect 7373 21387 7439 21390
rect 9305 21387 9371 21390
rect 11237 21450 11303 21453
rect 16113 21450 16179 21453
rect 11237 21448 16179 21450
rect 11237 21392 11242 21448
rect 11298 21392 16118 21448
rect 16174 21392 16179 21448
rect 11237 21390 16179 21392
rect 11237 21387 11303 21390
rect 16113 21387 16179 21390
rect 7557 21314 7623 21317
rect 5030 21312 7623 21314
rect 5030 21256 7562 21312
rect 7618 21256 7623 21312
rect 5030 21254 7623 21256
rect 0 21224 160 21254
rect 933 21251 999 21254
rect 7557 21251 7623 21254
rect 12198 21252 12204 21316
rect 12268 21252 12274 21316
rect 14590 21252 14596 21316
rect 14660 21314 14666 21316
rect 14917 21314 14983 21317
rect 14660 21312 14983 21314
rect 14660 21256 14922 21312
rect 14978 21256 14983 21312
rect 14660 21254 14983 21256
rect 14660 21252 14666 21254
rect 3913 21248 4229 21249
rect 3913 21184 3919 21248
rect 3983 21184 3999 21248
rect 4063 21184 4079 21248
rect 4143 21184 4159 21248
rect 4223 21184 4229 21248
rect 3913 21183 4229 21184
rect 9847 21248 10163 21249
rect 9847 21184 9853 21248
rect 9917 21184 9933 21248
rect 9997 21184 10013 21248
rect 10077 21184 10093 21248
rect 10157 21184 10163 21248
rect 9847 21183 10163 21184
rect 5901 21178 5967 21181
rect 9305 21178 9371 21181
rect 5901 21176 9371 21178
rect 5901 21120 5906 21176
rect 5962 21120 9310 21176
rect 9366 21120 9371 21176
rect 5901 21118 9371 21120
rect 5901 21115 5967 21118
rect 9305 21115 9371 21118
rect 0 21042 160 21072
rect 1577 21042 1643 21045
rect 12206 21042 12266 21252
rect 14917 21251 14983 21254
rect 15781 21248 16097 21249
rect 15781 21184 15787 21248
rect 15851 21184 15867 21248
rect 15931 21184 15947 21248
rect 16011 21184 16027 21248
rect 16091 21184 16097 21248
rect 15781 21183 16097 21184
rect 21715 21248 22031 21249
rect 21715 21184 21721 21248
rect 21785 21184 21801 21248
rect 21865 21184 21881 21248
rect 21945 21184 21961 21248
rect 22025 21184 22031 21248
rect 21715 21183 22031 21184
rect 24158 21116 24164 21180
rect 24228 21178 24234 21180
rect 24301 21178 24367 21181
rect 24228 21176 24367 21178
rect 24228 21120 24306 21176
rect 24362 21120 24367 21176
rect 24228 21118 24367 21120
rect 24228 21116 24234 21118
rect 24301 21115 24367 21118
rect 0 21040 1643 21042
rect 0 20984 1582 21040
rect 1638 20984 1643 21040
rect 0 20982 1643 20984
rect 0 20952 160 20982
rect 1577 20979 1643 20982
rect 1902 20982 12266 21042
rect 12525 21042 12591 21045
rect 16389 21042 16455 21045
rect 18965 21042 19031 21045
rect 12525 21040 19031 21042
rect 12525 20984 12530 21040
rect 12586 20984 16394 21040
rect 16450 20984 18970 21040
rect 19026 20984 19031 21040
rect 12525 20982 19031 20984
rect 1342 20844 1348 20908
rect 1412 20906 1418 20908
rect 1902 20906 1962 20982
rect 12525 20979 12591 20982
rect 16389 20979 16455 20982
rect 18965 20979 19031 20982
rect 24393 21042 24459 21045
rect 25840 21042 26000 21072
rect 24393 21040 26000 21042
rect 24393 20984 24398 21040
rect 24454 20984 26000 21040
rect 24393 20982 26000 20984
rect 24393 20979 24459 20982
rect 25840 20952 26000 20982
rect 1412 20846 1962 20906
rect 2129 20906 2195 20909
rect 8201 20906 8267 20909
rect 2129 20904 8267 20906
rect 2129 20848 2134 20904
rect 2190 20848 8206 20904
rect 8262 20848 8267 20904
rect 2129 20846 8267 20848
rect 1412 20844 1418 20846
rect 2129 20843 2195 20846
rect 8201 20843 8267 20846
rect 8385 20906 8451 20909
rect 12566 20906 12572 20908
rect 8385 20904 12572 20906
rect 8385 20848 8390 20904
rect 8446 20848 12572 20904
rect 8385 20846 12572 20848
rect 8385 20843 8451 20846
rect 12566 20844 12572 20846
rect 12636 20844 12642 20908
rect 16113 20906 16179 20909
rect 16614 20906 16620 20908
rect 16113 20904 16620 20906
rect 16113 20848 16118 20904
rect 16174 20848 16620 20904
rect 16113 20846 16620 20848
rect 16113 20843 16179 20846
rect 16614 20844 16620 20846
rect 16684 20844 16690 20908
rect 18229 20906 18295 20909
rect 19057 20906 19123 20909
rect 18229 20904 19123 20906
rect 18229 20848 18234 20904
rect 18290 20848 19062 20904
rect 19118 20848 19123 20904
rect 18229 20846 19123 20848
rect 18229 20843 18295 20846
rect 19057 20843 19123 20846
rect 0 20770 160 20800
rect 1393 20770 1459 20773
rect 0 20768 1459 20770
rect 0 20712 1398 20768
rect 1454 20712 1459 20768
rect 0 20710 1459 20712
rect 0 20680 160 20710
rect 1393 20707 1459 20710
rect 15469 20770 15535 20773
rect 17217 20770 17283 20773
rect 15469 20768 17283 20770
rect 15469 20712 15474 20768
rect 15530 20712 17222 20768
rect 17278 20712 17283 20768
rect 15469 20710 17283 20712
rect 15469 20707 15535 20710
rect 17217 20707 17283 20710
rect 6880 20704 7196 20705
rect 6880 20640 6886 20704
rect 6950 20640 6966 20704
rect 7030 20640 7046 20704
rect 7110 20640 7126 20704
rect 7190 20640 7196 20704
rect 6880 20639 7196 20640
rect 12814 20704 13130 20705
rect 12814 20640 12820 20704
rect 12884 20640 12900 20704
rect 12964 20640 12980 20704
rect 13044 20640 13060 20704
rect 13124 20640 13130 20704
rect 12814 20639 13130 20640
rect 18748 20704 19064 20705
rect 18748 20640 18754 20704
rect 18818 20640 18834 20704
rect 18898 20640 18914 20704
rect 18978 20640 18994 20704
rect 19058 20640 19064 20704
rect 18748 20639 19064 20640
rect 24682 20704 24998 20705
rect 24682 20640 24688 20704
rect 24752 20640 24768 20704
rect 24832 20640 24848 20704
rect 24912 20640 24928 20704
rect 24992 20640 24998 20704
rect 24682 20639 24998 20640
rect 1485 20634 1551 20637
rect 798 20632 1551 20634
rect 798 20576 1490 20632
rect 1546 20576 1551 20632
rect 798 20574 1551 20576
rect 0 20498 160 20528
rect 798 20498 858 20574
rect 1485 20571 1551 20574
rect 23933 20634 23999 20637
rect 23933 20632 24594 20634
rect 23933 20576 23938 20632
rect 23994 20576 24594 20632
rect 23933 20574 24594 20576
rect 23933 20571 23999 20574
rect 0 20438 858 20498
rect 3785 20498 3851 20501
rect 8937 20498 9003 20501
rect 3785 20496 9003 20498
rect 3785 20440 3790 20496
rect 3846 20440 8942 20496
rect 8998 20440 9003 20496
rect 3785 20438 9003 20440
rect 0 20408 160 20438
rect 3785 20435 3851 20438
rect 8937 20435 9003 20438
rect 12893 20498 12959 20501
rect 16430 20498 16436 20500
rect 12893 20496 16436 20498
rect 12893 20440 12898 20496
rect 12954 20440 16436 20496
rect 12893 20438 16436 20440
rect 12893 20435 12959 20438
rect 16430 20436 16436 20438
rect 16500 20436 16506 20500
rect 17350 20436 17356 20500
rect 17420 20498 17426 20500
rect 17493 20498 17559 20501
rect 17420 20496 17559 20498
rect 17420 20440 17498 20496
rect 17554 20440 17559 20496
rect 17420 20438 17559 20440
rect 24534 20498 24594 20574
rect 25840 20498 26000 20528
rect 24534 20438 26000 20498
rect 17420 20436 17426 20438
rect 17493 20435 17559 20438
rect 25840 20408 26000 20438
rect 2221 20362 2287 20365
rect 3417 20362 3483 20365
rect 4245 20362 4311 20365
rect 2221 20360 2790 20362
rect 2221 20304 2226 20360
rect 2282 20304 2790 20360
rect 2221 20302 2790 20304
rect 2221 20299 2287 20302
rect 0 20226 160 20256
rect 1209 20226 1275 20229
rect 0 20224 1275 20226
rect 0 20168 1214 20224
rect 1270 20168 1275 20224
rect 0 20166 1275 20168
rect 0 20136 160 20166
rect 1209 20163 1275 20166
rect 0 19954 160 19984
rect 1301 19954 1367 19957
rect 0 19952 1367 19954
rect 0 19896 1306 19952
rect 1362 19896 1367 19952
rect 0 19894 1367 19896
rect 2730 19954 2790 20302
rect 3417 20360 4311 20362
rect 3417 20304 3422 20360
rect 3478 20304 4250 20360
rect 4306 20304 4311 20360
rect 3417 20302 4311 20304
rect 3417 20299 3483 20302
rect 4245 20299 4311 20302
rect 10409 20362 10475 20365
rect 10685 20362 10751 20365
rect 10409 20360 10751 20362
rect 10409 20304 10414 20360
rect 10470 20304 10690 20360
rect 10746 20304 10751 20360
rect 10409 20302 10751 20304
rect 10409 20299 10475 20302
rect 10685 20299 10751 20302
rect 11053 20362 11119 20365
rect 17677 20362 17743 20365
rect 11053 20360 17743 20362
rect 11053 20304 11058 20360
rect 11114 20304 17682 20360
rect 17738 20304 17743 20360
rect 11053 20302 17743 20304
rect 11053 20299 11119 20302
rect 17677 20299 17743 20302
rect 22870 20164 22876 20228
rect 22940 20226 22946 20228
rect 25773 20226 25839 20229
rect 22940 20224 25839 20226
rect 22940 20168 25778 20224
rect 25834 20168 25839 20224
rect 22940 20166 25839 20168
rect 22940 20164 22946 20166
rect 25773 20163 25839 20166
rect 3913 20160 4229 20161
rect 3913 20096 3919 20160
rect 3983 20096 3999 20160
rect 4063 20096 4079 20160
rect 4143 20096 4159 20160
rect 4223 20096 4229 20160
rect 3913 20095 4229 20096
rect 9847 20160 10163 20161
rect 9847 20096 9853 20160
rect 9917 20096 9933 20160
rect 9997 20096 10013 20160
rect 10077 20096 10093 20160
rect 10157 20096 10163 20160
rect 9847 20095 10163 20096
rect 15781 20160 16097 20161
rect 15781 20096 15787 20160
rect 15851 20096 15867 20160
rect 15931 20096 15947 20160
rect 16011 20096 16027 20160
rect 16091 20096 16097 20160
rect 15781 20095 16097 20096
rect 21715 20160 22031 20161
rect 21715 20096 21721 20160
rect 21785 20096 21801 20160
rect 21865 20096 21881 20160
rect 21945 20096 21961 20160
rect 22025 20096 22031 20160
rect 21715 20095 22031 20096
rect 4981 20090 5047 20093
rect 9029 20090 9095 20093
rect 4981 20088 9095 20090
rect 4981 20032 4986 20088
rect 5042 20032 9034 20088
rect 9090 20032 9095 20088
rect 4981 20030 9095 20032
rect 4981 20027 5047 20030
rect 9029 20027 9095 20030
rect 4429 19954 4495 19957
rect 2730 19952 4495 19954
rect 2730 19896 4434 19952
rect 4490 19896 4495 19952
rect 2730 19894 4495 19896
rect 0 19864 160 19894
rect 1301 19891 1367 19894
rect 4429 19891 4495 19894
rect 5206 19892 5212 19956
rect 5276 19954 5282 19956
rect 9949 19954 10015 19957
rect 14917 19954 14983 19957
rect 5276 19952 10015 19954
rect 5276 19896 9954 19952
rect 10010 19896 10015 19952
rect 5276 19894 10015 19896
rect 5276 19892 5282 19894
rect 9949 19891 10015 19894
rect 10366 19952 14983 19954
rect 10366 19896 14922 19952
rect 14978 19896 14983 19952
rect 10366 19894 14983 19896
rect 10366 19821 10426 19894
rect 14917 19891 14983 19894
rect 23749 19954 23815 19957
rect 25840 19954 26000 19984
rect 23749 19952 26000 19954
rect 23749 19896 23754 19952
rect 23810 19896 26000 19952
rect 23749 19894 26000 19896
rect 23749 19891 23815 19894
rect 25840 19864 26000 19894
rect 473 19818 539 19821
rect 6085 19818 6151 19821
rect 10317 19820 10426 19821
rect 473 19816 6151 19818
rect 473 19760 478 19816
rect 534 19760 6090 19816
rect 6146 19760 6151 19816
rect 473 19758 6151 19760
rect 473 19755 539 19758
rect 6085 19755 6151 19758
rect 6732 19758 9506 19818
rect 0 19682 160 19712
rect 3325 19682 3391 19685
rect 0 19680 3391 19682
rect 0 19624 3330 19680
rect 3386 19624 3391 19680
rect 0 19622 3391 19624
rect 0 19592 160 19622
rect 3325 19619 3391 19622
rect 3509 19684 3575 19685
rect 6085 19684 6151 19685
rect 3509 19680 3556 19684
rect 3620 19682 3626 19684
rect 6085 19682 6132 19684
rect 3509 19624 3514 19680
rect 3509 19620 3556 19624
rect 3620 19622 3666 19682
rect 6040 19680 6132 19682
rect 6196 19682 6202 19684
rect 6732 19682 6792 19758
rect 6040 19624 6090 19680
rect 6040 19622 6132 19624
rect 3620 19620 3626 19622
rect 6085 19620 6132 19622
rect 6196 19622 6792 19682
rect 9446 19685 9506 19758
rect 10317 19816 10364 19820
rect 10428 19818 10434 19820
rect 11605 19818 11671 19821
rect 16573 19818 16639 19821
rect 10317 19760 10322 19816
rect 10317 19756 10364 19760
rect 10428 19758 10474 19818
rect 11605 19816 16639 19818
rect 11605 19760 11610 19816
rect 11666 19760 16578 19816
rect 16634 19760 16639 19816
rect 11605 19758 16639 19760
rect 10428 19756 10434 19758
rect 10317 19755 10383 19756
rect 11605 19755 11671 19758
rect 16573 19755 16639 19758
rect 9446 19680 9555 19685
rect 9446 19624 9494 19680
rect 9550 19624 9555 19680
rect 9446 19622 9555 19624
rect 6196 19620 6202 19622
rect 3509 19619 3575 19620
rect 6085 19619 6151 19620
rect 9489 19619 9555 19622
rect 10910 19620 10916 19684
rect 10980 19682 10986 19684
rect 11973 19682 12039 19685
rect 10980 19680 12039 19682
rect 10980 19624 11978 19680
rect 12034 19624 12039 19680
rect 10980 19622 12039 19624
rect 10980 19620 10986 19622
rect 11973 19619 12039 19622
rect 6880 19616 7196 19617
rect 6880 19552 6886 19616
rect 6950 19552 6966 19616
rect 7030 19552 7046 19616
rect 7110 19552 7126 19616
rect 7190 19552 7196 19616
rect 6880 19551 7196 19552
rect 12814 19616 13130 19617
rect 12814 19552 12820 19616
rect 12884 19552 12900 19616
rect 12964 19552 12980 19616
rect 13044 19552 13060 19616
rect 13124 19552 13130 19616
rect 12814 19551 13130 19552
rect 18748 19616 19064 19617
rect 18748 19552 18754 19616
rect 18818 19552 18834 19616
rect 18898 19552 18914 19616
rect 18978 19552 18994 19616
rect 19058 19552 19064 19616
rect 18748 19551 19064 19552
rect 24682 19616 24998 19617
rect 24682 19552 24688 19616
rect 24752 19552 24768 19616
rect 24832 19552 24848 19616
rect 24912 19552 24928 19616
rect 24992 19552 24998 19616
rect 24682 19551 24998 19552
rect 933 19546 999 19549
rect 4245 19546 4311 19549
rect 5625 19546 5691 19549
rect 13721 19548 13787 19549
rect 13670 19546 13676 19548
rect 933 19544 4311 19546
rect 933 19488 938 19544
rect 994 19488 4250 19544
rect 4306 19488 4311 19544
rect 933 19486 4311 19488
rect 933 19483 999 19486
rect 4245 19483 4311 19486
rect 4478 19544 5691 19546
rect 4478 19488 5630 19544
rect 5686 19488 5691 19544
rect 4478 19486 5691 19488
rect 13594 19486 13676 19546
rect 13740 19546 13787 19548
rect 17585 19546 17651 19549
rect 13740 19544 17651 19546
rect 13782 19488 17590 19544
rect 17646 19488 17651 19544
rect 0 19410 160 19440
rect 1301 19410 1367 19413
rect 0 19408 1367 19410
rect 0 19352 1306 19408
rect 1362 19352 1367 19408
rect 0 19350 1367 19352
rect 0 19320 160 19350
rect 1301 19347 1367 19350
rect 1577 19410 1643 19413
rect 2589 19410 2655 19413
rect 1577 19408 2655 19410
rect 1577 19352 1582 19408
rect 1638 19352 2594 19408
rect 2650 19352 2655 19408
rect 1577 19350 2655 19352
rect 1577 19347 1643 19350
rect 2589 19347 2655 19350
rect 3049 19410 3115 19413
rect 3601 19410 3667 19413
rect 4478 19410 4538 19486
rect 5625 19483 5691 19486
rect 13670 19484 13676 19486
rect 13740 19486 17651 19488
rect 13740 19484 13787 19486
rect 13721 19483 13787 19484
rect 17585 19483 17651 19486
rect 3049 19408 4538 19410
rect 3049 19352 3054 19408
rect 3110 19352 3606 19408
rect 3662 19352 4538 19408
rect 3049 19350 4538 19352
rect 3049 19347 3115 19350
rect 3601 19347 3667 19350
rect 5206 19348 5212 19412
rect 5276 19410 5282 19412
rect 5349 19410 5415 19413
rect 5276 19408 5415 19410
rect 5276 19352 5354 19408
rect 5410 19352 5415 19408
rect 5276 19350 5415 19352
rect 5276 19348 5282 19350
rect 5349 19347 5415 19350
rect 7189 19410 7255 19413
rect 8845 19410 8911 19413
rect 7189 19408 8911 19410
rect 7189 19352 7194 19408
rect 7250 19352 8850 19408
rect 8906 19352 8911 19408
rect 7189 19350 8911 19352
rect 7189 19347 7255 19350
rect 8845 19347 8911 19350
rect 13854 19348 13860 19412
rect 13924 19410 13930 19412
rect 14457 19410 14523 19413
rect 13924 19408 14523 19410
rect 13924 19352 14462 19408
rect 14518 19352 14523 19408
rect 13924 19350 14523 19352
rect 13924 19348 13930 19350
rect 14457 19347 14523 19350
rect 24209 19410 24275 19413
rect 25840 19410 26000 19440
rect 24209 19408 26000 19410
rect 24209 19352 24214 19408
rect 24270 19352 26000 19408
rect 24209 19350 26000 19352
rect 24209 19347 24275 19350
rect 25840 19320 26000 19350
rect 3509 19274 3575 19277
rect 3509 19272 4354 19274
rect 3509 19216 3514 19272
rect 3570 19216 4354 19272
rect 3509 19214 4354 19216
rect 3509 19211 3575 19214
rect 0 19138 160 19168
rect 749 19138 815 19141
rect 0 19136 815 19138
rect 0 19080 754 19136
rect 810 19080 815 19136
rect 0 19078 815 19080
rect 0 19048 160 19078
rect 749 19075 815 19078
rect 3913 19072 4229 19073
rect 3913 19008 3919 19072
rect 3983 19008 3999 19072
rect 4063 19008 4079 19072
rect 4143 19008 4159 19072
rect 4223 19008 4229 19072
rect 3913 19007 4229 19008
rect 4294 19002 4354 19214
rect 4470 19212 4476 19276
rect 4540 19274 4546 19276
rect 8753 19274 8819 19277
rect 4540 19272 8819 19274
rect 4540 19216 8758 19272
rect 8814 19216 8819 19272
rect 4540 19214 8819 19216
rect 4540 19212 4546 19214
rect 8753 19211 8819 19214
rect 11145 19274 11211 19277
rect 15745 19274 15811 19277
rect 11145 19272 15811 19274
rect 11145 19216 11150 19272
rect 11206 19216 15750 19272
rect 15806 19216 15811 19272
rect 11145 19214 15811 19216
rect 11145 19211 11211 19214
rect 15745 19211 15811 19214
rect 9847 19072 10163 19073
rect 9847 19008 9853 19072
rect 9917 19008 9933 19072
rect 9997 19008 10013 19072
rect 10077 19008 10093 19072
rect 10157 19008 10163 19072
rect 9847 19007 10163 19008
rect 15781 19072 16097 19073
rect 15781 19008 15787 19072
rect 15851 19008 15867 19072
rect 15931 19008 15947 19072
rect 16011 19008 16027 19072
rect 16091 19008 16097 19072
rect 15781 19007 16097 19008
rect 21715 19072 22031 19073
rect 21715 19008 21721 19072
rect 21785 19008 21801 19072
rect 21865 19008 21881 19072
rect 21945 19008 21961 19072
rect 22025 19008 22031 19072
rect 21715 19007 22031 19008
rect 4613 19002 4679 19005
rect 8293 19002 8359 19005
rect 4294 19000 8359 19002
rect 4294 18944 4618 19000
rect 4674 18944 8298 19000
rect 8354 18944 8359 19000
rect 4294 18942 8359 18944
rect 4613 18939 4679 18942
rect 8293 18939 8359 18942
rect 0 18866 160 18896
rect 933 18866 999 18869
rect 0 18864 999 18866
rect 0 18808 938 18864
rect 994 18808 999 18864
rect 0 18806 999 18808
rect 0 18776 160 18806
rect 933 18803 999 18806
rect 1945 18866 2011 18869
rect 7189 18866 7255 18869
rect 1945 18864 7255 18866
rect 1945 18808 1950 18864
rect 2006 18808 7194 18864
rect 7250 18808 7255 18864
rect 1945 18806 7255 18808
rect 1945 18803 2011 18806
rect 7189 18803 7255 18806
rect 10542 18804 10548 18868
rect 10612 18866 10618 18868
rect 14733 18866 14799 18869
rect 10612 18864 14799 18866
rect 10612 18808 14738 18864
rect 14794 18808 14799 18864
rect 10612 18806 14799 18808
rect 10612 18804 10618 18806
rect 14733 18803 14799 18806
rect 24393 18866 24459 18869
rect 25840 18866 26000 18896
rect 24393 18864 26000 18866
rect 24393 18808 24398 18864
rect 24454 18808 26000 18864
rect 24393 18806 26000 18808
rect 24393 18803 24459 18806
rect 25840 18776 26000 18806
rect 1577 18730 1643 18733
rect 6729 18730 6795 18733
rect 1577 18728 6795 18730
rect 1577 18672 1582 18728
rect 1638 18672 6734 18728
rect 6790 18672 6795 18728
rect 1577 18670 6795 18672
rect 1577 18667 1643 18670
rect 6729 18667 6795 18670
rect 8661 18730 8727 18733
rect 20621 18730 20687 18733
rect 8661 18728 20687 18730
rect 8661 18672 8666 18728
rect 8722 18672 20626 18728
rect 20682 18672 20687 18728
rect 8661 18670 20687 18672
rect 8661 18667 8727 18670
rect 20621 18667 20687 18670
rect 0 18594 160 18624
rect 749 18594 815 18597
rect 2865 18594 2931 18597
rect 0 18592 815 18594
rect 0 18536 754 18592
rect 810 18536 815 18592
rect 0 18534 815 18536
rect 0 18504 160 18534
rect 749 18531 815 18534
rect 2730 18592 2931 18594
rect 2730 18536 2870 18592
rect 2926 18536 2931 18592
rect 2730 18534 2931 18536
rect 0 18322 160 18352
rect 2730 18322 2790 18534
rect 2865 18531 2931 18534
rect 6880 18528 7196 18529
rect 6880 18464 6886 18528
rect 6950 18464 6966 18528
rect 7030 18464 7046 18528
rect 7110 18464 7126 18528
rect 7190 18464 7196 18528
rect 6880 18463 7196 18464
rect 12814 18528 13130 18529
rect 12814 18464 12820 18528
rect 12884 18464 12900 18528
rect 12964 18464 12980 18528
rect 13044 18464 13060 18528
rect 13124 18464 13130 18528
rect 12814 18463 13130 18464
rect 18748 18528 19064 18529
rect 18748 18464 18754 18528
rect 18818 18464 18834 18528
rect 18898 18464 18914 18528
rect 18978 18464 18994 18528
rect 19058 18464 19064 18528
rect 18748 18463 19064 18464
rect 24682 18528 24998 18529
rect 24682 18464 24688 18528
rect 24752 18464 24768 18528
rect 24832 18464 24848 18528
rect 24912 18464 24928 18528
rect 24992 18464 24998 18528
rect 24682 18463 24998 18464
rect 3509 18322 3575 18325
rect 0 18262 2790 18322
rect 3006 18320 3575 18322
rect 3006 18264 3514 18320
rect 3570 18264 3575 18320
rect 3006 18262 3575 18264
rect 0 18232 160 18262
rect 1945 18186 2011 18189
rect 3006 18186 3066 18262
rect 3509 18259 3575 18262
rect 12065 18322 12131 18325
rect 17677 18322 17743 18325
rect 12065 18320 17743 18322
rect 12065 18264 12070 18320
rect 12126 18264 17682 18320
rect 17738 18264 17743 18320
rect 12065 18262 17743 18264
rect 12065 18259 12131 18262
rect 17677 18259 17743 18262
rect 24393 18322 24459 18325
rect 25840 18322 26000 18352
rect 24393 18320 26000 18322
rect 24393 18264 24398 18320
rect 24454 18264 26000 18320
rect 24393 18262 26000 18264
rect 24393 18259 24459 18262
rect 25840 18232 26000 18262
rect 1945 18184 3066 18186
rect 1945 18128 1950 18184
rect 2006 18128 3066 18184
rect 1945 18126 3066 18128
rect 1945 18123 2011 18126
rect 9622 18124 9628 18188
rect 9692 18186 9698 18188
rect 10685 18186 10751 18189
rect 9692 18184 10751 18186
rect 9692 18128 10690 18184
rect 10746 18128 10751 18184
rect 9692 18126 10751 18128
rect 9692 18124 9698 18126
rect 10685 18123 10751 18126
rect 10961 18186 11027 18189
rect 15929 18186 15995 18189
rect 10961 18184 15995 18186
rect 10961 18128 10966 18184
rect 11022 18128 15934 18184
rect 15990 18128 15995 18184
rect 10961 18126 15995 18128
rect 10961 18123 11027 18126
rect 15929 18123 15995 18126
rect 16113 18186 16179 18189
rect 16430 18186 16436 18188
rect 16113 18184 16436 18186
rect 16113 18128 16118 18184
rect 16174 18128 16436 18184
rect 16113 18126 16436 18128
rect 16113 18123 16179 18126
rect 16430 18124 16436 18126
rect 16500 18124 16506 18188
rect 0 18050 160 18080
rect 1393 18050 1459 18053
rect 21357 18052 21423 18053
rect 21357 18050 21404 18052
rect 0 18048 1459 18050
rect 0 17992 1398 18048
rect 1454 17992 1459 18048
rect 0 17990 1459 17992
rect 21312 18048 21404 18050
rect 21312 17992 21362 18048
rect 21312 17990 21404 17992
rect 0 17960 160 17990
rect 1393 17987 1459 17990
rect 21357 17988 21404 17990
rect 21468 17988 21474 18052
rect 21357 17987 21423 17988
rect 3913 17984 4229 17985
rect 3913 17920 3919 17984
rect 3983 17920 3999 17984
rect 4063 17920 4079 17984
rect 4143 17920 4159 17984
rect 4223 17920 4229 17984
rect 3913 17919 4229 17920
rect 9847 17984 10163 17985
rect 9847 17920 9853 17984
rect 9917 17920 9933 17984
rect 9997 17920 10013 17984
rect 10077 17920 10093 17984
rect 10157 17920 10163 17984
rect 9847 17919 10163 17920
rect 15781 17984 16097 17985
rect 15781 17920 15787 17984
rect 15851 17920 15867 17984
rect 15931 17920 15947 17984
rect 16011 17920 16027 17984
rect 16091 17920 16097 17984
rect 15781 17919 16097 17920
rect 21715 17984 22031 17985
rect 21715 17920 21721 17984
rect 21785 17920 21801 17984
rect 21865 17920 21881 17984
rect 21945 17920 21961 17984
rect 22025 17920 22031 17984
rect 21715 17919 22031 17920
rect 24117 17914 24183 17917
rect 24117 17912 24962 17914
rect 24117 17856 24122 17912
rect 24178 17856 24962 17912
rect 24117 17854 24962 17856
rect 24117 17851 24183 17854
rect 0 17778 160 17808
rect 1301 17778 1367 17781
rect 0 17776 1367 17778
rect 0 17720 1306 17776
rect 1362 17720 1367 17776
rect 0 17718 1367 17720
rect 0 17688 160 17718
rect 1301 17715 1367 17718
rect 1761 17778 1827 17781
rect 4245 17778 4311 17781
rect 1761 17776 4311 17778
rect 1761 17720 1766 17776
rect 1822 17720 4250 17776
rect 4306 17720 4311 17776
rect 1761 17718 4311 17720
rect 1761 17715 1827 17718
rect 4245 17715 4311 17718
rect 5993 17778 6059 17781
rect 11462 17778 11468 17780
rect 5993 17776 11468 17778
rect 5993 17720 5998 17776
rect 6054 17720 11468 17776
rect 5993 17718 11468 17720
rect 5993 17715 6059 17718
rect 11462 17716 11468 17718
rect 11532 17716 11538 17780
rect 13353 17778 13419 17781
rect 13486 17778 13492 17780
rect 13353 17776 13492 17778
rect 13353 17720 13358 17776
rect 13414 17720 13492 17776
rect 13353 17718 13492 17720
rect 13353 17715 13419 17718
rect 13486 17716 13492 17718
rect 13556 17716 13562 17780
rect 24902 17778 24962 17854
rect 25840 17778 26000 17808
rect 24902 17718 26000 17778
rect 25840 17688 26000 17718
rect 9673 17642 9739 17645
rect 10317 17642 10383 17645
rect 9673 17640 10383 17642
rect 9673 17584 9678 17640
rect 9734 17584 10322 17640
rect 10378 17584 10383 17640
rect 9673 17582 10383 17584
rect 9673 17579 9739 17582
rect 10317 17579 10383 17582
rect 11513 17642 11579 17645
rect 11646 17642 11652 17644
rect 11513 17640 11652 17642
rect 11513 17584 11518 17640
rect 11574 17584 11652 17640
rect 11513 17582 11652 17584
rect 11513 17579 11579 17582
rect 11646 17580 11652 17582
rect 11716 17580 11722 17644
rect 13486 17580 13492 17644
rect 13556 17642 13562 17644
rect 23105 17642 23171 17645
rect 13556 17640 23171 17642
rect 13556 17584 23110 17640
rect 23166 17584 23171 17640
rect 13556 17582 23171 17584
rect 13556 17580 13562 17582
rect 23105 17579 23171 17582
rect 0 17506 160 17536
rect 933 17506 999 17509
rect 0 17504 999 17506
rect 0 17448 938 17504
rect 994 17448 999 17504
rect 0 17446 999 17448
rect 0 17416 160 17446
rect 933 17443 999 17446
rect 6880 17440 7196 17441
rect 6880 17376 6886 17440
rect 6950 17376 6966 17440
rect 7030 17376 7046 17440
rect 7110 17376 7126 17440
rect 7190 17376 7196 17440
rect 6880 17375 7196 17376
rect 12814 17440 13130 17441
rect 12814 17376 12820 17440
rect 12884 17376 12900 17440
rect 12964 17376 12980 17440
rect 13044 17376 13060 17440
rect 13124 17376 13130 17440
rect 12814 17375 13130 17376
rect 18748 17440 19064 17441
rect 18748 17376 18754 17440
rect 18818 17376 18834 17440
rect 18898 17376 18914 17440
rect 18978 17376 18994 17440
rect 19058 17376 19064 17440
rect 18748 17375 19064 17376
rect 24682 17440 24998 17441
rect 24682 17376 24688 17440
rect 24752 17376 24768 17440
rect 24832 17376 24848 17440
rect 24912 17376 24928 17440
rect 24992 17376 24998 17440
rect 24682 17375 24998 17376
rect 19425 17370 19491 17373
rect 19742 17370 19748 17372
rect 19425 17368 19748 17370
rect 19425 17312 19430 17368
rect 19486 17312 19748 17368
rect 19425 17310 19748 17312
rect 19425 17307 19491 17310
rect 19742 17308 19748 17310
rect 19812 17308 19818 17372
rect 0 17234 160 17264
rect 1853 17234 1919 17237
rect 0 17232 1919 17234
rect 0 17176 1858 17232
rect 1914 17176 1919 17232
rect 0 17174 1919 17176
rect 0 17144 160 17174
rect 1853 17171 1919 17174
rect 2221 17234 2287 17237
rect 17125 17234 17191 17237
rect 2221 17232 17191 17234
rect 2221 17176 2226 17232
rect 2282 17176 17130 17232
rect 17186 17176 17191 17232
rect 2221 17174 17191 17176
rect 2221 17171 2287 17174
rect 17125 17171 17191 17174
rect 18321 17234 18387 17237
rect 19926 17234 19932 17236
rect 18321 17232 19932 17234
rect 18321 17176 18326 17232
rect 18382 17176 19932 17232
rect 18321 17174 19932 17176
rect 18321 17171 18387 17174
rect 19926 17172 19932 17174
rect 19996 17172 20002 17236
rect 24025 17234 24091 17237
rect 25840 17234 26000 17264
rect 24025 17232 26000 17234
rect 24025 17176 24030 17232
rect 24086 17176 26000 17232
rect 24025 17174 26000 17176
rect 24025 17171 24091 17174
rect 25840 17144 26000 17174
rect 9673 17098 9739 17101
rect 10961 17098 11027 17101
rect 9673 17096 11027 17098
rect 9673 17040 9678 17096
rect 9734 17040 10966 17096
rect 11022 17040 11027 17096
rect 9673 17038 11027 17040
rect 9673 17035 9739 17038
rect 10961 17035 11027 17038
rect 0 16962 160 16992
rect 1301 16962 1367 16965
rect 0 16960 1367 16962
rect 0 16904 1306 16960
rect 1362 16904 1367 16960
rect 0 16902 1367 16904
rect 0 16872 160 16902
rect 1301 16899 1367 16902
rect 1669 16960 1735 16965
rect 1669 16904 1674 16960
rect 1730 16904 1735 16960
rect 1669 16899 1735 16904
rect 0 16690 160 16720
rect 1672 16693 1732 16899
rect 3913 16896 4229 16897
rect 3913 16832 3919 16896
rect 3983 16832 3999 16896
rect 4063 16832 4079 16896
rect 4143 16832 4159 16896
rect 4223 16832 4229 16896
rect 3913 16831 4229 16832
rect 9847 16896 10163 16897
rect 9847 16832 9853 16896
rect 9917 16832 9933 16896
rect 9997 16832 10013 16896
rect 10077 16832 10093 16896
rect 10157 16832 10163 16896
rect 9847 16831 10163 16832
rect 15781 16896 16097 16897
rect 15781 16832 15787 16896
rect 15851 16832 15867 16896
rect 15931 16832 15947 16896
rect 16011 16832 16027 16896
rect 16091 16832 16097 16896
rect 15781 16831 16097 16832
rect 21715 16896 22031 16897
rect 21715 16832 21721 16896
rect 21785 16832 21801 16896
rect 21865 16832 21881 16896
rect 21945 16832 21961 16896
rect 22025 16832 22031 16896
rect 21715 16831 22031 16832
rect 1301 16690 1367 16693
rect 0 16688 1367 16690
rect 0 16632 1306 16688
rect 1362 16632 1367 16688
rect 0 16630 1367 16632
rect 0 16600 160 16630
rect 1301 16627 1367 16630
rect 1669 16688 1735 16693
rect 1669 16632 1674 16688
rect 1730 16632 1735 16688
rect 1669 16627 1735 16632
rect 4245 16690 4311 16693
rect 4654 16690 4660 16692
rect 4245 16688 4660 16690
rect 4245 16632 4250 16688
rect 4306 16632 4660 16688
rect 4245 16630 4660 16632
rect 4245 16627 4311 16630
rect 4654 16628 4660 16630
rect 4724 16628 4730 16692
rect 24393 16690 24459 16693
rect 25840 16690 26000 16720
rect 24393 16688 26000 16690
rect 24393 16632 24398 16688
rect 24454 16632 26000 16688
rect 24393 16630 26000 16632
rect 24393 16627 24459 16630
rect 25840 16600 26000 16630
rect 10685 16556 10751 16557
rect 10685 16554 10732 16556
rect 10640 16552 10732 16554
rect 10640 16496 10690 16552
rect 10640 16494 10732 16496
rect 10685 16492 10732 16494
rect 10796 16492 10802 16556
rect 13353 16554 13419 16557
rect 13854 16554 13860 16556
rect 13353 16552 13860 16554
rect 13353 16496 13358 16552
rect 13414 16496 13860 16552
rect 13353 16494 13860 16496
rect 10685 16491 10751 16492
rect 13353 16491 13419 16494
rect 13854 16492 13860 16494
rect 13924 16492 13930 16556
rect 23933 16554 23999 16557
rect 23933 16552 25146 16554
rect 23933 16496 23938 16552
rect 23994 16496 25146 16552
rect 23933 16494 25146 16496
rect 23933 16491 23999 16494
rect 0 16418 160 16448
rect 1761 16418 1827 16421
rect 0 16416 1827 16418
rect 0 16360 1766 16416
rect 1822 16360 1827 16416
rect 0 16358 1827 16360
rect 0 16328 160 16358
rect 1761 16355 1827 16358
rect 6880 16352 7196 16353
rect 6880 16288 6886 16352
rect 6950 16288 6966 16352
rect 7030 16288 7046 16352
rect 7110 16288 7126 16352
rect 7190 16288 7196 16352
rect 6880 16287 7196 16288
rect 12814 16352 13130 16353
rect 12814 16288 12820 16352
rect 12884 16288 12900 16352
rect 12964 16288 12980 16352
rect 13044 16288 13060 16352
rect 13124 16288 13130 16352
rect 12814 16287 13130 16288
rect 18748 16352 19064 16353
rect 18748 16288 18754 16352
rect 18818 16288 18834 16352
rect 18898 16288 18914 16352
rect 18978 16288 18994 16352
rect 19058 16288 19064 16352
rect 18748 16287 19064 16288
rect 24682 16352 24998 16353
rect 24682 16288 24688 16352
rect 24752 16288 24768 16352
rect 24832 16288 24848 16352
rect 24912 16288 24928 16352
rect 24992 16288 24998 16352
rect 24682 16287 24998 16288
rect 1117 16282 1183 16285
rect 1117 16280 1962 16282
rect 1117 16224 1122 16280
rect 1178 16224 1962 16280
rect 1117 16222 1962 16224
rect 1117 16219 1183 16222
rect 0 16146 160 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 160 16086
rect 1577 16083 1643 16086
rect 1902 16010 1962 16222
rect 2681 16146 2747 16149
rect 3182 16146 3188 16148
rect 2681 16144 3188 16146
rect 2681 16088 2686 16144
rect 2742 16088 3188 16144
rect 2681 16086 3188 16088
rect 2681 16083 2747 16086
rect 3182 16084 3188 16086
rect 3252 16084 3258 16148
rect 25086 16146 25146 16494
rect 25840 16146 26000 16176
rect 25086 16086 26000 16146
rect 25840 16056 26000 16086
rect 4613 16010 4679 16013
rect 1902 16008 4679 16010
rect 1902 15952 4618 16008
rect 4674 15952 4679 16008
rect 1902 15950 4679 15952
rect 4613 15947 4679 15950
rect 10910 15948 10916 16012
rect 10980 16010 10986 16012
rect 22318 16010 22324 16012
rect 10980 15950 22324 16010
rect 10980 15948 10986 15950
rect 22318 15948 22324 15950
rect 22388 15948 22394 16012
rect 0 15874 160 15904
rect 3693 15874 3759 15877
rect 0 15872 3759 15874
rect 0 15816 3698 15872
rect 3754 15816 3759 15872
rect 0 15814 3759 15816
rect 0 15784 160 15814
rect 3693 15811 3759 15814
rect 3913 15808 4229 15809
rect 3913 15744 3919 15808
rect 3983 15744 3999 15808
rect 4063 15744 4079 15808
rect 4143 15744 4159 15808
rect 4223 15744 4229 15808
rect 3913 15743 4229 15744
rect 9847 15808 10163 15809
rect 9847 15744 9853 15808
rect 9917 15744 9933 15808
rect 9997 15744 10013 15808
rect 10077 15744 10093 15808
rect 10157 15744 10163 15808
rect 9847 15743 10163 15744
rect 15781 15808 16097 15809
rect 15781 15744 15787 15808
rect 15851 15744 15867 15808
rect 15931 15744 15947 15808
rect 16011 15744 16027 15808
rect 16091 15744 16097 15808
rect 15781 15743 16097 15744
rect 21715 15808 22031 15809
rect 21715 15744 21721 15808
rect 21785 15744 21801 15808
rect 21865 15744 21881 15808
rect 21945 15744 21961 15808
rect 22025 15744 22031 15808
rect 21715 15743 22031 15744
rect 0 15602 160 15632
rect 2589 15602 2655 15605
rect 6821 15602 6887 15605
rect 0 15542 1042 15602
rect 0 15512 160 15542
rect 982 15466 1042 15542
rect 2589 15600 6887 15602
rect 2589 15544 2594 15600
rect 2650 15544 6826 15600
rect 6882 15544 6887 15600
rect 2589 15542 6887 15544
rect 2589 15539 2655 15542
rect 6821 15539 6887 15542
rect 23749 15602 23815 15605
rect 25840 15602 26000 15632
rect 23749 15600 26000 15602
rect 23749 15544 23754 15600
rect 23810 15544 26000 15600
rect 23749 15542 26000 15544
rect 23749 15539 23815 15542
rect 25840 15512 26000 15542
rect 1393 15466 1459 15469
rect 982 15464 1459 15466
rect 982 15408 1398 15464
rect 1454 15408 1459 15464
rect 982 15406 1459 15408
rect 1393 15403 1459 15406
rect 5257 15466 5323 15469
rect 11421 15466 11487 15469
rect 5257 15464 11487 15466
rect 5257 15408 5262 15464
rect 5318 15408 11426 15464
rect 11482 15408 11487 15464
rect 5257 15406 11487 15408
rect 5257 15403 5323 15406
rect 11421 15403 11487 15406
rect 11973 15466 12039 15469
rect 12709 15466 12775 15469
rect 14549 15466 14615 15469
rect 11973 15464 14615 15466
rect 11973 15408 11978 15464
rect 12034 15408 12714 15464
rect 12770 15408 14554 15464
rect 14610 15408 14615 15464
rect 11973 15406 14615 15408
rect 11973 15403 12039 15406
rect 12709 15403 12775 15406
rect 14549 15403 14615 15406
rect 0 15330 160 15360
rect 4061 15330 4127 15333
rect 0 15328 4127 15330
rect 0 15272 4066 15328
rect 4122 15272 4127 15328
rect 0 15270 4127 15272
rect 0 15240 160 15270
rect 4061 15267 4127 15270
rect 4613 15330 4679 15333
rect 6637 15330 6703 15333
rect 4613 15328 6703 15330
rect 4613 15272 4618 15328
rect 4674 15272 6642 15328
rect 6698 15272 6703 15328
rect 4613 15270 6703 15272
rect 4613 15267 4679 15270
rect 6637 15267 6703 15270
rect 6880 15264 7196 15265
rect 6880 15200 6886 15264
rect 6950 15200 6966 15264
rect 7030 15200 7046 15264
rect 7110 15200 7126 15264
rect 7190 15200 7196 15264
rect 6880 15199 7196 15200
rect 12814 15264 13130 15265
rect 12814 15200 12820 15264
rect 12884 15200 12900 15264
rect 12964 15200 12980 15264
rect 13044 15200 13060 15264
rect 13124 15200 13130 15264
rect 12814 15199 13130 15200
rect 18748 15264 19064 15265
rect 18748 15200 18754 15264
rect 18818 15200 18834 15264
rect 18898 15200 18914 15264
rect 18978 15200 18994 15264
rect 19058 15200 19064 15264
rect 18748 15199 19064 15200
rect 24682 15264 24998 15265
rect 24682 15200 24688 15264
rect 24752 15200 24768 15264
rect 24832 15200 24848 15264
rect 24912 15200 24928 15264
rect 24992 15200 24998 15264
rect 24682 15199 24998 15200
rect 18045 15194 18111 15197
rect 18270 15194 18276 15196
rect 18045 15192 18276 15194
rect 18045 15136 18050 15192
rect 18106 15136 18276 15192
rect 18045 15134 18276 15136
rect 18045 15131 18111 15134
rect 18270 15132 18276 15134
rect 18340 15132 18346 15196
rect 24117 15194 24183 15197
rect 24117 15192 24594 15194
rect 24117 15136 24122 15192
rect 24178 15136 24594 15192
rect 24117 15134 24594 15136
rect 24117 15131 24183 15134
rect 0 15058 160 15088
rect 1761 15058 1827 15061
rect 0 15056 1827 15058
rect 0 15000 1766 15056
rect 1822 15000 1827 15056
rect 0 14998 1827 15000
rect 24534 15058 24594 15134
rect 25840 15058 26000 15088
rect 24534 14998 26000 15058
rect 0 14968 160 14998
rect 1761 14995 1827 14998
rect 25840 14968 26000 14998
rect 17902 14860 17908 14924
rect 17972 14922 17978 14924
rect 19425 14922 19491 14925
rect 17972 14920 19491 14922
rect 17972 14864 19430 14920
rect 19486 14864 19491 14920
rect 17972 14862 19491 14864
rect 17972 14860 17978 14862
rect 19425 14859 19491 14862
rect 0 14786 160 14816
rect 1485 14786 1551 14789
rect 0 14784 1551 14786
rect 0 14728 1490 14784
rect 1546 14728 1551 14784
rect 0 14726 1551 14728
rect 0 14696 160 14726
rect 1485 14723 1551 14726
rect 3913 14720 4229 14721
rect 3913 14656 3919 14720
rect 3983 14656 3999 14720
rect 4063 14656 4079 14720
rect 4143 14656 4159 14720
rect 4223 14656 4229 14720
rect 3913 14655 4229 14656
rect 9847 14720 10163 14721
rect 9847 14656 9853 14720
rect 9917 14656 9933 14720
rect 9997 14656 10013 14720
rect 10077 14656 10093 14720
rect 10157 14656 10163 14720
rect 9847 14655 10163 14656
rect 15781 14720 16097 14721
rect 15781 14656 15787 14720
rect 15851 14656 15867 14720
rect 15931 14656 15947 14720
rect 16011 14656 16027 14720
rect 16091 14656 16097 14720
rect 15781 14655 16097 14656
rect 21715 14720 22031 14721
rect 21715 14656 21721 14720
rect 21785 14656 21801 14720
rect 21865 14656 21881 14720
rect 21945 14656 21961 14720
rect 22025 14656 22031 14720
rect 21715 14655 22031 14656
rect 0 14514 160 14544
rect 1301 14514 1367 14517
rect 0 14512 1367 14514
rect 0 14456 1306 14512
rect 1362 14456 1367 14512
rect 0 14454 1367 14456
rect 0 14424 160 14454
rect 1301 14451 1367 14454
rect 2221 14514 2287 14517
rect 15193 14514 15259 14517
rect 2221 14512 15259 14514
rect 2221 14456 2226 14512
rect 2282 14456 15198 14512
rect 15254 14456 15259 14512
rect 2221 14454 15259 14456
rect 2221 14451 2287 14454
rect 15193 14451 15259 14454
rect 24393 14514 24459 14517
rect 25840 14514 26000 14544
rect 24393 14512 26000 14514
rect 24393 14456 24398 14512
rect 24454 14456 26000 14512
rect 24393 14454 26000 14456
rect 24393 14451 24459 14454
rect 25840 14424 26000 14454
rect 0 14242 160 14272
rect 1669 14242 1735 14245
rect 0 14240 1735 14242
rect 0 14184 1674 14240
rect 1730 14184 1735 14240
rect 0 14182 1735 14184
rect 0 14152 160 14182
rect 1669 14179 1735 14182
rect 6880 14176 7196 14177
rect 6880 14112 6886 14176
rect 6950 14112 6966 14176
rect 7030 14112 7046 14176
rect 7110 14112 7126 14176
rect 7190 14112 7196 14176
rect 6880 14111 7196 14112
rect 12814 14176 13130 14177
rect 12814 14112 12820 14176
rect 12884 14112 12900 14176
rect 12964 14112 12980 14176
rect 13044 14112 13060 14176
rect 13124 14112 13130 14176
rect 12814 14111 13130 14112
rect 18748 14176 19064 14177
rect 18748 14112 18754 14176
rect 18818 14112 18834 14176
rect 18898 14112 18914 14176
rect 18978 14112 18994 14176
rect 19058 14112 19064 14176
rect 18748 14111 19064 14112
rect 24682 14176 24998 14177
rect 24682 14112 24688 14176
rect 24752 14112 24768 14176
rect 24832 14112 24848 14176
rect 24912 14112 24928 14176
rect 24992 14112 24998 14176
rect 24682 14111 24998 14112
rect 0 13970 160 14000
rect 1301 13970 1367 13973
rect 0 13968 1367 13970
rect 0 13912 1306 13968
rect 1362 13912 1367 13968
rect 0 13910 1367 13912
rect 0 13880 160 13910
rect 1301 13907 1367 13910
rect 2313 13970 2379 13973
rect 5441 13970 5507 13973
rect 14641 13972 14707 13973
rect 2313 13968 5507 13970
rect 2313 13912 2318 13968
rect 2374 13912 5446 13968
rect 5502 13912 5507 13968
rect 2313 13910 5507 13912
rect 2313 13907 2379 13910
rect 5441 13907 5507 13910
rect 14590 13908 14596 13972
rect 14660 13970 14707 13972
rect 24485 13970 24551 13973
rect 25840 13970 26000 14000
rect 14660 13968 14752 13970
rect 14702 13912 14752 13968
rect 14660 13910 14752 13912
rect 24485 13968 26000 13970
rect 24485 13912 24490 13968
rect 24546 13912 26000 13968
rect 24485 13910 26000 13912
rect 14660 13908 14707 13910
rect 14641 13907 14707 13908
rect 24485 13907 24551 13910
rect 25840 13880 26000 13910
rect 1301 13836 1367 13837
rect 1301 13834 1348 13836
rect 1256 13832 1348 13834
rect 1256 13776 1306 13832
rect 1256 13774 1348 13776
rect 1301 13772 1348 13774
rect 1412 13772 1418 13836
rect 1485 13834 1551 13837
rect 1853 13834 1919 13837
rect 3049 13836 3115 13837
rect 1485 13832 1919 13834
rect 1485 13776 1490 13832
rect 1546 13776 1858 13832
rect 1914 13776 1919 13832
rect 1485 13774 1919 13776
rect 1301 13771 1367 13772
rect 1485 13771 1551 13774
rect 1853 13771 1919 13774
rect 2998 13772 3004 13836
rect 3068 13834 3115 13836
rect 3068 13832 3160 13834
rect 3110 13776 3160 13832
rect 3068 13774 3160 13776
rect 3068 13772 3115 13774
rect 3049 13771 3115 13772
rect 0 13698 160 13728
rect 3509 13698 3575 13701
rect 0 13696 3575 13698
rect 0 13640 3514 13696
rect 3570 13640 3575 13696
rect 0 13638 3575 13640
rect 0 13608 160 13638
rect 3509 13635 3575 13638
rect 6494 13636 6500 13700
rect 6564 13698 6570 13700
rect 7741 13698 7807 13701
rect 8569 13698 8635 13701
rect 6564 13696 7807 13698
rect 6564 13640 7746 13696
rect 7802 13640 7807 13696
rect 6564 13638 7807 13640
rect 6564 13636 6570 13638
rect 7741 13635 7807 13638
rect 7974 13696 8635 13698
rect 7974 13640 8574 13696
rect 8630 13640 8635 13696
rect 7974 13638 8635 13640
rect 3913 13632 4229 13633
rect 3913 13568 3919 13632
rect 3983 13568 3999 13632
rect 4063 13568 4079 13632
rect 4143 13568 4159 13632
rect 4223 13568 4229 13632
rect 3913 13567 4229 13568
rect 2313 13562 2379 13565
rect 7974 13562 8034 13638
rect 8569 13635 8635 13638
rect 12198 13636 12204 13700
rect 12268 13698 12274 13700
rect 12341 13698 12407 13701
rect 12268 13696 12407 13698
rect 12268 13640 12346 13696
rect 12402 13640 12407 13696
rect 12268 13638 12407 13640
rect 12268 13636 12274 13638
rect 12341 13635 12407 13638
rect 13854 13636 13860 13700
rect 13924 13698 13930 13700
rect 13997 13698 14063 13701
rect 13924 13696 14063 13698
rect 13924 13640 14002 13696
rect 14058 13640 14063 13696
rect 13924 13638 14063 13640
rect 13924 13636 13930 13638
rect 13997 13635 14063 13638
rect 9847 13632 10163 13633
rect 9847 13568 9853 13632
rect 9917 13568 9933 13632
rect 9997 13568 10013 13632
rect 10077 13568 10093 13632
rect 10157 13568 10163 13632
rect 9847 13567 10163 13568
rect 15781 13632 16097 13633
rect 15781 13568 15787 13632
rect 15851 13568 15867 13632
rect 15931 13568 15947 13632
rect 16011 13568 16027 13632
rect 16091 13568 16097 13632
rect 15781 13567 16097 13568
rect 21715 13632 22031 13633
rect 21715 13568 21721 13632
rect 21785 13568 21801 13632
rect 21865 13568 21881 13632
rect 21945 13568 21961 13632
rect 22025 13568 22031 13632
rect 21715 13567 22031 13568
rect 1166 13560 2379 13562
rect 1166 13504 2318 13560
rect 2374 13504 2379 13560
rect 1166 13502 2379 13504
rect 0 13426 160 13456
rect 1166 13426 1226 13502
rect 2313 13499 2379 13502
rect 4846 13502 8034 13562
rect 0 13366 1226 13426
rect 1301 13426 1367 13429
rect 1710 13426 1716 13428
rect 1301 13424 1716 13426
rect 1301 13368 1306 13424
rect 1362 13368 1716 13424
rect 1301 13366 1716 13368
rect 0 13336 160 13366
rect 1301 13363 1367 13366
rect 1710 13364 1716 13366
rect 1780 13364 1786 13428
rect 2078 13364 2084 13428
rect 2148 13426 2154 13428
rect 2589 13426 2655 13429
rect 2148 13424 2655 13426
rect 2148 13368 2594 13424
rect 2650 13368 2655 13424
rect 2148 13366 2655 13368
rect 2148 13364 2154 13366
rect 2589 13363 2655 13366
rect 2078 13228 2084 13292
rect 2148 13290 2154 13292
rect 4846 13290 4906 13502
rect 5022 13364 5028 13428
rect 5092 13426 5098 13428
rect 10317 13426 10383 13429
rect 5092 13424 10383 13426
rect 5092 13368 10322 13424
rect 10378 13368 10383 13424
rect 5092 13366 10383 13368
rect 5092 13364 5098 13366
rect 10317 13363 10383 13366
rect 24669 13426 24735 13429
rect 25840 13426 26000 13456
rect 24669 13424 26000 13426
rect 24669 13368 24674 13424
rect 24730 13368 26000 13424
rect 24669 13366 26000 13368
rect 24669 13363 24735 13366
rect 25840 13336 26000 13366
rect 2148 13230 4906 13290
rect 2148 13228 2154 13230
rect 0 13154 160 13184
rect 3509 13154 3575 13157
rect 0 13152 3575 13154
rect 0 13096 3514 13152
rect 3570 13096 3575 13152
rect 0 13094 3575 13096
rect 0 13064 160 13094
rect 3509 13091 3575 13094
rect 6880 13088 7196 13089
rect 6880 13024 6886 13088
rect 6950 13024 6966 13088
rect 7030 13024 7046 13088
rect 7110 13024 7126 13088
rect 7190 13024 7196 13088
rect 6880 13023 7196 13024
rect 12814 13088 13130 13089
rect 12814 13024 12820 13088
rect 12884 13024 12900 13088
rect 12964 13024 12980 13088
rect 13044 13024 13060 13088
rect 13124 13024 13130 13088
rect 12814 13023 13130 13024
rect 18748 13088 19064 13089
rect 18748 13024 18754 13088
rect 18818 13024 18834 13088
rect 18898 13024 18914 13088
rect 18978 13024 18994 13088
rect 19058 13024 19064 13088
rect 18748 13023 19064 13024
rect 24682 13088 24998 13089
rect 24682 13024 24688 13088
rect 24752 13024 24768 13088
rect 24832 13024 24848 13088
rect 24912 13024 24928 13088
rect 24992 13024 24998 13088
rect 24682 13023 24998 13024
rect 3233 13018 3299 13021
rect 3969 13018 4035 13021
rect 3233 13016 4035 13018
rect 3233 12960 3238 13016
rect 3294 12960 3974 13016
rect 4030 12960 4035 13016
rect 3233 12958 4035 12960
rect 3233 12955 3299 12958
rect 3969 12955 4035 12958
rect 0 12882 160 12912
rect 1577 12882 1643 12885
rect 0 12880 1643 12882
rect 0 12824 1582 12880
rect 1638 12824 1643 12880
rect 0 12822 1643 12824
rect 0 12792 160 12822
rect 1577 12819 1643 12822
rect 4613 12882 4679 12885
rect 7373 12882 7439 12885
rect 10542 12882 10548 12884
rect 4613 12880 10548 12882
rect 4613 12824 4618 12880
rect 4674 12824 7378 12880
rect 7434 12824 10548 12880
rect 4613 12822 10548 12824
rect 4613 12819 4679 12822
rect 7373 12819 7439 12822
rect 10542 12820 10548 12822
rect 10612 12820 10618 12884
rect 14365 12882 14431 12885
rect 20621 12882 20687 12885
rect 14365 12880 20687 12882
rect 14365 12824 14370 12880
rect 14426 12824 20626 12880
rect 20682 12824 20687 12880
rect 14365 12822 20687 12824
rect 14365 12819 14431 12822
rect 20621 12819 20687 12822
rect 24025 12882 24091 12885
rect 25840 12882 26000 12912
rect 24025 12880 26000 12882
rect 24025 12824 24030 12880
rect 24086 12824 26000 12880
rect 24025 12822 26000 12824
rect 24025 12819 24091 12822
rect 25840 12792 26000 12822
rect 2446 12684 2452 12748
rect 2516 12746 2522 12748
rect 5533 12746 5599 12749
rect 7465 12746 7531 12749
rect 2516 12744 7531 12746
rect 2516 12688 5538 12744
rect 5594 12688 7470 12744
rect 7526 12688 7531 12744
rect 2516 12686 7531 12688
rect 2516 12684 2522 12686
rect 5533 12683 5599 12686
rect 7465 12683 7531 12686
rect 10409 12746 10475 12749
rect 13629 12746 13695 12749
rect 10409 12744 13695 12746
rect 10409 12688 10414 12744
rect 10470 12688 13634 12744
rect 13690 12688 13695 12744
rect 10409 12686 13695 12688
rect 10409 12683 10475 12686
rect 13629 12683 13695 12686
rect 0 12610 160 12640
rect 1669 12610 1735 12613
rect 0 12608 1735 12610
rect 0 12552 1674 12608
rect 1730 12552 1735 12608
rect 0 12550 1735 12552
rect 0 12520 160 12550
rect 1669 12547 1735 12550
rect 3417 12610 3483 12613
rect 3785 12610 3851 12613
rect 3417 12608 3851 12610
rect 3417 12552 3422 12608
rect 3478 12552 3790 12608
rect 3846 12552 3851 12608
rect 3417 12550 3851 12552
rect 3417 12547 3483 12550
rect 3785 12547 3851 12550
rect 3913 12544 4229 12545
rect 3913 12480 3919 12544
rect 3983 12480 3999 12544
rect 4063 12480 4079 12544
rect 4143 12480 4159 12544
rect 4223 12480 4229 12544
rect 3913 12479 4229 12480
rect 9847 12544 10163 12545
rect 9847 12480 9853 12544
rect 9917 12480 9933 12544
rect 9997 12480 10013 12544
rect 10077 12480 10093 12544
rect 10157 12480 10163 12544
rect 9847 12479 10163 12480
rect 15781 12544 16097 12545
rect 15781 12480 15787 12544
rect 15851 12480 15867 12544
rect 15931 12480 15947 12544
rect 16011 12480 16027 12544
rect 16091 12480 16097 12544
rect 15781 12479 16097 12480
rect 21715 12544 22031 12545
rect 21715 12480 21721 12544
rect 21785 12480 21801 12544
rect 21865 12480 21881 12544
rect 21945 12480 21961 12544
rect 22025 12480 22031 12544
rect 21715 12479 22031 12480
rect 0 12338 160 12368
rect 2313 12338 2379 12341
rect 4613 12338 4679 12341
rect 0 12278 1410 12338
rect 0 12248 160 12278
rect 1350 12202 1410 12278
rect 2313 12336 4679 12338
rect 2313 12280 2318 12336
rect 2374 12280 4618 12336
rect 4674 12280 4679 12336
rect 2313 12278 4679 12280
rect 2313 12275 2379 12278
rect 4613 12275 4679 12278
rect 5165 12338 5231 12341
rect 6637 12338 6703 12341
rect 5165 12336 6703 12338
rect 5165 12280 5170 12336
rect 5226 12280 6642 12336
rect 6698 12280 6703 12336
rect 5165 12278 6703 12280
rect 5165 12275 5231 12278
rect 6637 12275 6703 12278
rect 12341 12338 12407 12341
rect 18321 12338 18387 12341
rect 12341 12336 18387 12338
rect 12341 12280 12346 12336
rect 12402 12280 18326 12336
rect 18382 12280 18387 12336
rect 12341 12278 18387 12280
rect 12341 12275 12407 12278
rect 18321 12275 18387 12278
rect 22502 12276 22508 12340
rect 22572 12338 22578 12340
rect 22645 12338 22711 12341
rect 22572 12336 22711 12338
rect 22572 12280 22650 12336
rect 22706 12280 22711 12336
rect 22572 12278 22711 12280
rect 22572 12276 22578 12278
rect 22645 12275 22711 12278
rect 23841 12338 23907 12341
rect 25840 12338 26000 12368
rect 23841 12336 26000 12338
rect 23841 12280 23846 12336
rect 23902 12280 26000 12336
rect 23841 12278 26000 12280
rect 23841 12275 23907 12278
rect 25840 12248 26000 12278
rect 2773 12202 2839 12205
rect 1350 12200 2839 12202
rect 1350 12144 2778 12200
rect 2834 12144 2839 12200
rect 1350 12142 2839 12144
rect 2773 12139 2839 12142
rect 3325 12202 3391 12205
rect 5901 12202 5967 12205
rect 3325 12200 5967 12202
rect 3325 12144 3330 12200
rect 3386 12144 5906 12200
rect 5962 12144 5967 12200
rect 3325 12142 5967 12144
rect 3325 12139 3391 12142
rect 5901 12139 5967 12142
rect 0 12066 160 12096
rect 1301 12066 1367 12069
rect 0 12064 1367 12066
rect 0 12008 1306 12064
rect 1362 12008 1367 12064
rect 0 12006 1367 12008
rect 0 11976 160 12006
rect 1301 12003 1367 12006
rect 6880 12000 7196 12001
rect 6880 11936 6886 12000
rect 6950 11936 6966 12000
rect 7030 11936 7046 12000
rect 7110 11936 7126 12000
rect 7190 11936 7196 12000
rect 6880 11935 7196 11936
rect 12814 12000 13130 12001
rect 12814 11936 12820 12000
rect 12884 11936 12900 12000
rect 12964 11936 12980 12000
rect 13044 11936 13060 12000
rect 13124 11936 13130 12000
rect 12814 11935 13130 11936
rect 18748 12000 19064 12001
rect 18748 11936 18754 12000
rect 18818 11936 18834 12000
rect 18898 11936 18914 12000
rect 18978 11936 18994 12000
rect 19058 11936 19064 12000
rect 18748 11935 19064 11936
rect 24682 12000 24998 12001
rect 24682 11936 24688 12000
rect 24752 11936 24768 12000
rect 24832 11936 24848 12000
rect 24912 11936 24928 12000
rect 24992 11936 24998 12000
rect 24682 11935 24998 11936
rect 0 11794 160 11824
rect 3969 11794 4035 11797
rect 17769 11794 17835 11797
rect 0 11792 4035 11794
rect 0 11736 3974 11792
rect 4030 11736 4035 11792
rect 0 11734 4035 11736
rect 0 11704 160 11734
rect 3969 11731 4035 11734
rect 12390 11792 17835 11794
rect 12390 11736 17774 11792
rect 17830 11736 17835 11792
rect 12390 11734 17835 11736
rect 2865 11658 2931 11661
rect 4061 11658 4127 11661
rect 12390 11658 12450 11734
rect 17769 11731 17835 11734
rect 21909 11794 21975 11797
rect 22369 11794 22435 11797
rect 22829 11794 22895 11797
rect 21909 11792 22895 11794
rect 21909 11736 21914 11792
rect 21970 11736 22374 11792
rect 22430 11736 22834 11792
rect 22890 11736 22895 11792
rect 21909 11734 22895 11736
rect 21909 11731 21975 11734
rect 22369 11731 22435 11734
rect 22829 11731 22895 11734
rect 24393 11794 24459 11797
rect 25840 11794 26000 11824
rect 24393 11792 26000 11794
rect 24393 11736 24398 11792
rect 24454 11736 26000 11792
rect 24393 11734 26000 11736
rect 24393 11731 24459 11734
rect 25840 11704 26000 11734
rect 2865 11656 12450 11658
rect 2865 11600 2870 11656
rect 2926 11600 4066 11656
rect 4122 11600 12450 11656
rect 2865 11598 12450 11600
rect 2865 11595 2931 11598
rect 4061 11595 4127 11598
rect 0 11522 160 11552
rect 3233 11522 3299 11525
rect 0 11520 3299 11522
rect 0 11464 3238 11520
rect 3294 11464 3299 11520
rect 0 11462 3299 11464
rect 0 11432 160 11462
rect 3233 11459 3299 11462
rect 3913 11456 4229 11457
rect 3913 11392 3919 11456
rect 3983 11392 3999 11456
rect 4063 11392 4079 11456
rect 4143 11392 4159 11456
rect 4223 11392 4229 11456
rect 3913 11391 4229 11392
rect 9847 11456 10163 11457
rect 9847 11392 9853 11456
rect 9917 11392 9933 11456
rect 9997 11392 10013 11456
rect 10077 11392 10093 11456
rect 10157 11392 10163 11456
rect 9847 11391 10163 11392
rect 15781 11456 16097 11457
rect 15781 11392 15787 11456
rect 15851 11392 15867 11456
rect 15931 11392 15947 11456
rect 16011 11392 16027 11456
rect 16091 11392 16097 11456
rect 15781 11391 16097 11392
rect 21715 11456 22031 11457
rect 21715 11392 21721 11456
rect 21785 11392 21801 11456
rect 21865 11392 21881 11456
rect 21945 11392 21961 11456
rect 22025 11392 22031 11456
rect 21715 11391 22031 11392
rect 0 11250 160 11280
rect 1761 11250 1827 11253
rect 0 11248 1827 11250
rect 0 11192 1766 11248
rect 1822 11192 1827 11248
rect 0 11190 1827 11192
rect 0 11160 160 11190
rect 1761 11187 1827 11190
rect 2681 11250 2747 11253
rect 4797 11250 4863 11253
rect 2681 11248 4863 11250
rect 2681 11192 2686 11248
rect 2742 11192 4802 11248
rect 4858 11192 4863 11248
rect 2681 11190 4863 11192
rect 2681 11187 2747 11190
rect 4797 11187 4863 11190
rect 16021 11250 16087 11253
rect 16614 11250 16620 11252
rect 16021 11248 16620 11250
rect 16021 11192 16026 11248
rect 16082 11192 16620 11248
rect 16021 11190 16620 11192
rect 16021 11187 16087 11190
rect 16614 11188 16620 11190
rect 16684 11188 16690 11252
rect 25037 11250 25103 11253
rect 25840 11250 26000 11280
rect 25037 11248 26000 11250
rect 25037 11192 25042 11248
rect 25098 11192 26000 11248
rect 25037 11190 26000 11192
rect 25037 11187 25103 11190
rect 25840 11160 26000 11190
rect 15009 11114 15075 11117
rect 17217 11114 17283 11117
rect 15009 11112 17283 11114
rect 15009 11056 15014 11112
rect 15070 11056 17222 11112
rect 17278 11056 17283 11112
rect 15009 11054 17283 11056
rect 15009 11051 15075 11054
rect 17217 11051 17283 11054
rect 0 10978 160 11008
rect 3325 10978 3391 10981
rect 0 10976 3391 10978
rect 0 10920 3330 10976
rect 3386 10920 3391 10976
rect 0 10918 3391 10920
rect 0 10888 160 10918
rect 3325 10915 3391 10918
rect 21030 10916 21036 10980
rect 21100 10978 21106 10980
rect 21173 10978 21239 10981
rect 21100 10976 21239 10978
rect 21100 10920 21178 10976
rect 21234 10920 21239 10976
rect 21100 10918 21239 10920
rect 21100 10916 21106 10918
rect 21173 10915 21239 10918
rect 6880 10912 7196 10913
rect 6880 10848 6886 10912
rect 6950 10848 6966 10912
rect 7030 10848 7046 10912
rect 7110 10848 7126 10912
rect 7190 10848 7196 10912
rect 6880 10847 7196 10848
rect 12814 10912 13130 10913
rect 12814 10848 12820 10912
rect 12884 10848 12900 10912
rect 12964 10848 12980 10912
rect 13044 10848 13060 10912
rect 13124 10848 13130 10912
rect 12814 10847 13130 10848
rect 18748 10912 19064 10913
rect 18748 10848 18754 10912
rect 18818 10848 18834 10912
rect 18898 10848 18914 10912
rect 18978 10848 18994 10912
rect 19058 10848 19064 10912
rect 18748 10847 19064 10848
rect 24682 10912 24998 10913
rect 24682 10848 24688 10912
rect 24752 10848 24768 10912
rect 24832 10848 24848 10912
rect 24912 10848 24928 10912
rect 24992 10848 24998 10912
rect 24682 10847 24998 10848
rect 0 10706 160 10736
rect 3141 10706 3207 10709
rect 0 10704 3207 10706
rect 0 10648 3146 10704
rect 3202 10648 3207 10704
rect 0 10646 3207 10648
rect 0 10616 160 10646
rect 3141 10643 3207 10646
rect 3969 10706 4035 10709
rect 6821 10706 6887 10709
rect 3969 10704 6887 10706
rect 3969 10648 3974 10704
rect 4030 10648 6826 10704
rect 6882 10648 6887 10704
rect 3969 10646 6887 10648
rect 3969 10643 4035 10646
rect 6821 10643 6887 10646
rect 24485 10706 24551 10709
rect 25840 10706 26000 10736
rect 24485 10704 26000 10706
rect 24485 10648 24490 10704
rect 24546 10648 26000 10704
rect 24485 10646 26000 10648
rect 24485 10643 24551 10646
rect 25840 10616 26000 10646
rect 7189 10570 7255 10573
rect 7649 10570 7715 10573
rect 7189 10568 7715 10570
rect 7189 10512 7194 10568
rect 7250 10512 7654 10568
rect 7710 10512 7715 10568
rect 7189 10510 7715 10512
rect 7189 10507 7255 10510
rect 7649 10507 7715 10510
rect 9121 10570 9187 10573
rect 15285 10570 15351 10573
rect 9121 10568 11898 10570
rect 9121 10512 9126 10568
rect 9182 10512 11898 10568
rect 9121 10510 11898 10512
rect 9121 10507 9187 10510
rect 0 10434 160 10464
rect 1485 10434 1551 10437
rect 0 10432 1551 10434
rect 0 10376 1490 10432
rect 1546 10376 1551 10432
rect 0 10374 1551 10376
rect 11838 10434 11898 10510
rect 12390 10568 15351 10570
rect 12390 10512 15290 10568
rect 15346 10512 15351 10568
rect 12390 10510 15351 10512
rect 12390 10434 12450 10510
rect 15285 10507 15351 10510
rect 11838 10374 12450 10434
rect 12801 10434 12867 10437
rect 14958 10434 14964 10436
rect 12801 10432 14964 10434
rect 12801 10376 12806 10432
rect 12862 10376 14964 10432
rect 12801 10374 14964 10376
rect 0 10344 160 10374
rect 1485 10371 1551 10374
rect 12801 10371 12867 10374
rect 14958 10372 14964 10374
rect 15028 10372 15034 10436
rect 3913 10368 4229 10369
rect 3913 10304 3919 10368
rect 3983 10304 3999 10368
rect 4063 10304 4079 10368
rect 4143 10304 4159 10368
rect 4223 10304 4229 10368
rect 3913 10303 4229 10304
rect 9847 10368 10163 10369
rect 9847 10304 9853 10368
rect 9917 10304 9933 10368
rect 9997 10304 10013 10368
rect 10077 10304 10093 10368
rect 10157 10304 10163 10368
rect 9847 10303 10163 10304
rect 15781 10368 16097 10369
rect 15781 10304 15787 10368
rect 15851 10304 15867 10368
rect 15931 10304 15947 10368
rect 16011 10304 16027 10368
rect 16091 10304 16097 10368
rect 15781 10303 16097 10304
rect 21715 10368 22031 10369
rect 21715 10304 21721 10368
rect 21785 10304 21801 10368
rect 21865 10304 21881 10368
rect 21945 10304 21961 10368
rect 22025 10304 22031 10368
rect 21715 10303 22031 10304
rect 6913 10298 6979 10301
rect 7557 10298 7623 10301
rect 6913 10296 7623 10298
rect 6913 10240 6918 10296
rect 6974 10240 7562 10296
rect 7618 10240 7623 10296
rect 6913 10238 7623 10240
rect 6913 10235 6979 10238
rect 7557 10235 7623 10238
rect 0 10162 160 10192
rect 2313 10162 2379 10165
rect 0 10160 2379 10162
rect 0 10104 2318 10160
rect 2374 10104 2379 10160
rect 0 10102 2379 10104
rect 0 10072 160 10102
rect 2313 10099 2379 10102
rect 4797 10164 4863 10165
rect 4797 10160 4844 10164
rect 4908 10162 4914 10164
rect 11697 10162 11763 10165
rect 12065 10162 12131 10165
rect 16665 10162 16731 10165
rect 4797 10104 4802 10160
rect 4797 10100 4844 10104
rect 4908 10102 4954 10162
rect 11697 10160 16731 10162
rect 11697 10104 11702 10160
rect 11758 10104 12070 10160
rect 12126 10104 16670 10160
rect 16726 10104 16731 10160
rect 11697 10102 16731 10104
rect 4908 10100 4914 10102
rect 4797 10099 4863 10100
rect 11697 10099 11763 10102
rect 12065 10099 12131 10102
rect 16665 10099 16731 10102
rect 23841 10162 23907 10165
rect 25840 10162 26000 10192
rect 23841 10160 26000 10162
rect 23841 10104 23846 10160
rect 23902 10104 26000 10160
rect 23841 10102 26000 10104
rect 23841 10099 23907 10102
rect 25840 10072 26000 10102
rect 11789 10026 11855 10029
rect 16573 10026 16639 10029
rect 11789 10024 16639 10026
rect 11789 9968 11794 10024
rect 11850 9968 16578 10024
rect 16634 9968 16639 10024
rect 11789 9966 16639 9968
rect 11789 9963 11855 9966
rect 16573 9963 16639 9966
rect 0 9890 160 9920
rect 1393 9890 1459 9893
rect 0 9888 1459 9890
rect 0 9832 1398 9888
rect 1454 9832 1459 9888
rect 0 9830 1459 9832
rect 0 9800 160 9830
rect 1393 9827 1459 9830
rect 6880 9824 7196 9825
rect 6880 9760 6886 9824
rect 6950 9760 6966 9824
rect 7030 9760 7046 9824
rect 7110 9760 7126 9824
rect 7190 9760 7196 9824
rect 6880 9759 7196 9760
rect 12814 9824 13130 9825
rect 12814 9760 12820 9824
rect 12884 9760 12900 9824
rect 12964 9760 12980 9824
rect 13044 9760 13060 9824
rect 13124 9760 13130 9824
rect 12814 9759 13130 9760
rect 18748 9824 19064 9825
rect 18748 9760 18754 9824
rect 18818 9760 18834 9824
rect 18898 9760 18914 9824
rect 18978 9760 18994 9824
rect 19058 9760 19064 9824
rect 18748 9759 19064 9760
rect 24682 9824 24998 9825
rect 24682 9760 24688 9824
rect 24752 9760 24768 9824
rect 24832 9760 24848 9824
rect 24912 9760 24928 9824
rect 24992 9760 24998 9824
rect 24682 9759 24998 9760
rect 17217 9754 17283 9757
rect 17350 9754 17356 9756
rect 17217 9752 17356 9754
rect 17217 9696 17222 9752
rect 17278 9696 17356 9752
rect 17217 9694 17356 9696
rect 17217 9691 17283 9694
rect 17350 9692 17356 9694
rect 17420 9692 17426 9756
rect 0 9618 160 9648
rect 2865 9618 2931 9621
rect 0 9616 2931 9618
rect 0 9560 2870 9616
rect 2926 9560 2931 9616
rect 0 9558 2931 9560
rect 0 9528 160 9558
rect 2865 9555 2931 9558
rect 5165 9618 5231 9621
rect 5533 9618 5599 9621
rect 5165 9616 5599 9618
rect 5165 9560 5170 9616
rect 5226 9560 5538 9616
rect 5594 9560 5599 9616
rect 5165 9558 5599 9560
rect 5165 9555 5231 9558
rect 5533 9555 5599 9558
rect 23933 9618 23999 9621
rect 25840 9618 26000 9648
rect 23933 9616 26000 9618
rect 23933 9560 23938 9616
rect 23994 9560 26000 9616
rect 23933 9558 26000 9560
rect 23933 9555 23999 9558
rect 25840 9528 26000 9558
rect 2129 9482 2195 9485
rect 9397 9482 9463 9485
rect 21633 9484 21699 9485
rect 2129 9480 9463 9482
rect 2129 9424 2134 9480
rect 2190 9424 9402 9480
rect 9458 9424 9463 9480
rect 2129 9422 9463 9424
rect 2129 9419 2195 9422
rect 9397 9419 9463 9422
rect 21582 9420 21588 9484
rect 21652 9482 21699 9484
rect 21652 9480 21744 9482
rect 21694 9424 21744 9480
rect 21652 9422 21744 9424
rect 21652 9420 21699 9422
rect 21633 9419 21699 9420
rect 0 9346 160 9376
rect 0 9286 1594 9346
rect 0 9256 160 9286
rect 0 9074 160 9104
rect 1301 9074 1367 9077
rect 0 9072 1367 9074
rect 0 9016 1306 9072
rect 1362 9016 1367 9072
rect 0 9014 1367 9016
rect 0 8984 160 9014
rect 1301 9011 1367 9014
rect 1534 8938 1594 9286
rect 3913 9280 4229 9281
rect 3913 9216 3919 9280
rect 3983 9216 3999 9280
rect 4063 9216 4079 9280
rect 4143 9216 4159 9280
rect 4223 9216 4229 9280
rect 3913 9215 4229 9216
rect 9847 9280 10163 9281
rect 9847 9216 9853 9280
rect 9917 9216 9933 9280
rect 9997 9216 10013 9280
rect 10077 9216 10093 9280
rect 10157 9216 10163 9280
rect 9847 9215 10163 9216
rect 15781 9280 16097 9281
rect 15781 9216 15787 9280
rect 15851 9216 15867 9280
rect 15931 9216 15947 9280
rect 16011 9216 16027 9280
rect 16091 9216 16097 9280
rect 15781 9215 16097 9216
rect 21715 9280 22031 9281
rect 21715 9216 21721 9280
rect 21785 9216 21801 9280
rect 21865 9216 21881 9280
rect 21945 9216 21961 9280
rect 22025 9216 22031 9280
rect 21715 9215 22031 9216
rect 5901 9210 5967 9213
rect 7373 9210 7439 9213
rect 5901 9208 7439 9210
rect 5901 9152 5906 9208
rect 5962 9152 7378 9208
rect 7434 9152 7439 9208
rect 5901 9150 7439 9152
rect 5901 9147 5967 9150
rect 7373 9147 7439 9150
rect 6913 9074 6979 9077
rect 7465 9074 7531 9077
rect 8385 9074 8451 9077
rect 6913 9072 8451 9074
rect 6913 9016 6918 9072
rect 6974 9016 7470 9072
rect 7526 9016 8390 9072
rect 8446 9016 8451 9072
rect 6913 9014 8451 9016
rect 6913 9011 6979 9014
rect 7465 9011 7531 9014
rect 8385 9011 8451 9014
rect 12157 9074 12223 9077
rect 18321 9074 18387 9077
rect 12157 9072 18387 9074
rect 12157 9016 12162 9072
rect 12218 9016 18326 9072
rect 18382 9016 18387 9072
rect 12157 9014 18387 9016
rect 12157 9011 12223 9014
rect 18321 9011 18387 9014
rect 23841 9074 23907 9077
rect 25840 9074 26000 9104
rect 23841 9072 26000 9074
rect 23841 9016 23846 9072
rect 23902 9016 26000 9072
rect 23841 9014 26000 9016
rect 23841 9011 23907 9014
rect 25840 8984 26000 9014
rect 1853 8938 1919 8941
rect 1534 8936 1919 8938
rect 1534 8880 1858 8936
rect 1914 8880 1919 8936
rect 1534 8878 1919 8880
rect 1853 8875 1919 8878
rect 2313 8938 2379 8941
rect 3417 8938 3483 8941
rect 24485 8938 24551 8941
rect 2313 8936 24551 8938
rect 2313 8880 2318 8936
rect 2374 8880 3422 8936
rect 3478 8880 24490 8936
rect 24546 8880 24551 8936
rect 2313 8878 24551 8880
rect 2313 8875 2379 8878
rect 3417 8875 3483 8878
rect 24485 8875 24551 8878
rect 0 8802 160 8832
rect 2865 8802 2931 8805
rect 0 8800 2931 8802
rect 0 8744 2870 8800
rect 2926 8744 2931 8800
rect 0 8742 2931 8744
rect 0 8712 160 8742
rect 2865 8739 2931 8742
rect 13445 8802 13511 8805
rect 17493 8802 17559 8805
rect 13445 8800 17559 8802
rect 13445 8744 13450 8800
rect 13506 8744 17498 8800
rect 17554 8744 17559 8800
rect 13445 8742 17559 8744
rect 13445 8739 13511 8742
rect 17493 8739 17559 8742
rect 6880 8736 7196 8737
rect 6880 8672 6886 8736
rect 6950 8672 6966 8736
rect 7030 8672 7046 8736
rect 7110 8672 7126 8736
rect 7190 8672 7196 8736
rect 6880 8671 7196 8672
rect 12814 8736 13130 8737
rect 12814 8672 12820 8736
rect 12884 8672 12900 8736
rect 12964 8672 12980 8736
rect 13044 8672 13060 8736
rect 13124 8672 13130 8736
rect 12814 8671 13130 8672
rect 18748 8736 19064 8737
rect 18748 8672 18754 8736
rect 18818 8672 18834 8736
rect 18898 8672 18914 8736
rect 18978 8672 18994 8736
rect 19058 8672 19064 8736
rect 18748 8671 19064 8672
rect 24682 8736 24998 8737
rect 24682 8672 24688 8736
rect 24752 8672 24768 8736
rect 24832 8672 24848 8736
rect 24912 8672 24928 8736
rect 24992 8672 24998 8736
rect 24682 8671 24998 8672
rect 606 8604 612 8668
rect 676 8666 682 8668
rect 4286 8666 4292 8668
rect 676 8606 4292 8666
rect 676 8604 682 8606
rect 4286 8604 4292 8606
rect 4356 8604 4362 8668
rect 17350 8604 17356 8668
rect 17420 8604 17426 8668
rect 0 8530 160 8560
rect 1577 8530 1643 8533
rect 0 8528 1643 8530
rect 0 8472 1582 8528
rect 1638 8472 1643 8528
rect 0 8470 1643 8472
rect 0 8440 160 8470
rect 1577 8467 1643 8470
rect 3325 8530 3391 8533
rect 3785 8530 3851 8533
rect 3325 8528 3851 8530
rect 3325 8472 3330 8528
rect 3386 8472 3790 8528
rect 3846 8472 3851 8528
rect 3325 8470 3851 8472
rect 3325 8467 3391 8470
rect 3785 8467 3851 8470
rect 3969 8530 4035 8533
rect 7649 8530 7715 8533
rect 3969 8528 7715 8530
rect 3969 8472 3974 8528
rect 4030 8472 7654 8528
rect 7710 8472 7715 8528
rect 3969 8470 7715 8472
rect 3969 8467 4035 8470
rect 7649 8467 7715 8470
rect 17358 8397 17418 8604
rect 23933 8530 23999 8533
rect 25840 8530 26000 8560
rect 23933 8528 26000 8530
rect 23933 8472 23938 8528
rect 23994 8472 26000 8528
rect 23933 8470 26000 8472
rect 23933 8467 23999 8470
rect 25840 8440 26000 8470
rect 3785 8394 3851 8397
rect 5390 8394 5396 8396
rect 3785 8392 5396 8394
rect 3785 8336 3790 8392
rect 3846 8336 5396 8392
rect 3785 8334 5396 8336
rect 3785 8331 3851 8334
rect 5390 8332 5396 8334
rect 5460 8332 5466 8396
rect 6545 8394 6611 8397
rect 7925 8394 7991 8397
rect 6545 8392 7991 8394
rect 6545 8336 6550 8392
rect 6606 8336 7930 8392
rect 7986 8336 7991 8392
rect 6545 8334 7991 8336
rect 17358 8392 17467 8397
rect 17358 8336 17406 8392
rect 17462 8336 17467 8392
rect 17358 8334 17467 8336
rect 6545 8331 6611 8334
rect 7925 8331 7991 8334
rect 17401 8331 17467 8334
rect 0 8258 160 8288
rect 0 8198 1042 8258
rect 0 8168 160 8198
rect 982 8122 1042 8198
rect 3913 8192 4229 8193
rect 3913 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4229 8192
rect 3913 8127 4229 8128
rect 9847 8192 10163 8193
rect 9847 8128 9853 8192
rect 9917 8128 9933 8192
rect 9997 8128 10013 8192
rect 10077 8128 10093 8192
rect 10157 8128 10163 8192
rect 9847 8127 10163 8128
rect 15781 8192 16097 8193
rect 15781 8128 15787 8192
rect 15851 8128 15867 8192
rect 15931 8128 15947 8192
rect 16011 8128 16027 8192
rect 16091 8128 16097 8192
rect 15781 8127 16097 8128
rect 21715 8192 22031 8193
rect 21715 8128 21721 8192
rect 21785 8128 21801 8192
rect 21865 8128 21881 8192
rect 21945 8128 21961 8192
rect 22025 8128 22031 8192
rect 21715 8127 22031 8128
rect 1761 8122 1827 8125
rect 982 8120 1827 8122
rect 982 8064 1766 8120
rect 1822 8064 1827 8120
rect 982 8062 1827 8064
rect 1761 8059 1827 8062
rect 0 7986 160 8016
rect 3049 7986 3115 7989
rect 0 7984 3115 7986
rect 0 7928 3054 7984
rect 3110 7928 3115 7984
rect 0 7926 3115 7928
rect 0 7896 160 7926
rect 3049 7923 3115 7926
rect 16849 7986 16915 7989
rect 19558 7986 19564 7988
rect 16849 7984 19564 7986
rect 16849 7928 16854 7984
rect 16910 7928 19564 7984
rect 16849 7926 19564 7928
rect 16849 7923 16915 7926
rect 19558 7924 19564 7926
rect 19628 7924 19634 7988
rect 25313 7986 25379 7989
rect 25840 7986 26000 8016
rect 25313 7984 26000 7986
rect 25313 7928 25318 7984
rect 25374 7928 26000 7984
rect 25313 7926 26000 7928
rect 25313 7923 25379 7926
rect 25840 7896 26000 7926
rect 2129 7850 2195 7853
rect 7465 7850 7531 7853
rect 2129 7848 7531 7850
rect 2129 7792 2134 7848
rect 2190 7792 7470 7848
rect 7526 7792 7531 7848
rect 2129 7790 7531 7792
rect 2129 7787 2195 7790
rect 7465 7787 7531 7790
rect 0 7714 160 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 160 7654
rect 1301 7651 1367 7654
rect 6880 7648 7196 7649
rect 6880 7584 6886 7648
rect 6950 7584 6966 7648
rect 7030 7584 7046 7648
rect 7110 7584 7126 7648
rect 7190 7584 7196 7648
rect 6880 7583 7196 7584
rect 12814 7648 13130 7649
rect 12814 7584 12820 7648
rect 12884 7584 12900 7648
rect 12964 7584 12980 7648
rect 13044 7584 13060 7648
rect 13124 7584 13130 7648
rect 12814 7583 13130 7584
rect 18748 7648 19064 7649
rect 18748 7584 18754 7648
rect 18818 7584 18834 7648
rect 18898 7584 18914 7648
rect 18978 7584 18994 7648
rect 19058 7584 19064 7648
rect 18748 7583 19064 7584
rect 24682 7648 24998 7649
rect 24682 7584 24688 7648
rect 24752 7584 24768 7648
rect 24832 7584 24848 7648
rect 24912 7584 24928 7648
rect 24992 7584 24998 7648
rect 24682 7583 24998 7584
rect 0 7442 160 7472
rect 24209 7442 24275 7445
rect 25840 7442 26000 7472
rect 0 7382 858 7442
rect 0 7352 160 7382
rect 798 7306 858 7382
rect 24209 7440 26000 7442
rect 24209 7384 24214 7440
rect 24270 7384 26000 7440
rect 24209 7382 26000 7384
rect 24209 7379 24275 7382
rect 25840 7352 26000 7382
rect 1393 7306 1459 7309
rect 798 7304 1459 7306
rect 798 7248 1398 7304
rect 1454 7248 1459 7304
rect 798 7246 1459 7248
rect 1393 7243 1459 7246
rect 13721 7306 13787 7309
rect 20110 7306 20116 7308
rect 13721 7304 20116 7306
rect 13721 7248 13726 7304
rect 13782 7248 20116 7304
rect 13721 7246 20116 7248
rect 13721 7243 13787 7246
rect 20110 7244 20116 7246
rect 20180 7244 20186 7308
rect 21081 7306 21147 7309
rect 24209 7306 24275 7309
rect 21081 7304 24275 7306
rect 21081 7248 21086 7304
rect 21142 7248 24214 7304
rect 24270 7248 24275 7304
rect 21081 7246 24275 7248
rect 21081 7243 21147 7246
rect 24209 7243 24275 7246
rect 0 7170 160 7200
rect 1301 7170 1367 7173
rect 0 7168 1367 7170
rect 0 7112 1306 7168
rect 1362 7112 1367 7168
rect 0 7110 1367 7112
rect 0 7080 160 7110
rect 1301 7107 1367 7110
rect 16665 7170 16731 7173
rect 18413 7170 18479 7173
rect 16665 7168 18479 7170
rect 16665 7112 16670 7168
rect 16726 7112 18418 7168
rect 18474 7112 18479 7168
rect 16665 7110 18479 7112
rect 16665 7107 16731 7110
rect 18413 7107 18479 7110
rect 3913 7104 4229 7105
rect 3913 7040 3919 7104
rect 3983 7040 3999 7104
rect 4063 7040 4079 7104
rect 4143 7040 4159 7104
rect 4223 7040 4229 7104
rect 3913 7039 4229 7040
rect 9847 7104 10163 7105
rect 9847 7040 9853 7104
rect 9917 7040 9933 7104
rect 9997 7040 10013 7104
rect 10077 7040 10093 7104
rect 10157 7040 10163 7104
rect 9847 7039 10163 7040
rect 15781 7104 16097 7105
rect 15781 7040 15787 7104
rect 15851 7040 15867 7104
rect 15931 7040 15947 7104
rect 16011 7040 16027 7104
rect 16091 7040 16097 7104
rect 15781 7039 16097 7040
rect 21715 7104 22031 7105
rect 21715 7040 21721 7104
rect 21785 7040 21801 7104
rect 21865 7040 21881 7104
rect 21945 7040 21961 7104
rect 22025 7040 22031 7104
rect 21715 7039 22031 7040
rect 0 6898 160 6928
rect 3325 6898 3391 6901
rect 0 6896 3391 6898
rect 0 6840 3330 6896
rect 3386 6840 3391 6896
rect 0 6838 3391 6840
rect 0 6808 160 6838
rect 3325 6835 3391 6838
rect 6729 6898 6795 6901
rect 9581 6898 9647 6901
rect 11881 6898 11947 6901
rect 6729 6896 11947 6898
rect 6729 6840 6734 6896
rect 6790 6840 9586 6896
rect 9642 6840 11886 6896
rect 11942 6840 11947 6896
rect 6729 6838 11947 6840
rect 6729 6835 6795 6838
rect 9581 6835 9647 6838
rect 11881 6835 11947 6838
rect 23473 6898 23539 6901
rect 25840 6898 26000 6928
rect 23473 6896 26000 6898
rect 23473 6840 23478 6896
rect 23534 6840 26000 6896
rect 23473 6838 26000 6840
rect 23473 6835 23539 6838
rect 25840 6808 26000 6838
rect 9029 6762 9095 6765
rect 9765 6762 9831 6765
rect 12249 6762 12315 6765
rect 16481 6762 16547 6765
rect 6686 6702 7482 6762
rect 0 6626 160 6656
rect 2129 6626 2195 6629
rect 0 6624 2195 6626
rect 0 6568 2134 6624
rect 2190 6568 2195 6624
rect 0 6566 2195 6568
rect 0 6536 160 6566
rect 2129 6563 2195 6566
rect 3693 6626 3759 6629
rect 6686 6626 6746 6702
rect 3693 6624 6746 6626
rect 3693 6568 3698 6624
rect 3754 6568 6746 6624
rect 3693 6566 6746 6568
rect 7422 6626 7482 6702
rect 9029 6760 9138 6762
rect 9029 6704 9034 6760
rect 9090 6704 9138 6760
rect 9029 6699 9138 6704
rect 9765 6760 12315 6762
rect 9765 6704 9770 6760
rect 9826 6704 12254 6760
rect 12310 6704 12315 6760
rect 9765 6702 12315 6704
rect 9765 6699 9831 6702
rect 12249 6699 12315 6702
rect 12620 6760 16547 6762
rect 12620 6704 16486 6760
rect 16542 6704 16547 6760
rect 12620 6702 16547 6704
rect 9078 6626 9138 6699
rect 12620 6626 12680 6702
rect 16481 6699 16547 6702
rect 20713 6762 20779 6765
rect 22553 6762 22619 6765
rect 23381 6762 23447 6765
rect 20713 6760 23447 6762
rect 20713 6704 20718 6760
rect 20774 6704 22558 6760
rect 22614 6704 23386 6760
rect 23442 6704 23447 6760
rect 20713 6702 23447 6704
rect 20713 6699 20779 6702
rect 22553 6699 22619 6702
rect 23381 6699 23447 6702
rect 7422 6566 12680 6626
rect 3693 6563 3759 6566
rect 6880 6560 7196 6561
rect 6880 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7196 6560
rect 6880 6495 7196 6496
rect 12814 6560 13130 6561
rect 12814 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13130 6560
rect 12814 6495 13130 6496
rect 18748 6560 19064 6561
rect 18748 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19064 6560
rect 18748 6495 19064 6496
rect 24682 6560 24998 6561
rect 24682 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 24998 6560
rect 24682 6495 24998 6496
rect 3325 6490 3391 6493
rect 4613 6490 4679 6493
rect 3325 6488 4679 6490
rect 3325 6432 3330 6488
rect 3386 6432 4618 6488
rect 4674 6432 4679 6488
rect 3325 6430 4679 6432
rect 3325 6427 3391 6430
rect 4613 6427 4679 6430
rect 0 6354 160 6384
rect 1209 6354 1275 6357
rect 0 6352 1275 6354
rect 0 6296 1214 6352
rect 1270 6296 1275 6352
rect 0 6294 1275 6296
rect 0 6264 160 6294
rect 1209 6291 1275 6294
rect 5441 6354 5507 6357
rect 16297 6354 16363 6357
rect 5441 6352 16363 6354
rect 5441 6296 5446 6352
rect 5502 6296 16302 6352
rect 16358 6296 16363 6352
rect 5441 6294 16363 6296
rect 5441 6291 5507 6294
rect 16297 6291 16363 6294
rect 23197 6354 23263 6357
rect 25840 6354 26000 6384
rect 23197 6352 26000 6354
rect 23197 6296 23202 6352
rect 23258 6296 26000 6352
rect 23197 6294 26000 6296
rect 23197 6291 23263 6294
rect 25840 6264 26000 6294
rect 933 6218 999 6221
rect 3693 6218 3759 6221
rect 933 6216 3759 6218
rect 933 6160 938 6216
rect 994 6160 3698 6216
rect 3754 6160 3759 6216
rect 933 6158 3759 6160
rect 933 6155 999 6158
rect 3693 6155 3759 6158
rect 4613 6218 4679 6221
rect 5257 6218 5323 6221
rect 4613 6216 5323 6218
rect 4613 6160 4618 6216
rect 4674 6160 5262 6216
rect 5318 6160 5323 6216
rect 4613 6158 5323 6160
rect 4613 6155 4679 6158
rect 5257 6155 5323 6158
rect 8569 6218 8635 6221
rect 13261 6218 13327 6221
rect 22645 6218 22711 6221
rect 8569 6216 13327 6218
rect 8569 6160 8574 6216
rect 8630 6160 13266 6216
rect 13322 6160 13327 6216
rect 8569 6158 13327 6160
rect 8569 6155 8635 6158
rect 13261 6155 13327 6158
rect 15518 6216 22711 6218
rect 15518 6160 22650 6216
rect 22706 6160 22711 6216
rect 15518 6158 22711 6160
rect 0 6082 160 6112
rect 1577 6082 1643 6085
rect 0 6080 1643 6082
rect 0 6024 1582 6080
rect 1638 6024 1643 6080
rect 0 6022 1643 6024
rect 0 5992 160 6022
rect 1577 6019 1643 6022
rect 10409 6082 10475 6085
rect 15518 6082 15578 6158
rect 22645 6155 22711 6158
rect 10409 6080 15578 6082
rect 10409 6024 10414 6080
rect 10470 6024 15578 6080
rect 10409 6022 15578 6024
rect 10409 6019 10475 6022
rect 3913 6016 4229 6017
rect 3913 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4229 6016
rect 3913 5951 4229 5952
rect 9847 6016 10163 6017
rect 9847 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10163 6016
rect 9847 5951 10163 5952
rect 15781 6016 16097 6017
rect 15781 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16097 6016
rect 15781 5951 16097 5952
rect 21715 6016 22031 6017
rect 21715 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22031 6016
rect 21715 5951 22031 5952
rect 10869 5946 10935 5949
rect 13813 5946 13879 5949
rect 10869 5944 13879 5946
rect 10869 5888 10874 5944
rect 10930 5888 13818 5944
rect 13874 5888 13879 5944
rect 10869 5886 13879 5888
rect 10869 5883 10935 5886
rect 13813 5883 13879 5886
rect 22326 5886 23628 5946
rect 0 5810 160 5840
rect 2773 5810 2839 5813
rect 0 5808 2839 5810
rect 0 5752 2778 5808
rect 2834 5752 2839 5808
rect 0 5750 2839 5752
rect 0 5720 160 5750
rect 2773 5747 2839 5750
rect 11237 5810 11303 5813
rect 14641 5810 14707 5813
rect 11237 5808 14707 5810
rect 11237 5752 11242 5808
rect 11298 5752 14646 5808
rect 14702 5752 14707 5808
rect 11237 5750 14707 5752
rect 11237 5747 11303 5750
rect 14641 5747 14707 5750
rect 21265 5810 21331 5813
rect 22326 5810 22386 5886
rect 21265 5808 22386 5810
rect 21265 5752 21270 5808
rect 21326 5752 22386 5808
rect 21265 5750 22386 5752
rect 22553 5810 22619 5813
rect 23381 5810 23447 5813
rect 22553 5808 23447 5810
rect 22553 5752 22558 5808
rect 22614 5752 23386 5808
rect 23442 5752 23447 5808
rect 22553 5750 23447 5752
rect 23568 5810 23628 5886
rect 25840 5810 26000 5840
rect 23568 5750 26000 5810
rect 21265 5747 21331 5750
rect 22553 5747 22619 5750
rect 23381 5747 23447 5750
rect 25840 5720 26000 5750
rect 1669 5674 1735 5677
rect 12341 5674 12407 5677
rect 1669 5672 12407 5674
rect 1669 5616 1674 5672
rect 1730 5616 12346 5672
rect 12402 5616 12407 5672
rect 1669 5614 12407 5616
rect 1669 5611 1735 5614
rect 12341 5611 12407 5614
rect 21633 5674 21699 5677
rect 23841 5674 23907 5677
rect 21633 5672 23907 5674
rect 21633 5616 21638 5672
rect 21694 5616 23846 5672
rect 23902 5616 23907 5672
rect 21633 5614 23907 5616
rect 21633 5611 21699 5614
rect 23841 5611 23907 5614
rect 0 5538 160 5568
rect 1117 5538 1183 5541
rect 0 5536 1183 5538
rect 0 5480 1122 5536
rect 1178 5480 1183 5536
rect 0 5478 1183 5480
rect 0 5448 160 5478
rect 1117 5475 1183 5478
rect 2497 5538 2563 5541
rect 2630 5538 2636 5540
rect 2497 5536 2636 5538
rect 2497 5480 2502 5536
rect 2558 5480 2636 5536
rect 2497 5478 2636 5480
rect 2497 5475 2563 5478
rect 2630 5476 2636 5478
rect 2700 5476 2706 5540
rect 20713 5538 20779 5541
rect 22277 5538 22343 5541
rect 20713 5536 22343 5538
rect 20713 5480 20718 5536
rect 20774 5480 22282 5536
rect 22338 5480 22343 5536
rect 20713 5478 22343 5480
rect 20713 5475 20779 5478
rect 22277 5475 22343 5478
rect 22553 5538 22619 5541
rect 22686 5538 22692 5540
rect 22553 5536 22692 5538
rect 22553 5480 22558 5536
rect 22614 5480 22692 5536
rect 22553 5478 22692 5480
rect 22553 5475 22619 5478
rect 22686 5476 22692 5478
rect 22756 5476 22762 5540
rect 6880 5472 7196 5473
rect 6880 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7196 5472
rect 6880 5407 7196 5408
rect 12814 5472 13130 5473
rect 12814 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13130 5472
rect 12814 5407 13130 5408
rect 18748 5472 19064 5473
rect 18748 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19064 5472
rect 18748 5407 19064 5408
rect 24682 5472 24998 5473
rect 24682 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 24998 5472
rect 24682 5407 24998 5408
rect 9581 5402 9647 5405
rect 12617 5402 12683 5405
rect 9581 5400 12683 5402
rect 9581 5344 9586 5400
rect 9642 5344 12622 5400
rect 12678 5344 12683 5400
rect 9581 5342 12683 5344
rect 9581 5339 9647 5342
rect 12617 5339 12683 5342
rect 13261 5404 13327 5405
rect 13261 5400 13308 5404
rect 13372 5402 13378 5404
rect 20713 5402 20779 5405
rect 23565 5402 23631 5405
rect 13261 5344 13266 5400
rect 13261 5340 13308 5344
rect 13372 5342 13418 5402
rect 20713 5400 23631 5402
rect 20713 5344 20718 5400
rect 20774 5344 23570 5400
rect 23626 5344 23631 5400
rect 20713 5342 23631 5344
rect 13372 5340 13378 5342
rect 13261 5339 13327 5340
rect 20713 5339 20779 5342
rect 23565 5339 23631 5342
rect 0 5266 160 5296
rect 0 5206 306 5266
rect 0 5176 160 5206
rect 246 4994 306 5206
rect 11830 5204 11836 5268
rect 11900 5266 11906 5268
rect 13537 5266 13603 5269
rect 11900 5264 13603 5266
rect 11900 5208 13542 5264
rect 13598 5208 13603 5264
rect 11900 5206 13603 5208
rect 11900 5204 11906 5206
rect 13537 5203 13603 5206
rect 14365 5266 14431 5269
rect 14590 5266 14596 5268
rect 14365 5264 14596 5266
rect 14365 5208 14370 5264
rect 14426 5208 14596 5264
rect 14365 5206 14596 5208
rect 14365 5203 14431 5206
rect 14590 5204 14596 5206
rect 14660 5204 14666 5268
rect 19701 5266 19767 5269
rect 21909 5266 21975 5269
rect 19701 5264 21975 5266
rect 19701 5208 19706 5264
rect 19762 5208 21914 5264
rect 21970 5208 21975 5264
rect 19701 5206 21975 5208
rect 19701 5203 19767 5206
rect 21909 5203 21975 5206
rect 22093 5266 22159 5269
rect 25840 5266 26000 5296
rect 22093 5264 26000 5266
rect 22093 5208 22098 5264
rect 22154 5208 26000 5264
rect 22093 5206 26000 5208
rect 22093 5203 22159 5206
rect 25840 5176 26000 5206
rect 8845 5130 8911 5133
rect 23473 5130 23539 5133
rect 8845 5128 23539 5130
rect 8845 5072 8850 5128
rect 8906 5072 23478 5128
rect 23534 5072 23539 5128
rect 8845 5070 23539 5072
rect 8845 5067 8911 5070
rect 23473 5067 23539 5070
rect 62 4934 306 4994
rect 23933 4994 23999 4997
rect 23933 4992 24962 4994
rect 23933 4936 23938 4992
rect 23994 4936 24962 4992
rect 23933 4934 24962 4936
rect 62 4314 122 4934
rect 23933 4931 23999 4934
rect 3913 4928 4229 4929
rect 3913 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4229 4928
rect 3913 4863 4229 4864
rect 9847 4928 10163 4929
rect 9847 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10163 4928
rect 9847 4863 10163 4864
rect 15781 4928 16097 4929
rect 15781 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16097 4928
rect 15781 4863 16097 4864
rect 21715 4928 22031 4929
rect 21715 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22031 4928
rect 21715 4863 22031 4864
rect 2957 4724 3023 4725
rect 2957 4722 3004 4724
rect 2912 4720 3004 4722
rect 3068 4722 3074 4724
rect 4061 4722 4127 4725
rect 3068 4720 4127 4722
rect 2912 4664 2962 4720
rect 3068 4664 4066 4720
rect 4122 4664 4127 4720
rect 2912 4662 3004 4664
rect 2957 4660 3004 4662
rect 3068 4662 4127 4664
rect 3068 4660 3074 4662
rect 2957 4659 3023 4660
rect 4061 4659 4127 4662
rect 10041 4722 10107 4725
rect 11329 4722 11395 4725
rect 12341 4722 12407 4725
rect 10041 4720 12407 4722
rect 10041 4664 10046 4720
rect 10102 4664 11334 4720
rect 11390 4664 12346 4720
rect 12402 4664 12407 4720
rect 10041 4662 12407 4664
rect 24902 4722 24962 4934
rect 25840 4722 26000 4752
rect 24902 4662 26000 4722
rect 10041 4659 10107 4662
rect 11329 4659 11395 4662
rect 12341 4659 12407 4662
rect 25840 4632 26000 4662
rect 3417 4586 3483 4589
rect 9397 4586 9463 4589
rect 3417 4584 9463 4586
rect 3417 4528 3422 4584
rect 3478 4528 9402 4584
rect 9458 4528 9463 4584
rect 3417 4526 9463 4528
rect 3417 4523 3483 4526
rect 9397 4523 9463 4526
rect 16297 4586 16363 4589
rect 22737 4586 22803 4589
rect 16297 4584 22803 4586
rect 16297 4528 16302 4584
rect 16358 4528 22742 4584
rect 22798 4528 22803 4584
rect 16297 4526 22803 4528
rect 16297 4523 16363 4526
rect 22737 4523 22803 4526
rect 20161 4450 20227 4453
rect 20713 4450 20779 4453
rect 20161 4448 20779 4450
rect 20161 4392 20166 4448
rect 20222 4392 20718 4448
rect 20774 4392 20779 4448
rect 20161 4390 20779 4392
rect 20161 4387 20227 4390
rect 20713 4387 20779 4390
rect 21357 4450 21423 4453
rect 21357 4448 22110 4450
rect 21357 4392 21362 4448
rect 21418 4392 22110 4448
rect 21357 4390 22110 4392
rect 21357 4387 21423 4390
rect 6880 4384 7196 4385
rect 6880 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7196 4384
rect 6880 4319 7196 4320
rect 12814 4384 13130 4385
rect 12814 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13130 4384
rect 12814 4319 13130 4320
rect 18748 4384 19064 4385
rect 18748 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19064 4384
rect 18748 4319 19064 4320
rect 1577 4314 1643 4317
rect 62 4312 1643 4314
rect 62 4256 1582 4312
rect 1638 4256 1643 4312
rect 62 4254 1643 4256
rect 1577 4251 1643 4254
rect 19517 4314 19583 4317
rect 21909 4314 21975 4317
rect 19517 4312 21975 4314
rect 19517 4256 19522 4312
rect 19578 4256 21914 4312
rect 21970 4256 21975 4312
rect 19517 4254 21975 4256
rect 19517 4251 19583 4254
rect 21909 4251 21975 4254
rect 12617 4178 12683 4181
rect 13854 4178 13860 4180
rect 4110 4118 4906 4178
rect 2589 4042 2655 4045
rect 4110 4042 4170 4118
rect 2589 4040 4170 4042
rect 2589 3984 2594 4040
rect 2650 3984 4170 4040
rect 2589 3982 4170 3984
rect 2589 3979 2655 3982
rect 4286 3980 4292 4044
rect 4356 4042 4362 4044
rect 4613 4042 4679 4045
rect 4356 4040 4679 4042
rect 4356 3984 4618 4040
rect 4674 3984 4679 4040
rect 4356 3982 4679 3984
rect 4846 4042 4906 4118
rect 12617 4176 13860 4178
rect 12617 4120 12622 4176
rect 12678 4120 13860 4176
rect 12617 4118 13860 4120
rect 12617 4115 12683 4118
rect 13854 4116 13860 4118
rect 13924 4116 13930 4180
rect 19333 4178 19399 4181
rect 19742 4178 19748 4180
rect 19333 4176 19748 4178
rect 19333 4120 19338 4176
rect 19394 4120 19748 4176
rect 19333 4118 19748 4120
rect 19333 4115 19399 4118
rect 19742 4116 19748 4118
rect 19812 4116 19818 4180
rect 22050 4178 22110 4390
rect 24682 4384 24998 4385
rect 24682 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 24998 4384
rect 24682 4319 24998 4320
rect 25840 4178 26000 4208
rect 22050 4118 26000 4178
rect 25840 4088 26000 4118
rect 7649 4042 7715 4045
rect 4846 4040 7715 4042
rect 4846 3984 7654 4040
rect 7710 3984 7715 4040
rect 4846 3982 7715 3984
rect 4356 3980 4362 3982
rect 4613 3979 4679 3982
rect 7649 3979 7715 3982
rect 12157 4044 12223 4045
rect 17677 4044 17743 4045
rect 12157 4040 12204 4044
rect 12268 4042 12274 4044
rect 12157 3984 12162 4040
rect 12157 3980 12204 3984
rect 12268 3982 12314 4042
rect 17677 4040 17724 4044
rect 17788 4042 17794 4044
rect 19885 4042 19951 4045
rect 25313 4042 25379 4045
rect 17677 3984 17682 4040
rect 12268 3980 12274 3982
rect 17677 3980 17724 3984
rect 17788 3982 17834 4042
rect 19885 4040 25379 4042
rect 19885 3984 19890 4040
rect 19946 3984 25318 4040
rect 25374 3984 25379 4040
rect 19885 3982 25379 3984
rect 17788 3980 17794 3982
rect 12157 3979 12223 3980
rect 17677 3979 17743 3980
rect 19885 3979 19951 3982
rect 25313 3979 25379 3982
rect 19517 3908 19583 3909
rect 19517 3906 19564 3908
rect 19472 3904 19564 3906
rect 19472 3848 19522 3904
rect 19472 3846 19564 3848
rect 19517 3844 19564 3846
rect 19628 3844 19634 3908
rect 19701 3906 19767 3909
rect 20437 3906 20503 3909
rect 21173 3908 21239 3909
rect 21449 3908 21515 3909
rect 21173 3906 21220 3908
rect 19701 3904 20503 3906
rect 19701 3848 19706 3904
rect 19762 3848 20442 3904
rect 20498 3848 20503 3904
rect 19701 3846 20503 3848
rect 21128 3904 21220 3906
rect 21128 3848 21178 3904
rect 21128 3846 21220 3848
rect 19517 3843 19583 3844
rect 19701 3843 19767 3846
rect 20437 3843 20503 3846
rect 21173 3844 21220 3846
rect 21284 3844 21290 3908
rect 21398 3844 21404 3908
rect 21468 3906 21515 3908
rect 21468 3904 21560 3906
rect 21510 3848 21560 3904
rect 21468 3846 21560 3848
rect 21468 3844 21515 3846
rect 21173 3843 21239 3844
rect 21449 3843 21515 3844
rect 3913 3840 4229 3841
rect 3913 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4229 3840
rect 3913 3775 4229 3776
rect 9847 3840 10163 3841
rect 9847 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10163 3840
rect 9847 3775 10163 3776
rect 15781 3840 16097 3841
rect 15781 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16097 3840
rect 15781 3775 16097 3776
rect 21715 3840 22031 3841
rect 21715 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22031 3840
rect 21715 3775 22031 3776
rect 19241 3770 19307 3773
rect 21173 3770 21239 3773
rect 19241 3768 21239 3770
rect 19241 3712 19246 3768
rect 19302 3712 21178 3768
rect 21234 3712 21239 3768
rect 19241 3710 21239 3712
rect 19241 3707 19307 3710
rect 21173 3707 21239 3710
rect 1761 3634 1827 3637
rect 20713 3634 20779 3637
rect 1761 3632 20779 3634
rect 1761 3576 1766 3632
rect 1822 3576 20718 3632
rect 20774 3576 20779 3632
rect 1761 3574 20779 3576
rect 1761 3571 1827 3574
rect 20713 3571 20779 3574
rect 23105 3634 23171 3637
rect 25840 3634 26000 3664
rect 23105 3632 26000 3634
rect 23105 3576 23110 3632
rect 23166 3576 26000 3632
rect 23105 3574 26000 3576
rect 23105 3571 23171 3574
rect 25840 3544 26000 3574
rect 2865 3498 2931 3501
rect 9673 3498 9739 3501
rect 2865 3496 9739 3498
rect 2865 3440 2870 3496
rect 2926 3440 9678 3496
rect 9734 3440 9739 3496
rect 2865 3438 9739 3440
rect 2865 3435 2931 3438
rect 9673 3435 9739 3438
rect 10133 3498 10199 3501
rect 10910 3498 10916 3500
rect 10133 3496 10916 3498
rect 10133 3440 10138 3496
rect 10194 3440 10916 3496
rect 10133 3438 10916 3440
rect 10133 3435 10199 3438
rect 10910 3436 10916 3438
rect 10980 3436 10986 3500
rect 17861 3498 17927 3501
rect 22093 3498 22159 3501
rect 17861 3496 22159 3498
rect 17861 3440 17866 3496
rect 17922 3440 22098 3496
rect 22154 3440 22159 3496
rect 17861 3438 22159 3440
rect 17861 3435 17927 3438
rect 22093 3435 22159 3438
rect 790 3300 796 3364
rect 860 3362 866 3364
rect 5533 3362 5599 3365
rect 19517 3362 19583 3365
rect 860 3360 5599 3362
rect 860 3304 5538 3360
rect 5594 3304 5599 3360
rect 860 3302 5599 3304
rect 860 3300 866 3302
rect 5533 3299 5599 3302
rect 19382 3360 19583 3362
rect 19382 3304 19522 3360
rect 19578 3304 19583 3360
rect 19382 3302 19583 3304
rect 6880 3296 7196 3297
rect 6880 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7196 3296
rect 6880 3231 7196 3232
rect 12814 3296 13130 3297
rect 12814 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13130 3296
rect 12814 3231 13130 3232
rect 18748 3296 19064 3297
rect 18748 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19064 3296
rect 18748 3231 19064 3232
rect 8385 3090 8451 3093
rect 11789 3090 11855 3093
rect 8385 3088 11855 3090
rect 8385 3032 8390 3088
rect 8446 3032 11794 3088
rect 11850 3032 11855 3088
rect 8385 3030 11855 3032
rect 8385 3027 8451 3030
rect 11789 3027 11855 3030
rect 4337 2954 4403 2957
rect 9397 2954 9463 2957
rect 4337 2952 9463 2954
rect 4337 2896 4342 2952
rect 4398 2896 9402 2952
rect 9458 2896 9463 2952
rect 4337 2894 9463 2896
rect 4337 2891 4403 2894
rect 9397 2891 9463 2894
rect 19382 2821 19442 3302
rect 19517 3299 19583 3302
rect 24682 3296 24998 3297
rect 24682 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 24998 3296
rect 24682 3231 24998 3232
rect 19517 3090 19583 3093
rect 20529 3090 20595 3093
rect 19517 3088 20595 3090
rect 19517 3032 19522 3088
rect 19578 3032 20534 3088
rect 20590 3032 20595 3088
rect 19517 3030 20595 3032
rect 19517 3027 19583 3030
rect 20529 3027 20595 3030
rect 22369 3090 22435 3093
rect 25840 3090 26000 3120
rect 22369 3088 26000 3090
rect 22369 3032 22374 3088
rect 22430 3032 26000 3088
rect 22369 3030 26000 3032
rect 22369 3027 22435 3030
rect 25840 3000 26000 3030
rect 4797 2818 4863 2821
rect 5901 2818 5967 2821
rect 4797 2816 5967 2818
rect 4797 2760 4802 2816
rect 4858 2760 5906 2816
rect 5962 2760 5967 2816
rect 4797 2758 5967 2760
rect 4797 2755 4863 2758
rect 5901 2755 5967 2758
rect 19333 2816 19442 2821
rect 19333 2760 19338 2816
rect 19394 2760 19442 2816
rect 19333 2758 19442 2760
rect 19333 2755 19399 2758
rect 3913 2752 4229 2753
rect 3913 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4229 2752
rect 3913 2687 4229 2688
rect 9847 2752 10163 2753
rect 9847 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10163 2752
rect 9847 2687 10163 2688
rect 15781 2752 16097 2753
rect 15781 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16097 2752
rect 15781 2687 16097 2688
rect 21715 2752 22031 2753
rect 21715 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22031 2752
rect 21715 2687 22031 2688
rect 9397 2684 9463 2685
rect 11973 2684 12039 2685
rect 14825 2684 14891 2685
rect 9397 2682 9444 2684
rect 9352 2680 9444 2682
rect 9352 2624 9402 2680
rect 9352 2622 9444 2624
rect 9397 2620 9444 2622
rect 9508 2620 9514 2684
rect 11973 2680 12020 2684
rect 12084 2682 12090 2684
rect 14774 2682 14780 2684
rect 11973 2624 11978 2680
rect 11973 2620 12020 2624
rect 12084 2622 12130 2682
rect 14734 2622 14780 2682
rect 14844 2680 14891 2684
rect 14886 2624 14891 2680
rect 12084 2620 12090 2622
rect 14774 2620 14780 2622
rect 14844 2620 14891 2624
rect 9397 2619 9463 2620
rect 11973 2619 12039 2620
rect 14825 2619 14891 2620
rect 15469 2684 15535 2685
rect 17493 2684 17559 2685
rect 15469 2680 15516 2684
rect 15580 2682 15586 2684
rect 15469 2624 15474 2680
rect 15469 2620 15516 2624
rect 15580 2622 15626 2682
rect 17493 2680 17540 2684
rect 17604 2682 17610 2684
rect 17493 2624 17498 2680
rect 15580 2620 15586 2622
rect 17493 2620 17540 2624
rect 17604 2622 17650 2682
rect 17604 2620 17610 2622
rect 18454 2620 18460 2684
rect 18524 2682 18530 2684
rect 18873 2682 18939 2685
rect 19241 2682 19307 2685
rect 18524 2680 18939 2682
rect 18524 2624 18878 2680
rect 18934 2624 18939 2680
rect 18524 2622 18939 2624
rect 18524 2620 18530 2622
rect 15469 2619 15535 2620
rect 17493 2619 17559 2620
rect 18873 2619 18939 2622
rect 19198 2680 19307 2682
rect 19198 2624 19246 2680
rect 19302 2624 19307 2680
rect 19198 2619 19307 2624
rect 19517 2682 19583 2685
rect 19742 2682 19748 2684
rect 19517 2680 19748 2682
rect 19517 2624 19522 2680
rect 19578 2624 19748 2680
rect 19517 2622 19748 2624
rect 19517 2619 19583 2622
rect 19742 2620 19748 2622
rect 19812 2620 19818 2684
rect 5717 2546 5783 2549
rect 5717 2544 9506 2546
rect 5717 2488 5722 2544
rect 5778 2488 9506 2544
rect 5717 2486 9506 2488
rect 5717 2483 5783 2486
rect 4429 2410 4495 2413
rect 9446 2410 9506 2486
rect 9622 2484 9628 2548
rect 9692 2546 9698 2548
rect 9765 2546 9831 2549
rect 13486 2546 13492 2548
rect 9692 2544 9831 2546
rect 9692 2488 9770 2544
rect 9826 2488 9831 2544
rect 9692 2486 9831 2488
rect 9692 2484 9698 2486
rect 9765 2483 9831 2486
rect 9998 2486 13492 2546
rect 9998 2410 10058 2486
rect 13486 2484 13492 2486
rect 13556 2484 13562 2548
rect 14733 2546 14799 2549
rect 16021 2546 16087 2549
rect 16941 2548 17007 2549
rect 16246 2546 16252 2548
rect 14733 2544 15946 2546
rect 14733 2488 14738 2544
rect 14794 2488 15946 2544
rect 14733 2486 15946 2488
rect 14733 2483 14799 2486
rect 4429 2408 9138 2410
rect 4429 2352 4434 2408
rect 4490 2352 9138 2408
rect 4429 2350 9138 2352
rect 9446 2350 10058 2410
rect 10133 2410 10199 2413
rect 10777 2410 10843 2413
rect 13629 2410 13695 2413
rect 10133 2408 10843 2410
rect 10133 2352 10138 2408
rect 10194 2352 10782 2408
rect 10838 2352 10843 2408
rect 10133 2350 10843 2352
rect 4429 2347 4495 2350
rect 3969 2274 4035 2277
rect 7741 2276 7807 2277
rect 8109 2276 8175 2277
rect 8477 2276 8543 2277
rect 8845 2276 8911 2277
rect 5022 2274 5028 2276
rect 3969 2272 5028 2274
rect 3969 2216 3974 2272
rect 4030 2216 5028 2272
rect 3969 2214 5028 2216
rect 3969 2211 4035 2214
rect 5022 2212 5028 2214
rect 5092 2212 5098 2276
rect 7741 2274 7788 2276
rect 7696 2272 7788 2274
rect 7696 2216 7746 2272
rect 7696 2214 7788 2216
rect 7741 2212 7788 2214
rect 7852 2212 7858 2276
rect 8109 2274 8156 2276
rect 8064 2272 8156 2274
rect 8064 2216 8114 2272
rect 8064 2214 8156 2216
rect 8109 2212 8156 2214
rect 8220 2212 8226 2276
rect 8477 2274 8524 2276
rect 8432 2272 8524 2274
rect 8432 2216 8482 2272
rect 8432 2214 8524 2216
rect 8477 2212 8524 2214
rect 8588 2212 8594 2276
rect 8845 2274 8892 2276
rect 8800 2272 8892 2274
rect 8800 2216 8850 2272
rect 8800 2214 8892 2216
rect 8845 2212 8892 2214
rect 8956 2212 8962 2276
rect 9078 2274 9138 2350
rect 10133 2347 10199 2350
rect 10777 2347 10843 2350
rect 11286 2408 13695 2410
rect 11286 2352 13634 2408
rect 13690 2352 13695 2408
rect 11286 2350 13695 2352
rect 15886 2410 15946 2486
rect 16021 2544 16252 2546
rect 16021 2488 16026 2544
rect 16082 2488 16252 2544
rect 16021 2486 16252 2488
rect 16021 2483 16087 2486
rect 16246 2484 16252 2486
rect 16316 2484 16322 2548
rect 16941 2546 16988 2548
rect 16896 2544 16988 2546
rect 16896 2488 16946 2544
rect 16896 2486 16988 2488
rect 16941 2484 16988 2486
rect 17052 2484 17058 2548
rect 18505 2546 18571 2549
rect 19198 2546 19258 2619
rect 18505 2544 19258 2546
rect 18505 2488 18510 2544
rect 18566 2488 19258 2544
rect 18505 2486 19258 2488
rect 16941 2483 17007 2484
rect 18505 2483 18571 2486
rect 21582 2484 21588 2548
rect 21652 2546 21658 2548
rect 21909 2546 21975 2549
rect 21652 2544 21975 2546
rect 21652 2488 21914 2544
rect 21970 2488 21975 2544
rect 21652 2486 21975 2488
rect 21652 2484 21658 2486
rect 21909 2483 21975 2486
rect 24025 2546 24091 2549
rect 25840 2546 26000 2576
rect 24025 2544 26000 2546
rect 24025 2488 24030 2544
rect 24086 2488 26000 2544
rect 24025 2486 26000 2488
rect 24025 2483 24091 2486
rect 25840 2456 26000 2486
rect 19609 2412 19675 2413
rect 19374 2410 19380 2412
rect 15886 2350 19380 2410
rect 11286 2274 11346 2350
rect 13629 2347 13695 2350
rect 19374 2348 19380 2350
rect 19444 2348 19450 2412
rect 19558 2348 19564 2412
rect 19628 2410 19675 2412
rect 20069 2410 20135 2413
rect 20805 2410 20871 2413
rect 19628 2408 19720 2410
rect 19670 2352 19720 2408
rect 19628 2350 19720 2352
rect 20069 2408 20871 2410
rect 20069 2352 20074 2408
rect 20130 2352 20810 2408
rect 20866 2352 20871 2408
rect 20069 2350 20871 2352
rect 19628 2348 19675 2350
rect 19609 2347 19675 2348
rect 20069 2347 20135 2350
rect 20805 2347 20871 2350
rect 9078 2214 11346 2274
rect 7741 2211 7807 2212
rect 8109 2211 8175 2212
rect 8477 2211 8543 2212
rect 8845 2211 8911 2212
rect 6880 2208 7196 2209
rect 6880 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7196 2208
rect 6880 2143 7196 2144
rect 12814 2208 13130 2209
rect 12814 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13130 2208
rect 12814 2143 13130 2144
rect 18748 2208 19064 2209
rect 18748 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19064 2208
rect 18748 2143 19064 2144
rect 24682 2208 24998 2209
rect 24682 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 24998 2208
rect 24682 2143 24998 2144
rect 2730 2078 5826 2138
rect 1158 1940 1164 2004
rect 1228 2002 1234 2004
rect 2730 2002 2790 2078
rect 1228 1942 2790 2002
rect 5533 2004 5599 2005
rect 5533 2000 5580 2004
rect 5644 2002 5650 2004
rect 5766 2002 5826 2078
rect 5993 2002 6059 2005
rect 5533 1944 5538 2000
rect 1228 1940 1234 1942
rect 5533 1940 5580 1944
rect 5644 1942 5690 2002
rect 5766 2000 6059 2002
rect 5766 1944 5998 2000
rect 6054 1944 6059 2000
rect 5766 1942 6059 1944
rect 5644 1940 5650 1942
rect 5533 1939 5599 1940
rect 5993 1939 6059 1942
rect 6310 1940 6316 2004
rect 6380 2002 6386 2004
rect 7005 2002 7071 2005
rect 6380 2000 7071 2002
rect 6380 1944 7010 2000
rect 7066 1944 7071 2000
rect 6380 1942 7071 1944
rect 6380 1940 6386 1942
rect 7005 1939 7071 1942
rect 13721 2002 13787 2005
rect 21173 2002 21239 2005
rect 25840 2002 26000 2032
rect 13721 2000 14474 2002
rect 13721 1944 13726 2000
rect 13782 1944 14474 2000
rect 13721 1942 14474 1944
rect 13721 1939 13787 1942
rect 13 1866 79 1869
rect 14273 1866 14339 1869
rect 13 1864 14339 1866
rect 13 1808 18 1864
rect 74 1808 14278 1864
rect 14334 1808 14339 1864
rect 13 1806 14339 1808
rect 14414 1866 14474 1942
rect 21173 2000 26000 2002
rect 21173 1944 21178 2000
rect 21234 1944 26000 2000
rect 21173 1942 26000 1944
rect 21173 1939 21239 1942
rect 25840 1912 26000 1942
rect 25405 1866 25471 1869
rect 14414 1864 25471 1866
rect 14414 1808 25410 1864
rect 25466 1808 25471 1864
rect 14414 1806 25471 1808
rect 13 1803 79 1806
rect 14273 1803 14339 1806
rect 25405 1803 25471 1806
rect 4429 1730 4495 1733
rect 9397 1730 9463 1733
rect 4429 1728 9463 1730
rect 4429 1672 4434 1728
rect 4490 1672 9402 1728
rect 9458 1672 9463 1728
rect 4429 1670 9463 1672
rect 4429 1667 4495 1670
rect 9397 1667 9463 1670
rect 3913 1664 4229 1665
rect 3913 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4229 1664
rect 3913 1599 4229 1600
rect 9847 1664 10163 1665
rect 9847 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10163 1664
rect 9847 1599 10163 1600
rect 15781 1664 16097 1665
rect 15781 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16097 1664
rect 15781 1599 16097 1600
rect 21715 1664 22031 1665
rect 21715 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22031 1664
rect 21715 1599 22031 1600
rect 4797 1594 4863 1597
rect 6913 1594 6979 1597
rect 4797 1592 6979 1594
rect 4797 1536 4802 1592
rect 4858 1536 6918 1592
rect 6974 1536 6979 1592
rect 4797 1534 6979 1536
rect 4797 1531 4863 1534
rect 6913 1531 6979 1534
rect 381 1458 447 1461
rect 9121 1458 9187 1461
rect 381 1456 9187 1458
rect 381 1400 386 1456
rect 442 1400 9126 1456
rect 9182 1400 9187 1456
rect 381 1398 9187 1400
rect 381 1395 447 1398
rect 9121 1395 9187 1398
rect 22553 1458 22619 1461
rect 25840 1458 26000 1488
rect 22553 1456 26000 1458
rect 22553 1400 22558 1456
rect 22614 1400 26000 1456
rect 22553 1398 26000 1400
rect 22553 1395 22619 1398
rect 25840 1368 26000 1398
rect 1669 1324 1735 1325
rect 2037 1324 2103 1325
rect 4429 1324 4495 1325
rect 1669 1322 1716 1324
rect 1624 1320 1716 1322
rect 1624 1264 1674 1320
rect 1624 1262 1716 1264
rect 1669 1260 1716 1262
rect 1780 1260 1786 1324
rect 2037 1322 2084 1324
rect 1992 1320 2084 1322
rect 1992 1264 2042 1320
rect 1992 1262 2084 1264
rect 2037 1260 2084 1262
rect 2148 1260 2154 1324
rect 4429 1320 4476 1324
rect 4540 1322 4546 1324
rect 6913 1322 6979 1325
rect 16481 1324 16547 1325
rect 16430 1322 16436 1324
rect 4429 1264 4434 1320
rect 4429 1260 4476 1264
rect 4540 1262 4586 1322
rect 5030 1320 6979 1322
rect 5030 1264 6918 1320
rect 6974 1264 6979 1320
rect 5030 1262 6979 1264
rect 16390 1262 16436 1322
rect 16500 1320 16547 1324
rect 16542 1264 16547 1320
rect 4540 1260 4546 1262
rect 1669 1259 1735 1260
rect 2037 1259 2103 1260
rect 4429 1259 4495 1260
rect 974 1124 980 1188
rect 1044 1186 1050 1188
rect 5030 1186 5090 1262
rect 6913 1259 6979 1262
rect 16430 1260 16436 1262
rect 16500 1260 16547 1264
rect 18086 1260 18092 1324
rect 18156 1322 18162 1324
rect 18505 1322 18571 1325
rect 18156 1320 18571 1322
rect 18156 1264 18510 1320
rect 18566 1264 18571 1320
rect 18156 1262 18571 1264
rect 18156 1260 18162 1262
rect 16481 1259 16547 1260
rect 18505 1259 18571 1262
rect 19926 1260 19932 1324
rect 19996 1322 20002 1324
rect 20989 1322 21055 1325
rect 19996 1320 21055 1322
rect 19996 1264 20994 1320
rect 21050 1264 21055 1320
rect 19996 1262 21055 1264
rect 19996 1260 20002 1262
rect 20989 1259 21055 1262
rect 1044 1126 5090 1186
rect 1044 1124 1050 1126
rect 6880 1120 7196 1121
rect 6880 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7196 1120
rect 6880 1055 7196 1056
rect 12814 1120 13130 1121
rect 12814 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13130 1120
rect 12814 1055 13130 1056
rect 18748 1120 19064 1121
rect 18748 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19064 1120
rect 18748 1055 19064 1056
rect 24682 1120 24998 1121
rect 24682 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 24998 1120
rect 24682 1055 24998 1056
rect 7925 914 7991 917
rect 17902 914 17908 916
rect 7925 912 17908 914
rect 7925 856 7930 912
rect 7986 856 17908 912
rect 7925 854 17908 856
rect 7925 851 7991 854
rect 17902 852 17908 854
rect 17972 852 17978 916
rect 21081 914 21147 917
rect 25840 914 26000 944
rect 21081 912 26000 914
rect 21081 856 21086 912
rect 21142 856 26000 912
rect 21081 854 26000 856
rect 21081 851 21147 854
rect 25840 824 26000 854
rect 6085 778 6151 781
rect 8702 778 8708 780
rect 6085 776 8708 778
rect 6085 720 6090 776
rect 6146 720 8708 776
rect 6085 718 8708 720
rect 6085 715 6151 718
rect 8702 716 8708 718
rect 8772 716 8778 780
<< via3 >>
rect 6886 43548 6950 43552
rect 6886 43492 6890 43548
rect 6890 43492 6946 43548
rect 6946 43492 6950 43548
rect 6886 43488 6950 43492
rect 6966 43548 7030 43552
rect 6966 43492 6970 43548
rect 6970 43492 7026 43548
rect 7026 43492 7030 43548
rect 6966 43488 7030 43492
rect 7046 43548 7110 43552
rect 7046 43492 7050 43548
rect 7050 43492 7106 43548
rect 7106 43492 7110 43548
rect 7046 43488 7110 43492
rect 7126 43548 7190 43552
rect 7126 43492 7130 43548
rect 7130 43492 7186 43548
rect 7186 43492 7190 43548
rect 7126 43488 7190 43492
rect 12820 43548 12884 43552
rect 12820 43492 12824 43548
rect 12824 43492 12880 43548
rect 12880 43492 12884 43548
rect 12820 43488 12884 43492
rect 12900 43548 12964 43552
rect 12900 43492 12904 43548
rect 12904 43492 12960 43548
rect 12960 43492 12964 43548
rect 12900 43488 12964 43492
rect 12980 43548 13044 43552
rect 12980 43492 12984 43548
rect 12984 43492 13040 43548
rect 13040 43492 13044 43548
rect 12980 43488 13044 43492
rect 13060 43548 13124 43552
rect 13060 43492 13064 43548
rect 13064 43492 13120 43548
rect 13120 43492 13124 43548
rect 13060 43488 13124 43492
rect 18754 43548 18818 43552
rect 18754 43492 18758 43548
rect 18758 43492 18814 43548
rect 18814 43492 18818 43548
rect 18754 43488 18818 43492
rect 18834 43548 18898 43552
rect 18834 43492 18838 43548
rect 18838 43492 18894 43548
rect 18894 43492 18898 43548
rect 18834 43488 18898 43492
rect 18914 43548 18978 43552
rect 18914 43492 18918 43548
rect 18918 43492 18974 43548
rect 18974 43492 18978 43548
rect 18914 43488 18978 43492
rect 18994 43548 19058 43552
rect 18994 43492 18998 43548
rect 18998 43492 19054 43548
rect 19054 43492 19058 43548
rect 18994 43488 19058 43492
rect 24688 43548 24752 43552
rect 24688 43492 24692 43548
rect 24692 43492 24748 43548
rect 24748 43492 24752 43548
rect 24688 43488 24752 43492
rect 24768 43548 24832 43552
rect 24768 43492 24772 43548
rect 24772 43492 24828 43548
rect 24828 43492 24832 43548
rect 24768 43488 24832 43492
rect 24848 43548 24912 43552
rect 24848 43492 24852 43548
rect 24852 43492 24908 43548
rect 24908 43492 24912 43548
rect 24848 43488 24912 43492
rect 24928 43548 24992 43552
rect 24928 43492 24932 43548
rect 24932 43492 24988 43548
rect 24988 43492 24992 43548
rect 24928 43488 24992 43492
rect 20668 43148 20732 43212
rect 11468 43012 11532 43076
rect 13676 43012 13740 43076
rect 3919 43004 3983 43008
rect 3919 42948 3923 43004
rect 3923 42948 3979 43004
rect 3979 42948 3983 43004
rect 3919 42944 3983 42948
rect 3999 43004 4063 43008
rect 3999 42948 4003 43004
rect 4003 42948 4059 43004
rect 4059 42948 4063 43004
rect 3999 42944 4063 42948
rect 4079 43004 4143 43008
rect 4079 42948 4083 43004
rect 4083 42948 4139 43004
rect 4139 42948 4143 43004
rect 4079 42944 4143 42948
rect 4159 43004 4223 43008
rect 4159 42948 4163 43004
rect 4163 42948 4219 43004
rect 4219 42948 4223 43004
rect 4159 42944 4223 42948
rect 9853 43004 9917 43008
rect 9853 42948 9857 43004
rect 9857 42948 9913 43004
rect 9913 42948 9917 43004
rect 9853 42944 9917 42948
rect 9933 43004 9997 43008
rect 9933 42948 9937 43004
rect 9937 42948 9993 43004
rect 9993 42948 9997 43004
rect 9933 42944 9997 42948
rect 10013 43004 10077 43008
rect 10013 42948 10017 43004
rect 10017 42948 10073 43004
rect 10073 42948 10077 43004
rect 10013 42944 10077 42948
rect 10093 43004 10157 43008
rect 10093 42948 10097 43004
rect 10097 42948 10153 43004
rect 10153 42948 10157 43004
rect 10093 42944 10157 42948
rect 15787 43004 15851 43008
rect 15787 42948 15791 43004
rect 15791 42948 15847 43004
rect 15847 42948 15851 43004
rect 15787 42944 15851 42948
rect 15867 43004 15931 43008
rect 15867 42948 15871 43004
rect 15871 42948 15927 43004
rect 15927 42948 15931 43004
rect 15867 42944 15931 42948
rect 15947 43004 16011 43008
rect 15947 42948 15951 43004
rect 15951 42948 16007 43004
rect 16007 42948 16011 43004
rect 15947 42944 16011 42948
rect 16027 43004 16091 43008
rect 16027 42948 16031 43004
rect 16031 42948 16087 43004
rect 16087 42948 16091 43004
rect 16027 42944 16091 42948
rect 21721 43004 21785 43008
rect 21721 42948 21725 43004
rect 21725 42948 21781 43004
rect 21781 42948 21785 43004
rect 21721 42944 21785 42948
rect 21801 43004 21865 43008
rect 21801 42948 21805 43004
rect 21805 42948 21861 43004
rect 21861 42948 21865 43004
rect 21801 42944 21865 42948
rect 21881 43004 21945 43008
rect 21881 42948 21885 43004
rect 21885 42948 21941 43004
rect 21941 42948 21945 43004
rect 21881 42944 21945 42948
rect 21961 43004 22025 43008
rect 21961 42948 21965 43004
rect 21965 42948 22021 43004
rect 22021 42948 22025 43004
rect 21961 42944 22025 42948
rect 11652 42876 11716 42940
rect 12204 42936 12268 42940
rect 12204 42880 12254 42936
rect 12254 42880 12268 42936
rect 12204 42876 12268 42880
rect 13308 42876 13372 42940
rect 14412 42876 14476 42940
rect 14964 42936 15028 42940
rect 14964 42880 14978 42936
rect 14978 42880 15028 42936
rect 14964 42876 15028 42880
rect 15332 42936 15396 42940
rect 15332 42880 15346 42936
rect 15346 42880 15396 42936
rect 15332 42876 15396 42880
rect 6886 42460 6950 42464
rect 6886 42404 6890 42460
rect 6890 42404 6946 42460
rect 6946 42404 6950 42460
rect 6886 42400 6950 42404
rect 6966 42460 7030 42464
rect 6966 42404 6970 42460
rect 6970 42404 7026 42460
rect 7026 42404 7030 42460
rect 6966 42400 7030 42404
rect 7046 42460 7110 42464
rect 7046 42404 7050 42460
rect 7050 42404 7106 42460
rect 7106 42404 7110 42460
rect 7046 42400 7110 42404
rect 7126 42460 7190 42464
rect 7126 42404 7130 42460
rect 7130 42404 7186 42460
rect 7186 42404 7190 42460
rect 7126 42400 7190 42404
rect 12820 42460 12884 42464
rect 12820 42404 12824 42460
rect 12824 42404 12880 42460
rect 12880 42404 12884 42460
rect 12820 42400 12884 42404
rect 12900 42460 12964 42464
rect 12900 42404 12904 42460
rect 12904 42404 12960 42460
rect 12960 42404 12964 42460
rect 12900 42400 12964 42404
rect 12980 42460 13044 42464
rect 12980 42404 12984 42460
rect 12984 42404 13040 42460
rect 13040 42404 13044 42460
rect 12980 42400 13044 42404
rect 13060 42460 13124 42464
rect 13060 42404 13064 42460
rect 13064 42404 13120 42460
rect 13120 42404 13124 42460
rect 13060 42400 13124 42404
rect 18754 42460 18818 42464
rect 18754 42404 18758 42460
rect 18758 42404 18814 42460
rect 18814 42404 18818 42460
rect 18754 42400 18818 42404
rect 18834 42460 18898 42464
rect 18834 42404 18838 42460
rect 18838 42404 18894 42460
rect 18894 42404 18898 42460
rect 18834 42400 18898 42404
rect 18914 42460 18978 42464
rect 18914 42404 18918 42460
rect 18918 42404 18974 42460
rect 18974 42404 18978 42460
rect 18914 42400 18978 42404
rect 18994 42460 19058 42464
rect 18994 42404 18998 42460
rect 18998 42404 19054 42460
rect 19054 42404 19058 42460
rect 18994 42400 19058 42404
rect 24688 42460 24752 42464
rect 24688 42404 24692 42460
rect 24692 42404 24748 42460
rect 24748 42404 24752 42460
rect 24688 42400 24752 42404
rect 24768 42460 24832 42464
rect 24768 42404 24772 42460
rect 24772 42404 24828 42460
rect 24828 42404 24832 42460
rect 24768 42400 24832 42404
rect 24848 42460 24912 42464
rect 24848 42404 24852 42460
rect 24852 42404 24908 42460
rect 24908 42404 24912 42460
rect 24848 42400 24912 42404
rect 24928 42460 24992 42464
rect 24928 42404 24932 42460
rect 24932 42404 24988 42460
rect 24988 42404 24992 42460
rect 24928 42400 24992 42404
rect 3919 41916 3983 41920
rect 3919 41860 3923 41916
rect 3923 41860 3979 41916
rect 3979 41860 3983 41916
rect 3919 41856 3983 41860
rect 3999 41916 4063 41920
rect 3999 41860 4003 41916
rect 4003 41860 4059 41916
rect 4059 41860 4063 41916
rect 3999 41856 4063 41860
rect 4079 41916 4143 41920
rect 4079 41860 4083 41916
rect 4083 41860 4139 41916
rect 4139 41860 4143 41916
rect 4079 41856 4143 41860
rect 4159 41916 4223 41920
rect 4159 41860 4163 41916
rect 4163 41860 4219 41916
rect 4219 41860 4223 41916
rect 4159 41856 4223 41860
rect 6316 41788 6380 41852
rect 6500 41788 6564 41852
rect 8156 42120 8220 42124
rect 8156 42064 8170 42120
rect 8170 42064 8220 42120
rect 8156 42060 8220 42064
rect 21036 42060 21100 42124
rect 9853 41916 9917 41920
rect 9853 41860 9857 41916
rect 9857 41860 9913 41916
rect 9913 41860 9917 41916
rect 9853 41856 9917 41860
rect 9933 41916 9997 41920
rect 9933 41860 9937 41916
rect 9937 41860 9993 41916
rect 9993 41860 9997 41916
rect 9933 41856 9997 41860
rect 10013 41916 10077 41920
rect 10013 41860 10017 41916
rect 10017 41860 10073 41916
rect 10073 41860 10077 41916
rect 10013 41856 10077 41860
rect 10093 41916 10157 41920
rect 10093 41860 10097 41916
rect 10097 41860 10153 41916
rect 10153 41860 10157 41916
rect 10093 41856 10157 41860
rect 15787 41916 15851 41920
rect 15787 41860 15791 41916
rect 15791 41860 15847 41916
rect 15847 41860 15851 41916
rect 15787 41856 15851 41860
rect 15867 41916 15931 41920
rect 15867 41860 15871 41916
rect 15871 41860 15927 41916
rect 15927 41860 15931 41916
rect 15867 41856 15931 41860
rect 15947 41916 16011 41920
rect 15947 41860 15951 41916
rect 15951 41860 16007 41916
rect 16007 41860 16011 41916
rect 15947 41856 16011 41860
rect 16027 41916 16091 41920
rect 16027 41860 16031 41916
rect 16031 41860 16087 41916
rect 16087 41860 16091 41916
rect 16027 41856 16091 41860
rect 7972 41788 8036 41852
rect 14596 41652 14660 41716
rect 21721 41916 21785 41920
rect 21721 41860 21725 41916
rect 21725 41860 21781 41916
rect 21781 41860 21785 41916
rect 21721 41856 21785 41860
rect 21801 41916 21865 41920
rect 21801 41860 21805 41916
rect 21805 41860 21861 41916
rect 21861 41860 21865 41916
rect 21801 41856 21865 41860
rect 21881 41916 21945 41920
rect 21881 41860 21885 41916
rect 21885 41860 21941 41916
rect 21941 41860 21945 41916
rect 21881 41856 21945 41860
rect 21961 41916 22025 41920
rect 21961 41860 21965 41916
rect 21965 41860 22021 41916
rect 22021 41860 22025 41916
rect 21961 41856 22025 41860
rect 17724 41788 17788 41852
rect 18276 41788 18340 41852
rect 17540 41712 17604 41716
rect 17540 41656 17590 41712
rect 17590 41656 17604 41712
rect 17540 41652 17604 41656
rect 1164 41516 1228 41580
rect 4844 41516 4908 41580
rect 14780 41516 14844 41580
rect 19196 41516 19260 41580
rect 9260 41380 9324 41444
rect 16252 41440 16316 41444
rect 16252 41384 16266 41440
rect 16266 41384 16316 41440
rect 16252 41380 16316 41384
rect 6886 41372 6950 41376
rect 6886 41316 6890 41372
rect 6890 41316 6946 41372
rect 6946 41316 6950 41372
rect 6886 41312 6950 41316
rect 6966 41372 7030 41376
rect 6966 41316 6970 41372
rect 6970 41316 7026 41372
rect 7026 41316 7030 41372
rect 6966 41312 7030 41316
rect 7046 41372 7110 41376
rect 7046 41316 7050 41372
rect 7050 41316 7106 41372
rect 7106 41316 7110 41372
rect 7046 41312 7110 41316
rect 7126 41372 7190 41376
rect 7126 41316 7130 41372
rect 7130 41316 7186 41372
rect 7186 41316 7190 41372
rect 7126 41312 7190 41316
rect 12820 41372 12884 41376
rect 12820 41316 12824 41372
rect 12824 41316 12880 41372
rect 12880 41316 12884 41372
rect 12820 41312 12884 41316
rect 12900 41372 12964 41376
rect 12900 41316 12904 41372
rect 12904 41316 12960 41372
rect 12960 41316 12964 41372
rect 12900 41312 12964 41316
rect 12980 41372 13044 41376
rect 12980 41316 12984 41372
rect 12984 41316 13040 41372
rect 13040 41316 13044 41372
rect 12980 41312 13044 41316
rect 13060 41372 13124 41376
rect 13060 41316 13064 41372
rect 13064 41316 13120 41372
rect 13120 41316 13124 41372
rect 13060 41312 13124 41316
rect 18754 41372 18818 41376
rect 18754 41316 18758 41372
rect 18758 41316 18814 41372
rect 18814 41316 18818 41372
rect 18754 41312 18818 41316
rect 18834 41372 18898 41376
rect 18834 41316 18838 41372
rect 18838 41316 18894 41372
rect 18894 41316 18898 41372
rect 18834 41312 18898 41316
rect 18914 41372 18978 41376
rect 18914 41316 18918 41372
rect 18918 41316 18974 41372
rect 18974 41316 18978 41372
rect 18914 41312 18978 41316
rect 18994 41372 19058 41376
rect 18994 41316 18998 41372
rect 18998 41316 19054 41372
rect 19054 41316 19058 41372
rect 18994 41312 19058 41316
rect 24688 41372 24752 41376
rect 24688 41316 24692 41372
rect 24692 41316 24748 41372
rect 24748 41316 24752 41372
rect 24688 41312 24752 41316
rect 24768 41372 24832 41376
rect 24768 41316 24772 41372
rect 24772 41316 24828 41372
rect 24828 41316 24832 41372
rect 24768 41312 24832 41316
rect 24848 41372 24912 41376
rect 24848 41316 24852 41372
rect 24852 41316 24908 41372
rect 24908 41316 24912 41372
rect 24848 41312 24912 41316
rect 24928 41372 24992 41376
rect 24928 41316 24932 41372
rect 24932 41316 24988 41372
rect 24988 41316 24992 41372
rect 24928 41312 24992 41316
rect 13492 40972 13556 41036
rect 3919 40828 3983 40832
rect 3919 40772 3923 40828
rect 3923 40772 3979 40828
rect 3979 40772 3983 40828
rect 3919 40768 3983 40772
rect 3999 40828 4063 40832
rect 3999 40772 4003 40828
rect 4003 40772 4059 40828
rect 4059 40772 4063 40828
rect 3999 40768 4063 40772
rect 4079 40828 4143 40832
rect 4079 40772 4083 40828
rect 4083 40772 4139 40828
rect 4139 40772 4143 40828
rect 4079 40768 4143 40772
rect 4159 40828 4223 40832
rect 4159 40772 4163 40828
rect 4163 40772 4219 40828
rect 4219 40772 4223 40828
rect 4159 40768 4223 40772
rect 9853 40828 9917 40832
rect 9853 40772 9857 40828
rect 9857 40772 9913 40828
rect 9913 40772 9917 40828
rect 9853 40768 9917 40772
rect 9933 40828 9997 40832
rect 9933 40772 9937 40828
rect 9937 40772 9993 40828
rect 9993 40772 9997 40828
rect 9933 40768 9997 40772
rect 10013 40828 10077 40832
rect 10013 40772 10017 40828
rect 10017 40772 10073 40828
rect 10073 40772 10077 40828
rect 10013 40768 10077 40772
rect 10093 40828 10157 40832
rect 10093 40772 10097 40828
rect 10097 40772 10153 40828
rect 10153 40772 10157 40828
rect 10093 40768 10157 40772
rect 15787 40828 15851 40832
rect 15787 40772 15791 40828
rect 15791 40772 15847 40828
rect 15847 40772 15851 40828
rect 15787 40768 15851 40772
rect 15867 40828 15931 40832
rect 15867 40772 15871 40828
rect 15871 40772 15927 40828
rect 15927 40772 15931 40828
rect 15867 40768 15931 40772
rect 15947 40828 16011 40832
rect 15947 40772 15951 40828
rect 15951 40772 16007 40828
rect 16007 40772 16011 40828
rect 15947 40768 16011 40772
rect 16027 40828 16091 40832
rect 16027 40772 16031 40828
rect 16031 40772 16087 40828
rect 16087 40772 16091 40828
rect 16027 40768 16091 40772
rect 21721 40828 21785 40832
rect 21721 40772 21725 40828
rect 21725 40772 21781 40828
rect 21781 40772 21785 40828
rect 21721 40768 21785 40772
rect 21801 40828 21865 40832
rect 21801 40772 21805 40828
rect 21805 40772 21861 40828
rect 21861 40772 21865 40828
rect 21801 40768 21865 40772
rect 21881 40828 21945 40832
rect 21881 40772 21885 40828
rect 21885 40772 21941 40828
rect 21941 40772 21945 40828
rect 21881 40768 21945 40772
rect 21961 40828 22025 40832
rect 21961 40772 21965 40828
rect 21965 40772 22021 40828
rect 22021 40772 22025 40828
rect 21961 40768 22025 40772
rect 20668 40564 20732 40628
rect 2084 40428 2148 40492
rect 1716 40292 1780 40356
rect 6886 40284 6950 40288
rect 6886 40228 6890 40284
rect 6890 40228 6946 40284
rect 6946 40228 6950 40284
rect 6886 40224 6950 40228
rect 6966 40284 7030 40288
rect 6966 40228 6970 40284
rect 6970 40228 7026 40284
rect 7026 40228 7030 40284
rect 6966 40224 7030 40228
rect 7046 40284 7110 40288
rect 7046 40228 7050 40284
rect 7050 40228 7106 40284
rect 7106 40228 7110 40284
rect 7046 40224 7110 40228
rect 7126 40284 7190 40288
rect 7126 40228 7130 40284
rect 7130 40228 7186 40284
rect 7186 40228 7190 40284
rect 7126 40224 7190 40228
rect 12820 40284 12884 40288
rect 12820 40228 12824 40284
rect 12824 40228 12880 40284
rect 12880 40228 12884 40284
rect 12820 40224 12884 40228
rect 12900 40284 12964 40288
rect 12900 40228 12904 40284
rect 12904 40228 12960 40284
rect 12960 40228 12964 40284
rect 12900 40224 12964 40228
rect 12980 40284 13044 40288
rect 12980 40228 12984 40284
rect 12984 40228 13040 40284
rect 13040 40228 13044 40284
rect 12980 40224 13044 40228
rect 13060 40284 13124 40288
rect 13060 40228 13064 40284
rect 13064 40228 13120 40284
rect 13120 40228 13124 40284
rect 13060 40224 13124 40228
rect 18754 40284 18818 40288
rect 18754 40228 18758 40284
rect 18758 40228 18814 40284
rect 18814 40228 18818 40284
rect 18754 40224 18818 40228
rect 18834 40284 18898 40288
rect 18834 40228 18838 40284
rect 18838 40228 18894 40284
rect 18894 40228 18898 40284
rect 18834 40224 18898 40228
rect 18914 40284 18978 40288
rect 18914 40228 18918 40284
rect 18918 40228 18974 40284
rect 18974 40228 18978 40284
rect 18914 40224 18978 40228
rect 18994 40284 19058 40288
rect 18994 40228 18998 40284
rect 18998 40228 19054 40284
rect 19054 40228 19058 40284
rect 18994 40224 19058 40228
rect 7788 40020 7852 40084
rect 9628 40080 9692 40084
rect 9628 40024 9678 40080
rect 9678 40024 9692 40080
rect 9628 40020 9692 40024
rect 24688 40284 24752 40288
rect 24688 40228 24692 40284
rect 24692 40228 24748 40284
rect 24748 40228 24752 40284
rect 24688 40224 24752 40228
rect 24768 40284 24832 40288
rect 24768 40228 24772 40284
rect 24772 40228 24828 40284
rect 24828 40228 24832 40284
rect 24768 40224 24832 40228
rect 24848 40284 24912 40288
rect 24848 40228 24852 40284
rect 24852 40228 24908 40284
rect 24908 40228 24912 40284
rect 24848 40224 24912 40228
rect 24928 40284 24992 40288
rect 24928 40228 24932 40284
rect 24932 40228 24988 40284
rect 24988 40228 24992 40284
rect 24928 40224 24992 40228
rect 19564 40020 19628 40084
rect 10548 39884 10612 39948
rect 3919 39740 3983 39744
rect 3919 39684 3923 39740
rect 3923 39684 3979 39740
rect 3979 39684 3983 39740
rect 3919 39680 3983 39684
rect 3999 39740 4063 39744
rect 3999 39684 4003 39740
rect 4003 39684 4059 39740
rect 4059 39684 4063 39740
rect 3999 39680 4063 39684
rect 4079 39740 4143 39744
rect 4079 39684 4083 39740
rect 4083 39684 4139 39740
rect 4139 39684 4143 39740
rect 4079 39680 4143 39684
rect 4159 39740 4223 39744
rect 4159 39684 4163 39740
rect 4163 39684 4219 39740
rect 4219 39684 4223 39740
rect 4159 39680 4223 39684
rect 9853 39740 9917 39744
rect 9853 39684 9857 39740
rect 9857 39684 9913 39740
rect 9913 39684 9917 39740
rect 9853 39680 9917 39684
rect 9933 39740 9997 39744
rect 9933 39684 9937 39740
rect 9937 39684 9993 39740
rect 9993 39684 9997 39740
rect 9933 39680 9997 39684
rect 10013 39740 10077 39744
rect 10013 39684 10017 39740
rect 10017 39684 10073 39740
rect 10073 39684 10077 39740
rect 10013 39680 10077 39684
rect 10093 39740 10157 39744
rect 10093 39684 10097 39740
rect 10097 39684 10153 39740
rect 10153 39684 10157 39740
rect 10093 39680 10157 39684
rect 15787 39740 15851 39744
rect 15787 39684 15791 39740
rect 15791 39684 15847 39740
rect 15847 39684 15851 39740
rect 15787 39680 15851 39684
rect 15867 39740 15931 39744
rect 15867 39684 15871 39740
rect 15871 39684 15927 39740
rect 15927 39684 15931 39740
rect 15867 39680 15931 39684
rect 15947 39740 16011 39744
rect 15947 39684 15951 39740
rect 15951 39684 16007 39740
rect 16007 39684 16011 39740
rect 15947 39680 16011 39684
rect 16027 39740 16091 39744
rect 16027 39684 16031 39740
rect 16031 39684 16087 39740
rect 16087 39684 16091 39740
rect 16027 39680 16091 39684
rect 21721 39740 21785 39744
rect 21721 39684 21725 39740
rect 21725 39684 21781 39740
rect 21781 39684 21785 39740
rect 21721 39680 21785 39684
rect 21801 39740 21865 39744
rect 21801 39684 21805 39740
rect 21805 39684 21861 39740
rect 21861 39684 21865 39740
rect 21801 39680 21865 39684
rect 21881 39740 21945 39744
rect 21881 39684 21885 39740
rect 21885 39684 21941 39740
rect 21941 39684 21945 39740
rect 21881 39680 21945 39684
rect 21961 39740 22025 39744
rect 21961 39684 21965 39740
rect 21965 39684 22021 39740
rect 22021 39684 22025 39740
rect 21961 39680 22025 39684
rect 7972 39340 8036 39404
rect 19748 39340 19812 39404
rect 6886 39196 6950 39200
rect 6886 39140 6890 39196
rect 6890 39140 6946 39196
rect 6946 39140 6950 39196
rect 6886 39136 6950 39140
rect 6966 39196 7030 39200
rect 6966 39140 6970 39196
rect 6970 39140 7026 39196
rect 7026 39140 7030 39196
rect 6966 39136 7030 39140
rect 7046 39196 7110 39200
rect 7046 39140 7050 39196
rect 7050 39140 7106 39196
rect 7106 39140 7110 39196
rect 7046 39136 7110 39140
rect 7126 39196 7190 39200
rect 7126 39140 7130 39196
rect 7130 39140 7186 39196
rect 7186 39140 7190 39196
rect 7126 39136 7190 39140
rect 12820 39196 12884 39200
rect 12820 39140 12824 39196
rect 12824 39140 12880 39196
rect 12880 39140 12884 39196
rect 12820 39136 12884 39140
rect 12900 39196 12964 39200
rect 12900 39140 12904 39196
rect 12904 39140 12960 39196
rect 12960 39140 12964 39196
rect 12900 39136 12964 39140
rect 12980 39196 13044 39200
rect 12980 39140 12984 39196
rect 12984 39140 13040 39196
rect 13040 39140 13044 39196
rect 12980 39136 13044 39140
rect 13060 39196 13124 39200
rect 13060 39140 13064 39196
rect 13064 39140 13120 39196
rect 13120 39140 13124 39196
rect 13060 39136 13124 39140
rect 18754 39196 18818 39200
rect 18754 39140 18758 39196
rect 18758 39140 18814 39196
rect 18814 39140 18818 39196
rect 18754 39136 18818 39140
rect 18834 39196 18898 39200
rect 18834 39140 18838 39196
rect 18838 39140 18894 39196
rect 18894 39140 18898 39196
rect 18834 39136 18898 39140
rect 18914 39196 18978 39200
rect 18914 39140 18918 39196
rect 18918 39140 18974 39196
rect 18974 39140 18978 39196
rect 18914 39136 18978 39140
rect 18994 39196 19058 39200
rect 18994 39140 18998 39196
rect 18998 39140 19054 39196
rect 19054 39140 19058 39196
rect 18994 39136 19058 39140
rect 24688 39196 24752 39200
rect 24688 39140 24692 39196
rect 24692 39140 24748 39196
rect 24748 39140 24752 39196
rect 24688 39136 24752 39140
rect 24768 39196 24832 39200
rect 24768 39140 24772 39196
rect 24772 39140 24828 39196
rect 24828 39140 24832 39196
rect 24768 39136 24832 39140
rect 24848 39196 24912 39200
rect 24848 39140 24852 39196
rect 24852 39140 24908 39196
rect 24908 39140 24912 39196
rect 24848 39136 24912 39140
rect 24928 39196 24992 39200
rect 24928 39140 24932 39196
rect 24932 39140 24988 39196
rect 24988 39140 24992 39196
rect 24928 39136 24992 39140
rect 13676 38932 13740 38996
rect 22508 38932 22572 38996
rect 1900 38720 1964 38724
rect 1900 38664 1950 38720
rect 1950 38664 1964 38720
rect 1900 38660 1964 38664
rect 612 38524 676 38588
rect 3919 38652 3983 38656
rect 3919 38596 3923 38652
rect 3923 38596 3979 38652
rect 3979 38596 3983 38652
rect 3919 38592 3983 38596
rect 3999 38652 4063 38656
rect 3999 38596 4003 38652
rect 4003 38596 4059 38652
rect 4059 38596 4063 38652
rect 3999 38592 4063 38596
rect 4079 38652 4143 38656
rect 4079 38596 4083 38652
rect 4083 38596 4139 38652
rect 4139 38596 4143 38652
rect 4079 38592 4143 38596
rect 4159 38652 4223 38656
rect 4159 38596 4163 38652
rect 4163 38596 4219 38652
rect 4219 38596 4223 38652
rect 4159 38592 4223 38596
rect 22324 38796 22388 38860
rect 19196 38660 19260 38724
rect 21404 38660 21468 38724
rect 9853 38652 9917 38656
rect 9853 38596 9857 38652
rect 9857 38596 9913 38652
rect 9913 38596 9917 38652
rect 9853 38592 9917 38596
rect 9933 38652 9997 38656
rect 9933 38596 9937 38652
rect 9937 38596 9993 38652
rect 9993 38596 9997 38652
rect 9933 38592 9997 38596
rect 10013 38652 10077 38656
rect 10013 38596 10017 38652
rect 10017 38596 10073 38652
rect 10073 38596 10077 38652
rect 10013 38592 10077 38596
rect 10093 38652 10157 38656
rect 10093 38596 10097 38652
rect 10097 38596 10153 38652
rect 10153 38596 10157 38652
rect 10093 38592 10157 38596
rect 15787 38652 15851 38656
rect 15787 38596 15791 38652
rect 15791 38596 15847 38652
rect 15847 38596 15851 38652
rect 15787 38592 15851 38596
rect 15867 38652 15931 38656
rect 15867 38596 15871 38652
rect 15871 38596 15927 38652
rect 15927 38596 15931 38652
rect 15867 38592 15931 38596
rect 15947 38652 16011 38656
rect 15947 38596 15951 38652
rect 15951 38596 16007 38652
rect 16007 38596 16011 38652
rect 15947 38592 16011 38596
rect 16027 38652 16091 38656
rect 16027 38596 16031 38652
rect 16031 38596 16087 38652
rect 16087 38596 16091 38652
rect 16027 38592 16091 38596
rect 21721 38652 21785 38656
rect 21721 38596 21725 38652
rect 21725 38596 21781 38652
rect 21781 38596 21785 38652
rect 21721 38592 21785 38596
rect 21801 38652 21865 38656
rect 21801 38596 21805 38652
rect 21805 38596 21861 38652
rect 21861 38596 21865 38652
rect 21801 38592 21865 38596
rect 21881 38652 21945 38656
rect 21881 38596 21885 38652
rect 21885 38596 21941 38652
rect 21941 38596 21945 38652
rect 21881 38592 21945 38596
rect 21961 38652 22025 38656
rect 21961 38596 21965 38652
rect 21965 38596 22021 38652
rect 22021 38596 22025 38652
rect 21961 38592 22025 38596
rect 12572 38388 12636 38452
rect 3004 38252 3068 38316
rect 6886 38108 6950 38112
rect 6886 38052 6890 38108
rect 6890 38052 6946 38108
rect 6946 38052 6950 38108
rect 6886 38048 6950 38052
rect 6966 38108 7030 38112
rect 6966 38052 6970 38108
rect 6970 38052 7026 38108
rect 7026 38052 7030 38108
rect 6966 38048 7030 38052
rect 7046 38108 7110 38112
rect 7046 38052 7050 38108
rect 7050 38052 7106 38108
rect 7106 38052 7110 38108
rect 7046 38048 7110 38052
rect 7126 38108 7190 38112
rect 7126 38052 7130 38108
rect 7130 38052 7186 38108
rect 7186 38052 7190 38108
rect 7126 38048 7190 38052
rect 12820 38108 12884 38112
rect 12820 38052 12824 38108
rect 12824 38052 12880 38108
rect 12880 38052 12884 38108
rect 12820 38048 12884 38052
rect 12900 38108 12964 38112
rect 12900 38052 12904 38108
rect 12904 38052 12960 38108
rect 12960 38052 12964 38108
rect 12900 38048 12964 38052
rect 12980 38108 13044 38112
rect 12980 38052 12984 38108
rect 12984 38052 13040 38108
rect 13040 38052 13044 38108
rect 12980 38048 13044 38052
rect 13060 38108 13124 38112
rect 13060 38052 13064 38108
rect 13064 38052 13120 38108
rect 13120 38052 13124 38108
rect 13060 38048 13124 38052
rect 18754 38108 18818 38112
rect 18754 38052 18758 38108
rect 18758 38052 18814 38108
rect 18814 38052 18818 38108
rect 18754 38048 18818 38052
rect 18834 38108 18898 38112
rect 18834 38052 18838 38108
rect 18838 38052 18894 38108
rect 18894 38052 18898 38108
rect 18834 38048 18898 38052
rect 18914 38108 18978 38112
rect 18914 38052 18918 38108
rect 18918 38052 18974 38108
rect 18974 38052 18978 38108
rect 18914 38048 18978 38052
rect 18994 38108 19058 38112
rect 18994 38052 18998 38108
rect 18998 38052 19054 38108
rect 19054 38052 19058 38108
rect 18994 38048 19058 38052
rect 24688 38108 24752 38112
rect 24688 38052 24692 38108
rect 24692 38052 24748 38108
rect 24748 38052 24752 38108
rect 24688 38048 24752 38052
rect 24768 38108 24832 38112
rect 24768 38052 24772 38108
rect 24772 38052 24828 38108
rect 24828 38052 24832 38108
rect 24768 38048 24832 38052
rect 24848 38108 24912 38112
rect 24848 38052 24852 38108
rect 24852 38052 24908 38108
rect 24908 38052 24912 38108
rect 24848 38048 24912 38052
rect 24928 38108 24992 38112
rect 24928 38052 24932 38108
rect 24932 38052 24988 38108
rect 24988 38052 24992 38108
rect 24928 38048 24992 38052
rect 980 37980 1044 38044
rect 3556 37844 3620 37908
rect 16620 37844 16684 37908
rect 4660 37708 4724 37772
rect 8892 37708 8956 37772
rect 3919 37564 3983 37568
rect 3919 37508 3923 37564
rect 3923 37508 3979 37564
rect 3979 37508 3983 37564
rect 3919 37504 3983 37508
rect 3999 37564 4063 37568
rect 3999 37508 4003 37564
rect 4003 37508 4059 37564
rect 4059 37508 4063 37564
rect 3999 37504 4063 37508
rect 4079 37564 4143 37568
rect 4079 37508 4083 37564
rect 4083 37508 4139 37564
rect 4139 37508 4143 37564
rect 4079 37504 4143 37508
rect 4159 37564 4223 37568
rect 4159 37508 4163 37564
rect 4163 37508 4219 37564
rect 4219 37508 4223 37564
rect 4159 37504 4223 37508
rect 9853 37564 9917 37568
rect 9853 37508 9857 37564
rect 9857 37508 9913 37564
rect 9913 37508 9917 37564
rect 9853 37504 9917 37508
rect 9933 37564 9997 37568
rect 9933 37508 9937 37564
rect 9937 37508 9993 37564
rect 9993 37508 9997 37564
rect 9933 37504 9997 37508
rect 10013 37564 10077 37568
rect 10013 37508 10017 37564
rect 10017 37508 10073 37564
rect 10073 37508 10077 37564
rect 10013 37504 10077 37508
rect 10093 37564 10157 37568
rect 10093 37508 10097 37564
rect 10097 37508 10153 37564
rect 10153 37508 10157 37564
rect 10093 37504 10157 37508
rect 15787 37564 15851 37568
rect 15787 37508 15791 37564
rect 15791 37508 15847 37564
rect 15847 37508 15851 37564
rect 15787 37504 15851 37508
rect 15867 37564 15931 37568
rect 15867 37508 15871 37564
rect 15871 37508 15927 37564
rect 15927 37508 15931 37564
rect 15867 37504 15931 37508
rect 15947 37564 16011 37568
rect 15947 37508 15951 37564
rect 15951 37508 16007 37564
rect 16007 37508 16011 37564
rect 15947 37504 16011 37508
rect 16027 37564 16091 37568
rect 16027 37508 16031 37564
rect 16031 37508 16087 37564
rect 16087 37508 16091 37564
rect 16027 37504 16091 37508
rect 21721 37564 21785 37568
rect 21721 37508 21725 37564
rect 21725 37508 21781 37564
rect 21781 37508 21785 37564
rect 21721 37504 21785 37508
rect 21801 37564 21865 37568
rect 21801 37508 21805 37564
rect 21805 37508 21861 37564
rect 21861 37508 21865 37564
rect 21801 37504 21865 37508
rect 21881 37564 21945 37568
rect 21881 37508 21885 37564
rect 21885 37508 21941 37564
rect 21941 37508 21945 37564
rect 21881 37504 21945 37508
rect 21961 37564 22025 37568
rect 21961 37508 21965 37564
rect 21965 37508 22021 37564
rect 22021 37508 22025 37564
rect 21961 37504 22025 37508
rect 8524 37300 8588 37364
rect 6886 37020 6950 37024
rect 6886 36964 6890 37020
rect 6890 36964 6946 37020
rect 6946 36964 6950 37020
rect 6886 36960 6950 36964
rect 6966 37020 7030 37024
rect 6966 36964 6970 37020
rect 6970 36964 7026 37020
rect 7026 36964 7030 37020
rect 6966 36960 7030 36964
rect 7046 37020 7110 37024
rect 7046 36964 7050 37020
rect 7050 36964 7106 37020
rect 7106 36964 7110 37020
rect 7046 36960 7110 36964
rect 7126 37020 7190 37024
rect 7126 36964 7130 37020
rect 7130 36964 7186 37020
rect 7186 36964 7190 37020
rect 7126 36960 7190 36964
rect 12820 37020 12884 37024
rect 12820 36964 12824 37020
rect 12824 36964 12880 37020
rect 12880 36964 12884 37020
rect 12820 36960 12884 36964
rect 12900 37020 12964 37024
rect 12900 36964 12904 37020
rect 12904 36964 12960 37020
rect 12960 36964 12964 37020
rect 12900 36960 12964 36964
rect 12980 37020 13044 37024
rect 12980 36964 12984 37020
rect 12984 36964 13040 37020
rect 13040 36964 13044 37020
rect 12980 36960 13044 36964
rect 13060 37020 13124 37024
rect 13060 36964 13064 37020
rect 13064 36964 13120 37020
rect 13120 36964 13124 37020
rect 13060 36960 13124 36964
rect 18754 37020 18818 37024
rect 18754 36964 18758 37020
rect 18758 36964 18814 37020
rect 18814 36964 18818 37020
rect 18754 36960 18818 36964
rect 18834 37020 18898 37024
rect 18834 36964 18838 37020
rect 18838 36964 18894 37020
rect 18894 36964 18898 37020
rect 18834 36960 18898 36964
rect 18914 37020 18978 37024
rect 18914 36964 18918 37020
rect 18918 36964 18974 37020
rect 18974 36964 18978 37020
rect 18914 36960 18978 36964
rect 18994 37020 19058 37024
rect 18994 36964 18998 37020
rect 18998 36964 19054 37020
rect 19054 36964 19058 37020
rect 18994 36960 19058 36964
rect 24688 37020 24752 37024
rect 24688 36964 24692 37020
rect 24692 36964 24748 37020
rect 24748 36964 24752 37020
rect 24688 36960 24752 36964
rect 24768 37020 24832 37024
rect 24768 36964 24772 37020
rect 24772 36964 24828 37020
rect 24828 36964 24832 37020
rect 24768 36960 24832 36964
rect 24848 37020 24912 37024
rect 24848 36964 24852 37020
rect 24852 36964 24908 37020
rect 24908 36964 24912 37020
rect 24848 36960 24912 36964
rect 24928 37020 24992 37024
rect 24928 36964 24932 37020
rect 24932 36964 24988 37020
rect 24988 36964 24992 37020
rect 24928 36960 24992 36964
rect 796 36620 860 36684
rect 3919 36476 3983 36480
rect 3919 36420 3923 36476
rect 3923 36420 3979 36476
rect 3979 36420 3983 36476
rect 3919 36416 3983 36420
rect 3999 36476 4063 36480
rect 3999 36420 4003 36476
rect 4003 36420 4059 36476
rect 4059 36420 4063 36476
rect 3999 36416 4063 36420
rect 4079 36476 4143 36480
rect 4079 36420 4083 36476
rect 4083 36420 4139 36476
rect 4139 36420 4143 36476
rect 4079 36416 4143 36420
rect 4159 36476 4223 36480
rect 4159 36420 4163 36476
rect 4163 36420 4219 36476
rect 4219 36420 4223 36476
rect 4159 36416 4223 36420
rect 9853 36476 9917 36480
rect 9853 36420 9857 36476
rect 9857 36420 9913 36476
rect 9913 36420 9917 36476
rect 9853 36416 9917 36420
rect 9933 36476 9997 36480
rect 9933 36420 9937 36476
rect 9937 36420 9993 36476
rect 9993 36420 9997 36476
rect 9933 36416 9997 36420
rect 10013 36476 10077 36480
rect 10013 36420 10017 36476
rect 10017 36420 10073 36476
rect 10073 36420 10077 36476
rect 10013 36416 10077 36420
rect 10093 36476 10157 36480
rect 10093 36420 10097 36476
rect 10097 36420 10153 36476
rect 10153 36420 10157 36476
rect 10093 36416 10157 36420
rect 15787 36476 15851 36480
rect 15787 36420 15791 36476
rect 15791 36420 15847 36476
rect 15847 36420 15851 36476
rect 15787 36416 15851 36420
rect 15867 36476 15931 36480
rect 15867 36420 15871 36476
rect 15871 36420 15927 36476
rect 15927 36420 15931 36476
rect 15867 36416 15931 36420
rect 15947 36476 16011 36480
rect 15947 36420 15951 36476
rect 15951 36420 16007 36476
rect 16007 36420 16011 36476
rect 15947 36416 16011 36420
rect 16027 36476 16091 36480
rect 16027 36420 16031 36476
rect 16031 36420 16087 36476
rect 16087 36420 16091 36476
rect 16027 36416 16091 36420
rect 21721 36476 21785 36480
rect 21721 36420 21725 36476
rect 21725 36420 21781 36476
rect 21781 36420 21785 36476
rect 21721 36416 21785 36420
rect 21801 36476 21865 36480
rect 21801 36420 21805 36476
rect 21805 36420 21861 36476
rect 21861 36420 21865 36476
rect 21801 36416 21865 36420
rect 21881 36476 21945 36480
rect 21881 36420 21885 36476
rect 21885 36420 21941 36476
rect 21941 36420 21945 36476
rect 21881 36416 21945 36420
rect 21961 36476 22025 36480
rect 21961 36420 21965 36476
rect 21965 36420 22021 36476
rect 22021 36420 22025 36476
rect 21961 36416 22025 36420
rect 21220 36076 21284 36140
rect 10364 35940 10428 36004
rect 6886 35932 6950 35936
rect 6886 35876 6890 35932
rect 6890 35876 6946 35932
rect 6946 35876 6950 35932
rect 6886 35872 6950 35876
rect 6966 35932 7030 35936
rect 6966 35876 6970 35932
rect 6970 35876 7026 35932
rect 7026 35876 7030 35932
rect 6966 35872 7030 35876
rect 7046 35932 7110 35936
rect 7046 35876 7050 35932
rect 7050 35876 7106 35932
rect 7106 35876 7110 35932
rect 7046 35872 7110 35876
rect 7126 35932 7190 35936
rect 7126 35876 7130 35932
rect 7130 35876 7186 35932
rect 7186 35876 7190 35932
rect 7126 35872 7190 35876
rect 12820 35932 12884 35936
rect 12820 35876 12824 35932
rect 12824 35876 12880 35932
rect 12880 35876 12884 35932
rect 12820 35872 12884 35876
rect 12900 35932 12964 35936
rect 12900 35876 12904 35932
rect 12904 35876 12960 35932
rect 12960 35876 12964 35932
rect 12900 35872 12964 35876
rect 12980 35932 13044 35936
rect 12980 35876 12984 35932
rect 12984 35876 13040 35932
rect 13040 35876 13044 35932
rect 12980 35872 13044 35876
rect 13060 35932 13124 35936
rect 13060 35876 13064 35932
rect 13064 35876 13120 35932
rect 13120 35876 13124 35932
rect 13060 35872 13124 35876
rect 18754 35932 18818 35936
rect 18754 35876 18758 35932
rect 18758 35876 18814 35932
rect 18814 35876 18818 35932
rect 18754 35872 18818 35876
rect 18834 35932 18898 35936
rect 18834 35876 18838 35932
rect 18838 35876 18894 35932
rect 18894 35876 18898 35932
rect 18834 35872 18898 35876
rect 18914 35932 18978 35936
rect 18914 35876 18918 35932
rect 18918 35876 18974 35932
rect 18974 35876 18978 35932
rect 18914 35872 18978 35876
rect 18994 35932 19058 35936
rect 18994 35876 18998 35932
rect 18998 35876 19054 35932
rect 19054 35876 19058 35932
rect 18994 35872 19058 35876
rect 24688 35932 24752 35936
rect 24688 35876 24692 35932
rect 24692 35876 24748 35932
rect 24748 35876 24752 35932
rect 24688 35872 24752 35876
rect 24768 35932 24832 35936
rect 24768 35876 24772 35932
rect 24772 35876 24828 35932
rect 24828 35876 24832 35932
rect 24768 35872 24832 35876
rect 24848 35932 24912 35936
rect 24848 35876 24852 35932
rect 24852 35876 24908 35932
rect 24908 35876 24912 35932
rect 24848 35872 24912 35876
rect 24928 35932 24992 35936
rect 24928 35876 24932 35932
rect 24932 35876 24988 35932
rect 24988 35876 24992 35932
rect 24928 35872 24992 35876
rect 3188 35804 3252 35868
rect 3188 35124 3252 35188
rect 8708 35592 8772 35596
rect 8708 35536 8758 35592
rect 8758 35536 8772 35592
rect 8708 35532 8772 35536
rect 3919 35388 3983 35392
rect 3919 35332 3923 35388
rect 3923 35332 3979 35388
rect 3979 35332 3983 35388
rect 3919 35328 3983 35332
rect 3999 35388 4063 35392
rect 3999 35332 4003 35388
rect 4003 35332 4059 35388
rect 4059 35332 4063 35388
rect 3999 35328 4063 35332
rect 4079 35388 4143 35392
rect 4079 35332 4083 35388
rect 4083 35332 4139 35388
rect 4139 35332 4143 35388
rect 4079 35328 4143 35332
rect 4159 35388 4223 35392
rect 4159 35332 4163 35388
rect 4163 35332 4219 35388
rect 4219 35332 4223 35388
rect 4159 35328 4223 35332
rect 9853 35388 9917 35392
rect 9853 35332 9857 35388
rect 9857 35332 9913 35388
rect 9913 35332 9917 35388
rect 9853 35328 9917 35332
rect 9933 35388 9997 35392
rect 9933 35332 9937 35388
rect 9937 35332 9993 35388
rect 9993 35332 9997 35388
rect 9933 35328 9997 35332
rect 10013 35388 10077 35392
rect 10013 35332 10017 35388
rect 10017 35332 10073 35388
rect 10073 35332 10077 35388
rect 10013 35328 10077 35332
rect 10093 35388 10157 35392
rect 10093 35332 10097 35388
rect 10097 35332 10153 35388
rect 10153 35332 10157 35388
rect 10093 35328 10157 35332
rect 15787 35388 15851 35392
rect 15787 35332 15791 35388
rect 15791 35332 15847 35388
rect 15847 35332 15851 35388
rect 15787 35328 15851 35332
rect 15867 35388 15931 35392
rect 15867 35332 15871 35388
rect 15871 35332 15927 35388
rect 15927 35332 15931 35388
rect 15867 35328 15931 35332
rect 15947 35388 16011 35392
rect 15947 35332 15951 35388
rect 15951 35332 16007 35388
rect 16007 35332 16011 35388
rect 15947 35328 16011 35332
rect 16027 35388 16091 35392
rect 16027 35332 16031 35388
rect 16031 35332 16087 35388
rect 16087 35332 16091 35388
rect 16027 35328 16091 35332
rect 21721 35388 21785 35392
rect 21721 35332 21725 35388
rect 21725 35332 21781 35388
rect 21781 35332 21785 35388
rect 21721 35328 21785 35332
rect 21801 35388 21865 35392
rect 21801 35332 21805 35388
rect 21805 35332 21861 35388
rect 21861 35332 21865 35388
rect 21801 35328 21865 35332
rect 21881 35388 21945 35392
rect 21881 35332 21885 35388
rect 21885 35332 21941 35388
rect 21941 35332 21945 35388
rect 21881 35328 21945 35332
rect 21961 35388 22025 35392
rect 21961 35332 21965 35388
rect 21965 35332 22021 35388
rect 22021 35332 22025 35388
rect 21961 35328 22025 35332
rect 5580 34852 5644 34916
rect 6886 34844 6950 34848
rect 6886 34788 6890 34844
rect 6890 34788 6946 34844
rect 6946 34788 6950 34844
rect 6886 34784 6950 34788
rect 6966 34844 7030 34848
rect 6966 34788 6970 34844
rect 6970 34788 7026 34844
rect 7026 34788 7030 34844
rect 6966 34784 7030 34788
rect 7046 34844 7110 34848
rect 7046 34788 7050 34844
rect 7050 34788 7106 34844
rect 7106 34788 7110 34844
rect 7046 34784 7110 34788
rect 7126 34844 7190 34848
rect 7126 34788 7130 34844
rect 7130 34788 7186 34844
rect 7186 34788 7190 34844
rect 7126 34784 7190 34788
rect 12820 34844 12884 34848
rect 12820 34788 12824 34844
rect 12824 34788 12880 34844
rect 12880 34788 12884 34844
rect 12820 34784 12884 34788
rect 12900 34844 12964 34848
rect 12900 34788 12904 34844
rect 12904 34788 12960 34844
rect 12960 34788 12964 34844
rect 12900 34784 12964 34788
rect 12980 34844 13044 34848
rect 12980 34788 12984 34844
rect 12984 34788 13040 34844
rect 13040 34788 13044 34844
rect 12980 34784 13044 34788
rect 13060 34844 13124 34848
rect 13060 34788 13064 34844
rect 13064 34788 13120 34844
rect 13120 34788 13124 34844
rect 13060 34784 13124 34788
rect 18754 34844 18818 34848
rect 18754 34788 18758 34844
rect 18758 34788 18814 34844
rect 18814 34788 18818 34844
rect 18754 34784 18818 34788
rect 18834 34844 18898 34848
rect 18834 34788 18838 34844
rect 18838 34788 18894 34844
rect 18894 34788 18898 34844
rect 18834 34784 18898 34788
rect 18914 34844 18978 34848
rect 18914 34788 18918 34844
rect 18918 34788 18974 34844
rect 18974 34788 18978 34844
rect 18914 34784 18978 34788
rect 18994 34844 19058 34848
rect 18994 34788 18998 34844
rect 18998 34788 19054 34844
rect 19054 34788 19058 34844
rect 18994 34784 19058 34788
rect 24688 34844 24752 34848
rect 24688 34788 24692 34844
rect 24692 34788 24748 34844
rect 24748 34788 24752 34844
rect 24688 34784 24752 34788
rect 24768 34844 24832 34848
rect 24768 34788 24772 34844
rect 24772 34788 24828 34844
rect 24828 34788 24832 34844
rect 24768 34784 24832 34788
rect 24848 34844 24912 34848
rect 24848 34788 24852 34844
rect 24852 34788 24908 34844
rect 24908 34788 24912 34844
rect 24848 34784 24912 34788
rect 24928 34844 24992 34848
rect 24928 34788 24932 34844
rect 24932 34788 24988 34844
rect 24988 34788 24992 34844
rect 24928 34784 24992 34788
rect 3919 34300 3983 34304
rect 3919 34244 3923 34300
rect 3923 34244 3979 34300
rect 3979 34244 3983 34300
rect 3919 34240 3983 34244
rect 3999 34300 4063 34304
rect 3999 34244 4003 34300
rect 4003 34244 4059 34300
rect 4059 34244 4063 34300
rect 3999 34240 4063 34244
rect 4079 34300 4143 34304
rect 4079 34244 4083 34300
rect 4083 34244 4139 34300
rect 4139 34244 4143 34300
rect 4079 34240 4143 34244
rect 4159 34300 4223 34304
rect 4159 34244 4163 34300
rect 4163 34244 4219 34300
rect 4219 34244 4223 34300
rect 4159 34240 4223 34244
rect 9853 34300 9917 34304
rect 9853 34244 9857 34300
rect 9857 34244 9913 34300
rect 9913 34244 9917 34300
rect 9853 34240 9917 34244
rect 9933 34300 9997 34304
rect 9933 34244 9937 34300
rect 9937 34244 9993 34300
rect 9993 34244 9997 34300
rect 9933 34240 9997 34244
rect 10013 34300 10077 34304
rect 10013 34244 10017 34300
rect 10017 34244 10073 34300
rect 10073 34244 10077 34300
rect 10013 34240 10077 34244
rect 10093 34300 10157 34304
rect 10093 34244 10097 34300
rect 10097 34244 10153 34300
rect 10153 34244 10157 34300
rect 10093 34240 10157 34244
rect 15787 34300 15851 34304
rect 15787 34244 15791 34300
rect 15791 34244 15847 34300
rect 15847 34244 15851 34300
rect 15787 34240 15851 34244
rect 15867 34300 15931 34304
rect 15867 34244 15871 34300
rect 15871 34244 15927 34300
rect 15927 34244 15931 34300
rect 15867 34240 15931 34244
rect 15947 34300 16011 34304
rect 15947 34244 15951 34300
rect 15951 34244 16007 34300
rect 16007 34244 16011 34300
rect 15947 34240 16011 34244
rect 16027 34300 16091 34304
rect 16027 34244 16031 34300
rect 16031 34244 16087 34300
rect 16087 34244 16091 34300
rect 16027 34240 16091 34244
rect 21721 34300 21785 34304
rect 21721 34244 21725 34300
rect 21725 34244 21781 34300
rect 21781 34244 21785 34300
rect 21721 34240 21785 34244
rect 21801 34300 21865 34304
rect 21801 34244 21805 34300
rect 21805 34244 21861 34300
rect 21861 34244 21865 34300
rect 21801 34240 21865 34244
rect 21881 34300 21945 34304
rect 21881 34244 21885 34300
rect 21885 34244 21941 34300
rect 21941 34244 21945 34300
rect 21881 34240 21945 34244
rect 21961 34300 22025 34304
rect 21961 34244 21965 34300
rect 21965 34244 22021 34300
rect 22021 34244 22025 34300
rect 21961 34240 22025 34244
rect 7604 33900 7668 33964
rect 14596 33900 14660 33964
rect 22876 33900 22940 33964
rect 6886 33756 6950 33760
rect 6886 33700 6890 33756
rect 6890 33700 6946 33756
rect 6946 33700 6950 33756
rect 6886 33696 6950 33700
rect 6966 33756 7030 33760
rect 6966 33700 6970 33756
rect 6970 33700 7026 33756
rect 7026 33700 7030 33756
rect 6966 33696 7030 33700
rect 7046 33756 7110 33760
rect 7046 33700 7050 33756
rect 7050 33700 7106 33756
rect 7106 33700 7110 33756
rect 7046 33696 7110 33700
rect 7126 33756 7190 33760
rect 7126 33700 7130 33756
rect 7130 33700 7186 33756
rect 7186 33700 7190 33756
rect 7126 33696 7190 33700
rect 12820 33756 12884 33760
rect 12820 33700 12824 33756
rect 12824 33700 12880 33756
rect 12880 33700 12884 33756
rect 12820 33696 12884 33700
rect 12900 33756 12964 33760
rect 12900 33700 12904 33756
rect 12904 33700 12960 33756
rect 12960 33700 12964 33756
rect 12900 33696 12964 33700
rect 12980 33756 13044 33760
rect 12980 33700 12984 33756
rect 12984 33700 13040 33756
rect 13040 33700 13044 33756
rect 12980 33696 13044 33700
rect 13060 33756 13124 33760
rect 13060 33700 13064 33756
rect 13064 33700 13120 33756
rect 13120 33700 13124 33756
rect 13060 33696 13124 33700
rect 18754 33756 18818 33760
rect 18754 33700 18758 33756
rect 18758 33700 18814 33756
rect 18814 33700 18818 33756
rect 18754 33696 18818 33700
rect 18834 33756 18898 33760
rect 18834 33700 18838 33756
rect 18838 33700 18894 33756
rect 18894 33700 18898 33756
rect 18834 33696 18898 33700
rect 18914 33756 18978 33760
rect 18914 33700 18918 33756
rect 18918 33700 18974 33756
rect 18974 33700 18978 33756
rect 18914 33696 18978 33700
rect 18994 33756 19058 33760
rect 18994 33700 18998 33756
rect 18998 33700 19054 33756
rect 19054 33700 19058 33756
rect 18994 33696 19058 33700
rect 24688 33756 24752 33760
rect 24688 33700 24692 33756
rect 24692 33700 24748 33756
rect 24748 33700 24752 33756
rect 24688 33696 24752 33700
rect 24768 33756 24832 33760
rect 24768 33700 24772 33756
rect 24772 33700 24828 33756
rect 24828 33700 24832 33756
rect 24768 33696 24832 33700
rect 24848 33756 24912 33760
rect 24848 33700 24852 33756
rect 24852 33700 24908 33756
rect 24908 33700 24912 33756
rect 24848 33696 24912 33700
rect 24928 33756 24992 33760
rect 24928 33700 24932 33756
rect 24932 33700 24988 33756
rect 24988 33700 24992 33756
rect 24928 33696 24992 33700
rect 1900 33628 1964 33692
rect 7972 33416 8036 33420
rect 7972 33360 7986 33416
rect 7986 33360 8036 33416
rect 7972 33356 8036 33360
rect 3919 33212 3983 33216
rect 3919 33156 3923 33212
rect 3923 33156 3979 33212
rect 3979 33156 3983 33212
rect 3919 33152 3983 33156
rect 3999 33212 4063 33216
rect 3999 33156 4003 33212
rect 4003 33156 4059 33212
rect 4059 33156 4063 33212
rect 3999 33152 4063 33156
rect 4079 33212 4143 33216
rect 4079 33156 4083 33212
rect 4083 33156 4139 33212
rect 4139 33156 4143 33212
rect 4079 33152 4143 33156
rect 4159 33212 4223 33216
rect 4159 33156 4163 33212
rect 4163 33156 4219 33212
rect 4219 33156 4223 33212
rect 4159 33152 4223 33156
rect 9853 33212 9917 33216
rect 9853 33156 9857 33212
rect 9857 33156 9913 33212
rect 9913 33156 9917 33212
rect 9853 33152 9917 33156
rect 9933 33212 9997 33216
rect 9933 33156 9937 33212
rect 9937 33156 9993 33212
rect 9993 33156 9997 33212
rect 9933 33152 9997 33156
rect 10013 33212 10077 33216
rect 10013 33156 10017 33212
rect 10017 33156 10073 33212
rect 10073 33156 10077 33212
rect 10013 33152 10077 33156
rect 10093 33212 10157 33216
rect 10093 33156 10097 33212
rect 10097 33156 10153 33212
rect 10153 33156 10157 33212
rect 10093 33152 10157 33156
rect 15787 33212 15851 33216
rect 15787 33156 15791 33212
rect 15791 33156 15847 33212
rect 15847 33156 15851 33212
rect 15787 33152 15851 33156
rect 15867 33212 15931 33216
rect 15867 33156 15871 33212
rect 15871 33156 15927 33212
rect 15927 33156 15931 33212
rect 15867 33152 15931 33156
rect 15947 33212 16011 33216
rect 15947 33156 15951 33212
rect 15951 33156 16007 33212
rect 16007 33156 16011 33212
rect 15947 33152 16011 33156
rect 16027 33212 16091 33216
rect 16027 33156 16031 33212
rect 16031 33156 16087 33212
rect 16087 33156 16091 33212
rect 16027 33152 16091 33156
rect 21721 33212 21785 33216
rect 21721 33156 21725 33212
rect 21725 33156 21781 33212
rect 21781 33156 21785 33212
rect 21721 33152 21785 33156
rect 21801 33212 21865 33216
rect 21801 33156 21805 33212
rect 21805 33156 21861 33212
rect 21861 33156 21865 33212
rect 21801 33152 21865 33156
rect 21881 33212 21945 33216
rect 21881 33156 21885 33212
rect 21885 33156 21941 33212
rect 21941 33156 21945 33212
rect 21881 33152 21945 33156
rect 21961 33212 22025 33216
rect 21961 33156 21965 33212
rect 21965 33156 22021 33212
rect 22021 33156 22025 33212
rect 21961 33152 22025 33156
rect 4476 33084 4540 33148
rect 21036 33084 21100 33148
rect 7420 32948 7484 33012
rect 3004 32812 3068 32876
rect 3556 32812 3620 32876
rect 4292 32812 4356 32876
rect 6886 32668 6950 32672
rect 6886 32612 6890 32668
rect 6890 32612 6946 32668
rect 6946 32612 6950 32668
rect 6886 32608 6950 32612
rect 6966 32668 7030 32672
rect 6966 32612 6970 32668
rect 6970 32612 7026 32668
rect 7026 32612 7030 32668
rect 6966 32608 7030 32612
rect 7046 32668 7110 32672
rect 7046 32612 7050 32668
rect 7050 32612 7106 32668
rect 7106 32612 7110 32668
rect 7046 32608 7110 32612
rect 7126 32668 7190 32672
rect 7126 32612 7130 32668
rect 7130 32612 7186 32668
rect 7186 32612 7190 32668
rect 7126 32608 7190 32612
rect 12820 32668 12884 32672
rect 12820 32612 12824 32668
rect 12824 32612 12880 32668
rect 12880 32612 12884 32668
rect 12820 32608 12884 32612
rect 12900 32668 12964 32672
rect 12900 32612 12904 32668
rect 12904 32612 12960 32668
rect 12960 32612 12964 32668
rect 12900 32608 12964 32612
rect 12980 32668 13044 32672
rect 12980 32612 12984 32668
rect 12984 32612 13040 32668
rect 13040 32612 13044 32668
rect 12980 32608 13044 32612
rect 13060 32668 13124 32672
rect 13060 32612 13064 32668
rect 13064 32612 13120 32668
rect 13120 32612 13124 32668
rect 13060 32608 13124 32612
rect 18754 32668 18818 32672
rect 18754 32612 18758 32668
rect 18758 32612 18814 32668
rect 18814 32612 18818 32668
rect 18754 32608 18818 32612
rect 18834 32668 18898 32672
rect 18834 32612 18838 32668
rect 18838 32612 18894 32668
rect 18894 32612 18898 32668
rect 18834 32608 18898 32612
rect 18914 32668 18978 32672
rect 18914 32612 18918 32668
rect 18918 32612 18974 32668
rect 18974 32612 18978 32668
rect 18914 32608 18978 32612
rect 18994 32668 19058 32672
rect 18994 32612 18998 32668
rect 18998 32612 19054 32668
rect 19054 32612 19058 32668
rect 18994 32608 19058 32612
rect 24688 32668 24752 32672
rect 24688 32612 24692 32668
rect 24692 32612 24748 32668
rect 24748 32612 24752 32668
rect 24688 32608 24752 32612
rect 24768 32668 24832 32672
rect 24768 32612 24772 32668
rect 24772 32612 24828 32668
rect 24828 32612 24832 32668
rect 24768 32608 24832 32612
rect 24848 32668 24912 32672
rect 24848 32612 24852 32668
rect 24852 32612 24908 32668
rect 24908 32612 24912 32668
rect 24848 32608 24912 32612
rect 24928 32668 24992 32672
rect 24928 32612 24932 32668
rect 24932 32612 24988 32668
rect 24988 32612 24992 32668
rect 24928 32608 24992 32612
rect 19380 32268 19444 32332
rect 3919 32124 3983 32128
rect 3919 32068 3923 32124
rect 3923 32068 3979 32124
rect 3979 32068 3983 32124
rect 3919 32064 3983 32068
rect 3999 32124 4063 32128
rect 3999 32068 4003 32124
rect 4003 32068 4059 32124
rect 4059 32068 4063 32124
rect 3999 32064 4063 32068
rect 4079 32124 4143 32128
rect 4079 32068 4083 32124
rect 4083 32068 4139 32124
rect 4139 32068 4143 32124
rect 4079 32064 4143 32068
rect 4159 32124 4223 32128
rect 4159 32068 4163 32124
rect 4163 32068 4219 32124
rect 4219 32068 4223 32124
rect 4159 32064 4223 32068
rect 9853 32124 9917 32128
rect 9853 32068 9857 32124
rect 9857 32068 9913 32124
rect 9913 32068 9917 32124
rect 9853 32064 9917 32068
rect 9933 32124 9997 32128
rect 9933 32068 9937 32124
rect 9937 32068 9993 32124
rect 9993 32068 9997 32124
rect 9933 32064 9997 32068
rect 10013 32124 10077 32128
rect 10013 32068 10017 32124
rect 10017 32068 10073 32124
rect 10073 32068 10077 32124
rect 10013 32064 10077 32068
rect 10093 32124 10157 32128
rect 10093 32068 10097 32124
rect 10097 32068 10153 32124
rect 10153 32068 10157 32124
rect 10093 32064 10157 32068
rect 15787 32124 15851 32128
rect 15787 32068 15791 32124
rect 15791 32068 15847 32124
rect 15847 32068 15851 32124
rect 15787 32064 15851 32068
rect 15867 32124 15931 32128
rect 15867 32068 15871 32124
rect 15871 32068 15927 32124
rect 15927 32068 15931 32124
rect 15867 32064 15931 32068
rect 15947 32124 16011 32128
rect 15947 32068 15951 32124
rect 15951 32068 16007 32124
rect 16007 32068 16011 32124
rect 15947 32064 16011 32068
rect 16027 32124 16091 32128
rect 16027 32068 16031 32124
rect 16031 32068 16087 32124
rect 16087 32068 16091 32124
rect 16027 32064 16091 32068
rect 21721 32124 21785 32128
rect 21721 32068 21725 32124
rect 21725 32068 21781 32124
rect 21781 32068 21785 32124
rect 21721 32064 21785 32068
rect 21801 32124 21865 32128
rect 21801 32068 21805 32124
rect 21805 32068 21861 32124
rect 21861 32068 21865 32124
rect 21801 32064 21865 32068
rect 21881 32124 21945 32128
rect 21881 32068 21885 32124
rect 21885 32068 21941 32124
rect 21941 32068 21945 32124
rect 21881 32064 21945 32068
rect 21961 32124 22025 32128
rect 21961 32068 21965 32124
rect 21965 32068 22021 32124
rect 22021 32068 22025 32124
rect 21961 32064 22025 32068
rect 12388 31996 12452 32060
rect 13492 31996 13556 32060
rect 15516 32056 15580 32060
rect 15516 32000 15566 32056
rect 15566 32000 15580 32056
rect 15516 31996 15580 32000
rect 4476 31860 4540 31924
rect 3556 31724 3620 31788
rect 7604 31724 7668 31788
rect 12388 31588 12452 31652
rect 6886 31580 6950 31584
rect 6886 31524 6890 31580
rect 6890 31524 6946 31580
rect 6946 31524 6950 31580
rect 6886 31520 6950 31524
rect 6966 31580 7030 31584
rect 6966 31524 6970 31580
rect 6970 31524 7026 31580
rect 7026 31524 7030 31580
rect 6966 31520 7030 31524
rect 7046 31580 7110 31584
rect 7046 31524 7050 31580
rect 7050 31524 7106 31580
rect 7106 31524 7110 31580
rect 7046 31520 7110 31524
rect 7126 31580 7190 31584
rect 7126 31524 7130 31580
rect 7130 31524 7186 31580
rect 7186 31524 7190 31580
rect 7126 31520 7190 31524
rect 3188 31180 3252 31244
rect 4660 31316 4724 31380
rect 12820 31580 12884 31584
rect 12820 31524 12824 31580
rect 12824 31524 12880 31580
rect 12880 31524 12884 31580
rect 12820 31520 12884 31524
rect 12900 31580 12964 31584
rect 12900 31524 12904 31580
rect 12904 31524 12960 31580
rect 12960 31524 12964 31580
rect 12900 31520 12964 31524
rect 12980 31580 13044 31584
rect 12980 31524 12984 31580
rect 12984 31524 13040 31580
rect 13040 31524 13044 31580
rect 12980 31520 13044 31524
rect 13060 31580 13124 31584
rect 13060 31524 13064 31580
rect 13064 31524 13120 31580
rect 13120 31524 13124 31580
rect 13060 31520 13124 31524
rect 18754 31580 18818 31584
rect 18754 31524 18758 31580
rect 18758 31524 18814 31580
rect 18814 31524 18818 31580
rect 18754 31520 18818 31524
rect 18834 31580 18898 31584
rect 18834 31524 18838 31580
rect 18838 31524 18894 31580
rect 18894 31524 18898 31580
rect 18834 31520 18898 31524
rect 18914 31580 18978 31584
rect 18914 31524 18918 31580
rect 18918 31524 18974 31580
rect 18974 31524 18978 31580
rect 18914 31520 18978 31524
rect 18994 31580 19058 31584
rect 18994 31524 18998 31580
rect 18998 31524 19054 31580
rect 19054 31524 19058 31580
rect 18994 31520 19058 31524
rect 13492 31316 13556 31380
rect 24688 31580 24752 31584
rect 24688 31524 24692 31580
rect 24692 31524 24748 31580
rect 24748 31524 24752 31580
rect 24688 31520 24752 31524
rect 24768 31580 24832 31584
rect 24768 31524 24772 31580
rect 24772 31524 24828 31580
rect 24828 31524 24832 31580
rect 24768 31520 24832 31524
rect 24848 31580 24912 31584
rect 24848 31524 24852 31580
rect 24852 31524 24908 31580
rect 24908 31524 24912 31580
rect 24848 31520 24912 31524
rect 24928 31580 24992 31584
rect 24928 31524 24932 31580
rect 24932 31524 24988 31580
rect 24988 31524 24992 31580
rect 24928 31520 24992 31524
rect 3919 31036 3983 31040
rect 3919 30980 3923 31036
rect 3923 30980 3979 31036
rect 3979 30980 3983 31036
rect 3919 30976 3983 30980
rect 3999 31036 4063 31040
rect 3999 30980 4003 31036
rect 4003 30980 4059 31036
rect 4059 30980 4063 31036
rect 3999 30976 4063 30980
rect 4079 31036 4143 31040
rect 4079 30980 4083 31036
rect 4083 30980 4139 31036
rect 4139 30980 4143 31036
rect 4079 30976 4143 30980
rect 4159 31036 4223 31040
rect 4159 30980 4163 31036
rect 4163 30980 4219 31036
rect 4219 30980 4223 31036
rect 4159 30976 4223 30980
rect 9853 31036 9917 31040
rect 9853 30980 9857 31036
rect 9857 30980 9913 31036
rect 9913 30980 9917 31036
rect 9853 30976 9917 30980
rect 9933 31036 9997 31040
rect 9933 30980 9937 31036
rect 9937 30980 9993 31036
rect 9993 30980 9997 31036
rect 9933 30976 9997 30980
rect 10013 31036 10077 31040
rect 10013 30980 10017 31036
rect 10017 30980 10073 31036
rect 10073 30980 10077 31036
rect 10013 30976 10077 30980
rect 10093 31036 10157 31040
rect 10093 30980 10097 31036
rect 10097 30980 10153 31036
rect 10153 30980 10157 31036
rect 10093 30976 10157 30980
rect 15787 31036 15851 31040
rect 15787 30980 15791 31036
rect 15791 30980 15847 31036
rect 15847 30980 15851 31036
rect 15787 30976 15851 30980
rect 15867 31036 15931 31040
rect 15867 30980 15871 31036
rect 15871 30980 15927 31036
rect 15927 30980 15931 31036
rect 15867 30976 15931 30980
rect 15947 31036 16011 31040
rect 15947 30980 15951 31036
rect 15951 30980 16007 31036
rect 16007 30980 16011 31036
rect 15947 30976 16011 30980
rect 16027 31036 16091 31040
rect 16027 30980 16031 31036
rect 16031 30980 16087 31036
rect 16087 30980 16091 31036
rect 16027 30976 16091 30980
rect 21721 31036 21785 31040
rect 21721 30980 21725 31036
rect 21725 30980 21781 31036
rect 21781 30980 21785 31036
rect 21721 30976 21785 30980
rect 21801 31036 21865 31040
rect 21801 30980 21805 31036
rect 21805 30980 21861 31036
rect 21861 30980 21865 31036
rect 21801 30976 21865 30980
rect 21881 31036 21945 31040
rect 21881 30980 21885 31036
rect 21885 30980 21941 31036
rect 21941 30980 21945 31036
rect 21881 30976 21945 30980
rect 21961 31036 22025 31040
rect 21961 30980 21965 31036
rect 21965 30980 22021 31036
rect 22021 30980 22025 31036
rect 21961 30976 22025 30980
rect 14044 30500 14108 30564
rect 6886 30492 6950 30496
rect 6886 30436 6890 30492
rect 6890 30436 6946 30492
rect 6946 30436 6950 30492
rect 6886 30432 6950 30436
rect 6966 30492 7030 30496
rect 6966 30436 6970 30492
rect 6970 30436 7026 30492
rect 7026 30436 7030 30492
rect 6966 30432 7030 30436
rect 7046 30492 7110 30496
rect 7046 30436 7050 30492
rect 7050 30436 7106 30492
rect 7106 30436 7110 30492
rect 7046 30432 7110 30436
rect 7126 30492 7190 30496
rect 7126 30436 7130 30492
rect 7130 30436 7186 30492
rect 7186 30436 7190 30492
rect 7126 30432 7190 30436
rect 12820 30492 12884 30496
rect 12820 30436 12824 30492
rect 12824 30436 12880 30492
rect 12880 30436 12884 30492
rect 12820 30432 12884 30436
rect 12900 30492 12964 30496
rect 12900 30436 12904 30492
rect 12904 30436 12960 30492
rect 12960 30436 12964 30492
rect 12900 30432 12964 30436
rect 12980 30492 13044 30496
rect 12980 30436 12984 30492
rect 12984 30436 13040 30492
rect 13040 30436 13044 30492
rect 12980 30432 13044 30436
rect 13060 30492 13124 30496
rect 13060 30436 13064 30492
rect 13064 30436 13120 30492
rect 13120 30436 13124 30492
rect 13060 30432 13124 30436
rect 18754 30492 18818 30496
rect 18754 30436 18758 30492
rect 18758 30436 18814 30492
rect 18814 30436 18818 30492
rect 18754 30432 18818 30436
rect 18834 30492 18898 30496
rect 18834 30436 18838 30492
rect 18838 30436 18894 30492
rect 18894 30436 18898 30492
rect 18834 30432 18898 30436
rect 18914 30492 18978 30496
rect 18914 30436 18918 30492
rect 18918 30436 18974 30492
rect 18974 30436 18978 30492
rect 18914 30432 18978 30436
rect 18994 30492 19058 30496
rect 18994 30436 18998 30492
rect 18998 30436 19054 30492
rect 19054 30436 19058 30492
rect 18994 30432 19058 30436
rect 24688 30492 24752 30496
rect 24688 30436 24692 30492
rect 24692 30436 24748 30492
rect 24748 30436 24752 30492
rect 24688 30432 24752 30436
rect 24768 30492 24832 30496
rect 24768 30436 24772 30492
rect 24772 30436 24828 30492
rect 24828 30436 24832 30492
rect 24768 30432 24832 30436
rect 24848 30492 24912 30496
rect 24848 30436 24852 30492
rect 24852 30436 24908 30492
rect 24908 30436 24912 30492
rect 24848 30432 24912 30436
rect 24928 30492 24992 30496
rect 24928 30436 24932 30492
rect 24932 30436 24988 30492
rect 24988 30436 24992 30492
rect 24928 30432 24992 30436
rect 4844 30288 4908 30292
rect 4844 30232 4858 30288
rect 4858 30232 4908 30288
rect 4844 30228 4908 30232
rect 12020 30364 12084 30428
rect 14412 30364 14476 30428
rect 3188 29956 3252 30020
rect 5212 30016 5276 30020
rect 6132 30092 6196 30156
rect 10364 30092 10428 30156
rect 5212 29960 5226 30016
rect 5226 29960 5276 30016
rect 5212 29956 5276 29960
rect 10364 30016 10428 30020
rect 10364 29960 10414 30016
rect 10414 29960 10428 30016
rect 10364 29956 10428 29960
rect 3919 29948 3983 29952
rect 3919 29892 3923 29948
rect 3923 29892 3979 29948
rect 3979 29892 3983 29948
rect 3919 29888 3983 29892
rect 3999 29948 4063 29952
rect 3999 29892 4003 29948
rect 4003 29892 4059 29948
rect 4059 29892 4063 29948
rect 3999 29888 4063 29892
rect 4079 29948 4143 29952
rect 4079 29892 4083 29948
rect 4083 29892 4139 29948
rect 4139 29892 4143 29948
rect 4079 29888 4143 29892
rect 4159 29948 4223 29952
rect 4159 29892 4163 29948
rect 4163 29892 4219 29948
rect 4219 29892 4223 29948
rect 4159 29888 4223 29892
rect 9853 29948 9917 29952
rect 9853 29892 9857 29948
rect 9857 29892 9913 29948
rect 9913 29892 9917 29948
rect 9853 29888 9917 29892
rect 9933 29948 9997 29952
rect 9933 29892 9937 29948
rect 9937 29892 9993 29948
rect 9993 29892 9997 29948
rect 9933 29888 9997 29892
rect 10013 29948 10077 29952
rect 10013 29892 10017 29948
rect 10017 29892 10073 29948
rect 10073 29892 10077 29948
rect 10013 29888 10077 29892
rect 10093 29948 10157 29952
rect 10093 29892 10097 29948
rect 10097 29892 10153 29948
rect 10153 29892 10157 29948
rect 10093 29888 10157 29892
rect 15787 29948 15851 29952
rect 15787 29892 15791 29948
rect 15791 29892 15847 29948
rect 15847 29892 15851 29948
rect 15787 29888 15851 29892
rect 15867 29948 15931 29952
rect 15867 29892 15871 29948
rect 15871 29892 15927 29948
rect 15927 29892 15931 29948
rect 15867 29888 15931 29892
rect 15947 29948 16011 29952
rect 15947 29892 15951 29948
rect 15951 29892 16007 29948
rect 16007 29892 16011 29948
rect 15947 29888 16011 29892
rect 16027 29948 16091 29952
rect 16027 29892 16031 29948
rect 16031 29892 16087 29948
rect 16087 29892 16091 29948
rect 16027 29888 16091 29892
rect 21721 29948 21785 29952
rect 21721 29892 21725 29948
rect 21725 29892 21781 29948
rect 21781 29892 21785 29948
rect 21721 29888 21785 29892
rect 21801 29948 21865 29952
rect 21801 29892 21805 29948
rect 21805 29892 21861 29948
rect 21861 29892 21865 29948
rect 21801 29888 21865 29892
rect 21881 29948 21945 29952
rect 21881 29892 21885 29948
rect 21885 29892 21941 29948
rect 21941 29892 21945 29948
rect 21881 29888 21945 29892
rect 21961 29948 22025 29952
rect 21961 29892 21965 29948
rect 21965 29892 22021 29948
rect 22021 29892 22025 29948
rect 21961 29888 22025 29892
rect 7972 29820 8036 29884
rect 2452 29548 2516 29612
rect 2084 29472 2148 29476
rect 2084 29416 2134 29472
rect 2134 29416 2148 29472
rect 2084 29412 2148 29416
rect 6886 29404 6950 29408
rect 6886 29348 6890 29404
rect 6890 29348 6946 29404
rect 6946 29348 6950 29404
rect 6886 29344 6950 29348
rect 6966 29404 7030 29408
rect 6966 29348 6970 29404
rect 6970 29348 7026 29404
rect 7026 29348 7030 29404
rect 6966 29344 7030 29348
rect 7046 29404 7110 29408
rect 7046 29348 7050 29404
rect 7050 29348 7106 29404
rect 7106 29348 7110 29404
rect 7046 29344 7110 29348
rect 7126 29404 7190 29408
rect 7126 29348 7130 29404
rect 7130 29348 7186 29404
rect 7186 29348 7190 29404
rect 7126 29344 7190 29348
rect 12820 29404 12884 29408
rect 12820 29348 12824 29404
rect 12824 29348 12880 29404
rect 12880 29348 12884 29404
rect 12820 29344 12884 29348
rect 12900 29404 12964 29408
rect 12900 29348 12904 29404
rect 12904 29348 12960 29404
rect 12960 29348 12964 29404
rect 12900 29344 12964 29348
rect 12980 29404 13044 29408
rect 12980 29348 12984 29404
rect 12984 29348 13040 29404
rect 13040 29348 13044 29404
rect 12980 29344 13044 29348
rect 13060 29404 13124 29408
rect 13060 29348 13064 29404
rect 13064 29348 13120 29404
rect 13120 29348 13124 29404
rect 13060 29344 13124 29348
rect 18754 29404 18818 29408
rect 18754 29348 18758 29404
rect 18758 29348 18814 29404
rect 18814 29348 18818 29404
rect 18754 29344 18818 29348
rect 18834 29404 18898 29408
rect 18834 29348 18838 29404
rect 18838 29348 18894 29404
rect 18894 29348 18898 29404
rect 18834 29344 18898 29348
rect 18914 29404 18978 29408
rect 18914 29348 18918 29404
rect 18918 29348 18974 29404
rect 18974 29348 18978 29404
rect 18914 29344 18978 29348
rect 18994 29404 19058 29408
rect 18994 29348 18998 29404
rect 18998 29348 19054 29404
rect 19054 29348 19058 29404
rect 18994 29344 19058 29348
rect 24688 29404 24752 29408
rect 24688 29348 24692 29404
rect 24692 29348 24748 29404
rect 24748 29348 24752 29404
rect 24688 29344 24752 29348
rect 24768 29404 24832 29408
rect 24768 29348 24772 29404
rect 24772 29348 24828 29404
rect 24828 29348 24832 29404
rect 24768 29344 24832 29348
rect 24848 29404 24912 29408
rect 24848 29348 24852 29404
rect 24852 29348 24908 29404
rect 24908 29348 24912 29404
rect 24848 29344 24912 29348
rect 24928 29404 24992 29408
rect 24928 29348 24932 29404
rect 24932 29348 24988 29404
rect 24988 29348 24992 29404
rect 24928 29344 24992 29348
rect 4292 29276 4356 29340
rect 14780 29004 14844 29068
rect 18460 29004 18524 29068
rect 3919 28860 3983 28864
rect 3919 28804 3923 28860
rect 3923 28804 3979 28860
rect 3979 28804 3983 28860
rect 3919 28800 3983 28804
rect 3999 28860 4063 28864
rect 3999 28804 4003 28860
rect 4003 28804 4059 28860
rect 4059 28804 4063 28860
rect 3999 28800 4063 28804
rect 4079 28860 4143 28864
rect 4079 28804 4083 28860
rect 4083 28804 4139 28860
rect 4139 28804 4143 28860
rect 4079 28800 4143 28804
rect 4159 28860 4223 28864
rect 4159 28804 4163 28860
rect 4163 28804 4219 28860
rect 4219 28804 4223 28860
rect 4159 28800 4223 28804
rect 9853 28860 9917 28864
rect 9853 28804 9857 28860
rect 9857 28804 9913 28860
rect 9913 28804 9917 28860
rect 9853 28800 9917 28804
rect 9933 28860 9997 28864
rect 9933 28804 9937 28860
rect 9937 28804 9993 28860
rect 9993 28804 9997 28860
rect 9933 28800 9997 28804
rect 10013 28860 10077 28864
rect 10013 28804 10017 28860
rect 10017 28804 10073 28860
rect 10073 28804 10077 28860
rect 10013 28800 10077 28804
rect 10093 28860 10157 28864
rect 10093 28804 10097 28860
rect 10097 28804 10153 28860
rect 10153 28804 10157 28860
rect 10093 28800 10157 28804
rect 15787 28860 15851 28864
rect 15787 28804 15791 28860
rect 15791 28804 15847 28860
rect 15847 28804 15851 28860
rect 15787 28800 15851 28804
rect 15867 28860 15931 28864
rect 15867 28804 15871 28860
rect 15871 28804 15927 28860
rect 15927 28804 15931 28860
rect 15867 28800 15931 28804
rect 15947 28860 16011 28864
rect 15947 28804 15951 28860
rect 15951 28804 16007 28860
rect 16007 28804 16011 28860
rect 15947 28800 16011 28804
rect 16027 28860 16091 28864
rect 16027 28804 16031 28860
rect 16031 28804 16087 28860
rect 16087 28804 16091 28860
rect 16027 28800 16091 28804
rect 9628 28792 9692 28796
rect 9628 28736 9678 28792
rect 9678 28736 9692 28792
rect 9628 28732 9692 28736
rect 21721 28860 21785 28864
rect 21721 28804 21725 28860
rect 21725 28804 21781 28860
rect 21781 28804 21785 28860
rect 21721 28800 21785 28804
rect 21801 28860 21865 28864
rect 21801 28804 21805 28860
rect 21805 28804 21861 28860
rect 21861 28804 21865 28860
rect 21801 28800 21865 28804
rect 21881 28860 21945 28864
rect 21881 28804 21885 28860
rect 21885 28804 21941 28860
rect 21941 28804 21945 28860
rect 21881 28800 21945 28804
rect 21961 28860 22025 28864
rect 21961 28804 21965 28860
rect 21965 28804 22021 28860
rect 22021 28804 22025 28860
rect 21961 28800 22025 28804
rect 2084 28460 2148 28524
rect 19196 28596 19260 28660
rect 6886 28316 6950 28320
rect 6886 28260 6890 28316
rect 6890 28260 6946 28316
rect 6946 28260 6950 28316
rect 6886 28256 6950 28260
rect 6966 28316 7030 28320
rect 6966 28260 6970 28316
rect 6970 28260 7026 28316
rect 7026 28260 7030 28316
rect 6966 28256 7030 28260
rect 7046 28316 7110 28320
rect 7046 28260 7050 28316
rect 7050 28260 7106 28316
rect 7106 28260 7110 28316
rect 7046 28256 7110 28260
rect 7126 28316 7190 28320
rect 7126 28260 7130 28316
rect 7130 28260 7186 28316
rect 7186 28260 7190 28316
rect 7126 28256 7190 28260
rect 12820 28316 12884 28320
rect 12820 28260 12824 28316
rect 12824 28260 12880 28316
rect 12880 28260 12884 28316
rect 12820 28256 12884 28260
rect 12900 28316 12964 28320
rect 12900 28260 12904 28316
rect 12904 28260 12960 28316
rect 12960 28260 12964 28316
rect 12900 28256 12964 28260
rect 12980 28316 13044 28320
rect 12980 28260 12984 28316
rect 12984 28260 13040 28316
rect 13040 28260 13044 28316
rect 12980 28256 13044 28260
rect 13060 28316 13124 28320
rect 13060 28260 13064 28316
rect 13064 28260 13120 28316
rect 13120 28260 13124 28316
rect 13060 28256 13124 28260
rect 18754 28316 18818 28320
rect 18754 28260 18758 28316
rect 18758 28260 18814 28316
rect 18814 28260 18818 28316
rect 18754 28256 18818 28260
rect 18834 28316 18898 28320
rect 18834 28260 18838 28316
rect 18838 28260 18894 28316
rect 18894 28260 18898 28316
rect 18834 28256 18898 28260
rect 18914 28316 18978 28320
rect 18914 28260 18918 28316
rect 18918 28260 18974 28316
rect 18974 28260 18978 28316
rect 18914 28256 18978 28260
rect 18994 28316 19058 28320
rect 18994 28260 18998 28316
rect 18998 28260 19054 28316
rect 19054 28260 19058 28316
rect 18994 28256 19058 28260
rect 24688 28316 24752 28320
rect 24688 28260 24692 28316
rect 24692 28260 24748 28316
rect 24748 28260 24752 28316
rect 24688 28256 24752 28260
rect 24768 28316 24832 28320
rect 24768 28260 24772 28316
rect 24772 28260 24828 28316
rect 24828 28260 24832 28316
rect 24768 28256 24832 28260
rect 24848 28316 24912 28320
rect 24848 28260 24852 28316
rect 24852 28260 24908 28316
rect 24908 28260 24912 28316
rect 24848 28256 24912 28260
rect 24928 28316 24992 28320
rect 24928 28260 24932 28316
rect 24932 28260 24988 28316
rect 24988 28260 24992 28316
rect 24928 28256 24992 28260
rect 1716 27916 1780 27980
rect 10732 27780 10796 27844
rect 3919 27772 3983 27776
rect 3919 27716 3923 27772
rect 3923 27716 3979 27772
rect 3979 27716 3983 27772
rect 3919 27712 3983 27716
rect 3999 27772 4063 27776
rect 3999 27716 4003 27772
rect 4003 27716 4059 27772
rect 4059 27716 4063 27772
rect 3999 27712 4063 27716
rect 4079 27772 4143 27776
rect 4079 27716 4083 27772
rect 4083 27716 4139 27772
rect 4139 27716 4143 27772
rect 4079 27712 4143 27716
rect 4159 27772 4223 27776
rect 4159 27716 4163 27772
rect 4163 27716 4219 27772
rect 4219 27716 4223 27772
rect 4159 27712 4223 27716
rect 9853 27772 9917 27776
rect 9853 27716 9857 27772
rect 9857 27716 9913 27772
rect 9913 27716 9917 27772
rect 9853 27712 9917 27716
rect 9933 27772 9997 27776
rect 9933 27716 9937 27772
rect 9937 27716 9993 27772
rect 9993 27716 9997 27772
rect 9933 27712 9997 27716
rect 10013 27772 10077 27776
rect 10013 27716 10017 27772
rect 10017 27716 10073 27772
rect 10073 27716 10077 27772
rect 10013 27712 10077 27716
rect 10093 27772 10157 27776
rect 10093 27716 10097 27772
rect 10097 27716 10153 27772
rect 10153 27716 10157 27772
rect 10093 27712 10157 27716
rect 15787 27772 15851 27776
rect 15787 27716 15791 27772
rect 15791 27716 15847 27772
rect 15847 27716 15851 27772
rect 15787 27712 15851 27716
rect 15867 27772 15931 27776
rect 15867 27716 15871 27772
rect 15871 27716 15927 27772
rect 15927 27716 15931 27772
rect 15867 27712 15931 27716
rect 15947 27772 16011 27776
rect 15947 27716 15951 27772
rect 15951 27716 16007 27772
rect 16007 27716 16011 27772
rect 15947 27712 16011 27716
rect 16027 27772 16091 27776
rect 16027 27716 16031 27772
rect 16031 27716 16087 27772
rect 16087 27716 16091 27772
rect 16027 27712 16091 27716
rect 21721 27772 21785 27776
rect 21721 27716 21725 27772
rect 21725 27716 21781 27772
rect 21781 27716 21785 27772
rect 21721 27712 21785 27716
rect 21801 27772 21865 27776
rect 21801 27716 21805 27772
rect 21805 27716 21861 27772
rect 21861 27716 21865 27772
rect 21801 27712 21865 27716
rect 21881 27772 21945 27776
rect 21881 27716 21885 27772
rect 21885 27716 21941 27772
rect 21941 27716 21945 27772
rect 21881 27712 21945 27716
rect 21961 27772 22025 27776
rect 21961 27716 21965 27772
rect 21965 27716 22021 27772
rect 22021 27716 22025 27772
rect 21961 27712 22025 27716
rect 5396 27644 5460 27708
rect 10548 27568 10612 27572
rect 10548 27512 10562 27568
rect 10562 27512 10612 27568
rect 10548 27508 10612 27512
rect 6886 27228 6950 27232
rect 6886 27172 6890 27228
rect 6890 27172 6946 27228
rect 6946 27172 6950 27228
rect 6886 27168 6950 27172
rect 6966 27228 7030 27232
rect 6966 27172 6970 27228
rect 6970 27172 7026 27228
rect 7026 27172 7030 27228
rect 6966 27168 7030 27172
rect 7046 27228 7110 27232
rect 7046 27172 7050 27228
rect 7050 27172 7106 27228
rect 7106 27172 7110 27228
rect 7046 27168 7110 27172
rect 7126 27228 7190 27232
rect 7126 27172 7130 27228
rect 7130 27172 7186 27228
rect 7186 27172 7190 27228
rect 7126 27168 7190 27172
rect 12820 27228 12884 27232
rect 12820 27172 12824 27228
rect 12824 27172 12880 27228
rect 12880 27172 12884 27228
rect 12820 27168 12884 27172
rect 12900 27228 12964 27232
rect 12900 27172 12904 27228
rect 12904 27172 12960 27228
rect 12960 27172 12964 27228
rect 12900 27168 12964 27172
rect 12980 27228 13044 27232
rect 12980 27172 12984 27228
rect 12984 27172 13040 27228
rect 13040 27172 13044 27228
rect 12980 27168 13044 27172
rect 13060 27228 13124 27232
rect 13060 27172 13064 27228
rect 13064 27172 13120 27228
rect 13120 27172 13124 27228
rect 13060 27168 13124 27172
rect 18754 27228 18818 27232
rect 18754 27172 18758 27228
rect 18758 27172 18814 27228
rect 18814 27172 18818 27228
rect 18754 27168 18818 27172
rect 18834 27228 18898 27232
rect 18834 27172 18838 27228
rect 18838 27172 18894 27228
rect 18894 27172 18898 27228
rect 18834 27168 18898 27172
rect 18914 27228 18978 27232
rect 18914 27172 18918 27228
rect 18918 27172 18974 27228
rect 18974 27172 18978 27228
rect 18914 27168 18978 27172
rect 18994 27228 19058 27232
rect 18994 27172 18998 27228
rect 18998 27172 19054 27228
rect 19054 27172 19058 27228
rect 18994 27168 19058 27172
rect 24688 27228 24752 27232
rect 24688 27172 24692 27228
rect 24692 27172 24748 27228
rect 24748 27172 24752 27228
rect 24688 27168 24752 27172
rect 24768 27228 24832 27232
rect 24768 27172 24772 27228
rect 24772 27172 24828 27228
rect 24828 27172 24832 27228
rect 24768 27168 24832 27172
rect 24848 27228 24912 27232
rect 24848 27172 24852 27228
rect 24852 27172 24908 27228
rect 24908 27172 24912 27228
rect 24848 27168 24912 27172
rect 24928 27228 24992 27232
rect 24928 27172 24932 27228
rect 24932 27172 24988 27228
rect 24988 27172 24992 27228
rect 24928 27168 24992 27172
rect 2268 27100 2332 27164
rect 17356 26888 17420 26892
rect 17356 26832 17406 26888
rect 17406 26832 17420 26888
rect 17356 26828 17420 26832
rect 3919 26684 3983 26688
rect 3919 26628 3923 26684
rect 3923 26628 3979 26684
rect 3979 26628 3983 26684
rect 3919 26624 3983 26628
rect 3999 26684 4063 26688
rect 3999 26628 4003 26684
rect 4003 26628 4059 26684
rect 4059 26628 4063 26684
rect 3999 26624 4063 26628
rect 4079 26684 4143 26688
rect 4079 26628 4083 26684
rect 4083 26628 4139 26684
rect 4139 26628 4143 26684
rect 4079 26624 4143 26628
rect 4159 26684 4223 26688
rect 4159 26628 4163 26684
rect 4163 26628 4219 26684
rect 4219 26628 4223 26684
rect 4159 26624 4223 26628
rect 9853 26684 9917 26688
rect 9853 26628 9857 26684
rect 9857 26628 9913 26684
rect 9913 26628 9917 26684
rect 9853 26624 9917 26628
rect 9933 26684 9997 26688
rect 9933 26628 9937 26684
rect 9937 26628 9993 26684
rect 9993 26628 9997 26684
rect 9933 26624 9997 26628
rect 10013 26684 10077 26688
rect 10013 26628 10017 26684
rect 10017 26628 10073 26684
rect 10073 26628 10077 26684
rect 10013 26624 10077 26628
rect 10093 26684 10157 26688
rect 10093 26628 10097 26684
rect 10097 26628 10153 26684
rect 10153 26628 10157 26684
rect 10093 26624 10157 26628
rect 15787 26684 15851 26688
rect 15787 26628 15791 26684
rect 15791 26628 15847 26684
rect 15847 26628 15851 26684
rect 15787 26624 15851 26628
rect 15867 26684 15931 26688
rect 15867 26628 15871 26684
rect 15871 26628 15927 26684
rect 15927 26628 15931 26684
rect 15867 26624 15931 26628
rect 15947 26684 16011 26688
rect 15947 26628 15951 26684
rect 15951 26628 16007 26684
rect 16007 26628 16011 26684
rect 15947 26624 16011 26628
rect 16027 26684 16091 26688
rect 16027 26628 16031 26684
rect 16031 26628 16087 26684
rect 16087 26628 16091 26684
rect 16027 26624 16091 26628
rect 21721 26684 21785 26688
rect 21721 26628 21725 26684
rect 21725 26628 21781 26684
rect 21781 26628 21785 26684
rect 21721 26624 21785 26628
rect 21801 26684 21865 26688
rect 21801 26628 21805 26684
rect 21805 26628 21861 26684
rect 21861 26628 21865 26684
rect 21801 26624 21865 26628
rect 21881 26684 21945 26688
rect 21881 26628 21885 26684
rect 21885 26628 21941 26684
rect 21941 26628 21945 26684
rect 21881 26624 21945 26628
rect 21961 26684 22025 26688
rect 21961 26628 21965 26684
rect 21965 26628 22021 26684
rect 22021 26628 22025 26684
rect 21961 26624 22025 26628
rect 6684 26556 6748 26620
rect 13676 26420 13740 26484
rect 10732 26148 10796 26212
rect 15332 26148 15396 26212
rect 16436 26208 16500 26212
rect 16436 26152 16450 26208
rect 16450 26152 16500 26208
rect 16436 26148 16500 26152
rect 19196 26148 19260 26212
rect 20116 26148 20180 26212
rect 6886 26140 6950 26144
rect 6886 26084 6890 26140
rect 6890 26084 6946 26140
rect 6946 26084 6950 26140
rect 6886 26080 6950 26084
rect 6966 26140 7030 26144
rect 6966 26084 6970 26140
rect 6970 26084 7026 26140
rect 7026 26084 7030 26140
rect 6966 26080 7030 26084
rect 7046 26140 7110 26144
rect 7046 26084 7050 26140
rect 7050 26084 7106 26140
rect 7106 26084 7110 26140
rect 7046 26080 7110 26084
rect 7126 26140 7190 26144
rect 7126 26084 7130 26140
rect 7130 26084 7186 26140
rect 7186 26084 7190 26140
rect 7126 26080 7190 26084
rect 12820 26140 12884 26144
rect 12820 26084 12824 26140
rect 12824 26084 12880 26140
rect 12880 26084 12884 26140
rect 12820 26080 12884 26084
rect 12900 26140 12964 26144
rect 12900 26084 12904 26140
rect 12904 26084 12960 26140
rect 12960 26084 12964 26140
rect 12900 26080 12964 26084
rect 12980 26140 13044 26144
rect 12980 26084 12984 26140
rect 12984 26084 13040 26140
rect 13040 26084 13044 26140
rect 12980 26080 13044 26084
rect 13060 26140 13124 26144
rect 13060 26084 13064 26140
rect 13064 26084 13120 26140
rect 13120 26084 13124 26140
rect 13060 26080 13124 26084
rect 18754 26140 18818 26144
rect 18754 26084 18758 26140
rect 18758 26084 18814 26140
rect 18814 26084 18818 26140
rect 18754 26080 18818 26084
rect 18834 26140 18898 26144
rect 18834 26084 18838 26140
rect 18838 26084 18894 26140
rect 18894 26084 18898 26140
rect 18834 26080 18898 26084
rect 18914 26140 18978 26144
rect 18914 26084 18918 26140
rect 18918 26084 18974 26140
rect 18974 26084 18978 26140
rect 18914 26080 18978 26084
rect 18994 26140 19058 26144
rect 18994 26084 18998 26140
rect 18998 26084 19054 26140
rect 19054 26084 19058 26140
rect 18994 26080 19058 26084
rect 24688 26140 24752 26144
rect 24688 26084 24692 26140
rect 24692 26084 24748 26140
rect 24748 26084 24752 26140
rect 24688 26080 24752 26084
rect 24768 26140 24832 26144
rect 24768 26084 24772 26140
rect 24772 26084 24828 26140
rect 24828 26084 24832 26140
rect 24768 26080 24832 26084
rect 24848 26140 24912 26144
rect 24848 26084 24852 26140
rect 24852 26084 24908 26140
rect 24908 26084 24912 26140
rect 24848 26080 24912 26084
rect 24928 26140 24992 26144
rect 24928 26084 24932 26140
rect 24932 26084 24988 26140
rect 24988 26084 24992 26140
rect 24928 26080 24992 26084
rect 3919 25596 3983 25600
rect 3919 25540 3923 25596
rect 3923 25540 3979 25596
rect 3979 25540 3983 25596
rect 3919 25536 3983 25540
rect 3999 25596 4063 25600
rect 3999 25540 4003 25596
rect 4003 25540 4059 25596
rect 4059 25540 4063 25596
rect 3999 25536 4063 25540
rect 4079 25596 4143 25600
rect 4079 25540 4083 25596
rect 4083 25540 4139 25596
rect 4139 25540 4143 25596
rect 4079 25536 4143 25540
rect 4159 25596 4223 25600
rect 4159 25540 4163 25596
rect 4163 25540 4219 25596
rect 4219 25540 4223 25596
rect 4159 25536 4223 25540
rect 9853 25596 9917 25600
rect 9853 25540 9857 25596
rect 9857 25540 9913 25596
rect 9913 25540 9917 25596
rect 9853 25536 9917 25540
rect 9933 25596 9997 25600
rect 9933 25540 9937 25596
rect 9937 25540 9993 25596
rect 9993 25540 9997 25596
rect 9933 25536 9997 25540
rect 10013 25596 10077 25600
rect 10013 25540 10017 25596
rect 10017 25540 10073 25596
rect 10073 25540 10077 25596
rect 10013 25536 10077 25540
rect 10093 25596 10157 25600
rect 10093 25540 10097 25596
rect 10097 25540 10153 25596
rect 10153 25540 10157 25596
rect 10093 25536 10157 25540
rect 15787 25596 15851 25600
rect 15787 25540 15791 25596
rect 15791 25540 15847 25596
rect 15847 25540 15851 25596
rect 15787 25536 15851 25540
rect 15867 25596 15931 25600
rect 15867 25540 15871 25596
rect 15871 25540 15927 25596
rect 15927 25540 15931 25596
rect 15867 25536 15931 25540
rect 15947 25596 16011 25600
rect 15947 25540 15951 25596
rect 15951 25540 16007 25596
rect 16007 25540 16011 25596
rect 15947 25536 16011 25540
rect 16027 25596 16091 25600
rect 16027 25540 16031 25596
rect 16031 25540 16087 25596
rect 16087 25540 16091 25596
rect 16027 25536 16091 25540
rect 21721 25596 21785 25600
rect 21721 25540 21725 25596
rect 21725 25540 21781 25596
rect 21781 25540 21785 25596
rect 21721 25536 21785 25540
rect 21801 25596 21865 25600
rect 21801 25540 21805 25596
rect 21805 25540 21861 25596
rect 21861 25540 21865 25596
rect 21801 25536 21865 25540
rect 21881 25596 21945 25600
rect 21881 25540 21885 25596
rect 21885 25540 21941 25596
rect 21941 25540 21945 25596
rect 21881 25536 21945 25540
rect 21961 25596 22025 25600
rect 21961 25540 21965 25596
rect 21965 25540 22021 25596
rect 22021 25540 22025 25596
rect 21961 25536 22025 25540
rect 14780 25332 14844 25396
rect 4844 25196 4908 25260
rect 7604 25060 7668 25124
rect 6886 25052 6950 25056
rect 6886 24996 6890 25052
rect 6890 24996 6946 25052
rect 6946 24996 6950 25052
rect 6886 24992 6950 24996
rect 6966 25052 7030 25056
rect 6966 24996 6970 25052
rect 6970 24996 7026 25052
rect 7026 24996 7030 25052
rect 6966 24992 7030 24996
rect 7046 25052 7110 25056
rect 7046 24996 7050 25052
rect 7050 24996 7106 25052
rect 7106 24996 7110 25052
rect 7046 24992 7110 24996
rect 7126 25052 7190 25056
rect 7126 24996 7130 25052
rect 7130 24996 7186 25052
rect 7186 24996 7190 25052
rect 7126 24992 7190 24996
rect 12820 25052 12884 25056
rect 12820 24996 12824 25052
rect 12824 24996 12880 25052
rect 12880 24996 12884 25052
rect 12820 24992 12884 24996
rect 12900 25052 12964 25056
rect 12900 24996 12904 25052
rect 12904 24996 12960 25052
rect 12960 24996 12964 25052
rect 12900 24992 12964 24996
rect 12980 25052 13044 25056
rect 12980 24996 12984 25052
rect 12984 24996 13040 25052
rect 13040 24996 13044 25052
rect 12980 24992 13044 24996
rect 13060 25052 13124 25056
rect 13060 24996 13064 25052
rect 13064 24996 13120 25052
rect 13120 24996 13124 25052
rect 13060 24992 13124 24996
rect 18754 25052 18818 25056
rect 18754 24996 18758 25052
rect 18758 24996 18814 25052
rect 18814 24996 18818 25052
rect 18754 24992 18818 24996
rect 18834 25052 18898 25056
rect 18834 24996 18838 25052
rect 18838 24996 18894 25052
rect 18894 24996 18898 25052
rect 18834 24992 18898 24996
rect 18914 25052 18978 25056
rect 18914 24996 18918 25052
rect 18918 24996 18974 25052
rect 18974 24996 18978 25052
rect 18914 24992 18978 24996
rect 18994 25052 19058 25056
rect 18994 24996 18998 25052
rect 18998 24996 19054 25052
rect 19054 24996 19058 25052
rect 18994 24992 19058 24996
rect 24688 25052 24752 25056
rect 24688 24996 24692 25052
rect 24692 24996 24748 25052
rect 24748 24996 24752 25052
rect 24688 24992 24752 24996
rect 24768 25052 24832 25056
rect 24768 24996 24772 25052
rect 24772 24996 24828 25052
rect 24828 24996 24832 25052
rect 24768 24992 24832 24996
rect 24848 25052 24912 25056
rect 24848 24996 24852 25052
rect 24852 24996 24908 25052
rect 24908 24996 24912 25052
rect 24848 24992 24912 24996
rect 24928 25052 24992 25056
rect 24928 24996 24932 25052
rect 24932 24996 24988 25052
rect 24988 24996 24992 25052
rect 24928 24992 24992 24996
rect 9076 24924 9140 24988
rect 10364 24924 10428 24988
rect 2084 24788 2148 24852
rect 4660 24788 4724 24852
rect 3919 24508 3983 24512
rect 3919 24452 3923 24508
rect 3923 24452 3979 24508
rect 3979 24452 3983 24508
rect 3919 24448 3983 24452
rect 3999 24508 4063 24512
rect 3999 24452 4003 24508
rect 4003 24452 4059 24508
rect 4059 24452 4063 24508
rect 3999 24448 4063 24452
rect 4079 24508 4143 24512
rect 4079 24452 4083 24508
rect 4083 24452 4139 24508
rect 4139 24452 4143 24508
rect 4079 24448 4143 24452
rect 4159 24508 4223 24512
rect 4159 24452 4163 24508
rect 4163 24452 4219 24508
rect 4219 24452 4223 24508
rect 4159 24448 4223 24452
rect 9853 24508 9917 24512
rect 9853 24452 9857 24508
rect 9857 24452 9913 24508
rect 9913 24452 9917 24508
rect 9853 24448 9917 24452
rect 9933 24508 9997 24512
rect 9933 24452 9937 24508
rect 9937 24452 9993 24508
rect 9993 24452 9997 24508
rect 9933 24448 9997 24452
rect 10013 24508 10077 24512
rect 10013 24452 10017 24508
rect 10017 24452 10073 24508
rect 10073 24452 10077 24508
rect 10013 24448 10077 24452
rect 10093 24508 10157 24512
rect 10093 24452 10097 24508
rect 10097 24452 10153 24508
rect 10153 24452 10157 24508
rect 10093 24448 10157 24452
rect 15787 24508 15851 24512
rect 15787 24452 15791 24508
rect 15791 24452 15847 24508
rect 15847 24452 15851 24508
rect 15787 24448 15851 24452
rect 15867 24508 15931 24512
rect 15867 24452 15871 24508
rect 15871 24452 15927 24508
rect 15927 24452 15931 24508
rect 15867 24448 15931 24452
rect 15947 24508 16011 24512
rect 15947 24452 15951 24508
rect 15951 24452 16007 24508
rect 16007 24452 16011 24508
rect 15947 24448 16011 24452
rect 16027 24508 16091 24512
rect 16027 24452 16031 24508
rect 16031 24452 16087 24508
rect 16087 24452 16091 24508
rect 16027 24448 16091 24452
rect 21721 24508 21785 24512
rect 21721 24452 21725 24508
rect 21725 24452 21781 24508
rect 21781 24452 21785 24508
rect 21721 24448 21785 24452
rect 21801 24508 21865 24512
rect 21801 24452 21805 24508
rect 21805 24452 21861 24508
rect 21861 24452 21865 24508
rect 21801 24448 21865 24452
rect 21881 24508 21945 24512
rect 21881 24452 21885 24508
rect 21885 24452 21941 24508
rect 21941 24452 21945 24508
rect 21881 24448 21945 24452
rect 21961 24508 22025 24512
rect 21961 24452 21965 24508
rect 21965 24452 22021 24508
rect 22021 24452 22025 24508
rect 21961 24448 22025 24452
rect 10916 24380 10980 24444
rect 24164 24108 24228 24172
rect 6886 23964 6950 23968
rect 6886 23908 6890 23964
rect 6890 23908 6946 23964
rect 6946 23908 6950 23964
rect 6886 23904 6950 23908
rect 6966 23964 7030 23968
rect 6966 23908 6970 23964
rect 6970 23908 7026 23964
rect 7026 23908 7030 23964
rect 6966 23904 7030 23908
rect 7046 23964 7110 23968
rect 7046 23908 7050 23964
rect 7050 23908 7106 23964
rect 7106 23908 7110 23964
rect 7046 23904 7110 23908
rect 7126 23964 7190 23968
rect 7126 23908 7130 23964
rect 7130 23908 7186 23964
rect 7186 23908 7190 23964
rect 7126 23904 7190 23908
rect 12820 23964 12884 23968
rect 12820 23908 12824 23964
rect 12824 23908 12880 23964
rect 12880 23908 12884 23964
rect 12820 23904 12884 23908
rect 12900 23964 12964 23968
rect 12900 23908 12904 23964
rect 12904 23908 12960 23964
rect 12960 23908 12964 23964
rect 12900 23904 12964 23908
rect 12980 23964 13044 23968
rect 12980 23908 12984 23964
rect 12984 23908 13040 23964
rect 13040 23908 13044 23964
rect 12980 23904 13044 23908
rect 13060 23964 13124 23968
rect 13060 23908 13064 23964
rect 13064 23908 13120 23964
rect 13120 23908 13124 23964
rect 13060 23904 13124 23908
rect 18754 23964 18818 23968
rect 18754 23908 18758 23964
rect 18758 23908 18814 23964
rect 18814 23908 18818 23964
rect 18754 23904 18818 23908
rect 18834 23964 18898 23968
rect 18834 23908 18838 23964
rect 18838 23908 18894 23964
rect 18894 23908 18898 23964
rect 18834 23904 18898 23908
rect 18914 23964 18978 23968
rect 18914 23908 18918 23964
rect 18918 23908 18974 23964
rect 18974 23908 18978 23964
rect 18914 23904 18978 23908
rect 18994 23964 19058 23968
rect 18994 23908 18998 23964
rect 18998 23908 19054 23964
rect 19054 23908 19058 23964
rect 18994 23904 19058 23908
rect 24688 23964 24752 23968
rect 24688 23908 24692 23964
rect 24692 23908 24748 23964
rect 24748 23908 24752 23964
rect 24688 23904 24752 23908
rect 24768 23964 24832 23968
rect 24768 23908 24772 23964
rect 24772 23908 24828 23964
rect 24828 23908 24832 23964
rect 24768 23904 24832 23908
rect 24848 23964 24912 23968
rect 24848 23908 24852 23964
rect 24852 23908 24908 23964
rect 24908 23908 24912 23964
rect 24848 23904 24912 23908
rect 24928 23964 24992 23968
rect 24928 23908 24932 23964
rect 24932 23908 24988 23964
rect 24988 23908 24992 23964
rect 24928 23904 24992 23908
rect 7604 23896 7668 23900
rect 7604 23840 7618 23896
rect 7618 23840 7668 23896
rect 7604 23836 7668 23840
rect 4660 23428 4724 23492
rect 7420 23428 7484 23492
rect 12204 23428 12268 23492
rect 3919 23420 3983 23424
rect 3919 23364 3923 23420
rect 3923 23364 3979 23420
rect 3979 23364 3983 23420
rect 3919 23360 3983 23364
rect 3999 23420 4063 23424
rect 3999 23364 4003 23420
rect 4003 23364 4059 23420
rect 4059 23364 4063 23420
rect 3999 23360 4063 23364
rect 4079 23420 4143 23424
rect 4079 23364 4083 23420
rect 4083 23364 4139 23420
rect 4139 23364 4143 23420
rect 4079 23360 4143 23364
rect 4159 23420 4223 23424
rect 4159 23364 4163 23420
rect 4163 23364 4219 23420
rect 4219 23364 4223 23420
rect 4159 23360 4223 23364
rect 9853 23420 9917 23424
rect 9853 23364 9857 23420
rect 9857 23364 9913 23420
rect 9913 23364 9917 23420
rect 9853 23360 9917 23364
rect 9933 23420 9997 23424
rect 9933 23364 9937 23420
rect 9937 23364 9993 23420
rect 9993 23364 9997 23420
rect 9933 23360 9997 23364
rect 10013 23420 10077 23424
rect 10013 23364 10017 23420
rect 10017 23364 10073 23420
rect 10073 23364 10077 23420
rect 10013 23360 10077 23364
rect 10093 23420 10157 23424
rect 10093 23364 10097 23420
rect 10097 23364 10153 23420
rect 10153 23364 10157 23420
rect 10093 23360 10157 23364
rect 5396 23352 5460 23356
rect 5396 23296 5446 23352
rect 5446 23296 5460 23352
rect 5396 23292 5460 23296
rect 14044 23428 14108 23492
rect 16620 23488 16684 23492
rect 16620 23432 16670 23488
rect 16670 23432 16684 23488
rect 16620 23428 16684 23432
rect 16988 23428 17052 23492
rect 22508 23428 22572 23492
rect 15787 23420 15851 23424
rect 15787 23364 15791 23420
rect 15791 23364 15847 23420
rect 15847 23364 15851 23420
rect 15787 23360 15851 23364
rect 15867 23420 15931 23424
rect 15867 23364 15871 23420
rect 15871 23364 15927 23420
rect 15927 23364 15931 23420
rect 15867 23360 15931 23364
rect 15947 23420 16011 23424
rect 15947 23364 15951 23420
rect 15951 23364 16007 23420
rect 16007 23364 16011 23420
rect 15947 23360 16011 23364
rect 16027 23420 16091 23424
rect 16027 23364 16031 23420
rect 16031 23364 16087 23420
rect 16087 23364 16091 23420
rect 16027 23360 16091 23364
rect 21721 23420 21785 23424
rect 21721 23364 21725 23420
rect 21725 23364 21781 23420
rect 21781 23364 21785 23420
rect 21721 23360 21785 23364
rect 21801 23420 21865 23424
rect 21801 23364 21805 23420
rect 21805 23364 21861 23420
rect 21861 23364 21865 23420
rect 21801 23360 21865 23364
rect 21881 23420 21945 23424
rect 21881 23364 21885 23420
rect 21885 23364 21941 23420
rect 21941 23364 21945 23420
rect 21881 23360 21945 23364
rect 21961 23420 22025 23424
rect 21961 23364 21965 23420
rect 21965 23364 22021 23420
rect 22021 23364 22025 23420
rect 21961 23360 22025 23364
rect 6886 22876 6950 22880
rect 6886 22820 6890 22876
rect 6890 22820 6946 22876
rect 6946 22820 6950 22876
rect 6886 22816 6950 22820
rect 6966 22876 7030 22880
rect 6966 22820 6970 22876
rect 6970 22820 7026 22876
rect 7026 22820 7030 22876
rect 6966 22816 7030 22820
rect 7046 22876 7110 22880
rect 7046 22820 7050 22876
rect 7050 22820 7106 22876
rect 7106 22820 7110 22876
rect 7046 22816 7110 22820
rect 7126 22876 7190 22880
rect 7126 22820 7130 22876
rect 7130 22820 7186 22876
rect 7186 22820 7190 22876
rect 7126 22816 7190 22820
rect 12820 22876 12884 22880
rect 12820 22820 12824 22876
rect 12824 22820 12880 22876
rect 12880 22820 12884 22876
rect 12820 22816 12884 22820
rect 12900 22876 12964 22880
rect 12900 22820 12904 22876
rect 12904 22820 12960 22876
rect 12960 22820 12964 22876
rect 12900 22816 12964 22820
rect 12980 22876 13044 22880
rect 12980 22820 12984 22876
rect 12984 22820 13040 22876
rect 13040 22820 13044 22876
rect 12980 22816 13044 22820
rect 13060 22876 13124 22880
rect 13060 22820 13064 22876
rect 13064 22820 13120 22876
rect 13120 22820 13124 22876
rect 13060 22816 13124 22820
rect 18754 22876 18818 22880
rect 18754 22820 18758 22876
rect 18758 22820 18814 22876
rect 18814 22820 18818 22876
rect 18754 22816 18818 22820
rect 18834 22876 18898 22880
rect 18834 22820 18838 22876
rect 18838 22820 18894 22876
rect 18894 22820 18898 22876
rect 18834 22816 18898 22820
rect 18914 22876 18978 22880
rect 18914 22820 18918 22876
rect 18918 22820 18974 22876
rect 18974 22820 18978 22876
rect 18914 22816 18978 22820
rect 18994 22876 19058 22880
rect 18994 22820 18998 22876
rect 18998 22820 19054 22876
rect 19054 22820 19058 22876
rect 18994 22816 19058 22820
rect 24688 22876 24752 22880
rect 24688 22820 24692 22876
rect 24692 22820 24748 22876
rect 24748 22820 24752 22876
rect 24688 22816 24752 22820
rect 24768 22876 24832 22880
rect 24768 22820 24772 22876
rect 24772 22820 24828 22876
rect 24828 22820 24832 22876
rect 24768 22816 24832 22820
rect 24848 22876 24912 22880
rect 24848 22820 24852 22876
rect 24852 22820 24908 22876
rect 24908 22820 24912 22876
rect 24848 22816 24912 22820
rect 24928 22876 24992 22880
rect 24928 22820 24932 22876
rect 24932 22820 24988 22876
rect 24988 22820 24992 22876
rect 24928 22816 24992 22820
rect 10364 22748 10428 22812
rect 2636 22068 2700 22132
rect 22692 22612 22756 22676
rect 3919 22332 3983 22336
rect 3919 22276 3923 22332
rect 3923 22276 3979 22332
rect 3979 22276 3983 22332
rect 3919 22272 3983 22276
rect 3999 22332 4063 22336
rect 3999 22276 4003 22332
rect 4003 22276 4059 22332
rect 4059 22276 4063 22332
rect 3999 22272 4063 22276
rect 4079 22332 4143 22336
rect 4079 22276 4083 22332
rect 4083 22276 4139 22332
rect 4139 22276 4143 22332
rect 4079 22272 4143 22276
rect 4159 22332 4223 22336
rect 4159 22276 4163 22332
rect 4163 22276 4219 22332
rect 4219 22276 4223 22332
rect 4159 22272 4223 22276
rect 9853 22332 9917 22336
rect 9853 22276 9857 22332
rect 9857 22276 9913 22332
rect 9913 22276 9917 22332
rect 9853 22272 9917 22276
rect 9933 22332 9997 22336
rect 9933 22276 9937 22332
rect 9937 22276 9993 22332
rect 9993 22276 9997 22332
rect 9933 22272 9997 22276
rect 10013 22332 10077 22336
rect 10013 22276 10017 22332
rect 10017 22276 10073 22332
rect 10073 22276 10077 22332
rect 10013 22272 10077 22276
rect 10093 22332 10157 22336
rect 10093 22276 10097 22332
rect 10097 22276 10153 22332
rect 10153 22276 10157 22332
rect 10093 22272 10157 22276
rect 15787 22332 15851 22336
rect 15787 22276 15791 22332
rect 15791 22276 15847 22332
rect 15847 22276 15851 22332
rect 15787 22272 15851 22276
rect 15867 22332 15931 22336
rect 15867 22276 15871 22332
rect 15871 22276 15927 22332
rect 15927 22276 15931 22332
rect 15867 22272 15931 22276
rect 15947 22332 16011 22336
rect 15947 22276 15951 22332
rect 15951 22276 16007 22332
rect 16007 22276 16011 22332
rect 15947 22272 16011 22276
rect 16027 22332 16091 22336
rect 16027 22276 16031 22332
rect 16031 22276 16087 22332
rect 16087 22276 16091 22332
rect 16027 22272 16091 22276
rect 21721 22332 21785 22336
rect 21721 22276 21725 22332
rect 21725 22276 21781 22332
rect 21781 22276 21785 22332
rect 21721 22272 21785 22276
rect 21801 22332 21865 22336
rect 21801 22276 21805 22332
rect 21805 22276 21861 22332
rect 21861 22276 21865 22332
rect 21801 22272 21865 22276
rect 21881 22332 21945 22336
rect 21881 22276 21885 22332
rect 21885 22276 21941 22332
rect 21941 22276 21945 22332
rect 21881 22272 21945 22276
rect 21961 22332 22025 22336
rect 21961 22276 21965 22332
rect 21965 22276 22021 22332
rect 22021 22276 22025 22332
rect 21961 22272 22025 22276
rect 11836 22264 11900 22268
rect 11836 22208 11886 22264
rect 11886 22208 11900 22264
rect 11836 22204 11900 22208
rect 12388 22204 12452 22268
rect 13492 22204 13556 22268
rect 5396 22068 5460 22132
rect 18092 22068 18156 22132
rect 21404 22068 21468 22132
rect 22508 22068 22572 22132
rect 4476 21992 4540 21996
rect 4476 21936 4490 21992
rect 4490 21936 4540 21992
rect 4476 21932 4540 21936
rect 13492 21932 13556 21996
rect 6886 21788 6950 21792
rect 6886 21732 6890 21788
rect 6890 21732 6946 21788
rect 6946 21732 6950 21788
rect 6886 21728 6950 21732
rect 6966 21788 7030 21792
rect 6966 21732 6970 21788
rect 6970 21732 7026 21788
rect 7026 21732 7030 21788
rect 6966 21728 7030 21732
rect 7046 21788 7110 21792
rect 7046 21732 7050 21788
rect 7050 21732 7106 21788
rect 7106 21732 7110 21788
rect 7046 21728 7110 21732
rect 7126 21788 7190 21792
rect 7126 21732 7130 21788
rect 7130 21732 7186 21788
rect 7186 21732 7190 21788
rect 7126 21728 7190 21732
rect 12820 21788 12884 21792
rect 12820 21732 12824 21788
rect 12824 21732 12880 21788
rect 12880 21732 12884 21788
rect 12820 21728 12884 21732
rect 12900 21788 12964 21792
rect 12900 21732 12904 21788
rect 12904 21732 12960 21788
rect 12960 21732 12964 21788
rect 12900 21728 12964 21732
rect 12980 21788 13044 21792
rect 12980 21732 12984 21788
rect 12984 21732 13040 21788
rect 13040 21732 13044 21788
rect 12980 21728 13044 21732
rect 13060 21788 13124 21792
rect 13060 21732 13064 21788
rect 13064 21732 13120 21788
rect 13120 21732 13124 21788
rect 13060 21728 13124 21732
rect 18754 21788 18818 21792
rect 18754 21732 18758 21788
rect 18758 21732 18814 21788
rect 18814 21732 18818 21788
rect 18754 21728 18818 21732
rect 18834 21788 18898 21792
rect 18834 21732 18838 21788
rect 18838 21732 18894 21788
rect 18894 21732 18898 21788
rect 18834 21728 18898 21732
rect 18914 21788 18978 21792
rect 18914 21732 18918 21788
rect 18918 21732 18974 21788
rect 18974 21732 18978 21788
rect 18914 21728 18978 21732
rect 18994 21788 19058 21792
rect 18994 21732 18998 21788
rect 18998 21732 19054 21788
rect 19054 21732 19058 21788
rect 18994 21728 19058 21732
rect 24688 21788 24752 21792
rect 24688 21732 24692 21788
rect 24692 21732 24748 21788
rect 24748 21732 24752 21788
rect 24688 21728 24752 21732
rect 24768 21788 24832 21792
rect 24768 21732 24772 21788
rect 24772 21732 24828 21788
rect 24828 21732 24832 21788
rect 24768 21728 24832 21732
rect 24848 21788 24912 21792
rect 24848 21732 24852 21788
rect 24852 21732 24908 21788
rect 24908 21732 24912 21788
rect 24848 21728 24912 21732
rect 24928 21788 24992 21792
rect 24928 21732 24932 21788
rect 24932 21732 24988 21788
rect 24988 21732 24992 21788
rect 24928 21728 24992 21732
rect 9076 21524 9140 21588
rect 21036 21524 21100 21588
rect 6684 21388 6748 21452
rect 12204 21252 12268 21316
rect 14596 21252 14660 21316
rect 3919 21244 3983 21248
rect 3919 21188 3923 21244
rect 3923 21188 3979 21244
rect 3979 21188 3983 21244
rect 3919 21184 3983 21188
rect 3999 21244 4063 21248
rect 3999 21188 4003 21244
rect 4003 21188 4059 21244
rect 4059 21188 4063 21244
rect 3999 21184 4063 21188
rect 4079 21244 4143 21248
rect 4079 21188 4083 21244
rect 4083 21188 4139 21244
rect 4139 21188 4143 21244
rect 4079 21184 4143 21188
rect 4159 21244 4223 21248
rect 4159 21188 4163 21244
rect 4163 21188 4219 21244
rect 4219 21188 4223 21244
rect 4159 21184 4223 21188
rect 9853 21244 9917 21248
rect 9853 21188 9857 21244
rect 9857 21188 9913 21244
rect 9913 21188 9917 21244
rect 9853 21184 9917 21188
rect 9933 21244 9997 21248
rect 9933 21188 9937 21244
rect 9937 21188 9993 21244
rect 9993 21188 9997 21244
rect 9933 21184 9997 21188
rect 10013 21244 10077 21248
rect 10013 21188 10017 21244
rect 10017 21188 10073 21244
rect 10073 21188 10077 21244
rect 10013 21184 10077 21188
rect 10093 21244 10157 21248
rect 10093 21188 10097 21244
rect 10097 21188 10153 21244
rect 10153 21188 10157 21244
rect 10093 21184 10157 21188
rect 15787 21244 15851 21248
rect 15787 21188 15791 21244
rect 15791 21188 15847 21244
rect 15847 21188 15851 21244
rect 15787 21184 15851 21188
rect 15867 21244 15931 21248
rect 15867 21188 15871 21244
rect 15871 21188 15927 21244
rect 15927 21188 15931 21244
rect 15867 21184 15931 21188
rect 15947 21244 16011 21248
rect 15947 21188 15951 21244
rect 15951 21188 16007 21244
rect 16007 21188 16011 21244
rect 15947 21184 16011 21188
rect 16027 21244 16091 21248
rect 16027 21188 16031 21244
rect 16031 21188 16087 21244
rect 16087 21188 16091 21244
rect 16027 21184 16091 21188
rect 21721 21244 21785 21248
rect 21721 21188 21725 21244
rect 21725 21188 21781 21244
rect 21781 21188 21785 21244
rect 21721 21184 21785 21188
rect 21801 21244 21865 21248
rect 21801 21188 21805 21244
rect 21805 21188 21861 21244
rect 21861 21188 21865 21244
rect 21801 21184 21865 21188
rect 21881 21244 21945 21248
rect 21881 21188 21885 21244
rect 21885 21188 21941 21244
rect 21941 21188 21945 21244
rect 21881 21184 21945 21188
rect 21961 21244 22025 21248
rect 21961 21188 21965 21244
rect 21965 21188 22021 21244
rect 22021 21188 22025 21244
rect 21961 21184 22025 21188
rect 24164 21116 24228 21180
rect 1348 20844 1412 20908
rect 12572 20844 12636 20908
rect 16620 20844 16684 20908
rect 6886 20700 6950 20704
rect 6886 20644 6890 20700
rect 6890 20644 6946 20700
rect 6946 20644 6950 20700
rect 6886 20640 6950 20644
rect 6966 20700 7030 20704
rect 6966 20644 6970 20700
rect 6970 20644 7026 20700
rect 7026 20644 7030 20700
rect 6966 20640 7030 20644
rect 7046 20700 7110 20704
rect 7046 20644 7050 20700
rect 7050 20644 7106 20700
rect 7106 20644 7110 20700
rect 7046 20640 7110 20644
rect 7126 20700 7190 20704
rect 7126 20644 7130 20700
rect 7130 20644 7186 20700
rect 7186 20644 7190 20700
rect 7126 20640 7190 20644
rect 12820 20700 12884 20704
rect 12820 20644 12824 20700
rect 12824 20644 12880 20700
rect 12880 20644 12884 20700
rect 12820 20640 12884 20644
rect 12900 20700 12964 20704
rect 12900 20644 12904 20700
rect 12904 20644 12960 20700
rect 12960 20644 12964 20700
rect 12900 20640 12964 20644
rect 12980 20700 13044 20704
rect 12980 20644 12984 20700
rect 12984 20644 13040 20700
rect 13040 20644 13044 20700
rect 12980 20640 13044 20644
rect 13060 20700 13124 20704
rect 13060 20644 13064 20700
rect 13064 20644 13120 20700
rect 13120 20644 13124 20700
rect 13060 20640 13124 20644
rect 18754 20700 18818 20704
rect 18754 20644 18758 20700
rect 18758 20644 18814 20700
rect 18814 20644 18818 20700
rect 18754 20640 18818 20644
rect 18834 20700 18898 20704
rect 18834 20644 18838 20700
rect 18838 20644 18894 20700
rect 18894 20644 18898 20700
rect 18834 20640 18898 20644
rect 18914 20700 18978 20704
rect 18914 20644 18918 20700
rect 18918 20644 18974 20700
rect 18974 20644 18978 20700
rect 18914 20640 18978 20644
rect 18994 20700 19058 20704
rect 18994 20644 18998 20700
rect 18998 20644 19054 20700
rect 19054 20644 19058 20700
rect 18994 20640 19058 20644
rect 24688 20700 24752 20704
rect 24688 20644 24692 20700
rect 24692 20644 24748 20700
rect 24748 20644 24752 20700
rect 24688 20640 24752 20644
rect 24768 20700 24832 20704
rect 24768 20644 24772 20700
rect 24772 20644 24828 20700
rect 24828 20644 24832 20700
rect 24768 20640 24832 20644
rect 24848 20700 24912 20704
rect 24848 20644 24852 20700
rect 24852 20644 24908 20700
rect 24908 20644 24912 20700
rect 24848 20640 24912 20644
rect 24928 20700 24992 20704
rect 24928 20644 24932 20700
rect 24932 20644 24988 20700
rect 24988 20644 24992 20700
rect 24928 20640 24992 20644
rect 16436 20436 16500 20500
rect 17356 20436 17420 20500
rect 22876 20164 22940 20228
rect 3919 20156 3983 20160
rect 3919 20100 3923 20156
rect 3923 20100 3979 20156
rect 3979 20100 3983 20156
rect 3919 20096 3983 20100
rect 3999 20156 4063 20160
rect 3999 20100 4003 20156
rect 4003 20100 4059 20156
rect 4059 20100 4063 20156
rect 3999 20096 4063 20100
rect 4079 20156 4143 20160
rect 4079 20100 4083 20156
rect 4083 20100 4139 20156
rect 4139 20100 4143 20156
rect 4079 20096 4143 20100
rect 4159 20156 4223 20160
rect 4159 20100 4163 20156
rect 4163 20100 4219 20156
rect 4219 20100 4223 20156
rect 4159 20096 4223 20100
rect 9853 20156 9917 20160
rect 9853 20100 9857 20156
rect 9857 20100 9913 20156
rect 9913 20100 9917 20156
rect 9853 20096 9917 20100
rect 9933 20156 9997 20160
rect 9933 20100 9937 20156
rect 9937 20100 9993 20156
rect 9993 20100 9997 20156
rect 9933 20096 9997 20100
rect 10013 20156 10077 20160
rect 10013 20100 10017 20156
rect 10017 20100 10073 20156
rect 10073 20100 10077 20156
rect 10013 20096 10077 20100
rect 10093 20156 10157 20160
rect 10093 20100 10097 20156
rect 10097 20100 10153 20156
rect 10153 20100 10157 20156
rect 10093 20096 10157 20100
rect 15787 20156 15851 20160
rect 15787 20100 15791 20156
rect 15791 20100 15847 20156
rect 15847 20100 15851 20156
rect 15787 20096 15851 20100
rect 15867 20156 15931 20160
rect 15867 20100 15871 20156
rect 15871 20100 15927 20156
rect 15927 20100 15931 20156
rect 15867 20096 15931 20100
rect 15947 20156 16011 20160
rect 15947 20100 15951 20156
rect 15951 20100 16007 20156
rect 16007 20100 16011 20156
rect 15947 20096 16011 20100
rect 16027 20156 16091 20160
rect 16027 20100 16031 20156
rect 16031 20100 16087 20156
rect 16087 20100 16091 20156
rect 16027 20096 16091 20100
rect 21721 20156 21785 20160
rect 21721 20100 21725 20156
rect 21725 20100 21781 20156
rect 21781 20100 21785 20156
rect 21721 20096 21785 20100
rect 21801 20156 21865 20160
rect 21801 20100 21805 20156
rect 21805 20100 21861 20156
rect 21861 20100 21865 20156
rect 21801 20096 21865 20100
rect 21881 20156 21945 20160
rect 21881 20100 21885 20156
rect 21885 20100 21941 20156
rect 21941 20100 21945 20156
rect 21881 20096 21945 20100
rect 21961 20156 22025 20160
rect 21961 20100 21965 20156
rect 21965 20100 22021 20156
rect 22021 20100 22025 20156
rect 21961 20096 22025 20100
rect 5212 19892 5276 19956
rect 3556 19680 3620 19684
rect 3556 19624 3570 19680
rect 3570 19624 3620 19680
rect 3556 19620 3620 19624
rect 6132 19680 6196 19684
rect 6132 19624 6146 19680
rect 6146 19624 6196 19680
rect 6132 19620 6196 19624
rect 10364 19816 10428 19820
rect 10364 19760 10378 19816
rect 10378 19760 10428 19816
rect 10364 19756 10428 19760
rect 10916 19620 10980 19684
rect 6886 19612 6950 19616
rect 6886 19556 6890 19612
rect 6890 19556 6946 19612
rect 6946 19556 6950 19612
rect 6886 19552 6950 19556
rect 6966 19612 7030 19616
rect 6966 19556 6970 19612
rect 6970 19556 7026 19612
rect 7026 19556 7030 19612
rect 6966 19552 7030 19556
rect 7046 19612 7110 19616
rect 7046 19556 7050 19612
rect 7050 19556 7106 19612
rect 7106 19556 7110 19612
rect 7046 19552 7110 19556
rect 7126 19612 7190 19616
rect 7126 19556 7130 19612
rect 7130 19556 7186 19612
rect 7186 19556 7190 19612
rect 7126 19552 7190 19556
rect 12820 19612 12884 19616
rect 12820 19556 12824 19612
rect 12824 19556 12880 19612
rect 12880 19556 12884 19612
rect 12820 19552 12884 19556
rect 12900 19612 12964 19616
rect 12900 19556 12904 19612
rect 12904 19556 12960 19612
rect 12960 19556 12964 19612
rect 12900 19552 12964 19556
rect 12980 19612 13044 19616
rect 12980 19556 12984 19612
rect 12984 19556 13040 19612
rect 13040 19556 13044 19612
rect 12980 19552 13044 19556
rect 13060 19612 13124 19616
rect 13060 19556 13064 19612
rect 13064 19556 13120 19612
rect 13120 19556 13124 19612
rect 13060 19552 13124 19556
rect 18754 19612 18818 19616
rect 18754 19556 18758 19612
rect 18758 19556 18814 19612
rect 18814 19556 18818 19612
rect 18754 19552 18818 19556
rect 18834 19612 18898 19616
rect 18834 19556 18838 19612
rect 18838 19556 18894 19612
rect 18894 19556 18898 19612
rect 18834 19552 18898 19556
rect 18914 19612 18978 19616
rect 18914 19556 18918 19612
rect 18918 19556 18974 19612
rect 18974 19556 18978 19612
rect 18914 19552 18978 19556
rect 18994 19612 19058 19616
rect 18994 19556 18998 19612
rect 18998 19556 19054 19612
rect 19054 19556 19058 19612
rect 18994 19552 19058 19556
rect 24688 19612 24752 19616
rect 24688 19556 24692 19612
rect 24692 19556 24748 19612
rect 24748 19556 24752 19612
rect 24688 19552 24752 19556
rect 24768 19612 24832 19616
rect 24768 19556 24772 19612
rect 24772 19556 24828 19612
rect 24828 19556 24832 19612
rect 24768 19552 24832 19556
rect 24848 19612 24912 19616
rect 24848 19556 24852 19612
rect 24852 19556 24908 19612
rect 24908 19556 24912 19612
rect 24848 19552 24912 19556
rect 24928 19612 24992 19616
rect 24928 19556 24932 19612
rect 24932 19556 24988 19612
rect 24988 19556 24992 19612
rect 24928 19552 24992 19556
rect 13676 19544 13740 19548
rect 13676 19488 13726 19544
rect 13726 19488 13740 19544
rect 13676 19484 13740 19488
rect 5212 19348 5276 19412
rect 13860 19348 13924 19412
rect 3919 19068 3983 19072
rect 3919 19012 3923 19068
rect 3923 19012 3979 19068
rect 3979 19012 3983 19068
rect 3919 19008 3983 19012
rect 3999 19068 4063 19072
rect 3999 19012 4003 19068
rect 4003 19012 4059 19068
rect 4059 19012 4063 19068
rect 3999 19008 4063 19012
rect 4079 19068 4143 19072
rect 4079 19012 4083 19068
rect 4083 19012 4139 19068
rect 4139 19012 4143 19068
rect 4079 19008 4143 19012
rect 4159 19068 4223 19072
rect 4159 19012 4163 19068
rect 4163 19012 4219 19068
rect 4219 19012 4223 19068
rect 4159 19008 4223 19012
rect 4476 19212 4540 19276
rect 9853 19068 9917 19072
rect 9853 19012 9857 19068
rect 9857 19012 9913 19068
rect 9913 19012 9917 19068
rect 9853 19008 9917 19012
rect 9933 19068 9997 19072
rect 9933 19012 9937 19068
rect 9937 19012 9993 19068
rect 9993 19012 9997 19068
rect 9933 19008 9997 19012
rect 10013 19068 10077 19072
rect 10013 19012 10017 19068
rect 10017 19012 10073 19068
rect 10073 19012 10077 19068
rect 10013 19008 10077 19012
rect 10093 19068 10157 19072
rect 10093 19012 10097 19068
rect 10097 19012 10153 19068
rect 10153 19012 10157 19068
rect 10093 19008 10157 19012
rect 15787 19068 15851 19072
rect 15787 19012 15791 19068
rect 15791 19012 15847 19068
rect 15847 19012 15851 19068
rect 15787 19008 15851 19012
rect 15867 19068 15931 19072
rect 15867 19012 15871 19068
rect 15871 19012 15927 19068
rect 15927 19012 15931 19068
rect 15867 19008 15931 19012
rect 15947 19068 16011 19072
rect 15947 19012 15951 19068
rect 15951 19012 16007 19068
rect 16007 19012 16011 19068
rect 15947 19008 16011 19012
rect 16027 19068 16091 19072
rect 16027 19012 16031 19068
rect 16031 19012 16087 19068
rect 16087 19012 16091 19068
rect 16027 19008 16091 19012
rect 21721 19068 21785 19072
rect 21721 19012 21725 19068
rect 21725 19012 21781 19068
rect 21781 19012 21785 19068
rect 21721 19008 21785 19012
rect 21801 19068 21865 19072
rect 21801 19012 21805 19068
rect 21805 19012 21861 19068
rect 21861 19012 21865 19068
rect 21801 19008 21865 19012
rect 21881 19068 21945 19072
rect 21881 19012 21885 19068
rect 21885 19012 21941 19068
rect 21941 19012 21945 19068
rect 21881 19008 21945 19012
rect 21961 19068 22025 19072
rect 21961 19012 21965 19068
rect 21965 19012 22021 19068
rect 22021 19012 22025 19068
rect 21961 19008 22025 19012
rect 10548 18804 10612 18868
rect 6886 18524 6950 18528
rect 6886 18468 6890 18524
rect 6890 18468 6946 18524
rect 6946 18468 6950 18524
rect 6886 18464 6950 18468
rect 6966 18524 7030 18528
rect 6966 18468 6970 18524
rect 6970 18468 7026 18524
rect 7026 18468 7030 18524
rect 6966 18464 7030 18468
rect 7046 18524 7110 18528
rect 7046 18468 7050 18524
rect 7050 18468 7106 18524
rect 7106 18468 7110 18524
rect 7046 18464 7110 18468
rect 7126 18524 7190 18528
rect 7126 18468 7130 18524
rect 7130 18468 7186 18524
rect 7186 18468 7190 18524
rect 7126 18464 7190 18468
rect 12820 18524 12884 18528
rect 12820 18468 12824 18524
rect 12824 18468 12880 18524
rect 12880 18468 12884 18524
rect 12820 18464 12884 18468
rect 12900 18524 12964 18528
rect 12900 18468 12904 18524
rect 12904 18468 12960 18524
rect 12960 18468 12964 18524
rect 12900 18464 12964 18468
rect 12980 18524 13044 18528
rect 12980 18468 12984 18524
rect 12984 18468 13040 18524
rect 13040 18468 13044 18524
rect 12980 18464 13044 18468
rect 13060 18524 13124 18528
rect 13060 18468 13064 18524
rect 13064 18468 13120 18524
rect 13120 18468 13124 18524
rect 13060 18464 13124 18468
rect 18754 18524 18818 18528
rect 18754 18468 18758 18524
rect 18758 18468 18814 18524
rect 18814 18468 18818 18524
rect 18754 18464 18818 18468
rect 18834 18524 18898 18528
rect 18834 18468 18838 18524
rect 18838 18468 18894 18524
rect 18894 18468 18898 18524
rect 18834 18464 18898 18468
rect 18914 18524 18978 18528
rect 18914 18468 18918 18524
rect 18918 18468 18974 18524
rect 18974 18468 18978 18524
rect 18914 18464 18978 18468
rect 18994 18524 19058 18528
rect 18994 18468 18998 18524
rect 18998 18468 19054 18524
rect 19054 18468 19058 18524
rect 18994 18464 19058 18468
rect 24688 18524 24752 18528
rect 24688 18468 24692 18524
rect 24692 18468 24748 18524
rect 24748 18468 24752 18524
rect 24688 18464 24752 18468
rect 24768 18524 24832 18528
rect 24768 18468 24772 18524
rect 24772 18468 24828 18524
rect 24828 18468 24832 18524
rect 24768 18464 24832 18468
rect 24848 18524 24912 18528
rect 24848 18468 24852 18524
rect 24852 18468 24908 18524
rect 24908 18468 24912 18524
rect 24848 18464 24912 18468
rect 24928 18524 24992 18528
rect 24928 18468 24932 18524
rect 24932 18468 24988 18524
rect 24988 18468 24992 18524
rect 24928 18464 24992 18468
rect 9628 18124 9692 18188
rect 16436 18124 16500 18188
rect 21404 18048 21468 18052
rect 21404 17992 21418 18048
rect 21418 17992 21468 18048
rect 21404 17988 21468 17992
rect 3919 17980 3983 17984
rect 3919 17924 3923 17980
rect 3923 17924 3979 17980
rect 3979 17924 3983 17980
rect 3919 17920 3983 17924
rect 3999 17980 4063 17984
rect 3999 17924 4003 17980
rect 4003 17924 4059 17980
rect 4059 17924 4063 17980
rect 3999 17920 4063 17924
rect 4079 17980 4143 17984
rect 4079 17924 4083 17980
rect 4083 17924 4139 17980
rect 4139 17924 4143 17980
rect 4079 17920 4143 17924
rect 4159 17980 4223 17984
rect 4159 17924 4163 17980
rect 4163 17924 4219 17980
rect 4219 17924 4223 17980
rect 4159 17920 4223 17924
rect 9853 17980 9917 17984
rect 9853 17924 9857 17980
rect 9857 17924 9913 17980
rect 9913 17924 9917 17980
rect 9853 17920 9917 17924
rect 9933 17980 9997 17984
rect 9933 17924 9937 17980
rect 9937 17924 9993 17980
rect 9993 17924 9997 17980
rect 9933 17920 9997 17924
rect 10013 17980 10077 17984
rect 10013 17924 10017 17980
rect 10017 17924 10073 17980
rect 10073 17924 10077 17980
rect 10013 17920 10077 17924
rect 10093 17980 10157 17984
rect 10093 17924 10097 17980
rect 10097 17924 10153 17980
rect 10153 17924 10157 17980
rect 10093 17920 10157 17924
rect 15787 17980 15851 17984
rect 15787 17924 15791 17980
rect 15791 17924 15847 17980
rect 15847 17924 15851 17980
rect 15787 17920 15851 17924
rect 15867 17980 15931 17984
rect 15867 17924 15871 17980
rect 15871 17924 15927 17980
rect 15927 17924 15931 17980
rect 15867 17920 15931 17924
rect 15947 17980 16011 17984
rect 15947 17924 15951 17980
rect 15951 17924 16007 17980
rect 16007 17924 16011 17980
rect 15947 17920 16011 17924
rect 16027 17980 16091 17984
rect 16027 17924 16031 17980
rect 16031 17924 16087 17980
rect 16087 17924 16091 17980
rect 16027 17920 16091 17924
rect 21721 17980 21785 17984
rect 21721 17924 21725 17980
rect 21725 17924 21781 17980
rect 21781 17924 21785 17980
rect 21721 17920 21785 17924
rect 21801 17980 21865 17984
rect 21801 17924 21805 17980
rect 21805 17924 21861 17980
rect 21861 17924 21865 17980
rect 21801 17920 21865 17924
rect 21881 17980 21945 17984
rect 21881 17924 21885 17980
rect 21885 17924 21941 17980
rect 21941 17924 21945 17980
rect 21881 17920 21945 17924
rect 21961 17980 22025 17984
rect 21961 17924 21965 17980
rect 21965 17924 22021 17980
rect 22021 17924 22025 17980
rect 21961 17920 22025 17924
rect 11468 17716 11532 17780
rect 13492 17716 13556 17780
rect 11652 17580 11716 17644
rect 13492 17580 13556 17644
rect 6886 17436 6950 17440
rect 6886 17380 6890 17436
rect 6890 17380 6946 17436
rect 6946 17380 6950 17436
rect 6886 17376 6950 17380
rect 6966 17436 7030 17440
rect 6966 17380 6970 17436
rect 6970 17380 7026 17436
rect 7026 17380 7030 17436
rect 6966 17376 7030 17380
rect 7046 17436 7110 17440
rect 7046 17380 7050 17436
rect 7050 17380 7106 17436
rect 7106 17380 7110 17436
rect 7046 17376 7110 17380
rect 7126 17436 7190 17440
rect 7126 17380 7130 17436
rect 7130 17380 7186 17436
rect 7186 17380 7190 17436
rect 7126 17376 7190 17380
rect 12820 17436 12884 17440
rect 12820 17380 12824 17436
rect 12824 17380 12880 17436
rect 12880 17380 12884 17436
rect 12820 17376 12884 17380
rect 12900 17436 12964 17440
rect 12900 17380 12904 17436
rect 12904 17380 12960 17436
rect 12960 17380 12964 17436
rect 12900 17376 12964 17380
rect 12980 17436 13044 17440
rect 12980 17380 12984 17436
rect 12984 17380 13040 17436
rect 13040 17380 13044 17436
rect 12980 17376 13044 17380
rect 13060 17436 13124 17440
rect 13060 17380 13064 17436
rect 13064 17380 13120 17436
rect 13120 17380 13124 17436
rect 13060 17376 13124 17380
rect 18754 17436 18818 17440
rect 18754 17380 18758 17436
rect 18758 17380 18814 17436
rect 18814 17380 18818 17436
rect 18754 17376 18818 17380
rect 18834 17436 18898 17440
rect 18834 17380 18838 17436
rect 18838 17380 18894 17436
rect 18894 17380 18898 17436
rect 18834 17376 18898 17380
rect 18914 17436 18978 17440
rect 18914 17380 18918 17436
rect 18918 17380 18974 17436
rect 18974 17380 18978 17436
rect 18914 17376 18978 17380
rect 18994 17436 19058 17440
rect 18994 17380 18998 17436
rect 18998 17380 19054 17436
rect 19054 17380 19058 17436
rect 18994 17376 19058 17380
rect 24688 17436 24752 17440
rect 24688 17380 24692 17436
rect 24692 17380 24748 17436
rect 24748 17380 24752 17436
rect 24688 17376 24752 17380
rect 24768 17436 24832 17440
rect 24768 17380 24772 17436
rect 24772 17380 24828 17436
rect 24828 17380 24832 17436
rect 24768 17376 24832 17380
rect 24848 17436 24912 17440
rect 24848 17380 24852 17436
rect 24852 17380 24908 17436
rect 24908 17380 24912 17436
rect 24848 17376 24912 17380
rect 24928 17436 24992 17440
rect 24928 17380 24932 17436
rect 24932 17380 24988 17436
rect 24988 17380 24992 17436
rect 24928 17376 24992 17380
rect 19748 17308 19812 17372
rect 19932 17172 19996 17236
rect 3919 16892 3983 16896
rect 3919 16836 3923 16892
rect 3923 16836 3979 16892
rect 3979 16836 3983 16892
rect 3919 16832 3983 16836
rect 3999 16892 4063 16896
rect 3999 16836 4003 16892
rect 4003 16836 4059 16892
rect 4059 16836 4063 16892
rect 3999 16832 4063 16836
rect 4079 16892 4143 16896
rect 4079 16836 4083 16892
rect 4083 16836 4139 16892
rect 4139 16836 4143 16892
rect 4079 16832 4143 16836
rect 4159 16892 4223 16896
rect 4159 16836 4163 16892
rect 4163 16836 4219 16892
rect 4219 16836 4223 16892
rect 4159 16832 4223 16836
rect 9853 16892 9917 16896
rect 9853 16836 9857 16892
rect 9857 16836 9913 16892
rect 9913 16836 9917 16892
rect 9853 16832 9917 16836
rect 9933 16892 9997 16896
rect 9933 16836 9937 16892
rect 9937 16836 9993 16892
rect 9993 16836 9997 16892
rect 9933 16832 9997 16836
rect 10013 16892 10077 16896
rect 10013 16836 10017 16892
rect 10017 16836 10073 16892
rect 10073 16836 10077 16892
rect 10013 16832 10077 16836
rect 10093 16892 10157 16896
rect 10093 16836 10097 16892
rect 10097 16836 10153 16892
rect 10153 16836 10157 16892
rect 10093 16832 10157 16836
rect 15787 16892 15851 16896
rect 15787 16836 15791 16892
rect 15791 16836 15847 16892
rect 15847 16836 15851 16892
rect 15787 16832 15851 16836
rect 15867 16892 15931 16896
rect 15867 16836 15871 16892
rect 15871 16836 15927 16892
rect 15927 16836 15931 16892
rect 15867 16832 15931 16836
rect 15947 16892 16011 16896
rect 15947 16836 15951 16892
rect 15951 16836 16007 16892
rect 16007 16836 16011 16892
rect 15947 16832 16011 16836
rect 16027 16892 16091 16896
rect 16027 16836 16031 16892
rect 16031 16836 16087 16892
rect 16087 16836 16091 16892
rect 16027 16832 16091 16836
rect 21721 16892 21785 16896
rect 21721 16836 21725 16892
rect 21725 16836 21781 16892
rect 21781 16836 21785 16892
rect 21721 16832 21785 16836
rect 21801 16892 21865 16896
rect 21801 16836 21805 16892
rect 21805 16836 21861 16892
rect 21861 16836 21865 16892
rect 21801 16832 21865 16836
rect 21881 16892 21945 16896
rect 21881 16836 21885 16892
rect 21885 16836 21941 16892
rect 21941 16836 21945 16892
rect 21881 16832 21945 16836
rect 21961 16892 22025 16896
rect 21961 16836 21965 16892
rect 21965 16836 22021 16892
rect 22021 16836 22025 16892
rect 21961 16832 22025 16836
rect 4660 16628 4724 16692
rect 10732 16552 10796 16556
rect 10732 16496 10746 16552
rect 10746 16496 10796 16552
rect 10732 16492 10796 16496
rect 13860 16492 13924 16556
rect 6886 16348 6950 16352
rect 6886 16292 6890 16348
rect 6890 16292 6946 16348
rect 6946 16292 6950 16348
rect 6886 16288 6950 16292
rect 6966 16348 7030 16352
rect 6966 16292 6970 16348
rect 6970 16292 7026 16348
rect 7026 16292 7030 16348
rect 6966 16288 7030 16292
rect 7046 16348 7110 16352
rect 7046 16292 7050 16348
rect 7050 16292 7106 16348
rect 7106 16292 7110 16348
rect 7046 16288 7110 16292
rect 7126 16348 7190 16352
rect 7126 16292 7130 16348
rect 7130 16292 7186 16348
rect 7186 16292 7190 16348
rect 7126 16288 7190 16292
rect 12820 16348 12884 16352
rect 12820 16292 12824 16348
rect 12824 16292 12880 16348
rect 12880 16292 12884 16348
rect 12820 16288 12884 16292
rect 12900 16348 12964 16352
rect 12900 16292 12904 16348
rect 12904 16292 12960 16348
rect 12960 16292 12964 16348
rect 12900 16288 12964 16292
rect 12980 16348 13044 16352
rect 12980 16292 12984 16348
rect 12984 16292 13040 16348
rect 13040 16292 13044 16348
rect 12980 16288 13044 16292
rect 13060 16348 13124 16352
rect 13060 16292 13064 16348
rect 13064 16292 13120 16348
rect 13120 16292 13124 16348
rect 13060 16288 13124 16292
rect 18754 16348 18818 16352
rect 18754 16292 18758 16348
rect 18758 16292 18814 16348
rect 18814 16292 18818 16348
rect 18754 16288 18818 16292
rect 18834 16348 18898 16352
rect 18834 16292 18838 16348
rect 18838 16292 18894 16348
rect 18894 16292 18898 16348
rect 18834 16288 18898 16292
rect 18914 16348 18978 16352
rect 18914 16292 18918 16348
rect 18918 16292 18974 16348
rect 18974 16292 18978 16348
rect 18914 16288 18978 16292
rect 18994 16348 19058 16352
rect 18994 16292 18998 16348
rect 18998 16292 19054 16348
rect 19054 16292 19058 16348
rect 18994 16288 19058 16292
rect 24688 16348 24752 16352
rect 24688 16292 24692 16348
rect 24692 16292 24748 16348
rect 24748 16292 24752 16348
rect 24688 16288 24752 16292
rect 24768 16348 24832 16352
rect 24768 16292 24772 16348
rect 24772 16292 24828 16348
rect 24828 16292 24832 16348
rect 24768 16288 24832 16292
rect 24848 16348 24912 16352
rect 24848 16292 24852 16348
rect 24852 16292 24908 16348
rect 24908 16292 24912 16348
rect 24848 16288 24912 16292
rect 24928 16348 24992 16352
rect 24928 16292 24932 16348
rect 24932 16292 24988 16348
rect 24988 16292 24992 16348
rect 24928 16288 24992 16292
rect 3188 16084 3252 16148
rect 10916 15948 10980 16012
rect 22324 15948 22388 16012
rect 3919 15804 3983 15808
rect 3919 15748 3923 15804
rect 3923 15748 3979 15804
rect 3979 15748 3983 15804
rect 3919 15744 3983 15748
rect 3999 15804 4063 15808
rect 3999 15748 4003 15804
rect 4003 15748 4059 15804
rect 4059 15748 4063 15804
rect 3999 15744 4063 15748
rect 4079 15804 4143 15808
rect 4079 15748 4083 15804
rect 4083 15748 4139 15804
rect 4139 15748 4143 15804
rect 4079 15744 4143 15748
rect 4159 15804 4223 15808
rect 4159 15748 4163 15804
rect 4163 15748 4219 15804
rect 4219 15748 4223 15804
rect 4159 15744 4223 15748
rect 9853 15804 9917 15808
rect 9853 15748 9857 15804
rect 9857 15748 9913 15804
rect 9913 15748 9917 15804
rect 9853 15744 9917 15748
rect 9933 15804 9997 15808
rect 9933 15748 9937 15804
rect 9937 15748 9993 15804
rect 9993 15748 9997 15804
rect 9933 15744 9997 15748
rect 10013 15804 10077 15808
rect 10013 15748 10017 15804
rect 10017 15748 10073 15804
rect 10073 15748 10077 15804
rect 10013 15744 10077 15748
rect 10093 15804 10157 15808
rect 10093 15748 10097 15804
rect 10097 15748 10153 15804
rect 10153 15748 10157 15804
rect 10093 15744 10157 15748
rect 15787 15804 15851 15808
rect 15787 15748 15791 15804
rect 15791 15748 15847 15804
rect 15847 15748 15851 15804
rect 15787 15744 15851 15748
rect 15867 15804 15931 15808
rect 15867 15748 15871 15804
rect 15871 15748 15927 15804
rect 15927 15748 15931 15804
rect 15867 15744 15931 15748
rect 15947 15804 16011 15808
rect 15947 15748 15951 15804
rect 15951 15748 16007 15804
rect 16007 15748 16011 15804
rect 15947 15744 16011 15748
rect 16027 15804 16091 15808
rect 16027 15748 16031 15804
rect 16031 15748 16087 15804
rect 16087 15748 16091 15804
rect 16027 15744 16091 15748
rect 21721 15804 21785 15808
rect 21721 15748 21725 15804
rect 21725 15748 21781 15804
rect 21781 15748 21785 15804
rect 21721 15744 21785 15748
rect 21801 15804 21865 15808
rect 21801 15748 21805 15804
rect 21805 15748 21861 15804
rect 21861 15748 21865 15804
rect 21801 15744 21865 15748
rect 21881 15804 21945 15808
rect 21881 15748 21885 15804
rect 21885 15748 21941 15804
rect 21941 15748 21945 15804
rect 21881 15744 21945 15748
rect 21961 15804 22025 15808
rect 21961 15748 21965 15804
rect 21965 15748 22021 15804
rect 22021 15748 22025 15804
rect 21961 15744 22025 15748
rect 6886 15260 6950 15264
rect 6886 15204 6890 15260
rect 6890 15204 6946 15260
rect 6946 15204 6950 15260
rect 6886 15200 6950 15204
rect 6966 15260 7030 15264
rect 6966 15204 6970 15260
rect 6970 15204 7026 15260
rect 7026 15204 7030 15260
rect 6966 15200 7030 15204
rect 7046 15260 7110 15264
rect 7046 15204 7050 15260
rect 7050 15204 7106 15260
rect 7106 15204 7110 15260
rect 7046 15200 7110 15204
rect 7126 15260 7190 15264
rect 7126 15204 7130 15260
rect 7130 15204 7186 15260
rect 7186 15204 7190 15260
rect 7126 15200 7190 15204
rect 12820 15260 12884 15264
rect 12820 15204 12824 15260
rect 12824 15204 12880 15260
rect 12880 15204 12884 15260
rect 12820 15200 12884 15204
rect 12900 15260 12964 15264
rect 12900 15204 12904 15260
rect 12904 15204 12960 15260
rect 12960 15204 12964 15260
rect 12900 15200 12964 15204
rect 12980 15260 13044 15264
rect 12980 15204 12984 15260
rect 12984 15204 13040 15260
rect 13040 15204 13044 15260
rect 12980 15200 13044 15204
rect 13060 15260 13124 15264
rect 13060 15204 13064 15260
rect 13064 15204 13120 15260
rect 13120 15204 13124 15260
rect 13060 15200 13124 15204
rect 18754 15260 18818 15264
rect 18754 15204 18758 15260
rect 18758 15204 18814 15260
rect 18814 15204 18818 15260
rect 18754 15200 18818 15204
rect 18834 15260 18898 15264
rect 18834 15204 18838 15260
rect 18838 15204 18894 15260
rect 18894 15204 18898 15260
rect 18834 15200 18898 15204
rect 18914 15260 18978 15264
rect 18914 15204 18918 15260
rect 18918 15204 18974 15260
rect 18974 15204 18978 15260
rect 18914 15200 18978 15204
rect 18994 15260 19058 15264
rect 18994 15204 18998 15260
rect 18998 15204 19054 15260
rect 19054 15204 19058 15260
rect 18994 15200 19058 15204
rect 24688 15260 24752 15264
rect 24688 15204 24692 15260
rect 24692 15204 24748 15260
rect 24748 15204 24752 15260
rect 24688 15200 24752 15204
rect 24768 15260 24832 15264
rect 24768 15204 24772 15260
rect 24772 15204 24828 15260
rect 24828 15204 24832 15260
rect 24768 15200 24832 15204
rect 24848 15260 24912 15264
rect 24848 15204 24852 15260
rect 24852 15204 24908 15260
rect 24908 15204 24912 15260
rect 24848 15200 24912 15204
rect 24928 15260 24992 15264
rect 24928 15204 24932 15260
rect 24932 15204 24988 15260
rect 24988 15204 24992 15260
rect 24928 15200 24992 15204
rect 18276 15132 18340 15196
rect 17908 14860 17972 14924
rect 3919 14716 3983 14720
rect 3919 14660 3923 14716
rect 3923 14660 3979 14716
rect 3979 14660 3983 14716
rect 3919 14656 3983 14660
rect 3999 14716 4063 14720
rect 3999 14660 4003 14716
rect 4003 14660 4059 14716
rect 4059 14660 4063 14716
rect 3999 14656 4063 14660
rect 4079 14716 4143 14720
rect 4079 14660 4083 14716
rect 4083 14660 4139 14716
rect 4139 14660 4143 14716
rect 4079 14656 4143 14660
rect 4159 14716 4223 14720
rect 4159 14660 4163 14716
rect 4163 14660 4219 14716
rect 4219 14660 4223 14716
rect 4159 14656 4223 14660
rect 9853 14716 9917 14720
rect 9853 14660 9857 14716
rect 9857 14660 9913 14716
rect 9913 14660 9917 14716
rect 9853 14656 9917 14660
rect 9933 14716 9997 14720
rect 9933 14660 9937 14716
rect 9937 14660 9993 14716
rect 9993 14660 9997 14716
rect 9933 14656 9997 14660
rect 10013 14716 10077 14720
rect 10013 14660 10017 14716
rect 10017 14660 10073 14716
rect 10073 14660 10077 14716
rect 10013 14656 10077 14660
rect 10093 14716 10157 14720
rect 10093 14660 10097 14716
rect 10097 14660 10153 14716
rect 10153 14660 10157 14716
rect 10093 14656 10157 14660
rect 15787 14716 15851 14720
rect 15787 14660 15791 14716
rect 15791 14660 15847 14716
rect 15847 14660 15851 14716
rect 15787 14656 15851 14660
rect 15867 14716 15931 14720
rect 15867 14660 15871 14716
rect 15871 14660 15927 14716
rect 15927 14660 15931 14716
rect 15867 14656 15931 14660
rect 15947 14716 16011 14720
rect 15947 14660 15951 14716
rect 15951 14660 16007 14716
rect 16007 14660 16011 14716
rect 15947 14656 16011 14660
rect 16027 14716 16091 14720
rect 16027 14660 16031 14716
rect 16031 14660 16087 14716
rect 16087 14660 16091 14716
rect 16027 14656 16091 14660
rect 21721 14716 21785 14720
rect 21721 14660 21725 14716
rect 21725 14660 21781 14716
rect 21781 14660 21785 14716
rect 21721 14656 21785 14660
rect 21801 14716 21865 14720
rect 21801 14660 21805 14716
rect 21805 14660 21861 14716
rect 21861 14660 21865 14716
rect 21801 14656 21865 14660
rect 21881 14716 21945 14720
rect 21881 14660 21885 14716
rect 21885 14660 21941 14716
rect 21941 14660 21945 14716
rect 21881 14656 21945 14660
rect 21961 14716 22025 14720
rect 21961 14660 21965 14716
rect 21965 14660 22021 14716
rect 22021 14660 22025 14716
rect 21961 14656 22025 14660
rect 6886 14172 6950 14176
rect 6886 14116 6890 14172
rect 6890 14116 6946 14172
rect 6946 14116 6950 14172
rect 6886 14112 6950 14116
rect 6966 14172 7030 14176
rect 6966 14116 6970 14172
rect 6970 14116 7026 14172
rect 7026 14116 7030 14172
rect 6966 14112 7030 14116
rect 7046 14172 7110 14176
rect 7046 14116 7050 14172
rect 7050 14116 7106 14172
rect 7106 14116 7110 14172
rect 7046 14112 7110 14116
rect 7126 14172 7190 14176
rect 7126 14116 7130 14172
rect 7130 14116 7186 14172
rect 7186 14116 7190 14172
rect 7126 14112 7190 14116
rect 12820 14172 12884 14176
rect 12820 14116 12824 14172
rect 12824 14116 12880 14172
rect 12880 14116 12884 14172
rect 12820 14112 12884 14116
rect 12900 14172 12964 14176
rect 12900 14116 12904 14172
rect 12904 14116 12960 14172
rect 12960 14116 12964 14172
rect 12900 14112 12964 14116
rect 12980 14172 13044 14176
rect 12980 14116 12984 14172
rect 12984 14116 13040 14172
rect 13040 14116 13044 14172
rect 12980 14112 13044 14116
rect 13060 14172 13124 14176
rect 13060 14116 13064 14172
rect 13064 14116 13120 14172
rect 13120 14116 13124 14172
rect 13060 14112 13124 14116
rect 18754 14172 18818 14176
rect 18754 14116 18758 14172
rect 18758 14116 18814 14172
rect 18814 14116 18818 14172
rect 18754 14112 18818 14116
rect 18834 14172 18898 14176
rect 18834 14116 18838 14172
rect 18838 14116 18894 14172
rect 18894 14116 18898 14172
rect 18834 14112 18898 14116
rect 18914 14172 18978 14176
rect 18914 14116 18918 14172
rect 18918 14116 18974 14172
rect 18974 14116 18978 14172
rect 18914 14112 18978 14116
rect 18994 14172 19058 14176
rect 18994 14116 18998 14172
rect 18998 14116 19054 14172
rect 19054 14116 19058 14172
rect 18994 14112 19058 14116
rect 24688 14172 24752 14176
rect 24688 14116 24692 14172
rect 24692 14116 24748 14172
rect 24748 14116 24752 14172
rect 24688 14112 24752 14116
rect 24768 14172 24832 14176
rect 24768 14116 24772 14172
rect 24772 14116 24828 14172
rect 24828 14116 24832 14172
rect 24768 14112 24832 14116
rect 24848 14172 24912 14176
rect 24848 14116 24852 14172
rect 24852 14116 24908 14172
rect 24908 14116 24912 14172
rect 24848 14112 24912 14116
rect 24928 14172 24992 14176
rect 24928 14116 24932 14172
rect 24932 14116 24988 14172
rect 24988 14116 24992 14172
rect 24928 14112 24992 14116
rect 14596 13968 14660 13972
rect 14596 13912 14646 13968
rect 14646 13912 14660 13968
rect 14596 13908 14660 13912
rect 1348 13832 1412 13836
rect 1348 13776 1362 13832
rect 1362 13776 1412 13832
rect 1348 13772 1412 13776
rect 3004 13832 3068 13836
rect 3004 13776 3054 13832
rect 3054 13776 3068 13832
rect 3004 13772 3068 13776
rect 6500 13636 6564 13700
rect 3919 13628 3983 13632
rect 3919 13572 3923 13628
rect 3923 13572 3979 13628
rect 3979 13572 3983 13628
rect 3919 13568 3983 13572
rect 3999 13628 4063 13632
rect 3999 13572 4003 13628
rect 4003 13572 4059 13628
rect 4059 13572 4063 13628
rect 3999 13568 4063 13572
rect 4079 13628 4143 13632
rect 4079 13572 4083 13628
rect 4083 13572 4139 13628
rect 4139 13572 4143 13628
rect 4079 13568 4143 13572
rect 4159 13628 4223 13632
rect 4159 13572 4163 13628
rect 4163 13572 4219 13628
rect 4219 13572 4223 13628
rect 4159 13568 4223 13572
rect 12204 13636 12268 13700
rect 13860 13636 13924 13700
rect 9853 13628 9917 13632
rect 9853 13572 9857 13628
rect 9857 13572 9913 13628
rect 9913 13572 9917 13628
rect 9853 13568 9917 13572
rect 9933 13628 9997 13632
rect 9933 13572 9937 13628
rect 9937 13572 9993 13628
rect 9993 13572 9997 13628
rect 9933 13568 9997 13572
rect 10013 13628 10077 13632
rect 10013 13572 10017 13628
rect 10017 13572 10073 13628
rect 10073 13572 10077 13628
rect 10013 13568 10077 13572
rect 10093 13628 10157 13632
rect 10093 13572 10097 13628
rect 10097 13572 10153 13628
rect 10153 13572 10157 13628
rect 10093 13568 10157 13572
rect 15787 13628 15851 13632
rect 15787 13572 15791 13628
rect 15791 13572 15847 13628
rect 15847 13572 15851 13628
rect 15787 13568 15851 13572
rect 15867 13628 15931 13632
rect 15867 13572 15871 13628
rect 15871 13572 15927 13628
rect 15927 13572 15931 13628
rect 15867 13568 15931 13572
rect 15947 13628 16011 13632
rect 15947 13572 15951 13628
rect 15951 13572 16007 13628
rect 16007 13572 16011 13628
rect 15947 13568 16011 13572
rect 16027 13628 16091 13632
rect 16027 13572 16031 13628
rect 16031 13572 16087 13628
rect 16087 13572 16091 13628
rect 16027 13568 16091 13572
rect 21721 13628 21785 13632
rect 21721 13572 21725 13628
rect 21725 13572 21781 13628
rect 21781 13572 21785 13628
rect 21721 13568 21785 13572
rect 21801 13628 21865 13632
rect 21801 13572 21805 13628
rect 21805 13572 21861 13628
rect 21861 13572 21865 13628
rect 21801 13568 21865 13572
rect 21881 13628 21945 13632
rect 21881 13572 21885 13628
rect 21885 13572 21941 13628
rect 21941 13572 21945 13628
rect 21881 13568 21945 13572
rect 21961 13628 22025 13632
rect 21961 13572 21965 13628
rect 21965 13572 22021 13628
rect 22021 13572 22025 13628
rect 21961 13568 22025 13572
rect 1716 13364 1780 13428
rect 2084 13364 2148 13428
rect 2084 13228 2148 13292
rect 5028 13364 5092 13428
rect 6886 13084 6950 13088
rect 6886 13028 6890 13084
rect 6890 13028 6946 13084
rect 6946 13028 6950 13084
rect 6886 13024 6950 13028
rect 6966 13084 7030 13088
rect 6966 13028 6970 13084
rect 6970 13028 7026 13084
rect 7026 13028 7030 13084
rect 6966 13024 7030 13028
rect 7046 13084 7110 13088
rect 7046 13028 7050 13084
rect 7050 13028 7106 13084
rect 7106 13028 7110 13084
rect 7046 13024 7110 13028
rect 7126 13084 7190 13088
rect 7126 13028 7130 13084
rect 7130 13028 7186 13084
rect 7186 13028 7190 13084
rect 7126 13024 7190 13028
rect 12820 13084 12884 13088
rect 12820 13028 12824 13084
rect 12824 13028 12880 13084
rect 12880 13028 12884 13084
rect 12820 13024 12884 13028
rect 12900 13084 12964 13088
rect 12900 13028 12904 13084
rect 12904 13028 12960 13084
rect 12960 13028 12964 13084
rect 12900 13024 12964 13028
rect 12980 13084 13044 13088
rect 12980 13028 12984 13084
rect 12984 13028 13040 13084
rect 13040 13028 13044 13084
rect 12980 13024 13044 13028
rect 13060 13084 13124 13088
rect 13060 13028 13064 13084
rect 13064 13028 13120 13084
rect 13120 13028 13124 13084
rect 13060 13024 13124 13028
rect 18754 13084 18818 13088
rect 18754 13028 18758 13084
rect 18758 13028 18814 13084
rect 18814 13028 18818 13084
rect 18754 13024 18818 13028
rect 18834 13084 18898 13088
rect 18834 13028 18838 13084
rect 18838 13028 18894 13084
rect 18894 13028 18898 13084
rect 18834 13024 18898 13028
rect 18914 13084 18978 13088
rect 18914 13028 18918 13084
rect 18918 13028 18974 13084
rect 18974 13028 18978 13084
rect 18914 13024 18978 13028
rect 18994 13084 19058 13088
rect 18994 13028 18998 13084
rect 18998 13028 19054 13084
rect 19054 13028 19058 13084
rect 18994 13024 19058 13028
rect 24688 13084 24752 13088
rect 24688 13028 24692 13084
rect 24692 13028 24748 13084
rect 24748 13028 24752 13084
rect 24688 13024 24752 13028
rect 24768 13084 24832 13088
rect 24768 13028 24772 13084
rect 24772 13028 24828 13084
rect 24828 13028 24832 13084
rect 24768 13024 24832 13028
rect 24848 13084 24912 13088
rect 24848 13028 24852 13084
rect 24852 13028 24908 13084
rect 24908 13028 24912 13084
rect 24848 13024 24912 13028
rect 24928 13084 24992 13088
rect 24928 13028 24932 13084
rect 24932 13028 24988 13084
rect 24988 13028 24992 13084
rect 24928 13024 24992 13028
rect 10548 12820 10612 12884
rect 2452 12684 2516 12748
rect 3919 12540 3983 12544
rect 3919 12484 3923 12540
rect 3923 12484 3979 12540
rect 3979 12484 3983 12540
rect 3919 12480 3983 12484
rect 3999 12540 4063 12544
rect 3999 12484 4003 12540
rect 4003 12484 4059 12540
rect 4059 12484 4063 12540
rect 3999 12480 4063 12484
rect 4079 12540 4143 12544
rect 4079 12484 4083 12540
rect 4083 12484 4139 12540
rect 4139 12484 4143 12540
rect 4079 12480 4143 12484
rect 4159 12540 4223 12544
rect 4159 12484 4163 12540
rect 4163 12484 4219 12540
rect 4219 12484 4223 12540
rect 4159 12480 4223 12484
rect 9853 12540 9917 12544
rect 9853 12484 9857 12540
rect 9857 12484 9913 12540
rect 9913 12484 9917 12540
rect 9853 12480 9917 12484
rect 9933 12540 9997 12544
rect 9933 12484 9937 12540
rect 9937 12484 9993 12540
rect 9993 12484 9997 12540
rect 9933 12480 9997 12484
rect 10013 12540 10077 12544
rect 10013 12484 10017 12540
rect 10017 12484 10073 12540
rect 10073 12484 10077 12540
rect 10013 12480 10077 12484
rect 10093 12540 10157 12544
rect 10093 12484 10097 12540
rect 10097 12484 10153 12540
rect 10153 12484 10157 12540
rect 10093 12480 10157 12484
rect 15787 12540 15851 12544
rect 15787 12484 15791 12540
rect 15791 12484 15847 12540
rect 15847 12484 15851 12540
rect 15787 12480 15851 12484
rect 15867 12540 15931 12544
rect 15867 12484 15871 12540
rect 15871 12484 15927 12540
rect 15927 12484 15931 12540
rect 15867 12480 15931 12484
rect 15947 12540 16011 12544
rect 15947 12484 15951 12540
rect 15951 12484 16007 12540
rect 16007 12484 16011 12540
rect 15947 12480 16011 12484
rect 16027 12540 16091 12544
rect 16027 12484 16031 12540
rect 16031 12484 16087 12540
rect 16087 12484 16091 12540
rect 16027 12480 16091 12484
rect 21721 12540 21785 12544
rect 21721 12484 21725 12540
rect 21725 12484 21781 12540
rect 21781 12484 21785 12540
rect 21721 12480 21785 12484
rect 21801 12540 21865 12544
rect 21801 12484 21805 12540
rect 21805 12484 21861 12540
rect 21861 12484 21865 12540
rect 21801 12480 21865 12484
rect 21881 12540 21945 12544
rect 21881 12484 21885 12540
rect 21885 12484 21941 12540
rect 21941 12484 21945 12540
rect 21881 12480 21945 12484
rect 21961 12540 22025 12544
rect 21961 12484 21965 12540
rect 21965 12484 22021 12540
rect 22021 12484 22025 12540
rect 21961 12480 22025 12484
rect 22508 12276 22572 12340
rect 6886 11996 6950 12000
rect 6886 11940 6890 11996
rect 6890 11940 6946 11996
rect 6946 11940 6950 11996
rect 6886 11936 6950 11940
rect 6966 11996 7030 12000
rect 6966 11940 6970 11996
rect 6970 11940 7026 11996
rect 7026 11940 7030 11996
rect 6966 11936 7030 11940
rect 7046 11996 7110 12000
rect 7046 11940 7050 11996
rect 7050 11940 7106 11996
rect 7106 11940 7110 11996
rect 7046 11936 7110 11940
rect 7126 11996 7190 12000
rect 7126 11940 7130 11996
rect 7130 11940 7186 11996
rect 7186 11940 7190 11996
rect 7126 11936 7190 11940
rect 12820 11996 12884 12000
rect 12820 11940 12824 11996
rect 12824 11940 12880 11996
rect 12880 11940 12884 11996
rect 12820 11936 12884 11940
rect 12900 11996 12964 12000
rect 12900 11940 12904 11996
rect 12904 11940 12960 11996
rect 12960 11940 12964 11996
rect 12900 11936 12964 11940
rect 12980 11996 13044 12000
rect 12980 11940 12984 11996
rect 12984 11940 13040 11996
rect 13040 11940 13044 11996
rect 12980 11936 13044 11940
rect 13060 11996 13124 12000
rect 13060 11940 13064 11996
rect 13064 11940 13120 11996
rect 13120 11940 13124 11996
rect 13060 11936 13124 11940
rect 18754 11996 18818 12000
rect 18754 11940 18758 11996
rect 18758 11940 18814 11996
rect 18814 11940 18818 11996
rect 18754 11936 18818 11940
rect 18834 11996 18898 12000
rect 18834 11940 18838 11996
rect 18838 11940 18894 11996
rect 18894 11940 18898 11996
rect 18834 11936 18898 11940
rect 18914 11996 18978 12000
rect 18914 11940 18918 11996
rect 18918 11940 18974 11996
rect 18974 11940 18978 11996
rect 18914 11936 18978 11940
rect 18994 11996 19058 12000
rect 18994 11940 18998 11996
rect 18998 11940 19054 11996
rect 19054 11940 19058 11996
rect 18994 11936 19058 11940
rect 24688 11996 24752 12000
rect 24688 11940 24692 11996
rect 24692 11940 24748 11996
rect 24748 11940 24752 11996
rect 24688 11936 24752 11940
rect 24768 11996 24832 12000
rect 24768 11940 24772 11996
rect 24772 11940 24828 11996
rect 24828 11940 24832 11996
rect 24768 11936 24832 11940
rect 24848 11996 24912 12000
rect 24848 11940 24852 11996
rect 24852 11940 24908 11996
rect 24908 11940 24912 11996
rect 24848 11936 24912 11940
rect 24928 11996 24992 12000
rect 24928 11940 24932 11996
rect 24932 11940 24988 11996
rect 24988 11940 24992 11996
rect 24928 11936 24992 11940
rect 3919 11452 3983 11456
rect 3919 11396 3923 11452
rect 3923 11396 3979 11452
rect 3979 11396 3983 11452
rect 3919 11392 3983 11396
rect 3999 11452 4063 11456
rect 3999 11396 4003 11452
rect 4003 11396 4059 11452
rect 4059 11396 4063 11452
rect 3999 11392 4063 11396
rect 4079 11452 4143 11456
rect 4079 11396 4083 11452
rect 4083 11396 4139 11452
rect 4139 11396 4143 11452
rect 4079 11392 4143 11396
rect 4159 11452 4223 11456
rect 4159 11396 4163 11452
rect 4163 11396 4219 11452
rect 4219 11396 4223 11452
rect 4159 11392 4223 11396
rect 9853 11452 9917 11456
rect 9853 11396 9857 11452
rect 9857 11396 9913 11452
rect 9913 11396 9917 11452
rect 9853 11392 9917 11396
rect 9933 11452 9997 11456
rect 9933 11396 9937 11452
rect 9937 11396 9993 11452
rect 9993 11396 9997 11452
rect 9933 11392 9997 11396
rect 10013 11452 10077 11456
rect 10013 11396 10017 11452
rect 10017 11396 10073 11452
rect 10073 11396 10077 11452
rect 10013 11392 10077 11396
rect 10093 11452 10157 11456
rect 10093 11396 10097 11452
rect 10097 11396 10153 11452
rect 10153 11396 10157 11452
rect 10093 11392 10157 11396
rect 15787 11452 15851 11456
rect 15787 11396 15791 11452
rect 15791 11396 15847 11452
rect 15847 11396 15851 11452
rect 15787 11392 15851 11396
rect 15867 11452 15931 11456
rect 15867 11396 15871 11452
rect 15871 11396 15927 11452
rect 15927 11396 15931 11452
rect 15867 11392 15931 11396
rect 15947 11452 16011 11456
rect 15947 11396 15951 11452
rect 15951 11396 16007 11452
rect 16007 11396 16011 11452
rect 15947 11392 16011 11396
rect 16027 11452 16091 11456
rect 16027 11396 16031 11452
rect 16031 11396 16087 11452
rect 16087 11396 16091 11452
rect 16027 11392 16091 11396
rect 21721 11452 21785 11456
rect 21721 11396 21725 11452
rect 21725 11396 21781 11452
rect 21781 11396 21785 11452
rect 21721 11392 21785 11396
rect 21801 11452 21865 11456
rect 21801 11396 21805 11452
rect 21805 11396 21861 11452
rect 21861 11396 21865 11452
rect 21801 11392 21865 11396
rect 21881 11452 21945 11456
rect 21881 11396 21885 11452
rect 21885 11396 21941 11452
rect 21941 11396 21945 11452
rect 21881 11392 21945 11396
rect 21961 11452 22025 11456
rect 21961 11396 21965 11452
rect 21965 11396 22021 11452
rect 22021 11396 22025 11452
rect 21961 11392 22025 11396
rect 16620 11188 16684 11252
rect 21036 10916 21100 10980
rect 6886 10908 6950 10912
rect 6886 10852 6890 10908
rect 6890 10852 6946 10908
rect 6946 10852 6950 10908
rect 6886 10848 6950 10852
rect 6966 10908 7030 10912
rect 6966 10852 6970 10908
rect 6970 10852 7026 10908
rect 7026 10852 7030 10908
rect 6966 10848 7030 10852
rect 7046 10908 7110 10912
rect 7046 10852 7050 10908
rect 7050 10852 7106 10908
rect 7106 10852 7110 10908
rect 7046 10848 7110 10852
rect 7126 10908 7190 10912
rect 7126 10852 7130 10908
rect 7130 10852 7186 10908
rect 7186 10852 7190 10908
rect 7126 10848 7190 10852
rect 12820 10908 12884 10912
rect 12820 10852 12824 10908
rect 12824 10852 12880 10908
rect 12880 10852 12884 10908
rect 12820 10848 12884 10852
rect 12900 10908 12964 10912
rect 12900 10852 12904 10908
rect 12904 10852 12960 10908
rect 12960 10852 12964 10908
rect 12900 10848 12964 10852
rect 12980 10908 13044 10912
rect 12980 10852 12984 10908
rect 12984 10852 13040 10908
rect 13040 10852 13044 10908
rect 12980 10848 13044 10852
rect 13060 10908 13124 10912
rect 13060 10852 13064 10908
rect 13064 10852 13120 10908
rect 13120 10852 13124 10908
rect 13060 10848 13124 10852
rect 18754 10908 18818 10912
rect 18754 10852 18758 10908
rect 18758 10852 18814 10908
rect 18814 10852 18818 10908
rect 18754 10848 18818 10852
rect 18834 10908 18898 10912
rect 18834 10852 18838 10908
rect 18838 10852 18894 10908
rect 18894 10852 18898 10908
rect 18834 10848 18898 10852
rect 18914 10908 18978 10912
rect 18914 10852 18918 10908
rect 18918 10852 18974 10908
rect 18974 10852 18978 10908
rect 18914 10848 18978 10852
rect 18994 10908 19058 10912
rect 18994 10852 18998 10908
rect 18998 10852 19054 10908
rect 19054 10852 19058 10908
rect 18994 10848 19058 10852
rect 24688 10908 24752 10912
rect 24688 10852 24692 10908
rect 24692 10852 24748 10908
rect 24748 10852 24752 10908
rect 24688 10848 24752 10852
rect 24768 10908 24832 10912
rect 24768 10852 24772 10908
rect 24772 10852 24828 10908
rect 24828 10852 24832 10908
rect 24768 10848 24832 10852
rect 24848 10908 24912 10912
rect 24848 10852 24852 10908
rect 24852 10852 24908 10908
rect 24908 10852 24912 10908
rect 24848 10848 24912 10852
rect 24928 10908 24992 10912
rect 24928 10852 24932 10908
rect 24932 10852 24988 10908
rect 24988 10852 24992 10908
rect 24928 10848 24992 10852
rect 14964 10372 15028 10436
rect 3919 10364 3983 10368
rect 3919 10308 3923 10364
rect 3923 10308 3979 10364
rect 3979 10308 3983 10364
rect 3919 10304 3983 10308
rect 3999 10364 4063 10368
rect 3999 10308 4003 10364
rect 4003 10308 4059 10364
rect 4059 10308 4063 10364
rect 3999 10304 4063 10308
rect 4079 10364 4143 10368
rect 4079 10308 4083 10364
rect 4083 10308 4139 10364
rect 4139 10308 4143 10364
rect 4079 10304 4143 10308
rect 4159 10364 4223 10368
rect 4159 10308 4163 10364
rect 4163 10308 4219 10364
rect 4219 10308 4223 10364
rect 4159 10304 4223 10308
rect 9853 10364 9917 10368
rect 9853 10308 9857 10364
rect 9857 10308 9913 10364
rect 9913 10308 9917 10364
rect 9853 10304 9917 10308
rect 9933 10364 9997 10368
rect 9933 10308 9937 10364
rect 9937 10308 9993 10364
rect 9993 10308 9997 10364
rect 9933 10304 9997 10308
rect 10013 10364 10077 10368
rect 10013 10308 10017 10364
rect 10017 10308 10073 10364
rect 10073 10308 10077 10364
rect 10013 10304 10077 10308
rect 10093 10364 10157 10368
rect 10093 10308 10097 10364
rect 10097 10308 10153 10364
rect 10153 10308 10157 10364
rect 10093 10304 10157 10308
rect 15787 10364 15851 10368
rect 15787 10308 15791 10364
rect 15791 10308 15847 10364
rect 15847 10308 15851 10364
rect 15787 10304 15851 10308
rect 15867 10364 15931 10368
rect 15867 10308 15871 10364
rect 15871 10308 15927 10364
rect 15927 10308 15931 10364
rect 15867 10304 15931 10308
rect 15947 10364 16011 10368
rect 15947 10308 15951 10364
rect 15951 10308 16007 10364
rect 16007 10308 16011 10364
rect 15947 10304 16011 10308
rect 16027 10364 16091 10368
rect 16027 10308 16031 10364
rect 16031 10308 16087 10364
rect 16087 10308 16091 10364
rect 16027 10304 16091 10308
rect 21721 10364 21785 10368
rect 21721 10308 21725 10364
rect 21725 10308 21781 10364
rect 21781 10308 21785 10364
rect 21721 10304 21785 10308
rect 21801 10364 21865 10368
rect 21801 10308 21805 10364
rect 21805 10308 21861 10364
rect 21861 10308 21865 10364
rect 21801 10304 21865 10308
rect 21881 10364 21945 10368
rect 21881 10308 21885 10364
rect 21885 10308 21941 10364
rect 21941 10308 21945 10364
rect 21881 10304 21945 10308
rect 21961 10364 22025 10368
rect 21961 10308 21965 10364
rect 21965 10308 22021 10364
rect 22021 10308 22025 10364
rect 21961 10304 22025 10308
rect 4844 10160 4908 10164
rect 4844 10104 4858 10160
rect 4858 10104 4908 10160
rect 4844 10100 4908 10104
rect 6886 9820 6950 9824
rect 6886 9764 6890 9820
rect 6890 9764 6946 9820
rect 6946 9764 6950 9820
rect 6886 9760 6950 9764
rect 6966 9820 7030 9824
rect 6966 9764 6970 9820
rect 6970 9764 7026 9820
rect 7026 9764 7030 9820
rect 6966 9760 7030 9764
rect 7046 9820 7110 9824
rect 7046 9764 7050 9820
rect 7050 9764 7106 9820
rect 7106 9764 7110 9820
rect 7046 9760 7110 9764
rect 7126 9820 7190 9824
rect 7126 9764 7130 9820
rect 7130 9764 7186 9820
rect 7186 9764 7190 9820
rect 7126 9760 7190 9764
rect 12820 9820 12884 9824
rect 12820 9764 12824 9820
rect 12824 9764 12880 9820
rect 12880 9764 12884 9820
rect 12820 9760 12884 9764
rect 12900 9820 12964 9824
rect 12900 9764 12904 9820
rect 12904 9764 12960 9820
rect 12960 9764 12964 9820
rect 12900 9760 12964 9764
rect 12980 9820 13044 9824
rect 12980 9764 12984 9820
rect 12984 9764 13040 9820
rect 13040 9764 13044 9820
rect 12980 9760 13044 9764
rect 13060 9820 13124 9824
rect 13060 9764 13064 9820
rect 13064 9764 13120 9820
rect 13120 9764 13124 9820
rect 13060 9760 13124 9764
rect 18754 9820 18818 9824
rect 18754 9764 18758 9820
rect 18758 9764 18814 9820
rect 18814 9764 18818 9820
rect 18754 9760 18818 9764
rect 18834 9820 18898 9824
rect 18834 9764 18838 9820
rect 18838 9764 18894 9820
rect 18894 9764 18898 9820
rect 18834 9760 18898 9764
rect 18914 9820 18978 9824
rect 18914 9764 18918 9820
rect 18918 9764 18974 9820
rect 18974 9764 18978 9820
rect 18914 9760 18978 9764
rect 18994 9820 19058 9824
rect 18994 9764 18998 9820
rect 18998 9764 19054 9820
rect 19054 9764 19058 9820
rect 18994 9760 19058 9764
rect 24688 9820 24752 9824
rect 24688 9764 24692 9820
rect 24692 9764 24748 9820
rect 24748 9764 24752 9820
rect 24688 9760 24752 9764
rect 24768 9820 24832 9824
rect 24768 9764 24772 9820
rect 24772 9764 24828 9820
rect 24828 9764 24832 9820
rect 24768 9760 24832 9764
rect 24848 9820 24912 9824
rect 24848 9764 24852 9820
rect 24852 9764 24908 9820
rect 24908 9764 24912 9820
rect 24848 9760 24912 9764
rect 24928 9820 24992 9824
rect 24928 9764 24932 9820
rect 24932 9764 24988 9820
rect 24988 9764 24992 9820
rect 24928 9760 24992 9764
rect 17356 9692 17420 9756
rect 21588 9480 21652 9484
rect 21588 9424 21638 9480
rect 21638 9424 21652 9480
rect 21588 9420 21652 9424
rect 3919 9276 3983 9280
rect 3919 9220 3923 9276
rect 3923 9220 3979 9276
rect 3979 9220 3983 9276
rect 3919 9216 3983 9220
rect 3999 9276 4063 9280
rect 3999 9220 4003 9276
rect 4003 9220 4059 9276
rect 4059 9220 4063 9276
rect 3999 9216 4063 9220
rect 4079 9276 4143 9280
rect 4079 9220 4083 9276
rect 4083 9220 4139 9276
rect 4139 9220 4143 9276
rect 4079 9216 4143 9220
rect 4159 9276 4223 9280
rect 4159 9220 4163 9276
rect 4163 9220 4219 9276
rect 4219 9220 4223 9276
rect 4159 9216 4223 9220
rect 9853 9276 9917 9280
rect 9853 9220 9857 9276
rect 9857 9220 9913 9276
rect 9913 9220 9917 9276
rect 9853 9216 9917 9220
rect 9933 9276 9997 9280
rect 9933 9220 9937 9276
rect 9937 9220 9993 9276
rect 9993 9220 9997 9276
rect 9933 9216 9997 9220
rect 10013 9276 10077 9280
rect 10013 9220 10017 9276
rect 10017 9220 10073 9276
rect 10073 9220 10077 9276
rect 10013 9216 10077 9220
rect 10093 9276 10157 9280
rect 10093 9220 10097 9276
rect 10097 9220 10153 9276
rect 10153 9220 10157 9276
rect 10093 9216 10157 9220
rect 15787 9276 15851 9280
rect 15787 9220 15791 9276
rect 15791 9220 15847 9276
rect 15847 9220 15851 9276
rect 15787 9216 15851 9220
rect 15867 9276 15931 9280
rect 15867 9220 15871 9276
rect 15871 9220 15927 9276
rect 15927 9220 15931 9276
rect 15867 9216 15931 9220
rect 15947 9276 16011 9280
rect 15947 9220 15951 9276
rect 15951 9220 16007 9276
rect 16007 9220 16011 9276
rect 15947 9216 16011 9220
rect 16027 9276 16091 9280
rect 16027 9220 16031 9276
rect 16031 9220 16087 9276
rect 16087 9220 16091 9276
rect 16027 9216 16091 9220
rect 21721 9276 21785 9280
rect 21721 9220 21725 9276
rect 21725 9220 21781 9276
rect 21781 9220 21785 9276
rect 21721 9216 21785 9220
rect 21801 9276 21865 9280
rect 21801 9220 21805 9276
rect 21805 9220 21861 9276
rect 21861 9220 21865 9276
rect 21801 9216 21865 9220
rect 21881 9276 21945 9280
rect 21881 9220 21885 9276
rect 21885 9220 21941 9276
rect 21941 9220 21945 9276
rect 21881 9216 21945 9220
rect 21961 9276 22025 9280
rect 21961 9220 21965 9276
rect 21965 9220 22021 9276
rect 22021 9220 22025 9276
rect 21961 9216 22025 9220
rect 6886 8732 6950 8736
rect 6886 8676 6890 8732
rect 6890 8676 6946 8732
rect 6946 8676 6950 8732
rect 6886 8672 6950 8676
rect 6966 8732 7030 8736
rect 6966 8676 6970 8732
rect 6970 8676 7026 8732
rect 7026 8676 7030 8732
rect 6966 8672 7030 8676
rect 7046 8732 7110 8736
rect 7046 8676 7050 8732
rect 7050 8676 7106 8732
rect 7106 8676 7110 8732
rect 7046 8672 7110 8676
rect 7126 8732 7190 8736
rect 7126 8676 7130 8732
rect 7130 8676 7186 8732
rect 7186 8676 7190 8732
rect 7126 8672 7190 8676
rect 12820 8732 12884 8736
rect 12820 8676 12824 8732
rect 12824 8676 12880 8732
rect 12880 8676 12884 8732
rect 12820 8672 12884 8676
rect 12900 8732 12964 8736
rect 12900 8676 12904 8732
rect 12904 8676 12960 8732
rect 12960 8676 12964 8732
rect 12900 8672 12964 8676
rect 12980 8732 13044 8736
rect 12980 8676 12984 8732
rect 12984 8676 13040 8732
rect 13040 8676 13044 8732
rect 12980 8672 13044 8676
rect 13060 8732 13124 8736
rect 13060 8676 13064 8732
rect 13064 8676 13120 8732
rect 13120 8676 13124 8732
rect 13060 8672 13124 8676
rect 18754 8732 18818 8736
rect 18754 8676 18758 8732
rect 18758 8676 18814 8732
rect 18814 8676 18818 8732
rect 18754 8672 18818 8676
rect 18834 8732 18898 8736
rect 18834 8676 18838 8732
rect 18838 8676 18894 8732
rect 18894 8676 18898 8732
rect 18834 8672 18898 8676
rect 18914 8732 18978 8736
rect 18914 8676 18918 8732
rect 18918 8676 18974 8732
rect 18974 8676 18978 8732
rect 18914 8672 18978 8676
rect 18994 8732 19058 8736
rect 18994 8676 18998 8732
rect 18998 8676 19054 8732
rect 19054 8676 19058 8732
rect 18994 8672 19058 8676
rect 24688 8732 24752 8736
rect 24688 8676 24692 8732
rect 24692 8676 24748 8732
rect 24748 8676 24752 8732
rect 24688 8672 24752 8676
rect 24768 8732 24832 8736
rect 24768 8676 24772 8732
rect 24772 8676 24828 8732
rect 24828 8676 24832 8732
rect 24768 8672 24832 8676
rect 24848 8732 24912 8736
rect 24848 8676 24852 8732
rect 24852 8676 24908 8732
rect 24908 8676 24912 8732
rect 24848 8672 24912 8676
rect 24928 8732 24992 8736
rect 24928 8676 24932 8732
rect 24932 8676 24988 8732
rect 24988 8676 24992 8732
rect 24928 8672 24992 8676
rect 612 8604 676 8668
rect 4292 8604 4356 8668
rect 17356 8604 17420 8668
rect 5396 8332 5460 8396
rect 3919 8188 3983 8192
rect 3919 8132 3923 8188
rect 3923 8132 3979 8188
rect 3979 8132 3983 8188
rect 3919 8128 3983 8132
rect 3999 8188 4063 8192
rect 3999 8132 4003 8188
rect 4003 8132 4059 8188
rect 4059 8132 4063 8188
rect 3999 8128 4063 8132
rect 4079 8188 4143 8192
rect 4079 8132 4083 8188
rect 4083 8132 4139 8188
rect 4139 8132 4143 8188
rect 4079 8128 4143 8132
rect 4159 8188 4223 8192
rect 4159 8132 4163 8188
rect 4163 8132 4219 8188
rect 4219 8132 4223 8188
rect 4159 8128 4223 8132
rect 9853 8188 9917 8192
rect 9853 8132 9857 8188
rect 9857 8132 9913 8188
rect 9913 8132 9917 8188
rect 9853 8128 9917 8132
rect 9933 8188 9997 8192
rect 9933 8132 9937 8188
rect 9937 8132 9993 8188
rect 9993 8132 9997 8188
rect 9933 8128 9997 8132
rect 10013 8188 10077 8192
rect 10013 8132 10017 8188
rect 10017 8132 10073 8188
rect 10073 8132 10077 8188
rect 10013 8128 10077 8132
rect 10093 8188 10157 8192
rect 10093 8132 10097 8188
rect 10097 8132 10153 8188
rect 10153 8132 10157 8188
rect 10093 8128 10157 8132
rect 15787 8188 15851 8192
rect 15787 8132 15791 8188
rect 15791 8132 15847 8188
rect 15847 8132 15851 8188
rect 15787 8128 15851 8132
rect 15867 8188 15931 8192
rect 15867 8132 15871 8188
rect 15871 8132 15927 8188
rect 15927 8132 15931 8188
rect 15867 8128 15931 8132
rect 15947 8188 16011 8192
rect 15947 8132 15951 8188
rect 15951 8132 16007 8188
rect 16007 8132 16011 8188
rect 15947 8128 16011 8132
rect 16027 8188 16091 8192
rect 16027 8132 16031 8188
rect 16031 8132 16087 8188
rect 16087 8132 16091 8188
rect 16027 8128 16091 8132
rect 21721 8188 21785 8192
rect 21721 8132 21725 8188
rect 21725 8132 21781 8188
rect 21781 8132 21785 8188
rect 21721 8128 21785 8132
rect 21801 8188 21865 8192
rect 21801 8132 21805 8188
rect 21805 8132 21861 8188
rect 21861 8132 21865 8188
rect 21801 8128 21865 8132
rect 21881 8188 21945 8192
rect 21881 8132 21885 8188
rect 21885 8132 21941 8188
rect 21941 8132 21945 8188
rect 21881 8128 21945 8132
rect 21961 8188 22025 8192
rect 21961 8132 21965 8188
rect 21965 8132 22021 8188
rect 22021 8132 22025 8188
rect 21961 8128 22025 8132
rect 19564 7924 19628 7988
rect 6886 7644 6950 7648
rect 6886 7588 6890 7644
rect 6890 7588 6946 7644
rect 6946 7588 6950 7644
rect 6886 7584 6950 7588
rect 6966 7644 7030 7648
rect 6966 7588 6970 7644
rect 6970 7588 7026 7644
rect 7026 7588 7030 7644
rect 6966 7584 7030 7588
rect 7046 7644 7110 7648
rect 7046 7588 7050 7644
rect 7050 7588 7106 7644
rect 7106 7588 7110 7644
rect 7046 7584 7110 7588
rect 7126 7644 7190 7648
rect 7126 7588 7130 7644
rect 7130 7588 7186 7644
rect 7186 7588 7190 7644
rect 7126 7584 7190 7588
rect 12820 7644 12884 7648
rect 12820 7588 12824 7644
rect 12824 7588 12880 7644
rect 12880 7588 12884 7644
rect 12820 7584 12884 7588
rect 12900 7644 12964 7648
rect 12900 7588 12904 7644
rect 12904 7588 12960 7644
rect 12960 7588 12964 7644
rect 12900 7584 12964 7588
rect 12980 7644 13044 7648
rect 12980 7588 12984 7644
rect 12984 7588 13040 7644
rect 13040 7588 13044 7644
rect 12980 7584 13044 7588
rect 13060 7644 13124 7648
rect 13060 7588 13064 7644
rect 13064 7588 13120 7644
rect 13120 7588 13124 7644
rect 13060 7584 13124 7588
rect 18754 7644 18818 7648
rect 18754 7588 18758 7644
rect 18758 7588 18814 7644
rect 18814 7588 18818 7644
rect 18754 7584 18818 7588
rect 18834 7644 18898 7648
rect 18834 7588 18838 7644
rect 18838 7588 18894 7644
rect 18894 7588 18898 7644
rect 18834 7584 18898 7588
rect 18914 7644 18978 7648
rect 18914 7588 18918 7644
rect 18918 7588 18974 7644
rect 18974 7588 18978 7644
rect 18914 7584 18978 7588
rect 18994 7644 19058 7648
rect 18994 7588 18998 7644
rect 18998 7588 19054 7644
rect 19054 7588 19058 7644
rect 18994 7584 19058 7588
rect 24688 7644 24752 7648
rect 24688 7588 24692 7644
rect 24692 7588 24748 7644
rect 24748 7588 24752 7644
rect 24688 7584 24752 7588
rect 24768 7644 24832 7648
rect 24768 7588 24772 7644
rect 24772 7588 24828 7644
rect 24828 7588 24832 7644
rect 24768 7584 24832 7588
rect 24848 7644 24912 7648
rect 24848 7588 24852 7644
rect 24852 7588 24908 7644
rect 24908 7588 24912 7644
rect 24848 7584 24912 7588
rect 24928 7644 24992 7648
rect 24928 7588 24932 7644
rect 24932 7588 24988 7644
rect 24988 7588 24992 7644
rect 24928 7584 24992 7588
rect 20116 7244 20180 7308
rect 3919 7100 3983 7104
rect 3919 7044 3923 7100
rect 3923 7044 3979 7100
rect 3979 7044 3983 7100
rect 3919 7040 3983 7044
rect 3999 7100 4063 7104
rect 3999 7044 4003 7100
rect 4003 7044 4059 7100
rect 4059 7044 4063 7100
rect 3999 7040 4063 7044
rect 4079 7100 4143 7104
rect 4079 7044 4083 7100
rect 4083 7044 4139 7100
rect 4139 7044 4143 7100
rect 4079 7040 4143 7044
rect 4159 7100 4223 7104
rect 4159 7044 4163 7100
rect 4163 7044 4219 7100
rect 4219 7044 4223 7100
rect 4159 7040 4223 7044
rect 9853 7100 9917 7104
rect 9853 7044 9857 7100
rect 9857 7044 9913 7100
rect 9913 7044 9917 7100
rect 9853 7040 9917 7044
rect 9933 7100 9997 7104
rect 9933 7044 9937 7100
rect 9937 7044 9993 7100
rect 9993 7044 9997 7100
rect 9933 7040 9997 7044
rect 10013 7100 10077 7104
rect 10013 7044 10017 7100
rect 10017 7044 10073 7100
rect 10073 7044 10077 7100
rect 10013 7040 10077 7044
rect 10093 7100 10157 7104
rect 10093 7044 10097 7100
rect 10097 7044 10153 7100
rect 10153 7044 10157 7100
rect 10093 7040 10157 7044
rect 15787 7100 15851 7104
rect 15787 7044 15791 7100
rect 15791 7044 15847 7100
rect 15847 7044 15851 7100
rect 15787 7040 15851 7044
rect 15867 7100 15931 7104
rect 15867 7044 15871 7100
rect 15871 7044 15927 7100
rect 15927 7044 15931 7100
rect 15867 7040 15931 7044
rect 15947 7100 16011 7104
rect 15947 7044 15951 7100
rect 15951 7044 16007 7100
rect 16007 7044 16011 7100
rect 15947 7040 16011 7044
rect 16027 7100 16091 7104
rect 16027 7044 16031 7100
rect 16031 7044 16087 7100
rect 16087 7044 16091 7100
rect 16027 7040 16091 7044
rect 21721 7100 21785 7104
rect 21721 7044 21725 7100
rect 21725 7044 21781 7100
rect 21781 7044 21785 7100
rect 21721 7040 21785 7044
rect 21801 7100 21865 7104
rect 21801 7044 21805 7100
rect 21805 7044 21861 7100
rect 21861 7044 21865 7100
rect 21801 7040 21865 7044
rect 21881 7100 21945 7104
rect 21881 7044 21885 7100
rect 21885 7044 21941 7100
rect 21941 7044 21945 7100
rect 21881 7040 21945 7044
rect 21961 7100 22025 7104
rect 21961 7044 21965 7100
rect 21965 7044 22021 7100
rect 22021 7044 22025 7100
rect 21961 7040 22025 7044
rect 6886 6556 6950 6560
rect 6886 6500 6890 6556
rect 6890 6500 6946 6556
rect 6946 6500 6950 6556
rect 6886 6496 6950 6500
rect 6966 6556 7030 6560
rect 6966 6500 6970 6556
rect 6970 6500 7026 6556
rect 7026 6500 7030 6556
rect 6966 6496 7030 6500
rect 7046 6556 7110 6560
rect 7046 6500 7050 6556
rect 7050 6500 7106 6556
rect 7106 6500 7110 6556
rect 7046 6496 7110 6500
rect 7126 6556 7190 6560
rect 7126 6500 7130 6556
rect 7130 6500 7186 6556
rect 7186 6500 7190 6556
rect 7126 6496 7190 6500
rect 12820 6556 12884 6560
rect 12820 6500 12824 6556
rect 12824 6500 12880 6556
rect 12880 6500 12884 6556
rect 12820 6496 12884 6500
rect 12900 6556 12964 6560
rect 12900 6500 12904 6556
rect 12904 6500 12960 6556
rect 12960 6500 12964 6556
rect 12900 6496 12964 6500
rect 12980 6556 13044 6560
rect 12980 6500 12984 6556
rect 12984 6500 13040 6556
rect 13040 6500 13044 6556
rect 12980 6496 13044 6500
rect 13060 6556 13124 6560
rect 13060 6500 13064 6556
rect 13064 6500 13120 6556
rect 13120 6500 13124 6556
rect 13060 6496 13124 6500
rect 18754 6556 18818 6560
rect 18754 6500 18758 6556
rect 18758 6500 18814 6556
rect 18814 6500 18818 6556
rect 18754 6496 18818 6500
rect 18834 6556 18898 6560
rect 18834 6500 18838 6556
rect 18838 6500 18894 6556
rect 18894 6500 18898 6556
rect 18834 6496 18898 6500
rect 18914 6556 18978 6560
rect 18914 6500 18918 6556
rect 18918 6500 18974 6556
rect 18974 6500 18978 6556
rect 18914 6496 18978 6500
rect 18994 6556 19058 6560
rect 18994 6500 18998 6556
rect 18998 6500 19054 6556
rect 19054 6500 19058 6556
rect 18994 6496 19058 6500
rect 24688 6556 24752 6560
rect 24688 6500 24692 6556
rect 24692 6500 24748 6556
rect 24748 6500 24752 6556
rect 24688 6496 24752 6500
rect 24768 6556 24832 6560
rect 24768 6500 24772 6556
rect 24772 6500 24828 6556
rect 24828 6500 24832 6556
rect 24768 6496 24832 6500
rect 24848 6556 24912 6560
rect 24848 6500 24852 6556
rect 24852 6500 24908 6556
rect 24908 6500 24912 6556
rect 24848 6496 24912 6500
rect 24928 6556 24992 6560
rect 24928 6500 24932 6556
rect 24932 6500 24988 6556
rect 24988 6500 24992 6556
rect 24928 6496 24992 6500
rect 3919 6012 3983 6016
rect 3919 5956 3923 6012
rect 3923 5956 3979 6012
rect 3979 5956 3983 6012
rect 3919 5952 3983 5956
rect 3999 6012 4063 6016
rect 3999 5956 4003 6012
rect 4003 5956 4059 6012
rect 4059 5956 4063 6012
rect 3999 5952 4063 5956
rect 4079 6012 4143 6016
rect 4079 5956 4083 6012
rect 4083 5956 4139 6012
rect 4139 5956 4143 6012
rect 4079 5952 4143 5956
rect 4159 6012 4223 6016
rect 4159 5956 4163 6012
rect 4163 5956 4219 6012
rect 4219 5956 4223 6012
rect 4159 5952 4223 5956
rect 9853 6012 9917 6016
rect 9853 5956 9857 6012
rect 9857 5956 9913 6012
rect 9913 5956 9917 6012
rect 9853 5952 9917 5956
rect 9933 6012 9997 6016
rect 9933 5956 9937 6012
rect 9937 5956 9993 6012
rect 9993 5956 9997 6012
rect 9933 5952 9997 5956
rect 10013 6012 10077 6016
rect 10013 5956 10017 6012
rect 10017 5956 10073 6012
rect 10073 5956 10077 6012
rect 10013 5952 10077 5956
rect 10093 6012 10157 6016
rect 10093 5956 10097 6012
rect 10097 5956 10153 6012
rect 10153 5956 10157 6012
rect 10093 5952 10157 5956
rect 15787 6012 15851 6016
rect 15787 5956 15791 6012
rect 15791 5956 15847 6012
rect 15847 5956 15851 6012
rect 15787 5952 15851 5956
rect 15867 6012 15931 6016
rect 15867 5956 15871 6012
rect 15871 5956 15927 6012
rect 15927 5956 15931 6012
rect 15867 5952 15931 5956
rect 15947 6012 16011 6016
rect 15947 5956 15951 6012
rect 15951 5956 16007 6012
rect 16007 5956 16011 6012
rect 15947 5952 16011 5956
rect 16027 6012 16091 6016
rect 16027 5956 16031 6012
rect 16031 5956 16087 6012
rect 16087 5956 16091 6012
rect 16027 5952 16091 5956
rect 21721 6012 21785 6016
rect 21721 5956 21725 6012
rect 21725 5956 21781 6012
rect 21781 5956 21785 6012
rect 21721 5952 21785 5956
rect 21801 6012 21865 6016
rect 21801 5956 21805 6012
rect 21805 5956 21861 6012
rect 21861 5956 21865 6012
rect 21801 5952 21865 5956
rect 21881 6012 21945 6016
rect 21881 5956 21885 6012
rect 21885 5956 21941 6012
rect 21941 5956 21945 6012
rect 21881 5952 21945 5956
rect 21961 6012 22025 6016
rect 21961 5956 21965 6012
rect 21965 5956 22021 6012
rect 22021 5956 22025 6012
rect 21961 5952 22025 5956
rect 2636 5476 2700 5540
rect 22692 5476 22756 5540
rect 6886 5468 6950 5472
rect 6886 5412 6890 5468
rect 6890 5412 6946 5468
rect 6946 5412 6950 5468
rect 6886 5408 6950 5412
rect 6966 5468 7030 5472
rect 6966 5412 6970 5468
rect 6970 5412 7026 5468
rect 7026 5412 7030 5468
rect 6966 5408 7030 5412
rect 7046 5468 7110 5472
rect 7046 5412 7050 5468
rect 7050 5412 7106 5468
rect 7106 5412 7110 5468
rect 7046 5408 7110 5412
rect 7126 5468 7190 5472
rect 7126 5412 7130 5468
rect 7130 5412 7186 5468
rect 7186 5412 7190 5468
rect 7126 5408 7190 5412
rect 12820 5468 12884 5472
rect 12820 5412 12824 5468
rect 12824 5412 12880 5468
rect 12880 5412 12884 5468
rect 12820 5408 12884 5412
rect 12900 5468 12964 5472
rect 12900 5412 12904 5468
rect 12904 5412 12960 5468
rect 12960 5412 12964 5468
rect 12900 5408 12964 5412
rect 12980 5468 13044 5472
rect 12980 5412 12984 5468
rect 12984 5412 13040 5468
rect 13040 5412 13044 5468
rect 12980 5408 13044 5412
rect 13060 5468 13124 5472
rect 13060 5412 13064 5468
rect 13064 5412 13120 5468
rect 13120 5412 13124 5468
rect 13060 5408 13124 5412
rect 18754 5468 18818 5472
rect 18754 5412 18758 5468
rect 18758 5412 18814 5468
rect 18814 5412 18818 5468
rect 18754 5408 18818 5412
rect 18834 5468 18898 5472
rect 18834 5412 18838 5468
rect 18838 5412 18894 5468
rect 18894 5412 18898 5468
rect 18834 5408 18898 5412
rect 18914 5468 18978 5472
rect 18914 5412 18918 5468
rect 18918 5412 18974 5468
rect 18974 5412 18978 5468
rect 18914 5408 18978 5412
rect 18994 5468 19058 5472
rect 18994 5412 18998 5468
rect 18998 5412 19054 5468
rect 19054 5412 19058 5468
rect 18994 5408 19058 5412
rect 24688 5468 24752 5472
rect 24688 5412 24692 5468
rect 24692 5412 24748 5468
rect 24748 5412 24752 5468
rect 24688 5408 24752 5412
rect 24768 5468 24832 5472
rect 24768 5412 24772 5468
rect 24772 5412 24828 5468
rect 24828 5412 24832 5468
rect 24768 5408 24832 5412
rect 24848 5468 24912 5472
rect 24848 5412 24852 5468
rect 24852 5412 24908 5468
rect 24908 5412 24912 5468
rect 24848 5408 24912 5412
rect 24928 5468 24992 5472
rect 24928 5412 24932 5468
rect 24932 5412 24988 5468
rect 24988 5412 24992 5468
rect 24928 5408 24992 5412
rect 13308 5400 13372 5404
rect 13308 5344 13322 5400
rect 13322 5344 13372 5400
rect 13308 5340 13372 5344
rect 11836 5204 11900 5268
rect 14596 5204 14660 5268
rect 3919 4924 3983 4928
rect 3919 4868 3923 4924
rect 3923 4868 3979 4924
rect 3979 4868 3983 4924
rect 3919 4864 3983 4868
rect 3999 4924 4063 4928
rect 3999 4868 4003 4924
rect 4003 4868 4059 4924
rect 4059 4868 4063 4924
rect 3999 4864 4063 4868
rect 4079 4924 4143 4928
rect 4079 4868 4083 4924
rect 4083 4868 4139 4924
rect 4139 4868 4143 4924
rect 4079 4864 4143 4868
rect 4159 4924 4223 4928
rect 4159 4868 4163 4924
rect 4163 4868 4219 4924
rect 4219 4868 4223 4924
rect 4159 4864 4223 4868
rect 9853 4924 9917 4928
rect 9853 4868 9857 4924
rect 9857 4868 9913 4924
rect 9913 4868 9917 4924
rect 9853 4864 9917 4868
rect 9933 4924 9997 4928
rect 9933 4868 9937 4924
rect 9937 4868 9993 4924
rect 9993 4868 9997 4924
rect 9933 4864 9997 4868
rect 10013 4924 10077 4928
rect 10013 4868 10017 4924
rect 10017 4868 10073 4924
rect 10073 4868 10077 4924
rect 10013 4864 10077 4868
rect 10093 4924 10157 4928
rect 10093 4868 10097 4924
rect 10097 4868 10153 4924
rect 10153 4868 10157 4924
rect 10093 4864 10157 4868
rect 15787 4924 15851 4928
rect 15787 4868 15791 4924
rect 15791 4868 15847 4924
rect 15847 4868 15851 4924
rect 15787 4864 15851 4868
rect 15867 4924 15931 4928
rect 15867 4868 15871 4924
rect 15871 4868 15927 4924
rect 15927 4868 15931 4924
rect 15867 4864 15931 4868
rect 15947 4924 16011 4928
rect 15947 4868 15951 4924
rect 15951 4868 16007 4924
rect 16007 4868 16011 4924
rect 15947 4864 16011 4868
rect 16027 4924 16091 4928
rect 16027 4868 16031 4924
rect 16031 4868 16087 4924
rect 16087 4868 16091 4924
rect 16027 4864 16091 4868
rect 21721 4924 21785 4928
rect 21721 4868 21725 4924
rect 21725 4868 21781 4924
rect 21781 4868 21785 4924
rect 21721 4864 21785 4868
rect 21801 4924 21865 4928
rect 21801 4868 21805 4924
rect 21805 4868 21861 4924
rect 21861 4868 21865 4924
rect 21801 4864 21865 4868
rect 21881 4924 21945 4928
rect 21881 4868 21885 4924
rect 21885 4868 21941 4924
rect 21941 4868 21945 4924
rect 21881 4864 21945 4868
rect 21961 4924 22025 4928
rect 21961 4868 21965 4924
rect 21965 4868 22021 4924
rect 22021 4868 22025 4924
rect 21961 4864 22025 4868
rect 3004 4720 3068 4724
rect 3004 4664 3018 4720
rect 3018 4664 3068 4720
rect 3004 4660 3068 4664
rect 6886 4380 6950 4384
rect 6886 4324 6890 4380
rect 6890 4324 6946 4380
rect 6946 4324 6950 4380
rect 6886 4320 6950 4324
rect 6966 4380 7030 4384
rect 6966 4324 6970 4380
rect 6970 4324 7026 4380
rect 7026 4324 7030 4380
rect 6966 4320 7030 4324
rect 7046 4380 7110 4384
rect 7046 4324 7050 4380
rect 7050 4324 7106 4380
rect 7106 4324 7110 4380
rect 7046 4320 7110 4324
rect 7126 4380 7190 4384
rect 7126 4324 7130 4380
rect 7130 4324 7186 4380
rect 7186 4324 7190 4380
rect 7126 4320 7190 4324
rect 12820 4380 12884 4384
rect 12820 4324 12824 4380
rect 12824 4324 12880 4380
rect 12880 4324 12884 4380
rect 12820 4320 12884 4324
rect 12900 4380 12964 4384
rect 12900 4324 12904 4380
rect 12904 4324 12960 4380
rect 12960 4324 12964 4380
rect 12900 4320 12964 4324
rect 12980 4380 13044 4384
rect 12980 4324 12984 4380
rect 12984 4324 13040 4380
rect 13040 4324 13044 4380
rect 12980 4320 13044 4324
rect 13060 4380 13124 4384
rect 13060 4324 13064 4380
rect 13064 4324 13120 4380
rect 13120 4324 13124 4380
rect 13060 4320 13124 4324
rect 18754 4380 18818 4384
rect 18754 4324 18758 4380
rect 18758 4324 18814 4380
rect 18814 4324 18818 4380
rect 18754 4320 18818 4324
rect 18834 4380 18898 4384
rect 18834 4324 18838 4380
rect 18838 4324 18894 4380
rect 18894 4324 18898 4380
rect 18834 4320 18898 4324
rect 18914 4380 18978 4384
rect 18914 4324 18918 4380
rect 18918 4324 18974 4380
rect 18974 4324 18978 4380
rect 18914 4320 18978 4324
rect 18994 4380 19058 4384
rect 18994 4324 18998 4380
rect 18998 4324 19054 4380
rect 19054 4324 19058 4380
rect 18994 4320 19058 4324
rect 4292 3980 4356 4044
rect 13860 4116 13924 4180
rect 19748 4116 19812 4180
rect 24688 4380 24752 4384
rect 24688 4324 24692 4380
rect 24692 4324 24748 4380
rect 24748 4324 24752 4380
rect 24688 4320 24752 4324
rect 24768 4380 24832 4384
rect 24768 4324 24772 4380
rect 24772 4324 24828 4380
rect 24828 4324 24832 4380
rect 24768 4320 24832 4324
rect 24848 4380 24912 4384
rect 24848 4324 24852 4380
rect 24852 4324 24908 4380
rect 24908 4324 24912 4380
rect 24848 4320 24912 4324
rect 24928 4380 24992 4384
rect 24928 4324 24932 4380
rect 24932 4324 24988 4380
rect 24988 4324 24992 4380
rect 24928 4320 24992 4324
rect 12204 4040 12268 4044
rect 12204 3984 12218 4040
rect 12218 3984 12268 4040
rect 12204 3980 12268 3984
rect 17724 4040 17788 4044
rect 17724 3984 17738 4040
rect 17738 3984 17788 4040
rect 17724 3980 17788 3984
rect 19564 3904 19628 3908
rect 19564 3848 19578 3904
rect 19578 3848 19628 3904
rect 19564 3844 19628 3848
rect 21220 3904 21284 3908
rect 21220 3848 21234 3904
rect 21234 3848 21284 3904
rect 21220 3844 21284 3848
rect 21404 3904 21468 3908
rect 21404 3848 21454 3904
rect 21454 3848 21468 3904
rect 21404 3844 21468 3848
rect 3919 3836 3983 3840
rect 3919 3780 3923 3836
rect 3923 3780 3979 3836
rect 3979 3780 3983 3836
rect 3919 3776 3983 3780
rect 3999 3836 4063 3840
rect 3999 3780 4003 3836
rect 4003 3780 4059 3836
rect 4059 3780 4063 3836
rect 3999 3776 4063 3780
rect 4079 3836 4143 3840
rect 4079 3780 4083 3836
rect 4083 3780 4139 3836
rect 4139 3780 4143 3836
rect 4079 3776 4143 3780
rect 4159 3836 4223 3840
rect 4159 3780 4163 3836
rect 4163 3780 4219 3836
rect 4219 3780 4223 3836
rect 4159 3776 4223 3780
rect 9853 3836 9917 3840
rect 9853 3780 9857 3836
rect 9857 3780 9913 3836
rect 9913 3780 9917 3836
rect 9853 3776 9917 3780
rect 9933 3836 9997 3840
rect 9933 3780 9937 3836
rect 9937 3780 9993 3836
rect 9993 3780 9997 3836
rect 9933 3776 9997 3780
rect 10013 3836 10077 3840
rect 10013 3780 10017 3836
rect 10017 3780 10073 3836
rect 10073 3780 10077 3836
rect 10013 3776 10077 3780
rect 10093 3836 10157 3840
rect 10093 3780 10097 3836
rect 10097 3780 10153 3836
rect 10153 3780 10157 3836
rect 10093 3776 10157 3780
rect 15787 3836 15851 3840
rect 15787 3780 15791 3836
rect 15791 3780 15847 3836
rect 15847 3780 15851 3836
rect 15787 3776 15851 3780
rect 15867 3836 15931 3840
rect 15867 3780 15871 3836
rect 15871 3780 15927 3836
rect 15927 3780 15931 3836
rect 15867 3776 15931 3780
rect 15947 3836 16011 3840
rect 15947 3780 15951 3836
rect 15951 3780 16007 3836
rect 16007 3780 16011 3836
rect 15947 3776 16011 3780
rect 16027 3836 16091 3840
rect 16027 3780 16031 3836
rect 16031 3780 16087 3836
rect 16087 3780 16091 3836
rect 16027 3776 16091 3780
rect 21721 3836 21785 3840
rect 21721 3780 21725 3836
rect 21725 3780 21781 3836
rect 21781 3780 21785 3836
rect 21721 3776 21785 3780
rect 21801 3836 21865 3840
rect 21801 3780 21805 3836
rect 21805 3780 21861 3836
rect 21861 3780 21865 3836
rect 21801 3776 21865 3780
rect 21881 3836 21945 3840
rect 21881 3780 21885 3836
rect 21885 3780 21941 3836
rect 21941 3780 21945 3836
rect 21881 3776 21945 3780
rect 21961 3836 22025 3840
rect 21961 3780 21965 3836
rect 21965 3780 22021 3836
rect 22021 3780 22025 3836
rect 21961 3776 22025 3780
rect 10916 3436 10980 3500
rect 796 3300 860 3364
rect 6886 3292 6950 3296
rect 6886 3236 6890 3292
rect 6890 3236 6946 3292
rect 6946 3236 6950 3292
rect 6886 3232 6950 3236
rect 6966 3292 7030 3296
rect 6966 3236 6970 3292
rect 6970 3236 7026 3292
rect 7026 3236 7030 3292
rect 6966 3232 7030 3236
rect 7046 3292 7110 3296
rect 7046 3236 7050 3292
rect 7050 3236 7106 3292
rect 7106 3236 7110 3292
rect 7046 3232 7110 3236
rect 7126 3292 7190 3296
rect 7126 3236 7130 3292
rect 7130 3236 7186 3292
rect 7186 3236 7190 3292
rect 7126 3232 7190 3236
rect 12820 3292 12884 3296
rect 12820 3236 12824 3292
rect 12824 3236 12880 3292
rect 12880 3236 12884 3292
rect 12820 3232 12884 3236
rect 12900 3292 12964 3296
rect 12900 3236 12904 3292
rect 12904 3236 12960 3292
rect 12960 3236 12964 3292
rect 12900 3232 12964 3236
rect 12980 3292 13044 3296
rect 12980 3236 12984 3292
rect 12984 3236 13040 3292
rect 13040 3236 13044 3292
rect 12980 3232 13044 3236
rect 13060 3292 13124 3296
rect 13060 3236 13064 3292
rect 13064 3236 13120 3292
rect 13120 3236 13124 3292
rect 13060 3232 13124 3236
rect 18754 3292 18818 3296
rect 18754 3236 18758 3292
rect 18758 3236 18814 3292
rect 18814 3236 18818 3292
rect 18754 3232 18818 3236
rect 18834 3292 18898 3296
rect 18834 3236 18838 3292
rect 18838 3236 18894 3292
rect 18894 3236 18898 3292
rect 18834 3232 18898 3236
rect 18914 3292 18978 3296
rect 18914 3236 18918 3292
rect 18918 3236 18974 3292
rect 18974 3236 18978 3292
rect 18914 3232 18978 3236
rect 18994 3292 19058 3296
rect 18994 3236 18998 3292
rect 18998 3236 19054 3292
rect 19054 3236 19058 3292
rect 18994 3232 19058 3236
rect 24688 3292 24752 3296
rect 24688 3236 24692 3292
rect 24692 3236 24748 3292
rect 24748 3236 24752 3292
rect 24688 3232 24752 3236
rect 24768 3292 24832 3296
rect 24768 3236 24772 3292
rect 24772 3236 24828 3292
rect 24828 3236 24832 3292
rect 24768 3232 24832 3236
rect 24848 3292 24912 3296
rect 24848 3236 24852 3292
rect 24852 3236 24908 3292
rect 24908 3236 24912 3292
rect 24848 3232 24912 3236
rect 24928 3292 24992 3296
rect 24928 3236 24932 3292
rect 24932 3236 24988 3292
rect 24988 3236 24992 3292
rect 24928 3232 24992 3236
rect 3919 2748 3983 2752
rect 3919 2692 3923 2748
rect 3923 2692 3979 2748
rect 3979 2692 3983 2748
rect 3919 2688 3983 2692
rect 3999 2748 4063 2752
rect 3999 2692 4003 2748
rect 4003 2692 4059 2748
rect 4059 2692 4063 2748
rect 3999 2688 4063 2692
rect 4079 2748 4143 2752
rect 4079 2692 4083 2748
rect 4083 2692 4139 2748
rect 4139 2692 4143 2748
rect 4079 2688 4143 2692
rect 4159 2748 4223 2752
rect 4159 2692 4163 2748
rect 4163 2692 4219 2748
rect 4219 2692 4223 2748
rect 4159 2688 4223 2692
rect 9853 2748 9917 2752
rect 9853 2692 9857 2748
rect 9857 2692 9913 2748
rect 9913 2692 9917 2748
rect 9853 2688 9917 2692
rect 9933 2748 9997 2752
rect 9933 2692 9937 2748
rect 9937 2692 9993 2748
rect 9993 2692 9997 2748
rect 9933 2688 9997 2692
rect 10013 2748 10077 2752
rect 10013 2692 10017 2748
rect 10017 2692 10073 2748
rect 10073 2692 10077 2748
rect 10013 2688 10077 2692
rect 10093 2748 10157 2752
rect 10093 2692 10097 2748
rect 10097 2692 10153 2748
rect 10153 2692 10157 2748
rect 10093 2688 10157 2692
rect 15787 2748 15851 2752
rect 15787 2692 15791 2748
rect 15791 2692 15847 2748
rect 15847 2692 15851 2748
rect 15787 2688 15851 2692
rect 15867 2748 15931 2752
rect 15867 2692 15871 2748
rect 15871 2692 15927 2748
rect 15927 2692 15931 2748
rect 15867 2688 15931 2692
rect 15947 2748 16011 2752
rect 15947 2692 15951 2748
rect 15951 2692 16007 2748
rect 16007 2692 16011 2748
rect 15947 2688 16011 2692
rect 16027 2748 16091 2752
rect 16027 2692 16031 2748
rect 16031 2692 16087 2748
rect 16087 2692 16091 2748
rect 16027 2688 16091 2692
rect 21721 2748 21785 2752
rect 21721 2692 21725 2748
rect 21725 2692 21781 2748
rect 21781 2692 21785 2748
rect 21721 2688 21785 2692
rect 21801 2748 21865 2752
rect 21801 2692 21805 2748
rect 21805 2692 21861 2748
rect 21861 2692 21865 2748
rect 21801 2688 21865 2692
rect 21881 2748 21945 2752
rect 21881 2692 21885 2748
rect 21885 2692 21941 2748
rect 21941 2692 21945 2748
rect 21881 2688 21945 2692
rect 21961 2748 22025 2752
rect 21961 2692 21965 2748
rect 21965 2692 22021 2748
rect 22021 2692 22025 2748
rect 21961 2688 22025 2692
rect 9444 2680 9508 2684
rect 9444 2624 9458 2680
rect 9458 2624 9508 2680
rect 9444 2620 9508 2624
rect 12020 2680 12084 2684
rect 12020 2624 12034 2680
rect 12034 2624 12084 2680
rect 12020 2620 12084 2624
rect 14780 2680 14844 2684
rect 14780 2624 14830 2680
rect 14830 2624 14844 2680
rect 14780 2620 14844 2624
rect 15516 2680 15580 2684
rect 15516 2624 15530 2680
rect 15530 2624 15580 2680
rect 15516 2620 15580 2624
rect 17540 2680 17604 2684
rect 17540 2624 17554 2680
rect 17554 2624 17604 2680
rect 17540 2620 17604 2624
rect 18460 2620 18524 2684
rect 19748 2620 19812 2684
rect 9628 2484 9692 2548
rect 13492 2484 13556 2548
rect 5028 2212 5092 2276
rect 7788 2272 7852 2276
rect 7788 2216 7802 2272
rect 7802 2216 7852 2272
rect 7788 2212 7852 2216
rect 8156 2272 8220 2276
rect 8156 2216 8170 2272
rect 8170 2216 8220 2272
rect 8156 2212 8220 2216
rect 8524 2272 8588 2276
rect 8524 2216 8538 2272
rect 8538 2216 8588 2272
rect 8524 2212 8588 2216
rect 8892 2272 8956 2276
rect 8892 2216 8906 2272
rect 8906 2216 8956 2272
rect 8892 2212 8956 2216
rect 16252 2484 16316 2548
rect 16988 2544 17052 2548
rect 16988 2488 17002 2544
rect 17002 2488 17052 2544
rect 16988 2484 17052 2488
rect 21588 2484 21652 2548
rect 19380 2348 19444 2412
rect 19564 2408 19628 2412
rect 19564 2352 19614 2408
rect 19614 2352 19628 2408
rect 19564 2348 19628 2352
rect 6886 2204 6950 2208
rect 6886 2148 6890 2204
rect 6890 2148 6946 2204
rect 6946 2148 6950 2204
rect 6886 2144 6950 2148
rect 6966 2204 7030 2208
rect 6966 2148 6970 2204
rect 6970 2148 7026 2204
rect 7026 2148 7030 2204
rect 6966 2144 7030 2148
rect 7046 2204 7110 2208
rect 7046 2148 7050 2204
rect 7050 2148 7106 2204
rect 7106 2148 7110 2204
rect 7046 2144 7110 2148
rect 7126 2204 7190 2208
rect 7126 2148 7130 2204
rect 7130 2148 7186 2204
rect 7186 2148 7190 2204
rect 7126 2144 7190 2148
rect 12820 2204 12884 2208
rect 12820 2148 12824 2204
rect 12824 2148 12880 2204
rect 12880 2148 12884 2204
rect 12820 2144 12884 2148
rect 12900 2204 12964 2208
rect 12900 2148 12904 2204
rect 12904 2148 12960 2204
rect 12960 2148 12964 2204
rect 12900 2144 12964 2148
rect 12980 2204 13044 2208
rect 12980 2148 12984 2204
rect 12984 2148 13040 2204
rect 13040 2148 13044 2204
rect 12980 2144 13044 2148
rect 13060 2204 13124 2208
rect 13060 2148 13064 2204
rect 13064 2148 13120 2204
rect 13120 2148 13124 2204
rect 13060 2144 13124 2148
rect 18754 2204 18818 2208
rect 18754 2148 18758 2204
rect 18758 2148 18814 2204
rect 18814 2148 18818 2204
rect 18754 2144 18818 2148
rect 18834 2204 18898 2208
rect 18834 2148 18838 2204
rect 18838 2148 18894 2204
rect 18894 2148 18898 2204
rect 18834 2144 18898 2148
rect 18914 2204 18978 2208
rect 18914 2148 18918 2204
rect 18918 2148 18974 2204
rect 18974 2148 18978 2204
rect 18914 2144 18978 2148
rect 18994 2204 19058 2208
rect 18994 2148 18998 2204
rect 18998 2148 19054 2204
rect 19054 2148 19058 2204
rect 18994 2144 19058 2148
rect 24688 2204 24752 2208
rect 24688 2148 24692 2204
rect 24692 2148 24748 2204
rect 24748 2148 24752 2204
rect 24688 2144 24752 2148
rect 24768 2204 24832 2208
rect 24768 2148 24772 2204
rect 24772 2148 24828 2204
rect 24828 2148 24832 2204
rect 24768 2144 24832 2148
rect 24848 2204 24912 2208
rect 24848 2148 24852 2204
rect 24852 2148 24908 2204
rect 24908 2148 24912 2204
rect 24848 2144 24912 2148
rect 24928 2204 24992 2208
rect 24928 2148 24932 2204
rect 24932 2148 24988 2204
rect 24988 2148 24992 2204
rect 24928 2144 24992 2148
rect 1164 1940 1228 2004
rect 5580 2000 5644 2004
rect 5580 1944 5594 2000
rect 5594 1944 5644 2000
rect 5580 1940 5644 1944
rect 6316 1940 6380 2004
rect 3919 1660 3983 1664
rect 3919 1604 3923 1660
rect 3923 1604 3979 1660
rect 3979 1604 3983 1660
rect 3919 1600 3983 1604
rect 3999 1660 4063 1664
rect 3999 1604 4003 1660
rect 4003 1604 4059 1660
rect 4059 1604 4063 1660
rect 3999 1600 4063 1604
rect 4079 1660 4143 1664
rect 4079 1604 4083 1660
rect 4083 1604 4139 1660
rect 4139 1604 4143 1660
rect 4079 1600 4143 1604
rect 4159 1660 4223 1664
rect 4159 1604 4163 1660
rect 4163 1604 4219 1660
rect 4219 1604 4223 1660
rect 4159 1600 4223 1604
rect 9853 1660 9917 1664
rect 9853 1604 9857 1660
rect 9857 1604 9913 1660
rect 9913 1604 9917 1660
rect 9853 1600 9917 1604
rect 9933 1660 9997 1664
rect 9933 1604 9937 1660
rect 9937 1604 9993 1660
rect 9993 1604 9997 1660
rect 9933 1600 9997 1604
rect 10013 1660 10077 1664
rect 10013 1604 10017 1660
rect 10017 1604 10073 1660
rect 10073 1604 10077 1660
rect 10013 1600 10077 1604
rect 10093 1660 10157 1664
rect 10093 1604 10097 1660
rect 10097 1604 10153 1660
rect 10153 1604 10157 1660
rect 10093 1600 10157 1604
rect 15787 1660 15851 1664
rect 15787 1604 15791 1660
rect 15791 1604 15847 1660
rect 15847 1604 15851 1660
rect 15787 1600 15851 1604
rect 15867 1660 15931 1664
rect 15867 1604 15871 1660
rect 15871 1604 15927 1660
rect 15927 1604 15931 1660
rect 15867 1600 15931 1604
rect 15947 1660 16011 1664
rect 15947 1604 15951 1660
rect 15951 1604 16007 1660
rect 16007 1604 16011 1660
rect 15947 1600 16011 1604
rect 16027 1660 16091 1664
rect 16027 1604 16031 1660
rect 16031 1604 16087 1660
rect 16087 1604 16091 1660
rect 16027 1600 16091 1604
rect 21721 1660 21785 1664
rect 21721 1604 21725 1660
rect 21725 1604 21781 1660
rect 21781 1604 21785 1660
rect 21721 1600 21785 1604
rect 21801 1660 21865 1664
rect 21801 1604 21805 1660
rect 21805 1604 21861 1660
rect 21861 1604 21865 1660
rect 21801 1600 21865 1604
rect 21881 1660 21945 1664
rect 21881 1604 21885 1660
rect 21885 1604 21941 1660
rect 21941 1604 21945 1660
rect 21881 1600 21945 1604
rect 21961 1660 22025 1664
rect 21961 1604 21965 1660
rect 21965 1604 22021 1660
rect 22021 1604 22025 1660
rect 21961 1600 22025 1604
rect 1716 1320 1780 1324
rect 1716 1264 1730 1320
rect 1730 1264 1780 1320
rect 1716 1260 1780 1264
rect 2084 1320 2148 1324
rect 2084 1264 2098 1320
rect 2098 1264 2148 1320
rect 2084 1260 2148 1264
rect 4476 1320 4540 1324
rect 4476 1264 4490 1320
rect 4490 1264 4540 1320
rect 4476 1260 4540 1264
rect 16436 1320 16500 1324
rect 16436 1264 16486 1320
rect 16486 1264 16500 1320
rect 980 1124 1044 1188
rect 16436 1260 16500 1264
rect 18092 1260 18156 1324
rect 19932 1260 19996 1324
rect 6886 1116 6950 1120
rect 6886 1060 6890 1116
rect 6890 1060 6946 1116
rect 6946 1060 6950 1116
rect 6886 1056 6950 1060
rect 6966 1116 7030 1120
rect 6966 1060 6970 1116
rect 6970 1060 7026 1116
rect 7026 1060 7030 1116
rect 6966 1056 7030 1060
rect 7046 1116 7110 1120
rect 7046 1060 7050 1116
rect 7050 1060 7106 1116
rect 7106 1060 7110 1116
rect 7046 1056 7110 1060
rect 7126 1116 7190 1120
rect 7126 1060 7130 1116
rect 7130 1060 7186 1116
rect 7186 1060 7190 1116
rect 7126 1056 7190 1060
rect 12820 1116 12884 1120
rect 12820 1060 12824 1116
rect 12824 1060 12880 1116
rect 12880 1060 12884 1116
rect 12820 1056 12884 1060
rect 12900 1116 12964 1120
rect 12900 1060 12904 1116
rect 12904 1060 12960 1116
rect 12960 1060 12964 1116
rect 12900 1056 12964 1060
rect 12980 1116 13044 1120
rect 12980 1060 12984 1116
rect 12984 1060 13040 1116
rect 13040 1060 13044 1116
rect 12980 1056 13044 1060
rect 13060 1116 13124 1120
rect 13060 1060 13064 1116
rect 13064 1060 13120 1116
rect 13120 1060 13124 1116
rect 13060 1056 13124 1060
rect 18754 1116 18818 1120
rect 18754 1060 18758 1116
rect 18758 1060 18814 1116
rect 18814 1060 18818 1116
rect 18754 1056 18818 1060
rect 18834 1116 18898 1120
rect 18834 1060 18838 1116
rect 18838 1060 18894 1116
rect 18894 1060 18898 1116
rect 18834 1056 18898 1060
rect 18914 1116 18978 1120
rect 18914 1060 18918 1116
rect 18918 1060 18974 1116
rect 18974 1060 18978 1116
rect 18914 1056 18978 1060
rect 18994 1116 19058 1120
rect 18994 1060 18998 1116
rect 18998 1060 19054 1116
rect 19054 1060 19058 1116
rect 18994 1056 19058 1060
rect 24688 1116 24752 1120
rect 24688 1060 24692 1116
rect 24692 1060 24748 1116
rect 24748 1060 24752 1116
rect 24688 1056 24752 1060
rect 24768 1116 24832 1120
rect 24768 1060 24772 1116
rect 24772 1060 24828 1116
rect 24828 1060 24832 1116
rect 24768 1056 24832 1060
rect 24848 1116 24912 1120
rect 24848 1060 24852 1116
rect 24852 1060 24908 1116
rect 24908 1060 24912 1116
rect 24848 1056 24912 1060
rect 24928 1116 24992 1120
rect 24928 1060 24932 1116
rect 24932 1060 24988 1116
rect 24988 1060 24992 1116
rect 24928 1056 24992 1060
rect 17908 852 17972 916
rect 8708 716 8772 780
<< metal4 >>
rect 3911 43008 4231 43568
rect 3911 42944 3919 43008
rect 3983 42944 3999 43008
rect 4063 42944 4079 43008
rect 4143 42944 4159 43008
rect 4223 42944 4231 43008
rect 3911 41920 4231 42944
rect 3911 41856 3919 41920
rect 3983 41856 3999 41920
rect 4063 41856 4079 41920
rect 4143 41856 4159 41920
rect 4223 41856 4231 41920
rect 1163 41580 1229 41581
rect 1163 41516 1164 41580
rect 1228 41516 1229 41580
rect 1163 41515 1229 41516
rect 611 38588 677 38589
rect 611 38524 612 38588
rect 676 38524 677 38588
rect 611 38523 677 38524
rect 614 8669 674 38523
rect 979 38044 1045 38045
rect 979 37980 980 38044
rect 1044 37980 1045 38044
rect 979 37979 1045 37980
rect 795 36684 861 36685
rect 795 36620 796 36684
rect 860 36620 861 36684
rect 795 36619 861 36620
rect 611 8668 677 8669
rect 611 8604 612 8668
rect 676 8604 677 8668
rect 611 8603 677 8604
rect 798 3365 858 36619
rect 795 3364 861 3365
rect 795 3300 796 3364
rect 860 3300 861 3364
rect 795 3299 861 3300
rect 982 1189 1042 37979
rect 1166 2005 1226 41515
rect 3911 40832 4231 41856
rect 6878 43552 7198 43568
rect 6878 43488 6886 43552
rect 6950 43488 6966 43552
rect 7030 43488 7046 43552
rect 7110 43488 7126 43552
rect 7190 43488 7198 43552
rect 6878 42464 7198 43488
rect 6878 42400 6886 42464
rect 6950 42400 6966 42464
rect 7030 42400 7046 42464
rect 7110 42400 7126 42464
rect 7190 42400 7198 42464
rect 6315 41852 6381 41853
rect 6315 41788 6316 41852
rect 6380 41788 6381 41852
rect 6315 41787 6381 41788
rect 6499 41852 6565 41853
rect 6499 41788 6500 41852
rect 6564 41788 6565 41852
rect 6499 41787 6565 41788
rect 4843 41580 4909 41581
rect 4843 41516 4844 41580
rect 4908 41516 4909 41580
rect 4843 41515 4909 41516
rect 3911 40768 3919 40832
rect 3983 40768 3999 40832
rect 4063 40768 4079 40832
rect 4143 40768 4159 40832
rect 4223 40768 4231 40832
rect 2083 40492 2149 40493
rect 2083 40428 2084 40492
rect 2148 40428 2149 40492
rect 2083 40427 2149 40428
rect 1715 40356 1781 40357
rect 1715 40292 1716 40356
rect 1780 40292 1781 40356
rect 1715 40291 1781 40292
rect 1718 27981 1778 40291
rect 1899 38724 1965 38725
rect 1899 38660 1900 38724
rect 1964 38660 1965 38724
rect 1899 38659 1965 38660
rect 1902 33693 1962 38659
rect 1899 33692 1965 33693
rect 1899 33628 1900 33692
rect 1964 33628 1965 33692
rect 1899 33627 1965 33628
rect 2086 31770 2146 40427
rect 3911 39744 4231 40768
rect 3911 39680 3919 39744
rect 3983 39680 3999 39744
rect 4063 39680 4079 39744
rect 4143 39680 4159 39744
rect 4223 39680 4231 39744
rect 3911 38656 4231 39680
rect 3911 38592 3919 38656
rect 3983 38592 3999 38656
rect 4063 38592 4079 38656
rect 4143 38592 4159 38656
rect 4223 38592 4231 38656
rect 3003 38316 3069 38317
rect 3003 38252 3004 38316
rect 3068 38252 3069 38316
rect 3003 38251 3069 38252
rect 3006 32877 3066 38251
rect 3555 37908 3621 37909
rect 3555 37844 3556 37908
rect 3620 37844 3621 37908
rect 3555 37843 3621 37844
rect 3187 35868 3253 35869
rect 3187 35804 3188 35868
rect 3252 35804 3253 35868
rect 3187 35803 3253 35804
rect 3190 35189 3250 35803
rect 3187 35188 3253 35189
rect 3187 35124 3188 35188
rect 3252 35124 3253 35188
rect 3187 35123 3253 35124
rect 3558 32877 3618 37843
rect 3911 37568 4231 38592
rect 4659 37772 4725 37773
rect 4659 37708 4660 37772
rect 4724 37708 4725 37772
rect 4659 37707 4725 37708
rect 3911 37504 3919 37568
rect 3983 37504 3999 37568
rect 4063 37504 4079 37568
rect 4143 37504 4159 37568
rect 4223 37504 4231 37568
rect 3911 36480 4231 37504
rect 3911 36416 3919 36480
rect 3983 36416 3999 36480
rect 4063 36416 4079 36480
rect 4143 36416 4159 36480
rect 4223 36416 4231 36480
rect 3911 35392 4231 36416
rect 3911 35328 3919 35392
rect 3983 35328 3999 35392
rect 4063 35328 4079 35392
rect 4143 35328 4159 35392
rect 4223 35328 4231 35392
rect 3911 34304 4231 35328
rect 3911 34240 3919 34304
rect 3983 34240 3999 34304
rect 4063 34240 4079 34304
rect 4143 34240 4159 34304
rect 4223 34240 4231 34304
rect 3911 33216 4231 34240
rect 3911 33152 3919 33216
rect 3983 33152 3999 33216
rect 4063 33152 4079 33216
rect 4143 33152 4159 33216
rect 4223 33152 4231 33216
rect 3003 32876 3069 32877
rect 3003 32812 3004 32876
rect 3068 32812 3069 32876
rect 3003 32811 3069 32812
rect 3555 32876 3621 32877
rect 3555 32812 3556 32876
rect 3620 32812 3621 32876
rect 3555 32811 3621 32812
rect 3911 32128 4231 33152
rect 4475 33148 4541 33149
rect 4475 33084 4476 33148
rect 4540 33084 4541 33148
rect 4475 33083 4541 33084
rect 4291 32876 4357 32877
rect 4291 32812 4292 32876
rect 4356 32812 4357 32876
rect 4291 32811 4357 32812
rect 3911 32064 3919 32128
rect 3983 32064 3999 32128
rect 4063 32064 4079 32128
rect 4143 32064 4159 32128
rect 4223 32064 4231 32128
rect 3555 31788 3621 31789
rect 2086 31710 2330 31770
rect 3555 31724 3556 31788
rect 3620 31724 3621 31788
rect 3555 31723 3621 31724
rect 2083 29476 2149 29477
rect 2083 29412 2084 29476
rect 2148 29412 2149 29476
rect 2083 29411 2149 29412
rect 2086 28525 2146 29411
rect 2083 28524 2149 28525
rect 2083 28460 2084 28524
rect 2148 28460 2149 28524
rect 2083 28459 2149 28460
rect 1715 27980 1781 27981
rect 1715 27916 1716 27980
rect 1780 27916 1781 27980
rect 1715 27915 1781 27916
rect 2086 24853 2146 28459
rect 2270 27165 2330 31710
rect 3187 31244 3253 31245
rect 3187 31180 3188 31244
rect 3252 31180 3253 31244
rect 3187 31179 3253 31180
rect 3190 30021 3250 31179
rect 3187 30020 3253 30021
rect 3187 29956 3188 30020
rect 3252 29956 3253 30020
rect 3187 29955 3253 29956
rect 2451 29612 2517 29613
rect 2451 29548 2452 29612
rect 2516 29548 2517 29612
rect 2451 29547 2517 29548
rect 2267 27164 2333 27165
rect 2267 27100 2268 27164
rect 2332 27100 2333 27164
rect 2267 27099 2333 27100
rect 2083 24852 2149 24853
rect 2083 24788 2084 24852
rect 2148 24788 2149 24852
rect 2083 24787 2149 24788
rect 2270 22110 2330 27099
rect 2086 22050 2330 22110
rect 1347 20908 1413 20909
rect 1347 20844 1348 20908
rect 1412 20844 1413 20908
rect 1347 20843 1413 20844
rect 1350 13837 1410 20843
rect 1347 13836 1413 13837
rect 1347 13772 1348 13836
rect 1412 13772 1413 13836
rect 1347 13771 1413 13772
rect 2086 13429 2146 22050
rect 1715 13428 1781 13429
rect 1715 13364 1716 13428
rect 1780 13364 1781 13428
rect 1715 13363 1781 13364
rect 2083 13428 2149 13429
rect 2083 13364 2084 13428
rect 2148 13364 2149 13428
rect 2083 13363 2149 13364
rect 1163 2004 1229 2005
rect 1163 1940 1164 2004
rect 1228 1940 1229 2004
rect 1163 1939 1229 1940
rect 1718 1325 1778 13363
rect 2083 13292 2149 13293
rect 2083 13228 2084 13292
rect 2148 13228 2149 13292
rect 2083 13227 2149 13228
rect 2086 1325 2146 13227
rect 2454 12749 2514 29547
rect 2635 22132 2701 22133
rect 2635 22068 2636 22132
rect 2700 22068 2701 22132
rect 2635 22067 2701 22068
rect 2451 12748 2517 12749
rect 2451 12684 2452 12748
rect 2516 12684 2517 12748
rect 2451 12683 2517 12684
rect 2638 5541 2698 22067
rect 3190 16149 3250 29955
rect 3558 19685 3618 31723
rect 3911 31040 4231 32064
rect 3911 30976 3919 31040
rect 3983 30976 3999 31040
rect 4063 30976 4079 31040
rect 4143 30976 4159 31040
rect 4223 30976 4231 31040
rect 3911 29952 4231 30976
rect 3911 29888 3919 29952
rect 3983 29888 3999 29952
rect 4063 29888 4079 29952
rect 4143 29888 4159 29952
rect 4223 29888 4231 29952
rect 3911 28864 4231 29888
rect 4294 29341 4354 32811
rect 4478 31925 4538 33083
rect 4475 31924 4541 31925
rect 4475 31860 4476 31924
rect 4540 31860 4541 31924
rect 4475 31859 4541 31860
rect 4291 29340 4357 29341
rect 4291 29276 4292 29340
rect 4356 29276 4357 29340
rect 4291 29275 4357 29276
rect 3911 28800 3919 28864
rect 3983 28800 3999 28864
rect 4063 28800 4079 28864
rect 4143 28800 4159 28864
rect 4223 28800 4231 28864
rect 3911 27776 4231 28800
rect 3911 27712 3919 27776
rect 3983 27712 3999 27776
rect 4063 27712 4079 27776
rect 4143 27712 4159 27776
rect 4223 27712 4231 27776
rect 3911 26688 4231 27712
rect 3911 26624 3919 26688
rect 3983 26624 3999 26688
rect 4063 26624 4079 26688
rect 4143 26624 4159 26688
rect 4223 26624 4231 26688
rect 3911 25600 4231 26624
rect 3911 25536 3919 25600
rect 3983 25536 3999 25600
rect 4063 25536 4079 25600
rect 4143 25536 4159 25600
rect 4223 25536 4231 25600
rect 3911 24512 4231 25536
rect 3911 24448 3919 24512
rect 3983 24448 3999 24512
rect 4063 24448 4079 24512
rect 4143 24448 4159 24512
rect 4223 24448 4231 24512
rect 3911 23424 4231 24448
rect 3911 23360 3919 23424
rect 3983 23360 3999 23424
rect 4063 23360 4079 23424
rect 4143 23360 4159 23424
rect 4223 23360 4231 23424
rect 3911 22336 4231 23360
rect 3911 22272 3919 22336
rect 3983 22272 3999 22336
rect 4063 22272 4079 22336
rect 4143 22272 4159 22336
rect 4223 22272 4231 22336
rect 3911 21248 4231 22272
rect 4478 21997 4538 31859
rect 4662 31381 4722 37707
rect 4659 31380 4725 31381
rect 4659 31316 4660 31380
rect 4724 31316 4725 31380
rect 4659 31315 4725 31316
rect 4662 24853 4722 31315
rect 4846 30293 4906 41515
rect 5579 34916 5645 34917
rect 5579 34852 5580 34916
rect 5644 34852 5645 34916
rect 5579 34851 5645 34852
rect 4843 30292 4909 30293
rect 4843 30228 4844 30292
rect 4908 30228 4909 30292
rect 4843 30227 4909 30228
rect 5211 30020 5277 30021
rect 5211 29956 5212 30020
rect 5276 29956 5277 30020
rect 5211 29955 5277 29956
rect 4843 25260 4909 25261
rect 4843 25196 4844 25260
rect 4908 25196 4909 25260
rect 4843 25195 4909 25196
rect 4659 24852 4725 24853
rect 4659 24788 4660 24852
rect 4724 24788 4725 24852
rect 4659 24787 4725 24788
rect 4659 23492 4725 23493
rect 4659 23428 4660 23492
rect 4724 23428 4725 23492
rect 4659 23427 4725 23428
rect 4475 21996 4541 21997
rect 4475 21932 4476 21996
rect 4540 21932 4541 21996
rect 4475 21931 4541 21932
rect 3911 21184 3919 21248
rect 3983 21184 3999 21248
rect 4063 21184 4079 21248
rect 4143 21184 4159 21248
rect 4223 21184 4231 21248
rect 3911 20160 4231 21184
rect 3911 20096 3919 20160
rect 3983 20096 3999 20160
rect 4063 20096 4079 20160
rect 4143 20096 4159 20160
rect 4223 20096 4231 20160
rect 3555 19684 3621 19685
rect 3555 19620 3556 19684
rect 3620 19620 3621 19684
rect 3555 19619 3621 19620
rect 3911 19072 4231 20096
rect 4475 19276 4541 19277
rect 4475 19212 4476 19276
rect 4540 19212 4541 19276
rect 4475 19211 4541 19212
rect 3911 19008 3919 19072
rect 3983 19008 3999 19072
rect 4063 19008 4079 19072
rect 4143 19008 4159 19072
rect 4223 19008 4231 19072
rect 3911 17984 4231 19008
rect 3911 17920 3919 17984
rect 3983 17920 3999 17984
rect 4063 17920 4079 17984
rect 4143 17920 4159 17984
rect 4223 17920 4231 17984
rect 3911 16896 4231 17920
rect 3911 16832 3919 16896
rect 3983 16832 3999 16896
rect 4063 16832 4079 16896
rect 4143 16832 4159 16896
rect 4223 16832 4231 16896
rect 3187 16148 3253 16149
rect 3187 16084 3188 16148
rect 3252 16084 3253 16148
rect 3187 16083 3253 16084
rect 3911 15808 4231 16832
rect 3911 15744 3919 15808
rect 3983 15744 3999 15808
rect 4063 15744 4079 15808
rect 4143 15744 4159 15808
rect 4223 15744 4231 15808
rect 3911 14720 4231 15744
rect 3911 14656 3919 14720
rect 3983 14656 3999 14720
rect 4063 14656 4079 14720
rect 4143 14656 4159 14720
rect 4223 14656 4231 14720
rect 3003 13836 3069 13837
rect 3003 13772 3004 13836
rect 3068 13772 3069 13836
rect 3003 13771 3069 13772
rect 2635 5540 2701 5541
rect 2635 5476 2636 5540
rect 2700 5476 2701 5540
rect 2635 5475 2701 5476
rect 3006 4725 3066 13771
rect 3911 13632 4231 14656
rect 3911 13568 3919 13632
rect 3983 13568 3999 13632
rect 4063 13568 4079 13632
rect 4143 13568 4159 13632
rect 4223 13568 4231 13632
rect 3911 12544 4231 13568
rect 3911 12480 3919 12544
rect 3983 12480 3999 12544
rect 4063 12480 4079 12544
rect 4143 12480 4159 12544
rect 4223 12480 4231 12544
rect 3911 11456 4231 12480
rect 3911 11392 3919 11456
rect 3983 11392 3999 11456
rect 4063 11392 4079 11456
rect 4143 11392 4159 11456
rect 4223 11392 4231 11456
rect 3911 10368 4231 11392
rect 3911 10304 3919 10368
rect 3983 10304 3999 10368
rect 4063 10304 4079 10368
rect 4143 10304 4159 10368
rect 4223 10304 4231 10368
rect 3911 9280 4231 10304
rect 3911 9216 3919 9280
rect 3983 9216 3999 9280
rect 4063 9216 4079 9280
rect 4143 9216 4159 9280
rect 4223 9216 4231 9280
rect 3911 8192 4231 9216
rect 4291 8668 4357 8669
rect 4291 8604 4292 8668
rect 4356 8604 4357 8668
rect 4291 8603 4357 8604
rect 3911 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4231 8192
rect 3911 7104 4231 8128
rect 3911 7040 3919 7104
rect 3983 7040 3999 7104
rect 4063 7040 4079 7104
rect 4143 7040 4159 7104
rect 4223 7040 4231 7104
rect 3911 6016 4231 7040
rect 3911 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4231 6016
rect 3911 4928 4231 5952
rect 3911 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4231 4928
rect 3003 4724 3069 4725
rect 3003 4660 3004 4724
rect 3068 4660 3069 4724
rect 3003 4659 3069 4660
rect 3911 3840 4231 4864
rect 4294 4045 4354 8603
rect 4291 4044 4357 4045
rect 4291 3980 4292 4044
rect 4356 3980 4357 4044
rect 4291 3979 4357 3980
rect 3911 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4231 3840
rect 3911 2752 4231 3776
rect 3911 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4231 2752
rect 3911 1664 4231 2688
rect 3911 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4231 1664
rect 1715 1324 1781 1325
rect 1715 1260 1716 1324
rect 1780 1260 1781 1324
rect 1715 1259 1781 1260
rect 2083 1324 2149 1325
rect 2083 1260 2084 1324
rect 2148 1260 2149 1324
rect 2083 1259 2149 1260
rect 979 1188 1045 1189
rect 979 1124 980 1188
rect 1044 1124 1045 1188
rect 979 1123 1045 1124
rect 3911 1040 4231 1600
rect 4478 1325 4538 19211
rect 4662 16693 4722 23427
rect 4659 16692 4725 16693
rect 4659 16628 4660 16692
rect 4724 16628 4725 16692
rect 4659 16627 4725 16628
rect 4846 10165 4906 25195
rect 5214 19957 5274 29955
rect 5395 27708 5461 27709
rect 5395 27644 5396 27708
rect 5460 27644 5461 27708
rect 5395 27643 5461 27644
rect 5398 23357 5458 27643
rect 5395 23356 5461 23357
rect 5395 23292 5396 23356
rect 5460 23292 5461 23356
rect 5395 23291 5461 23292
rect 5395 22132 5461 22133
rect 5395 22068 5396 22132
rect 5460 22068 5461 22132
rect 5395 22067 5461 22068
rect 5211 19956 5277 19957
rect 5211 19892 5212 19956
rect 5276 19892 5277 19956
rect 5211 19891 5277 19892
rect 5214 19413 5274 19891
rect 5211 19412 5277 19413
rect 5211 19348 5212 19412
rect 5276 19348 5277 19412
rect 5211 19347 5277 19348
rect 5027 13428 5093 13429
rect 5027 13364 5028 13428
rect 5092 13364 5093 13428
rect 5027 13363 5093 13364
rect 4843 10164 4909 10165
rect 4843 10100 4844 10164
rect 4908 10100 4909 10164
rect 4843 10099 4909 10100
rect 5030 2277 5090 13363
rect 5398 8397 5458 22067
rect 5395 8396 5461 8397
rect 5395 8332 5396 8396
rect 5460 8332 5461 8396
rect 5395 8331 5461 8332
rect 5027 2276 5093 2277
rect 5027 2212 5028 2276
rect 5092 2212 5093 2276
rect 5027 2211 5093 2212
rect 5582 2005 5642 34851
rect 6131 30156 6197 30157
rect 6131 30092 6132 30156
rect 6196 30092 6197 30156
rect 6131 30091 6197 30092
rect 6134 19685 6194 30091
rect 6131 19684 6197 19685
rect 6131 19620 6132 19684
rect 6196 19620 6197 19684
rect 6131 19619 6197 19620
rect 6318 2005 6378 41787
rect 6502 13701 6562 41787
rect 6878 41376 7198 42400
rect 9845 43008 10165 43568
rect 12812 43552 13132 43568
rect 12812 43488 12820 43552
rect 12884 43488 12900 43552
rect 12964 43488 12980 43552
rect 13044 43488 13060 43552
rect 13124 43488 13132 43552
rect 11467 43076 11533 43077
rect 11467 43012 11468 43076
rect 11532 43012 11533 43076
rect 11467 43011 11533 43012
rect 9845 42944 9853 43008
rect 9917 42944 9933 43008
rect 9997 42944 10013 43008
rect 10077 42944 10093 43008
rect 10157 42944 10165 43008
rect 8155 42124 8221 42125
rect 8155 42060 8156 42124
rect 8220 42060 8221 42124
rect 8155 42059 8221 42060
rect 7971 41852 8037 41853
rect 7971 41788 7972 41852
rect 8036 41788 8037 41852
rect 7971 41787 8037 41788
rect 6878 41312 6886 41376
rect 6950 41312 6966 41376
rect 7030 41312 7046 41376
rect 7110 41312 7126 41376
rect 7190 41312 7198 41376
rect 6878 40288 7198 41312
rect 6878 40224 6886 40288
rect 6950 40224 6966 40288
rect 7030 40224 7046 40288
rect 7110 40224 7126 40288
rect 7190 40224 7198 40288
rect 6878 39200 7198 40224
rect 7787 40084 7853 40085
rect 7787 40020 7788 40084
rect 7852 40020 7853 40084
rect 7787 40019 7853 40020
rect 6878 39136 6886 39200
rect 6950 39136 6966 39200
rect 7030 39136 7046 39200
rect 7110 39136 7126 39200
rect 7190 39136 7198 39200
rect 6878 38112 7198 39136
rect 6878 38048 6886 38112
rect 6950 38048 6966 38112
rect 7030 38048 7046 38112
rect 7110 38048 7126 38112
rect 7190 38048 7198 38112
rect 6878 37024 7198 38048
rect 6878 36960 6886 37024
rect 6950 36960 6966 37024
rect 7030 36960 7046 37024
rect 7110 36960 7126 37024
rect 7190 36960 7198 37024
rect 6878 35936 7198 36960
rect 6878 35872 6886 35936
rect 6950 35872 6966 35936
rect 7030 35872 7046 35936
rect 7110 35872 7126 35936
rect 7190 35872 7198 35936
rect 6878 34848 7198 35872
rect 6878 34784 6886 34848
rect 6950 34784 6966 34848
rect 7030 34784 7046 34848
rect 7110 34784 7126 34848
rect 7190 34784 7198 34848
rect 6878 33760 7198 34784
rect 7603 33964 7669 33965
rect 7603 33900 7604 33964
rect 7668 33900 7669 33964
rect 7603 33899 7669 33900
rect 6878 33696 6886 33760
rect 6950 33696 6966 33760
rect 7030 33696 7046 33760
rect 7110 33696 7126 33760
rect 7190 33696 7198 33760
rect 6878 32672 7198 33696
rect 7419 33012 7485 33013
rect 7419 32948 7420 33012
rect 7484 32948 7485 33012
rect 7419 32947 7485 32948
rect 6878 32608 6886 32672
rect 6950 32608 6966 32672
rect 7030 32608 7046 32672
rect 7110 32608 7126 32672
rect 7190 32608 7198 32672
rect 6878 31584 7198 32608
rect 6878 31520 6886 31584
rect 6950 31520 6966 31584
rect 7030 31520 7046 31584
rect 7110 31520 7126 31584
rect 7190 31520 7198 31584
rect 6878 30496 7198 31520
rect 6878 30432 6886 30496
rect 6950 30432 6966 30496
rect 7030 30432 7046 30496
rect 7110 30432 7126 30496
rect 7190 30432 7198 30496
rect 6878 29408 7198 30432
rect 6878 29344 6886 29408
rect 6950 29344 6966 29408
rect 7030 29344 7046 29408
rect 7110 29344 7126 29408
rect 7190 29344 7198 29408
rect 6878 28320 7198 29344
rect 6878 28256 6886 28320
rect 6950 28256 6966 28320
rect 7030 28256 7046 28320
rect 7110 28256 7126 28320
rect 7190 28256 7198 28320
rect 6878 27232 7198 28256
rect 6878 27168 6886 27232
rect 6950 27168 6966 27232
rect 7030 27168 7046 27232
rect 7110 27168 7126 27232
rect 7190 27168 7198 27232
rect 6683 26620 6749 26621
rect 6683 26556 6684 26620
rect 6748 26556 6749 26620
rect 6683 26555 6749 26556
rect 6686 21453 6746 26555
rect 6878 26144 7198 27168
rect 6878 26080 6886 26144
rect 6950 26080 6966 26144
rect 7030 26080 7046 26144
rect 7110 26080 7126 26144
rect 7190 26080 7198 26144
rect 6878 25056 7198 26080
rect 6878 24992 6886 25056
rect 6950 24992 6966 25056
rect 7030 24992 7046 25056
rect 7110 24992 7126 25056
rect 7190 24992 7198 25056
rect 6878 23968 7198 24992
rect 6878 23904 6886 23968
rect 6950 23904 6966 23968
rect 7030 23904 7046 23968
rect 7110 23904 7126 23968
rect 7190 23904 7198 23968
rect 6878 22880 7198 23904
rect 7422 23493 7482 32947
rect 7606 31789 7666 33899
rect 7603 31788 7669 31789
rect 7603 31724 7604 31788
rect 7668 31724 7669 31788
rect 7603 31723 7669 31724
rect 7606 25125 7666 31723
rect 7603 25124 7669 25125
rect 7603 25060 7604 25124
rect 7668 25060 7669 25124
rect 7603 25059 7669 25060
rect 7606 23901 7666 25059
rect 7603 23900 7669 23901
rect 7603 23836 7604 23900
rect 7668 23836 7669 23900
rect 7603 23835 7669 23836
rect 7419 23492 7485 23493
rect 7419 23428 7420 23492
rect 7484 23428 7485 23492
rect 7419 23427 7485 23428
rect 6878 22816 6886 22880
rect 6950 22816 6966 22880
rect 7030 22816 7046 22880
rect 7110 22816 7126 22880
rect 7190 22816 7198 22880
rect 6878 21792 7198 22816
rect 6878 21728 6886 21792
rect 6950 21728 6966 21792
rect 7030 21728 7046 21792
rect 7110 21728 7126 21792
rect 7190 21728 7198 21792
rect 6683 21452 6749 21453
rect 6683 21388 6684 21452
rect 6748 21388 6749 21452
rect 6683 21387 6749 21388
rect 6878 20704 7198 21728
rect 6878 20640 6886 20704
rect 6950 20640 6966 20704
rect 7030 20640 7046 20704
rect 7110 20640 7126 20704
rect 7190 20640 7198 20704
rect 6878 19616 7198 20640
rect 6878 19552 6886 19616
rect 6950 19552 6966 19616
rect 7030 19552 7046 19616
rect 7110 19552 7126 19616
rect 7190 19552 7198 19616
rect 6878 18528 7198 19552
rect 6878 18464 6886 18528
rect 6950 18464 6966 18528
rect 7030 18464 7046 18528
rect 7110 18464 7126 18528
rect 7190 18464 7198 18528
rect 6878 17440 7198 18464
rect 6878 17376 6886 17440
rect 6950 17376 6966 17440
rect 7030 17376 7046 17440
rect 7110 17376 7126 17440
rect 7190 17376 7198 17440
rect 6878 16352 7198 17376
rect 6878 16288 6886 16352
rect 6950 16288 6966 16352
rect 7030 16288 7046 16352
rect 7110 16288 7126 16352
rect 7190 16288 7198 16352
rect 6878 15264 7198 16288
rect 6878 15200 6886 15264
rect 6950 15200 6966 15264
rect 7030 15200 7046 15264
rect 7110 15200 7126 15264
rect 7190 15200 7198 15264
rect 6878 14176 7198 15200
rect 6878 14112 6886 14176
rect 6950 14112 6966 14176
rect 7030 14112 7046 14176
rect 7110 14112 7126 14176
rect 7190 14112 7198 14176
rect 6499 13700 6565 13701
rect 6499 13636 6500 13700
rect 6564 13636 6565 13700
rect 6499 13635 6565 13636
rect 6878 13088 7198 14112
rect 6878 13024 6886 13088
rect 6950 13024 6966 13088
rect 7030 13024 7046 13088
rect 7110 13024 7126 13088
rect 7190 13024 7198 13088
rect 6878 12000 7198 13024
rect 6878 11936 6886 12000
rect 6950 11936 6966 12000
rect 7030 11936 7046 12000
rect 7110 11936 7126 12000
rect 7190 11936 7198 12000
rect 6878 10912 7198 11936
rect 6878 10848 6886 10912
rect 6950 10848 6966 10912
rect 7030 10848 7046 10912
rect 7110 10848 7126 10912
rect 7190 10848 7198 10912
rect 6878 9824 7198 10848
rect 6878 9760 6886 9824
rect 6950 9760 6966 9824
rect 7030 9760 7046 9824
rect 7110 9760 7126 9824
rect 7190 9760 7198 9824
rect 6878 8736 7198 9760
rect 6878 8672 6886 8736
rect 6950 8672 6966 8736
rect 7030 8672 7046 8736
rect 7110 8672 7126 8736
rect 7190 8672 7198 8736
rect 6878 7648 7198 8672
rect 6878 7584 6886 7648
rect 6950 7584 6966 7648
rect 7030 7584 7046 7648
rect 7110 7584 7126 7648
rect 7190 7584 7198 7648
rect 6878 6560 7198 7584
rect 6878 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7198 6560
rect 6878 5472 7198 6496
rect 6878 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7198 5472
rect 6878 4384 7198 5408
rect 6878 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7198 4384
rect 6878 3296 7198 4320
rect 6878 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7198 3296
rect 6878 2208 7198 3232
rect 7790 2277 7850 40019
rect 7974 39405 8034 41787
rect 7971 39404 8037 39405
rect 7971 39340 7972 39404
rect 8036 39340 8037 39404
rect 7971 39339 8037 39340
rect 7971 33420 8037 33421
rect 7971 33356 7972 33420
rect 8036 33356 8037 33420
rect 7971 33355 8037 33356
rect 7974 29885 8034 33355
rect 7971 29884 8037 29885
rect 7971 29820 7972 29884
rect 8036 29820 8037 29884
rect 7971 29819 8037 29820
rect 8158 2277 8218 42059
rect 9845 41920 10165 42944
rect 9845 41856 9853 41920
rect 9917 41856 9933 41920
rect 9997 41856 10013 41920
rect 10077 41856 10093 41920
rect 10157 41856 10165 41920
rect 9259 41444 9325 41445
rect 9259 41380 9260 41444
rect 9324 41380 9325 41444
rect 9259 41379 9325 41380
rect 8891 37772 8957 37773
rect 8891 37708 8892 37772
rect 8956 37708 8957 37772
rect 8891 37707 8957 37708
rect 8523 37364 8589 37365
rect 8523 37300 8524 37364
rect 8588 37300 8589 37364
rect 8523 37299 8589 37300
rect 8526 2277 8586 37299
rect 8707 35596 8773 35597
rect 8707 35532 8708 35596
rect 8772 35532 8773 35596
rect 8707 35531 8773 35532
rect 7787 2276 7853 2277
rect 7787 2212 7788 2276
rect 7852 2212 7853 2276
rect 7787 2211 7853 2212
rect 8155 2276 8221 2277
rect 8155 2212 8156 2276
rect 8220 2212 8221 2276
rect 8155 2211 8221 2212
rect 8523 2276 8589 2277
rect 8523 2212 8524 2276
rect 8588 2212 8589 2276
rect 8523 2211 8589 2212
rect 6878 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7198 2208
rect 5579 2004 5645 2005
rect 5579 1940 5580 2004
rect 5644 1940 5645 2004
rect 5579 1939 5645 1940
rect 6315 2004 6381 2005
rect 6315 1940 6316 2004
rect 6380 1940 6381 2004
rect 6315 1939 6381 1940
rect 4475 1324 4541 1325
rect 4475 1260 4476 1324
rect 4540 1260 4541 1324
rect 4475 1259 4541 1260
rect 6878 1120 7198 2144
rect 6878 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7198 1120
rect 6878 1040 7198 1056
rect 8710 781 8770 35531
rect 8894 2277 8954 37707
rect 9262 28250 9322 41379
rect 9845 40832 10165 41856
rect 9845 40768 9853 40832
rect 9917 40768 9933 40832
rect 9997 40768 10013 40832
rect 10077 40768 10093 40832
rect 10157 40768 10165 40832
rect 9627 40084 9693 40085
rect 9627 40020 9628 40084
rect 9692 40020 9693 40084
rect 9627 40019 9693 40020
rect 9630 28797 9690 40019
rect 9845 39744 10165 40768
rect 10547 39948 10613 39949
rect 10547 39884 10548 39948
rect 10612 39884 10613 39948
rect 10547 39883 10613 39884
rect 9845 39680 9853 39744
rect 9917 39680 9933 39744
rect 9997 39680 10013 39744
rect 10077 39680 10093 39744
rect 10157 39680 10165 39744
rect 9845 38656 10165 39680
rect 9845 38592 9853 38656
rect 9917 38592 9933 38656
rect 9997 38592 10013 38656
rect 10077 38592 10093 38656
rect 10157 38592 10165 38656
rect 9845 37568 10165 38592
rect 9845 37504 9853 37568
rect 9917 37504 9933 37568
rect 9997 37504 10013 37568
rect 10077 37504 10093 37568
rect 10157 37504 10165 37568
rect 9845 36480 10165 37504
rect 9845 36416 9853 36480
rect 9917 36416 9933 36480
rect 9997 36416 10013 36480
rect 10077 36416 10093 36480
rect 10157 36416 10165 36480
rect 9845 35392 10165 36416
rect 10363 36004 10429 36005
rect 10363 35940 10364 36004
rect 10428 35940 10429 36004
rect 10363 35939 10429 35940
rect 9845 35328 9853 35392
rect 9917 35328 9933 35392
rect 9997 35328 10013 35392
rect 10077 35328 10093 35392
rect 10157 35328 10165 35392
rect 9845 34304 10165 35328
rect 9845 34240 9853 34304
rect 9917 34240 9933 34304
rect 9997 34240 10013 34304
rect 10077 34240 10093 34304
rect 10157 34240 10165 34304
rect 9845 33216 10165 34240
rect 9845 33152 9853 33216
rect 9917 33152 9933 33216
rect 9997 33152 10013 33216
rect 10077 33152 10093 33216
rect 10157 33152 10165 33216
rect 9845 32128 10165 33152
rect 9845 32064 9853 32128
rect 9917 32064 9933 32128
rect 9997 32064 10013 32128
rect 10077 32064 10093 32128
rect 10157 32064 10165 32128
rect 9845 31040 10165 32064
rect 9845 30976 9853 31040
rect 9917 30976 9933 31040
rect 9997 30976 10013 31040
rect 10077 30976 10093 31040
rect 10157 30976 10165 31040
rect 9845 29952 10165 30976
rect 10366 30157 10426 35939
rect 10363 30156 10429 30157
rect 10363 30092 10364 30156
rect 10428 30092 10429 30156
rect 10363 30091 10429 30092
rect 10363 30020 10429 30021
rect 10363 29956 10364 30020
rect 10428 29956 10429 30020
rect 10363 29955 10429 29956
rect 9845 29888 9853 29952
rect 9917 29888 9933 29952
rect 9997 29888 10013 29952
rect 10077 29888 10093 29952
rect 10157 29888 10165 29952
rect 9845 28864 10165 29888
rect 9845 28800 9853 28864
rect 9917 28800 9933 28864
rect 9997 28800 10013 28864
rect 10077 28800 10093 28864
rect 10157 28800 10165 28864
rect 9627 28796 9693 28797
rect 9627 28732 9628 28796
rect 9692 28732 9693 28796
rect 9627 28731 9693 28732
rect 9262 28190 9690 28250
rect 9075 24988 9141 24989
rect 9075 24924 9076 24988
rect 9140 24924 9141 24988
rect 9075 24923 9141 24924
rect 9078 21589 9138 24923
rect 9630 22110 9690 28190
rect 9446 22050 9690 22110
rect 9845 27776 10165 28800
rect 9845 27712 9853 27776
rect 9917 27712 9933 27776
rect 9997 27712 10013 27776
rect 10077 27712 10093 27776
rect 10157 27712 10165 27776
rect 9845 26688 10165 27712
rect 9845 26624 9853 26688
rect 9917 26624 9933 26688
rect 9997 26624 10013 26688
rect 10077 26624 10093 26688
rect 10157 26624 10165 26688
rect 9845 25600 10165 26624
rect 9845 25536 9853 25600
rect 9917 25536 9933 25600
rect 9997 25536 10013 25600
rect 10077 25536 10093 25600
rect 10157 25536 10165 25600
rect 9845 24512 10165 25536
rect 10366 24989 10426 29955
rect 10550 27573 10610 39883
rect 10731 27844 10797 27845
rect 10731 27780 10732 27844
rect 10796 27780 10797 27844
rect 10731 27779 10797 27780
rect 10547 27572 10613 27573
rect 10547 27508 10548 27572
rect 10612 27508 10613 27572
rect 10547 27507 10613 27508
rect 10734 26890 10794 27779
rect 10550 26830 10794 26890
rect 10363 24988 10429 24989
rect 10363 24924 10364 24988
rect 10428 24924 10429 24988
rect 10363 24923 10429 24924
rect 9845 24448 9853 24512
rect 9917 24448 9933 24512
rect 9997 24448 10013 24512
rect 10077 24448 10093 24512
rect 10157 24448 10165 24512
rect 9845 23424 10165 24448
rect 9845 23360 9853 23424
rect 9917 23360 9933 23424
rect 9997 23360 10013 23424
rect 10077 23360 10093 23424
rect 10157 23360 10165 23424
rect 9845 22336 10165 23360
rect 10363 22812 10429 22813
rect 10363 22748 10364 22812
rect 10428 22748 10429 22812
rect 10363 22747 10429 22748
rect 9845 22272 9853 22336
rect 9917 22272 9933 22336
rect 9997 22272 10013 22336
rect 10077 22272 10093 22336
rect 10157 22272 10165 22336
rect 9075 21588 9141 21589
rect 9075 21524 9076 21588
rect 9140 21524 9141 21588
rect 9075 21523 9141 21524
rect 9446 2685 9506 22050
rect 9845 21248 10165 22272
rect 9845 21184 9853 21248
rect 9917 21184 9933 21248
rect 9997 21184 10013 21248
rect 10077 21184 10093 21248
rect 10157 21184 10165 21248
rect 9845 20160 10165 21184
rect 9845 20096 9853 20160
rect 9917 20096 9933 20160
rect 9997 20096 10013 20160
rect 10077 20096 10093 20160
rect 10157 20096 10165 20160
rect 9845 19072 10165 20096
rect 10366 19821 10426 22747
rect 10363 19820 10429 19821
rect 10363 19756 10364 19820
rect 10428 19756 10429 19820
rect 10363 19755 10429 19756
rect 9845 19008 9853 19072
rect 9917 19008 9933 19072
rect 9997 19008 10013 19072
rect 10077 19008 10093 19072
rect 10157 19008 10165 19072
rect 9627 18188 9693 18189
rect 9627 18124 9628 18188
rect 9692 18124 9693 18188
rect 9627 18123 9693 18124
rect 9443 2684 9509 2685
rect 9443 2620 9444 2684
rect 9508 2620 9509 2684
rect 9443 2619 9509 2620
rect 9630 2549 9690 18123
rect 9845 17984 10165 19008
rect 10550 18869 10610 26830
rect 10731 26212 10797 26213
rect 10731 26148 10732 26212
rect 10796 26148 10797 26212
rect 10731 26147 10797 26148
rect 10547 18868 10613 18869
rect 10547 18804 10548 18868
rect 10612 18804 10613 18868
rect 10547 18803 10613 18804
rect 9845 17920 9853 17984
rect 9917 17920 9933 17984
rect 9997 17920 10013 17984
rect 10077 17920 10093 17984
rect 10157 17920 10165 17984
rect 9845 16896 10165 17920
rect 9845 16832 9853 16896
rect 9917 16832 9933 16896
rect 9997 16832 10013 16896
rect 10077 16832 10093 16896
rect 10157 16832 10165 16896
rect 9845 15808 10165 16832
rect 9845 15744 9853 15808
rect 9917 15744 9933 15808
rect 9997 15744 10013 15808
rect 10077 15744 10093 15808
rect 10157 15744 10165 15808
rect 9845 14720 10165 15744
rect 9845 14656 9853 14720
rect 9917 14656 9933 14720
rect 9997 14656 10013 14720
rect 10077 14656 10093 14720
rect 10157 14656 10165 14720
rect 9845 13632 10165 14656
rect 9845 13568 9853 13632
rect 9917 13568 9933 13632
rect 9997 13568 10013 13632
rect 10077 13568 10093 13632
rect 10157 13568 10165 13632
rect 9845 12544 10165 13568
rect 10550 12885 10610 18803
rect 10734 16557 10794 26147
rect 10915 24444 10981 24445
rect 10915 24380 10916 24444
rect 10980 24380 10981 24444
rect 10915 24379 10981 24380
rect 10918 19685 10978 24379
rect 10915 19684 10981 19685
rect 10915 19620 10916 19684
rect 10980 19620 10981 19684
rect 10915 19619 10981 19620
rect 11470 17781 11530 43011
rect 11651 42940 11717 42941
rect 11651 42876 11652 42940
rect 11716 42876 11717 42940
rect 11651 42875 11717 42876
rect 12203 42940 12269 42941
rect 12203 42876 12204 42940
rect 12268 42876 12269 42940
rect 12203 42875 12269 42876
rect 11467 17780 11533 17781
rect 11467 17716 11468 17780
rect 11532 17716 11533 17780
rect 11467 17715 11533 17716
rect 11654 17645 11714 42875
rect 12019 30428 12085 30429
rect 12019 30364 12020 30428
rect 12084 30364 12085 30428
rect 12019 30363 12085 30364
rect 11835 22268 11901 22269
rect 11835 22204 11836 22268
rect 11900 22204 11901 22268
rect 11835 22203 11901 22204
rect 11651 17644 11717 17645
rect 11651 17580 11652 17644
rect 11716 17580 11717 17644
rect 11651 17579 11717 17580
rect 10731 16556 10797 16557
rect 10731 16492 10732 16556
rect 10796 16492 10797 16556
rect 10731 16491 10797 16492
rect 10915 16012 10981 16013
rect 10915 15948 10916 16012
rect 10980 15948 10981 16012
rect 10915 15947 10981 15948
rect 10547 12884 10613 12885
rect 10547 12820 10548 12884
rect 10612 12820 10613 12884
rect 10547 12819 10613 12820
rect 9845 12480 9853 12544
rect 9917 12480 9933 12544
rect 9997 12480 10013 12544
rect 10077 12480 10093 12544
rect 10157 12480 10165 12544
rect 9845 11456 10165 12480
rect 9845 11392 9853 11456
rect 9917 11392 9933 11456
rect 9997 11392 10013 11456
rect 10077 11392 10093 11456
rect 10157 11392 10165 11456
rect 9845 10368 10165 11392
rect 9845 10304 9853 10368
rect 9917 10304 9933 10368
rect 9997 10304 10013 10368
rect 10077 10304 10093 10368
rect 10157 10304 10165 10368
rect 9845 9280 10165 10304
rect 9845 9216 9853 9280
rect 9917 9216 9933 9280
rect 9997 9216 10013 9280
rect 10077 9216 10093 9280
rect 10157 9216 10165 9280
rect 9845 8192 10165 9216
rect 9845 8128 9853 8192
rect 9917 8128 9933 8192
rect 9997 8128 10013 8192
rect 10077 8128 10093 8192
rect 10157 8128 10165 8192
rect 9845 7104 10165 8128
rect 9845 7040 9853 7104
rect 9917 7040 9933 7104
rect 9997 7040 10013 7104
rect 10077 7040 10093 7104
rect 10157 7040 10165 7104
rect 9845 6016 10165 7040
rect 9845 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10165 6016
rect 9845 4928 10165 5952
rect 9845 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10165 4928
rect 9845 3840 10165 4864
rect 9845 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10165 3840
rect 9845 2752 10165 3776
rect 10918 3501 10978 15947
rect 11838 5269 11898 22203
rect 11835 5268 11901 5269
rect 11835 5204 11836 5268
rect 11900 5204 11901 5268
rect 11835 5203 11901 5204
rect 10915 3500 10981 3501
rect 10915 3436 10916 3500
rect 10980 3436 10981 3500
rect 10915 3435 10981 3436
rect 9845 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10165 2752
rect 9627 2548 9693 2549
rect 9627 2484 9628 2548
rect 9692 2484 9693 2548
rect 9627 2483 9693 2484
rect 8891 2276 8957 2277
rect 8891 2212 8892 2276
rect 8956 2212 8957 2276
rect 8891 2211 8957 2212
rect 9845 1664 10165 2688
rect 12022 2685 12082 30363
rect 12206 23493 12266 42875
rect 12812 42464 13132 43488
rect 13675 43076 13741 43077
rect 13675 43012 13676 43076
rect 13740 43012 13741 43076
rect 13675 43011 13741 43012
rect 13307 42940 13373 42941
rect 13307 42876 13308 42940
rect 13372 42876 13373 42940
rect 13307 42875 13373 42876
rect 12812 42400 12820 42464
rect 12884 42400 12900 42464
rect 12964 42400 12980 42464
rect 13044 42400 13060 42464
rect 13124 42400 13132 42464
rect 12812 41376 13132 42400
rect 12812 41312 12820 41376
rect 12884 41312 12900 41376
rect 12964 41312 12980 41376
rect 13044 41312 13060 41376
rect 13124 41312 13132 41376
rect 12812 40288 13132 41312
rect 12812 40224 12820 40288
rect 12884 40224 12900 40288
rect 12964 40224 12980 40288
rect 13044 40224 13060 40288
rect 13124 40224 13132 40288
rect 12812 39200 13132 40224
rect 12812 39136 12820 39200
rect 12884 39136 12900 39200
rect 12964 39136 12980 39200
rect 13044 39136 13060 39200
rect 13124 39136 13132 39200
rect 12571 38452 12637 38453
rect 12571 38388 12572 38452
rect 12636 38388 12637 38452
rect 12571 38387 12637 38388
rect 12387 32060 12453 32061
rect 12387 31996 12388 32060
rect 12452 31996 12453 32060
rect 12387 31995 12453 31996
rect 12390 31653 12450 31995
rect 12387 31652 12453 31653
rect 12387 31588 12388 31652
rect 12452 31588 12453 31652
rect 12387 31587 12453 31588
rect 12203 23492 12269 23493
rect 12203 23428 12204 23492
rect 12268 23428 12269 23492
rect 12203 23427 12269 23428
rect 12387 22268 12453 22269
rect 12387 22204 12388 22268
rect 12452 22204 12453 22268
rect 12387 22203 12453 22204
rect 12390 22130 12450 22203
rect 12206 22070 12450 22130
rect 12206 21317 12266 22070
rect 12203 21316 12269 21317
rect 12203 21252 12204 21316
rect 12268 21252 12269 21316
rect 12203 21251 12269 21252
rect 12574 20909 12634 38387
rect 12812 38112 13132 39136
rect 12812 38048 12820 38112
rect 12884 38048 12900 38112
rect 12964 38048 12980 38112
rect 13044 38048 13060 38112
rect 13124 38048 13132 38112
rect 12812 37024 13132 38048
rect 12812 36960 12820 37024
rect 12884 36960 12900 37024
rect 12964 36960 12980 37024
rect 13044 36960 13060 37024
rect 13124 36960 13132 37024
rect 12812 35936 13132 36960
rect 12812 35872 12820 35936
rect 12884 35872 12900 35936
rect 12964 35872 12980 35936
rect 13044 35872 13060 35936
rect 13124 35872 13132 35936
rect 12812 34848 13132 35872
rect 12812 34784 12820 34848
rect 12884 34784 12900 34848
rect 12964 34784 12980 34848
rect 13044 34784 13060 34848
rect 13124 34784 13132 34848
rect 12812 33760 13132 34784
rect 12812 33696 12820 33760
rect 12884 33696 12900 33760
rect 12964 33696 12980 33760
rect 13044 33696 13060 33760
rect 13124 33696 13132 33760
rect 12812 32672 13132 33696
rect 12812 32608 12820 32672
rect 12884 32608 12900 32672
rect 12964 32608 12980 32672
rect 13044 32608 13060 32672
rect 13124 32608 13132 32672
rect 12812 31584 13132 32608
rect 12812 31520 12820 31584
rect 12884 31520 12900 31584
rect 12964 31520 12980 31584
rect 13044 31520 13060 31584
rect 13124 31520 13132 31584
rect 12812 30496 13132 31520
rect 12812 30432 12820 30496
rect 12884 30432 12900 30496
rect 12964 30432 12980 30496
rect 13044 30432 13060 30496
rect 13124 30432 13132 30496
rect 12812 29408 13132 30432
rect 12812 29344 12820 29408
rect 12884 29344 12900 29408
rect 12964 29344 12980 29408
rect 13044 29344 13060 29408
rect 13124 29344 13132 29408
rect 12812 28320 13132 29344
rect 12812 28256 12820 28320
rect 12884 28256 12900 28320
rect 12964 28256 12980 28320
rect 13044 28256 13060 28320
rect 13124 28256 13132 28320
rect 12812 27232 13132 28256
rect 12812 27168 12820 27232
rect 12884 27168 12900 27232
rect 12964 27168 12980 27232
rect 13044 27168 13060 27232
rect 13124 27168 13132 27232
rect 12812 26144 13132 27168
rect 12812 26080 12820 26144
rect 12884 26080 12900 26144
rect 12964 26080 12980 26144
rect 13044 26080 13060 26144
rect 13124 26080 13132 26144
rect 12812 25056 13132 26080
rect 12812 24992 12820 25056
rect 12884 24992 12900 25056
rect 12964 24992 12980 25056
rect 13044 24992 13060 25056
rect 13124 24992 13132 25056
rect 12812 23968 13132 24992
rect 12812 23904 12820 23968
rect 12884 23904 12900 23968
rect 12964 23904 12980 23968
rect 13044 23904 13060 23968
rect 13124 23904 13132 23968
rect 12812 22880 13132 23904
rect 12812 22816 12820 22880
rect 12884 22816 12900 22880
rect 12964 22816 12980 22880
rect 13044 22816 13060 22880
rect 13124 22816 13132 22880
rect 12812 21792 13132 22816
rect 12812 21728 12820 21792
rect 12884 21728 12900 21792
rect 12964 21728 12980 21792
rect 13044 21728 13060 21792
rect 13124 21728 13132 21792
rect 12571 20908 12637 20909
rect 12571 20844 12572 20908
rect 12636 20844 12637 20908
rect 12571 20843 12637 20844
rect 12812 20704 13132 21728
rect 12812 20640 12820 20704
rect 12884 20640 12900 20704
rect 12964 20640 12980 20704
rect 13044 20640 13060 20704
rect 13124 20640 13132 20704
rect 12812 19616 13132 20640
rect 12812 19552 12820 19616
rect 12884 19552 12900 19616
rect 12964 19552 12980 19616
rect 13044 19552 13060 19616
rect 13124 19552 13132 19616
rect 12812 18528 13132 19552
rect 12812 18464 12820 18528
rect 12884 18464 12900 18528
rect 12964 18464 12980 18528
rect 13044 18464 13060 18528
rect 13124 18464 13132 18528
rect 12812 17440 13132 18464
rect 12812 17376 12820 17440
rect 12884 17376 12900 17440
rect 12964 17376 12980 17440
rect 13044 17376 13060 17440
rect 13124 17376 13132 17440
rect 12812 16352 13132 17376
rect 12812 16288 12820 16352
rect 12884 16288 12900 16352
rect 12964 16288 12980 16352
rect 13044 16288 13060 16352
rect 13124 16288 13132 16352
rect 12812 15264 13132 16288
rect 12812 15200 12820 15264
rect 12884 15200 12900 15264
rect 12964 15200 12980 15264
rect 13044 15200 13060 15264
rect 13124 15200 13132 15264
rect 12812 14176 13132 15200
rect 12812 14112 12820 14176
rect 12884 14112 12900 14176
rect 12964 14112 12980 14176
rect 13044 14112 13060 14176
rect 13124 14112 13132 14176
rect 12203 13700 12269 13701
rect 12203 13636 12204 13700
rect 12268 13636 12269 13700
rect 12203 13635 12269 13636
rect 12206 4045 12266 13635
rect 12812 13088 13132 14112
rect 12812 13024 12820 13088
rect 12884 13024 12900 13088
rect 12964 13024 12980 13088
rect 13044 13024 13060 13088
rect 13124 13024 13132 13088
rect 12812 12000 13132 13024
rect 12812 11936 12820 12000
rect 12884 11936 12900 12000
rect 12964 11936 12980 12000
rect 13044 11936 13060 12000
rect 13124 11936 13132 12000
rect 12812 10912 13132 11936
rect 12812 10848 12820 10912
rect 12884 10848 12900 10912
rect 12964 10848 12980 10912
rect 13044 10848 13060 10912
rect 13124 10848 13132 10912
rect 12812 9824 13132 10848
rect 12812 9760 12820 9824
rect 12884 9760 12900 9824
rect 12964 9760 12980 9824
rect 13044 9760 13060 9824
rect 13124 9760 13132 9824
rect 12812 8736 13132 9760
rect 12812 8672 12820 8736
rect 12884 8672 12900 8736
rect 12964 8672 12980 8736
rect 13044 8672 13060 8736
rect 13124 8672 13132 8736
rect 12812 7648 13132 8672
rect 12812 7584 12820 7648
rect 12884 7584 12900 7648
rect 12964 7584 12980 7648
rect 13044 7584 13060 7648
rect 13124 7584 13132 7648
rect 12812 6560 13132 7584
rect 12812 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13132 6560
rect 12812 5472 13132 6496
rect 12812 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13132 5472
rect 12812 4384 13132 5408
rect 13310 5405 13370 42875
rect 13491 41036 13557 41037
rect 13491 40972 13492 41036
rect 13556 40972 13557 41036
rect 13491 40971 13557 40972
rect 13494 32061 13554 40971
rect 13678 38997 13738 43011
rect 15779 43008 16099 43568
rect 15779 42944 15787 43008
rect 15851 42944 15867 43008
rect 15931 42944 15947 43008
rect 16011 42944 16027 43008
rect 16091 42944 16099 43008
rect 14411 42940 14477 42941
rect 14411 42876 14412 42940
rect 14476 42876 14477 42940
rect 14411 42875 14477 42876
rect 14963 42940 15029 42941
rect 14963 42876 14964 42940
rect 15028 42876 15029 42940
rect 14963 42875 15029 42876
rect 15331 42940 15397 42941
rect 15331 42876 15332 42940
rect 15396 42876 15397 42940
rect 15331 42875 15397 42876
rect 13675 38996 13741 38997
rect 13675 38932 13676 38996
rect 13740 38932 13741 38996
rect 13675 38931 13741 38932
rect 13491 32060 13557 32061
rect 13491 31996 13492 32060
rect 13556 31996 13557 32060
rect 13491 31995 13557 31996
rect 13491 31380 13557 31381
rect 13491 31316 13492 31380
rect 13556 31316 13557 31380
rect 13491 31315 13557 31316
rect 13494 22269 13554 31315
rect 14043 30564 14109 30565
rect 14043 30500 14044 30564
rect 14108 30500 14109 30564
rect 14043 30499 14109 30500
rect 13675 26484 13741 26485
rect 13675 26420 13676 26484
rect 13740 26420 13741 26484
rect 13675 26419 13741 26420
rect 13491 22268 13557 22269
rect 13491 22204 13492 22268
rect 13556 22204 13557 22268
rect 13491 22203 13557 22204
rect 13491 21996 13557 21997
rect 13491 21932 13492 21996
rect 13556 21932 13557 21996
rect 13491 21931 13557 21932
rect 13494 17781 13554 21931
rect 13678 19549 13738 26419
rect 14046 23493 14106 30499
rect 14414 30429 14474 42875
rect 14595 41716 14661 41717
rect 14595 41652 14596 41716
rect 14660 41652 14661 41716
rect 14595 41651 14661 41652
rect 14598 33965 14658 41651
rect 14779 41580 14845 41581
rect 14779 41516 14780 41580
rect 14844 41516 14845 41580
rect 14779 41515 14845 41516
rect 14595 33964 14661 33965
rect 14595 33900 14596 33964
rect 14660 33900 14661 33964
rect 14595 33899 14661 33900
rect 14411 30428 14477 30429
rect 14411 30364 14412 30428
rect 14476 30364 14477 30428
rect 14411 30363 14477 30364
rect 14782 29069 14842 41515
rect 14779 29068 14845 29069
rect 14779 29004 14780 29068
rect 14844 29004 14845 29068
rect 14779 29003 14845 29004
rect 14779 25396 14845 25397
rect 14779 25332 14780 25396
rect 14844 25332 14845 25396
rect 14779 25331 14845 25332
rect 14043 23492 14109 23493
rect 14043 23428 14044 23492
rect 14108 23428 14109 23492
rect 14043 23427 14109 23428
rect 14595 21316 14661 21317
rect 14595 21252 14596 21316
rect 14660 21252 14661 21316
rect 14595 21251 14661 21252
rect 13675 19548 13741 19549
rect 13675 19484 13676 19548
rect 13740 19484 13741 19548
rect 13675 19483 13741 19484
rect 13859 19412 13925 19413
rect 13859 19348 13860 19412
rect 13924 19348 13925 19412
rect 13859 19347 13925 19348
rect 13491 17780 13557 17781
rect 13491 17716 13492 17780
rect 13556 17716 13557 17780
rect 13491 17715 13557 17716
rect 13491 17644 13557 17645
rect 13491 17580 13492 17644
rect 13556 17580 13557 17644
rect 13491 17579 13557 17580
rect 13307 5404 13373 5405
rect 13307 5340 13308 5404
rect 13372 5340 13373 5404
rect 13307 5339 13373 5340
rect 12812 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13132 4384
rect 12203 4044 12269 4045
rect 12203 3980 12204 4044
rect 12268 3980 12269 4044
rect 12203 3979 12269 3980
rect 12812 3296 13132 4320
rect 12812 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13132 3296
rect 12019 2684 12085 2685
rect 12019 2620 12020 2684
rect 12084 2620 12085 2684
rect 12019 2619 12085 2620
rect 9845 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10165 1664
rect 9845 1040 10165 1600
rect 12812 2208 13132 3232
rect 13494 2549 13554 17579
rect 13862 16557 13922 19347
rect 13859 16556 13925 16557
rect 13859 16492 13860 16556
rect 13924 16492 13925 16556
rect 13859 16491 13925 16492
rect 14598 13973 14658 21251
rect 14595 13972 14661 13973
rect 14595 13908 14596 13972
rect 14660 13908 14661 13972
rect 14595 13907 14661 13908
rect 13859 13700 13925 13701
rect 13859 13636 13860 13700
rect 13924 13636 13925 13700
rect 13859 13635 13925 13636
rect 13862 4181 13922 13635
rect 14598 5269 14658 13907
rect 14595 5268 14661 5269
rect 14595 5204 14596 5268
rect 14660 5204 14661 5268
rect 14595 5203 14661 5204
rect 13859 4180 13925 4181
rect 13859 4116 13860 4180
rect 13924 4116 13925 4180
rect 13859 4115 13925 4116
rect 14782 2685 14842 25331
rect 14966 10437 15026 42875
rect 15334 26213 15394 42875
rect 15779 41920 16099 42944
rect 15779 41856 15787 41920
rect 15851 41856 15867 41920
rect 15931 41856 15947 41920
rect 16011 41856 16027 41920
rect 16091 41856 16099 41920
rect 15779 40832 16099 41856
rect 18746 43552 19066 43568
rect 18746 43488 18754 43552
rect 18818 43488 18834 43552
rect 18898 43488 18914 43552
rect 18978 43488 18994 43552
rect 19058 43488 19066 43552
rect 18746 42464 19066 43488
rect 20667 43212 20733 43213
rect 20667 43148 20668 43212
rect 20732 43148 20733 43212
rect 20667 43147 20733 43148
rect 18746 42400 18754 42464
rect 18818 42400 18834 42464
rect 18898 42400 18914 42464
rect 18978 42400 18994 42464
rect 19058 42400 19066 42464
rect 17723 41852 17789 41853
rect 17723 41788 17724 41852
rect 17788 41788 17789 41852
rect 17723 41787 17789 41788
rect 18275 41852 18341 41853
rect 18275 41788 18276 41852
rect 18340 41788 18341 41852
rect 18275 41787 18341 41788
rect 17539 41716 17605 41717
rect 17539 41652 17540 41716
rect 17604 41652 17605 41716
rect 17539 41651 17605 41652
rect 16251 41444 16317 41445
rect 16251 41380 16252 41444
rect 16316 41380 16317 41444
rect 16251 41379 16317 41380
rect 15779 40768 15787 40832
rect 15851 40768 15867 40832
rect 15931 40768 15947 40832
rect 16011 40768 16027 40832
rect 16091 40768 16099 40832
rect 15779 39744 16099 40768
rect 15779 39680 15787 39744
rect 15851 39680 15867 39744
rect 15931 39680 15947 39744
rect 16011 39680 16027 39744
rect 16091 39680 16099 39744
rect 15779 38656 16099 39680
rect 15779 38592 15787 38656
rect 15851 38592 15867 38656
rect 15931 38592 15947 38656
rect 16011 38592 16027 38656
rect 16091 38592 16099 38656
rect 15779 37568 16099 38592
rect 15779 37504 15787 37568
rect 15851 37504 15867 37568
rect 15931 37504 15947 37568
rect 16011 37504 16027 37568
rect 16091 37504 16099 37568
rect 15779 36480 16099 37504
rect 15779 36416 15787 36480
rect 15851 36416 15867 36480
rect 15931 36416 15947 36480
rect 16011 36416 16027 36480
rect 16091 36416 16099 36480
rect 15779 35392 16099 36416
rect 15779 35328 15787 35392
rect 15851 35328 15867 35392
rect 15931 35328 15947 35392
rect 16011 35328 16027 35392
rect 16091 35328 16099 35392
rect 15779 34304 16099 35328
rect 15779 34240 15787 34304
rect 15851 34240 15867 34304
rect 15931 34240 15947 34304
rect 16011 34240 16027 34304
rect 16091 34240 16099 34304
rect 15779 33216 16099 34240
rect 15779 33152 15787 33216
rect 15851 33152 15867 33216
rect 15931 33152 15947 33216
rect 16011 33152 16027 33216
rect 16091 33152 16099 33216
rect 15779 32128 16099 33152
rect 15779 32064 15787 32128
rect 15851 32064 15867 32128
rect 15931 32064 15947 32128
rect 16011 32064 16027 32128
rect 16091 32064 16099 32128
rect 15515 32060 15581 32061
rect 15515 31996 15516 32060
rect 15580 31996 15581 32060
rect 15515 31995 15581 31996
rect 15331 26212 15397 26213
rect 15331 26148 15332 26212
rect 15396 26148 15397 26212
rect 15331 26147 15397 26148
rect 14963 10436 15029 10437
rect 14963 10372 14964 10436
rect 15028 10372 15029 10436
rect 14963 10371 15029 10372
rect 15518 2685 15578 31995
rect 15779 31040 16099 32064
rect 15779 30976 15787 31040
rect 15851 30976 15867 31040
rect 15931 30976 15947 31040
rect 16011 30976 16027 31040
rect 16091 30976 16099 31040
rect 15779 29952 16099 30976
rect 15779 29888 15787 29952
rect 15851 29888 15867 29952
rect 15931 29888 15947 29952
rect 16011 29888 16027 29952
rect 16091 29888 16099 29952
rect 15779 28864 16099 29888
rect 15779 28800 15787 28864
rect 15851 28800 15867 28864
rect 15931 28800 15947 28864
rect 16011 28800 16027 28864
rect 16091 28800 16099 28864
rect 15779 27776 16099 28800
rect 15779 27712 15787 27776
rect 15851 27712 15867 27776
rect 15931 27712 15947 27776
rect 16011 27712 16027 27776
rect 16091 27712 16099 27776
rect 15779 26688 16099 27712
rect 15779 26624 15787 26688
rect 15851 26624 15867 26688
rect 15931 26624 15947 26688
rect 16011 26624 16027 26688
rect 16091 26624 16099 26688
rect 15779 25600 16099 26624
rect 15779 25536 15787 25600
rect 15851 25536 15867 25600
rect 15931 25536 15947 25600
rect 16011 25536 16027 25600
rect 16091 25536 16099 25600
rect 15779 24512 16099 25536
rect 15779 24448 15787 24512
rect 15851 24448 15867 24512
rect 15931 24448 15947 24512
rect 16011 24448 16027 24512
rect 16091 24448 16099 24512
rect 15779 23424 16099 24448
rect 15779 23360 15787 23424
rect 15851 23360 15867 23424
rect 15931 23360 15947 23424
rect 16011 23360 16027 23424
rect 16091 23360 16099 23424
rect 15779 22336 16099 23360
rect 15779 22272 15787 22336
rect 15851 22272 15867 22336
rect 15931 22272 15947 22336
rect 16011 22272 16027 22336
rect 16091 22272 16099 22336
rect 15779 21248 16099 22272
rect 15779 21184 15787 21248
rect 15851 21184 15867 21248
rect 15931 21184 15947 21248
rect 16011 21184 16027 21248
rect 16091 21184 16099 21248
rect 15779 20160 16099 21184
rect 15779 20096 15787 20160
rect 15851 20096 15867 20160
rect 15931 20096 15947 20160
rect 16011 20096 16027 20160
rect 16091 20096 16099 20160
rect 15779 19072 16099 20096
rect 15779 19008 15787 19072
rect 15851 19008 15867 19072
rect 15931 19008 15947 19072
rect 16011 19008 16027 19072
rect 16091 19008 16099 19072
rect 15779 17984 16099 19008
rect 15779 17920 15787 17984
rect 15851 17920 15867 17984
rect 15931 17920 15947 17984
rect 16011 17920 16027 17984
rect 16091 17920 16099 17984
rect 15779 16896 16099 17920
rect 15779 16832 15787 16896
rect 15851 16832 15867 16896
rect 15931 16832 15947 16896
rect 16011 16832 16027 16896
rect 16091 16832 16099 16896
rect 15779 15808 16099 16832
rect 15779 15744 15787 15808
rect 15851 15744 15867 15808
rect 15931 15744 15947 15808
rect 16011 15744 16027 15808
rect 16091 15744 16099 15808
rect 15779 14720 16099 15744
rect 15779 14656 15787 14720
rect 15851 14656 15867 14720
rect 15931 14656 15947 14720
rect 16011 14656 16027 14720
rect 16091 14656 16099 14720
rect 15779 13632 16099 14656
rect 15779 13568 15787 13632
rect 15851 13568 15867 13632
rect 15931 13568 15947 13632
rect 16011 13568 16027 13632
rect 16091 13568 16099 13632
rect 15779 12544 16099 13568
rect 15779 12480 15787 12544
rect 15851 12480 15867 12544
rect 15931 12480 15947 12544
rect 16011 12480 16027 12544
rect 16091 12480 16099 12544
rect 15779 11456 16099 12480
rect 15779 11392 15787 11456
rect 15851 11392 15867 11456
rect 15931 11392 15947 11456
rect 16011 11392 16027 11456
rect 16091 11392 16099 11456
rect 15779 10368 16099 11392
rect 15779 10304 15787 10368
rect 15851 10304 15867 10368
rect 15931 10304 15947 10368
rect 16011 10304 16027 10368
rect 16091 10304 16099 10368
rect 15779 9280 16099 10304
rect 15779 9216 15787 9280
rect 15851 9216 15867 9280
rect 15931 9216 15947 9280
rect 16011 9216 16027 9280
rect 16091 9216 16099 9280
rect 15779 8192 16099 9216
rect 15779 8128 15787 8192
rect 15851 8128 15867 8192
rect 15931 8128 15947 8192
rect 16011 8128 16027 8192
rect 16091 8128 16099 8192
rect 15779 7104 16099 8128
rect 15779 7040 15787 7104
rect 15851 7040 15867 7104
rect 15931 7040 15947 7104
rect 16011 7040 16027 7104
rect 16091 7040 16099 7104
rect 15779 6016 16099 7040
rect 15779 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16099 6016
rect 15779 4928 16099 5952
rect 15779 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16099 4928
rect 15779 3840 16099 4864
rect 15779 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16099 3840
rect 15779 2752 16099 3776
rect 15779 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16099 2752
rect 14779 2684 14845 2685
rect 14779 2620 14780 2684
rect 14844 2620 14845 2684
rect 14779 2619 14845 2620
rect 15515 2684 15581 2685
rect 15515 2620 15516 2684
rect 15580 2620 15581 2684
rect 15515 2619 15581 2620
rect 13491 2548 13557 2549
rect 13491 2484 13492 2548
rect 13556 2484 13557 2548
rect 13491 2483 13557 2484
rect 12812 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13132 2208
rect 12812 1120 13132 2144
rect 12812 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13132 1120
rect 12812 1040 13132 1056
rect 15779 1664 16099 2688
rect 16254 2549 16314 41379
rect 16619 37908 16685 37909
rect 16619 37844 16620 37908
rect 16684 37844 16685 37908
rect 16619 37843 16685 37844
rect 16435 26212 16501 26213
rect 16435 26148 16436 26212
rect 16500 26148 16501 26212
rect 16435 26147 16501 26148
rect 16438 20501 16498 26147
rect 16622 23493 16682 37843
rect 17355 26892 17421 26893
rect 17355 26828 17356 26892
rect 17420 26828 17421 26892
rect 17355 26827 17421 26828
rect 16619 23492 16685 23493
rect 16619 23428 16620 23492
rect 16684 23428 16685 23492
rect 16619 23427 16685 23428
rect 16987 23492 17053 23493
rect 16987 23428 16988 23492
rect 17052 23428 17053 23492
rect 16987 23427 17053 23428
rect 16619 20908 16685 20909
rect 16619 20844 16620 20908
rect 16684 20844 16685 20908
rect 16619 20843 16685 20844
rect 16435 20500 16501 20501
rect 16435 20436 16436 20500
rect 16500 20436 16501 20500
rect 16435 20435 16501 20436
rect 16435 18188 16501 18189
rect 16435 18124 16436 18188
rect 16500 18124 16501 18188
rect 16435 18123 16501 18124
rect 16251 2548 16317 2549
rect 16251 2484 16252 2548
rect 16316 2484 16317 2548
rect 16251 2483 16317 2484
rect 15779 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16099 1664
rect 15779 1040 16099 1600
rect 16438 1325 16498 18123
rect 16622 11253 16682 20843
rect 16619 11252 16685 11253
rect 16619 11188 16620 11252
rect 16684 11188 16685 11252
rect 16619 11187 16685 11188
rect 16990 2549 17050 23427
rect 17358 20501 17418 26827
rect 17355 20500 17421 20501
rect 17355 20436 17356 20500
rect 17420 20436 17421 20500
rect 17355 20435 17421 20436
rect 17355 9756 17421 9757
rect 17355 9692 17356 9756
rect 17420 9692 17421 9756
rect 17355 9691 17421 9692
rect 17358 8669 17418 9691
rect 17355 8668 17421 8669
rect 17355 8604 17356 8668
rect 17420 8604 17421 8668
rect 17355 8603 17421 8604
rect 17542 2685 17602 41651
rect 17726 4045 17786 41787
rect 18091 22132 18157 22133
rect 18091 22068 18092 22132
rect 18156 22068 18157 22132
rect 18091 22067 18157 22068
rect 17907 14924 17973 14925
rect 17907 14860 17908 14924
rect 17972 14860 17973 14924
rect 17907 14859 17973 14860
rect 17723 4044 17789 4045
rect 17723 3980 17724 4044
rect 17788 3980 17789 4044
rect 17723 3979 17789 3980
rect 17539 2684 17605 2685
rect 17539 2620 17540 2684
rect 17604 2620 17605 2684
rect 17539 2619 17605 2620
rect 16987 2548 17053 2549
rect 16987 2484 16988 2548
rect 17052 2484 17053 2548
rect 16987 2483 17053 2484
rect 16435 1324 16501 1325
rect 16435 1260 16436 1324
rect 16500 1260 16501 1324
rect 16435 1259 16501 1260
rect 17910 917 17970 14859
rect 18094 1325 18154 22067
rect 18278 15197 18338 41787
rect 18746 41376 19066 42400
rect 19195 41580 19261 41581
rect 19195 41516 19196 41580
rect 19260 41516 19261 41580
rect 19195 41515 19261 41516
rect 18746 41312 18754 41376
rect 18818 41312 18834 41376
rect 18898 41312 18914 41376
rect 18978 41312 18994 41376
rect 19058 41312 19066 41376
rect 18746 40288 19066 41312
rect 18746 40224 18754 40288
rect 18818 40224 18834 40288
rect 18898 40224 18914 40288
rect 18978 40224 18994 40288
rect 19058 40224 19066 40288
rect 18746 39200 19066 40224
rect 18746 39136 18754 39200
rect 18818 39136 18834 39200
rect 18898 39136 18914 39200
rect 18978 39136 18994 39200
rect 19058 39136 19066 39200
rect 18746 38112 19066 39136
rect 19198 38725 19258 41515
rect 20670 40629 20730 43147
rect 21713 43008 22033 43568
rect 21713 42944 21721 43008
rect 21785 42944 21801 43008
rect 21865 42944 21881 43008
rect 21945 42944 21961 43008
rect 22025 42944 22033 43008
rect 21035 42124 21101 42125
rect 21035 42060 21036 42124
rect 21100 42060 21101 42124
rect 21035 42059 21101 42060
rect 20667 40628 20733 40629
rect 20667 40564 20668 40628
rect 20732 40564 20733 40628
rect 20667 40563 20733 40564
rect 19563 40084 19629 40085
rect 19563 40020 19564 40084
rect 19628 40020 19629 40084
rect 19563 40019 19629 40020
rect 19195 38724 19261 38725
rect 19195 38660 19196 38724
rect 19260 38660 19261 38724
rect 19195 38659 19261 38660
rect 18746 38048 18754 38112
rect 18818 38048 18834 38112
rect 18898 38048 18914 38112
rect 18978 38048 18994 38112
rect 19058 38048 19066 38112
rect 18746 37024 19066 38048
rect 18746 36960 18754 37024
rect 18818 36960 18834 37024
rect 18898 36960 18914 37024
rect 18978 36960 18994 37024
rect 19058 36960 19066 37024
rect 18746 35936 19066 36960
rect 18746 35872 18754 35936
rect 18818 35872 18834 35936
rect 18898 35872 18914 35936
rect 18978 35872 18994 35936
rect 19058 35872 19066 35936
rect 18746 34848 19066 35872
rect 18746 34784 18754 34848
rect 18818 34784 18834 34848
rect 18898 34784 18914 34848
rect 18978 34784 18994 34848
rect 19058 34784 19066 34848
rect 18746 33760 19066 34784
rect 18746 33696 18754 33760
rect 18818 33696 18834 33760
rect 18898 33696 18914 33760
rect 18978 33696 18994 33760
rect 19058 33696 19066 33760
rect 18746 32672 19066 33696
rect 18746 32608 18754 32672
rect 18818 32608 18834 32672
rect 18898 32608 18914 32672
rect 18978 32608 18994 32672
rect 19058 32608 19066 32672
rect 18746 31584 19066 32608
rect 19379 32332 19445 32333
rect 19379 32268 19380 32332
rect 19444 32268 19445 32332
rect 19379 32267 19445 32268
rect 18746 31520 18754 31584
rect 18818 31520 18834 31584
rect 18898 31520 18914 31584
rect 18978 31520 18994 31584
rect 19058 31520 19066 31584
rect 18746 30496 19066 31520
rect 18746 30432 18754 30496
rect 18818 30432 18834 30496
rect 18898 30432 18914 30496
rect 18978 30432 18994 30496
rect 19058 30432 19066 30496
rect 18746 29408 19066 30432
rect 18746 29344 18754 29408
rect 18818 29344 18834 29408
rect 18898 29344 18914 29408
rect 18978 29344 18994 29408
rect 19058 29344 19066 29408
rect 18459 29068 18525 29069
rect 18459 29004 18460 29068
rect 18524 29004 18525 29068
rect 18459 29003 18525 29004
rect 18275 15196 18341 15197
rect 18275 15132 18276 15196
rect 18340 15132 18341 15196
rect 18275 15131 18341 15132
rect 18462 2685 18522 29003
rect 18746 28320 19066 29344
rect 19195 28660 19261 28661
rect 19195 28596 19196 28660
rect 19260 28596 19261 28660
rect 19195 28595 19261 28596
rect 18746 28256 18754 28320
rect 18818 28256 18834 28320
rect 18898 28256 18914 28320
rect 18978 28256 18994 28320
rect 19058 28256 19066 28320
rect 18746 27232 19066 28256
rect 18746 27168 18754 27232
rect 18818 27168 18834 27232
rect 18898 27168 18914 27232
rect 18978 27168 18994 27232
rect 19058 27168 19066 27232
rect 18746 26144 19066 27168
rect 19198 26213 19258 28595
rect 19195 26212 19261 26213
rect 19195 26148 19196 26212
rect 19260 26148 19261 26212
rect 19195 26147 19261 26148
rect 18746 26080 18754 26144
rect 18818 26080 18834 26144
rect 18898 26080 18914 26144
rect 18978 26080 18994 26144
rect 19058 26080 19066 26144
rect 18746 25056 19066 26080
rect 18746 24992 18754 25056
rect 18818 24992 18834 25056
rect 18898 24992 18914 25056
rect 18978 24992 18994 25056
rect 19058 24992 19066 25056
rect 18746 23968 19066 24992
rect 18746 23904 18754 23968
rect 18818 23904 18834 23968
rect 18898 23904 18914 23968
rect 18978 23904 18994 23968
rect 19058 23904 19066 23968
rect 18746 22880 19066 23904
rect 18746 22816 18754 22880
rect 18818 22816 18834 22880
rect 18898 22816 18914 22880
rect 18978 22816 18994 22880
rect 19058 22816 19066 22880
rect 18746 21792 19066 22816
rect 18746 21728 18754 21792
rect 18818 21728 18834 21792
rect 18898 21728 18914 21792
rect 18978 21728 18994 21792
rect 19058 21728 19066 21792
rect 18746 20704 19066 21728
rect 18746 20640 18754 20704
rect 18818 20640 18834 20704
rect 18898 20640 18914 20704
rect 18978 20640 18994 20704
rect 19058 20640 19066 20704
rect 18746 19616 19066 20640
rect 18746 19552 18754 19616
rect 18818 19552 18834 19616
rect 18898 19552 18914 19616
rect 18978 19552 18994 19616
rect 19058 19552 19066 19616
rect 18746 18528 19066 19552
rect 18746 18464 18754 18528
rect 18818 18464 18834 18528
rect 18898 18464 18914 18528
rect 18978 18464 18994 18528
rect 19058 18464 19066 18528
rect 18746 17440 19066 18464
rect 18746 17376 18754 17440
rect 18818 17376 18834 17440
rect 18898 17376 18914 17440
rect 18978 17376 18994 17440
rect 19058 17376 19066 17440
rect 18746 16352 19066 17376
rect 18746 16288 18754 16352
rect 18818 16288 18834 16352
rect 18898 16288 18914 16352
rect 18978 16288 18994 16352
rect 19058 16288 19066 16352
rect 18746 15264 19066 16288
rect 18746 15200 18754 15264
rect 18818 15200 18834 15264
rect 18898 15200 18914 15264
rect 18978 15200 18994 15264
rect 19058 15200 19066 15264
rect 18746 14176 19066 15200
rect 18746 14112 18754 14176
rect 18818 14112 18834 14176
rect 18898 14112 18914 14176
rect 18978 14112 18994 14176
rect 19058 14112 19066 14176
rect 18746 13088 19066 14112
rect 18746 13024 18754 13088
rect 18818 13024 18834 13088
rect 18898 13024 18914 13088
rect 18978 13024 18994 13088
rect 19058 13024 19066 13088
rect 18746 12000 19066 13024
rect 18746 11936 18754 12000
rect 18818 11936 18834 12000
rect 18898 11936 18914 12000
rect 18978 11936 18994 12000
rect 19058 11936 19066 12000
rect 18746 10912 19066 11936
rect 18746 10848 18754 10912
rect 18818 10848 18834 10912
rect 18898 10848 18914 10912
rect 18978 10848 18994 10912
rect 19058 10848 19066 10912
rect 18746 9824 19066 10848
rect 18746 9760 18754 9824
rect 18818 9760 18834 9824
rect 18898 9760 18914 9824
rect 18978 9760 18994 9824
rect 19058 9760 19066 9824
rect 18746 8736 19066 9760
rect 18746 8672 18754 8736
rect 18818 8672 18834 8736
rect 18898 8672 18914 8736
rect 18978 8672 18994 8736
rect 19058 8672 19066 8736
rect 18746 7648 19066 8672
rect 18746 7584 18754 7648
rect 18818 7584 18834 7648
rect 18898 7584 18914 7648
rect 18978 7584 18994 7648
rect 19058 7584 19066 7648
rect 18746 6560 19066 7584
rect 18746 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19066 6560
rect 18746 5472 19066 6496
rect 18746 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19066 5472
rect 18746 4384 19066 5408
rect 18746 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19066 4384
rect 18746 3296 19066 4320
rect 18746 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19066 3296
rect 18459 2684 18525 2685
rect 18459 2620 18460 2684
rect 18524 2620 18525 2684
rect 18459 2619 18525 2620
rect 18746 2208 19066 3232
rect 19382 2413 19442 32267
rect 19566 7989 19626 40019
rect 19747 39404 19813 39405
rect 19747 39340 19748 39404
rect 19812 39340 19813 39404
rect 19747 39339 19813 39340
rect 19750 17373 19810 39339
rect 21038 33149 21098 42059
rect 21713 41920 22033 42944
rect 21713 41856 21721 41920
rect 21785 41856 21801 41920
rect 21865 41856 21881 41920
rect 21945 41856 21961 41920
rect 22025 41856 22033 41920
rect 21713 40832 22033 41856
rect 21713 40768 21721 40832
rect 21785 40768 21801 40832
rect 21865 40768 21881 40832
rect 21945 40768 21961 40832
rect 22025 40768 22033 40832
rect 21713 39744 22033 40768
rect 21713 39680 21721 39744
rect 21785 39680 21801 39744
rect 21865 39680 21881 39744
rect 21945 39680 21961 39744
rect 22025 39680 22033 39744
rect 21403 38724 21469 38725
rect 21403 38660 21404 38724
rect 21468 38660 21469 38724
rect 21403 38659 21469 38660
rect 21219 36140 21285 36141
rect 21219 36076 21220 36140
rect 21284 36076 21285 36140
rect 21219 36075 21285 36076
rect 21035 33148 21101 33149
rect 21035 33084 21036 33148
rect 21100 33084 21101 33148
rect 21035 33083 21101 33084
rect 20115 26212 20181 26213
rect 20115 26148 20116 26212
rect 20180 26148 20181 26212
rect 20115 26147 20181 26148
rect 19747 17372 19813 17373
rect 19747 17308 19748 17372
rect 19812 17308 19813 17372
rect 19747 17307 19813 17308
rect 19931 17236 19997 17237
rect 19931 17172 19932 17236
rect 19996 17172 19997 17236
rect 19931 17171 19997 17172
rect 19563 7988 19629 7989
rect 19563 7924 19564 7988
rect 19628 7924 19629 7988
rect 19563 7923 19629 7924
rect 19747 4180 19813 4181
rect 19747 4116 19748 4180
rect 19812 4116 19813 4180
rect 19747 4115 19813 4116
rect 19563 3908 19629 3909
rect 19563 3844 19564 3908
rect 19628 3844 19629 3908
rect 19563 3843 19629 3844
rect 19566 2413 19626 3843
rect 19750 2685 19810 4115
rect 19747 2684 19813 2685
rect 19747 2620 19748 2684
rect 19812 2620 19813 2684
rect 19747 2619 19813 2620
rect 19379 2412 19445 2413
rect 19379 2348 19380 2412
rect 19444 2348 19445 2412
rect 19379 2347 19445 2348
rect 19563 2412 19629 2413
rect 19563 2348 19564 2412
rect 19628 2348 19629 2412
rect 19563 2347 19629 2348
rect 18746 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19066 2208
rect 18091 1324 18157 1325
rect 18091 1260 18092 1324
rect 18156 1260 18157 1324
rect 18091 1259 18157 1260
rect 18746 1120 19066 2144
rect 19934 1325 19994 17171
rect 20118 7309 20178 26147
rect 21035 21588 21101 21589
rect 21035 21524 21036 21588
rect 21100 21524 21101 21588
rect 21035 21523 21101 21524
rect 21038 10981 21098 21523
rect 21035 10980 21101 10981
rect 21035 10916 21036 10980
rect 21100 10916 21101 10980
rect 21035 10915 21101 10916
rect 20115 7308 20181 7309
rect 20115 7244 20116 7308
rect 20180 7244 20181 7308
rect 20115 7243 20181 7244
rect 21222 3909 21282 36075
rect 21406 22133 21466 38659
rect 21713 38656 22033 39680
rect 24680 43552 25000 43568
rect 24680 43488 24688 43552
rect 24752 43488 24768 43552
rect 24832 43488 24848 43552
rect 24912 43488 24928 43552
rect 24992 43488 25000 43552
rect 24680 42464 25000 43488
rect 24680 42400 24688 42464
rect 24752 42400 24768 42464
rect 24832 42400 24848 42464
rect 24912 42400 24928 42464
rect 24992 42400 25000 42464
rect 24680 41376 25000 42400
rect 24680 41312 24688 41376
rect 24752 41312 24768 41376
rect 24832 41312 24848 41376
rect 24912 41312 24928 41376
rect 24992 41312 25000 41376
rect 24680 40288 25000 41312
rect 24680 40224 24688 40288
rect 24752 40224 24768 40288
rect 24832 40224 24848 40288
rect 24912 40224 24928 40288
rect 24992 40224 25000 40288
rect 24680 39200 25000 40224
rect 24680 39136 24688 39200
rect 24752 39136 24768 39200
rect 24832 39136 24848 39200
rect 24912 39136 24928 39200
rect 24992 39136 25000 39200
rect 22507 38996 22573 38997
rect 22507 38932 22508 38996
rect 22572 38932 22573 38996
rect 22507 38931 22573 38932
rect 22323 38860 22389 38861
rect 22323 38796 22324 38860
rect 22388 38796 22389 38860
rect 22323 38795 22389 38796
rect 21713 38592 21721 38656
rect 21785 38592 21801 38656
rect 21865 38592 21881 38656
rect 21945 38592 21961 38656
rect 22025 38592 22033 38656
rect 21713 37568 22033 38592
rect 21713 37504 21721 37568
rect 21785 37504 21801 37568
rect 21865 37504 21881 37568
rect 21945 37504 21961 37568
rect 22025 37504 22033 37568
rect 21713 36480 22033 37504
rect 21713 36416 21721 36480
rect 21785 36416 21801 36480
rect 21865 36416 21881 36480
rect 21945 36416 21961 36480
rect 22025 36416 22033 36480
rect 21713 35392 22033 36416
rect 21713 35328 21721 35392
rect 21785 35328 21801 35392
rect 21865 35328 21881 35392
rect 21945 35328 21961 35392
rect 22025 35328 22033 35392
rect 21713 34304 22033 35328
rect 21713 34240 21721 34304
rect 21785 34240 21801 34304
rect 21865 34240 21881 34304
rect 21945 34240 21961 34304
rect 22025 34240 22033 34304
rect 21713 33216 22033 34240
rect 21713 33152 21721 33216
rect 21785 33152 21801 33216
rect 21865 33152 21881 33216
rect 21945 33152 21961 33216
rect 22025 33152 22033 33216
rect 21713 32128 22033 33152
rect 21713 32064 21721 32128
rect 21785 32064 21801 32128
rect 21865 32064 21881 32128
rect 21945 32064 21961 32128
rect 22025 32064 22033 32128
rect 21713 31040 22033 32064
rect 21713 30976 21721 31040
rect 21785 30976 21801 31040
rect 21865 30976 21881 31040
rect 21945 30976 21961 31040
rect 22025 30976 22033 31040
rect 21713 29952 22033 30976
rect 21713 29888 21721 29952
rect 21785 29888 21801 29952
rect 21865 29888 21881 29952
rect 21945 29888 21961 29952
rect 22025 29888 22033 29952
rect 21713 28864 22033 29888
rect 21713 28800 21721 28864
rect 21785 28800 21801 28864
rect 21865 28800 21881 28864
rect 21945 28800 21961 28864
rect 22025 28800 22033 28864
rect 21713 27776 22033 28800
rect 21713 27712 21721 27776
rect 21785 27712 21801 27776
rect 21865 27712 21881 27776
rect 21945 27712 21961 27776
rect 22025 27712 22033 27776
rect 21713 26688 22033 27712
rect 21713 26624 21721 26688
rect 21785 26624 21801 26688
rect 21865 26624 21881 26688
rect 21945 26624 21961 26688
rect 22025 26624 22033 26688
rect 21713 25600 22033 26624
rect 21713 25536 21721 25600
rect 21785 25536 21801 25600
rect 21865 25536 21881 25600
rect 21945 25536 21961 25600
rect 22025 25536 22033 25600
rect 21713 24512 22033 25536
rect 21713 24448 21721 24512
rect 21785 24448 21801 24512
rect 21865 24448 21881 24512
rect 21945 24448 21961 24512
rect 22025 24448 22033 24512
rect 21713 23424 22033 24448
rect 21713 23360 21721 23424
rect 21785 23360 21801 23424
rect 21865 23360 21881 23424
rect 21945 23360 21961 23424
rect 22025 23360 22033 23424
rect 21713 22336 22033 23360
rect 21713 22272 21721 22336
rect 21785 22272 21801 22336
rect 21865 22272 21881 22336
rect 21945 22272 21961 22336
rect 22025 22272 22033 22336
rect 21403 22132 21469 22133
rect 21403 22068 21404 22132
rect 21468 22068 21469 22132
rect 21403 22067 21469 22068
rect 21713 21248 22033 22272
rect 21713 21184 21721 21248
rect 21785 21184 21801 21248
rect 21865 21184 21881 21248
rect 21945 21184 21961 21248
rect 22025 21184 22033 21248
rect 21713 20160 22033 21184
rect 21713 20096 21721 20160
rect 21785 20096 21801 20160
rect 21865 20096 21881 20160
rect 21945 20096 21961 20160
rect 22025 20096 22033 20160
rect 21713 19072 22033 20096
rect 21713 19008 21721 19072
rect 21785 19008 21801 19072
rect 21865 19008 21881 19072
rect 21945 19008 21961 19072
rect 22025 19008 22033 19072
rect 21403 18052 21469 18053
rect 21403 17988 21404 18052
rect 21468 17988 21469 18052
rect 21403 17987 21469 17988
rect 21406 3909 21466 17987
rect 21713 17984 22033 19008
rect 21713 17920 21721 17984
rect 21785 17920 21801 17984
rect 21865 17920 21881 17984
rect 21945 17920 21961 17984
rect 22025 17920 22033 17984
rect 21713 16896 22033 17920
rect 21713 16832 21721 16896
rect 21785 16832 21801 16896
rect 21865 16832 21881 16896
rect 21945 16832 21961 16896
rect 22025 16832 22033 16896
rect 21713 15808 22033 16832
rect 22326 16013 22386 38795
rect 22510 23493 22570 38931
rect 24680 38112 25000 39136
rect 24680 38048 24688 38112
rect 24752 38048 24768 38112
rect 24832 38048 24848 38112
rect 24912 38048 24928 38112
rect 24992 38048 25000 38112
rect 24680 37024 25000 38048
rect 24680 36960 24688 37024
rect 24752 36960 24768 37024
rect 24832 36960 24848 37024
rect 24912 36960 24928 37024
rect 24992 36960 25000 37024
rect 24680 35936 25000 36960
rect 24680 35872 24688 35936
rect 24752 35872 24768 35936
rect 24832 35872 24848 35936
rect 24912 35872 24928 35936
rect 24992 35872 25000 35936
rect 24680 34848 25000 35872
rect 24680 34784 24688 34848
rect 24752 34784 24768 34848
rect 24832 34784 24848 34848
rect 24912 34784 24928 34848
rect 24992 34784 25000 34848
rect 22875 33964 22941 33965
rect 22875 33900 22876 33964
rect 22940 33900 22941 33964
rect 22875 33899 22941 33900
rect 22507 23492 22573 23493
rect 22507 23428 22508 23492
rect 22572 23428 22573 23492
rect 22507 23427 22573 23428
rect 22691 22676 22757 22677
rect 22691 22612 22692 22676
rect 22756 22612 22757 22676
rect 22691 22611 22757 22612
rect 22507 22132 22573 22133
rect 22507 22068 22508 22132
rect 22572 22068 22573 22132
rect 22507 22067 22573 22068
rect 22323 16012 22389 16013
rect 22323 15948 22324 16012
rect 22388 15948 22389 16012
rect 22323 15947 22389 15948
rect 21713 15744 21721 15808
rect 21785 15744 21801 15808
rect 21865 15744 21881 15808
rect 21945 15744 21961 15808
rect 22025 15744 22033 15808
rect 21713 14720 22033 15744
rect 21713 14656 21721 14720
rect 21785 14656 21801 14720
rect 21865 14656 21881 14720
rect 21945 14656 21961 14720
rect 22025 14656 22033 14720
rect 21713 13632 22033 14656
rect 21713 13568 21721 13632
rect 21785 13568 21801 13632
rect 21865 13568 21881 13632
rect 21945 13568 21961 13632
rect 22025 13568 22033 13632
rect 21713 12544 22033 13568
rect 21713 12480 21721 12544
rect 21785 12480 21801 12544
rect 21865 12480 21881 12544
rect 21945 12480 21961 12544
rect 22025 12480 22033 12544
rect 21713 11456 22033 12480
rect 22510 12341 22570 22067
rect 22507 12340 22573 12341
rect 22507 12276 22508 12340
rect 22572 12276 22573 12340
rect 22507 12275 22573 12276
rect 21713 11392 21721 11456
rect 21785 11392 21801 11456
rect 21865 11392 21881 11456
rect 21945 11392 21961 11456
rect 22025 11392 22033 11456
rect 21713 10368 22033 11392
rect 21713 10304 21721 10368
rect 21785 10304 21801 10368
rect 21865 10304 21881 10368
rect 21945 10304 21961 10368
rect 22025 10304 22033 10368
rect 21587 9484 21653 9485
rect 21587 9420 21588 9484
rect 21652 9420 21653 9484
rect 21587 9419 21653 9420
rect 21219 3908 21285 3909
rect 21219 3844 21220 3908
rect 21284 3844 21285 3908
rect 21219 3843 21285 3844
rect 21403 3908 21469 3909
rect 21403 3844 21404 3908
rect 21468 3844 21469 3908
rect 21403 3843 21469 3844
rect 21590 2549 21650 9419
rect 21713 9280 22033 10304
rect 21713 9216 21721 9280
rect 21785 9216 21801 9280
rect 21865 9216 21881 9280
rect 21945 9216 21961 9280
rect 22025 9216 22033 9280
rect 21713 8192 22033 9216
rect 21713 8128 21721 8192
rect 21785 8128 21801 8192
rect 21865 8128 21881 8192
rect 21945 8128 21961 8192
rect 22025 8128 22033 8192
rect 21713 7104 22033 8128
rect 21713 7040 21721 7104
rect 21785 7040 21801 7104
rect 21865 7040 21881 7104
rect 21945 7040 21961 7104
rect 22025 7040 22033 7104
rect 21713 6016 22033 7040
rect 21713 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22033 6016
rect 21713 4928 22033 5952
rect 22694 5541 22754 22611
rect 22878 20229 22938 33899
rect 24680 33760 25000 34784
rect 24680 33696 24688 33760
rect 24752 33696 24768 33760
rect 24832 33696 24848 33760
rect 24912 33696 24928 33760
rect 24992 33696 25000 33760
rect 24680 32672 25000 33696
rect 24680 32608 24688 32672
rect 24752 32608 24768 32672
rect 24832 32608 24848 32672
rect 24912 32608 24928 32672
rect 24992 32608 25000 32672
rect 24680 31584 25000 32608
rect 24680 31520 24688 31584
rect 24752 31520 24768 31584
rect 24832 31520 24848 31584
rect 24912 31520 24928 31584
rect 24992 31520 25000 31584
rect 24680 30496 25000 31520
rect 24680 30432 24688 30496
rect 24752 30432 24768 30496
rect 24832 30432 24848 30496
rect 24912 30432 24928 30496
rect 24992 30432 25000 30496
rect 24680 29408 25000 30432
rect 24680 29344 24688 29408
rect 24752 29344 24768 29408
rect 24832 29344 24848 29408
rect 24912 29344 24928 29408
rect 24992 29344 25000 29408
rect 24680 28320 25000 29344
rect 24680 28256 24688 28320
rect 24752 28256 24768 28320
rect 24832 28256 24848 28320
rect 24912 28256 24928 28320
rect 24992 28256 25000 28320
rect 24680 27232 25000 28256
rect 24680 27168 24688 27232
rect 24752 27168 24768 27232
rect 24832 27168 24848 27232
rect 24912 27168 24928 27232
rect 24992 27168 25000 27232
rect 24680 26144 25000 27168
rect 24680 26080 24688 26144
rect 24752 26080 24768 26144
rect 24832 26080 24848 26144
rect 24912 26080 24928 26144
rect 24992 26080 25000 26144
rect 24680 25056 25000 26080
rect 24680 24992 24688 25056
rect 24752 24992 24768 25056
rect 24832 24992 24848 25056
rect 24912 24992 24928 25056
rect 24992 24992 25000 25056
rect 24163 24172 24229 24173
rect 24163 24108 24164 24172
rect 24228 24108 24229 24172
rect 24163 24107 24229 24108
rect 24166 21181 24226 24107
rect 24680 23968 25000 24992
rect 24680 23904 24688 23968
rect 24752 23904 24768 23968
rect 24832 23904 24848 23968
rect 24912 23904 24928 23968
rect 24992 23904 25000 23968
rect 24680 22880 25000 23904
rect 24680 22816 24688 22880
rect 24752 22816 24768 22880
rect 24832 22816 24848 22880
rect 24912 22816 24928 22880
rect 24992 22816 25000 22880
rect 24680 21792 25000 22816
rect 24680 21728 24688 21792
rect 24752 21728 24768 21792
rect 24832 21728 24848 21792
rect 24912 21728 24928 21792
rect 24992 21728 25000 21792
rect 24163 21180 24229 21181
rect 24163 21116 24164 21180
rect 24228 21116 24229 21180
rect 24163 21115 24229 21116
rect 24680 20704 25000 21728
rect 24680 20640 24688 20704
rect 24752 20640 24768 20704
rect 24832 20640 24848 20704
rect 24912 20640 24928 20704
rect 24992 20640 25000 20704
rect 22875 20228 22941 20229
rect 22875 20164 22876 20228
rect 22940 20164 22941 20228
rect 22875 20163 22941 20164
rect 24680 19616 25000 20640
rect 24680 19552 24688 19616
rect 24752 19552 24768 19616
rect 24832 19552 24848 19616
rect 24912 19552 24928 19616
rect 24992 19552 25000 19616
rect 24680 18528 25000 19552
rect 24680 18464 24688 18528
rect 24752 18464 24768 18528
rect 24832 18464 24848 18528
rect 24912 18464 24928 18528
rect 24992 18464 25000 18528
rect 24680 17440 25000 18464
rect 24680 17376 24688 17440
rect 24752 17376 24768 17440
rect 24832 17376 24848 17440
rect 24912 17376 24928 17440
rect 24992 17376 25000 17440
rect 24680 16352 25000 17376
rect 24680 16288 24688 16352
rect 24752 16288 24768 16352
rect 24832 16288 24848 16352
rect 24912 16288 24928 16352
rect 24992 16288 25000 16352
rect 24680 15264 25000 16288
rect 24680 15200 24688 15264
rect 24752 15200 24768 15264
rect 24832 15200 24848 15264
rect 24912 15200 24928 15264
rect 24992 15200 25000 15264
rect 24680 14176 25000 15200
rect 24680 14112 24688 14176
rect 24752 14112 24768 14176
rect 24832 14112 24848 14176
rect 24912 14112 24928 14176
rect 24992 14112 25000 14176
rect 24680 13088 25000 14112
rect 24680 13024 24688 13088
rect 24752 13024 24768 13088
rect 24832 13024 24848 13088
rect 24912 13024 24928 13088
rect 24992 13024 25000 13088
rect 24680 12000 25000 13024
rect 24680 11936 24688 12000
rect 24752 11936 24768 12000
rect 24832 11936 24848 12000
rect 24912 11936 24928 12000
rect 24992 11936 25000 12000
rect 24680 10912 25000 11936
rect 24680 10848 24688 10912
rect 24752 10848 24768 10912
rect 24832 10848 24848 10912
rect 24912 10848 24928 10912
rect 24992 10848 25000 10912
rect 24680 9824 25000 10848
rect 24680 9760 24688 9824
rect 24752 9760 24768 9824
rect 24832 9760 24848 9824
rect 24912 9760 24928 9824
rect 24992 9760 25000 9824
rect 24680 8736 25000 9760
rect 24680 8672 24688 8736
rect 24752 8672 24768 8736
rect 24832 8672 24848 8736
rect 24912 8672 24928 8736
rect 24992 8672 25000 8736
rect 24680 7648 25000 8672
rect 24680 7584 24688 7648
rect 24752 7584 24768 7648
rect 24832 7584 24848 7648
rect 24912 7584 24928 7648
rect 24992 7584 25000 7648
rect 24680 6560 25000 7584
rect 24680 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 25000 6560
rect 22691 5540 22757 5541
rect 22691 5476 22692 5540
rect 22756 5476 22757 5540
rect 22691 5475 22757 5476
rect 21713 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22033 4928
rect 21713 3840 22033 4864
rect 21713 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22033 3840
rect 21713 2752 22033 3776
rect 21713 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22033 2752
rect 21587 2548 21653 2549
rect 21587 2484 21588 2548
rect 21652 2484 21653 2548
rect 21587 2483 21653 2484
rect 21713 1664 22033 2688
rect 21713 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22033 1664
rect 19931 1324 19997 1325
rect 19931 1260 19932 1324
rect 19996 1260 19997 1324
rect 19931 1259 19997 1260
rect 18746 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19066 1120
rect 18746 1040 19066 1056
rect 21713 1040 22033 1600
rect 24680 5472 25000 6496
rect 24680 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 25000 5472
rect 24680 4384 25000 5408
rect 24680 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 25000 4384
rect 24680 3296 25000 4320
rect 24680 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 25000 3296
rect 24680 2208 25000 3232
rect 24680 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 25000 2208
rect 24680 1120 25000 2144
rect 24680 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 25000 1120
rect 24680 1040 25000 1056
rect 17907 916 17973 917
rect 17907 852 17908 916
rect 17972 852 17973 916
rect 17907 851 17973 852
rect 8707 780 8773 781
rect 8707 716 8708 780
rect 8772 716 8773 780
rect 8707 715 8773 716
use sky130_fd_sc_hd__clkbuf_1  _000_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23644 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _001_
timestamp 1688980957
transform 1 0 23644 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _002_
timestamp 1688980957
transform 1 0 23644 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _003_
timestamp 1688980957
transform 1 0 21896 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _004_
timestamp 1688980957
transform 1 0 23460 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _005_
timestamp 1688980957
transform 1 0 22448 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _006_
timestamp 1688980957
transform 1 0 23276 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _007_
timestamp 1688980957
transform 1 0 23000 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _008_
timestamp 1688980957
transform 1 0 23460 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _009_
timestamp 1688980957
transform 1 0 23552 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _010_
timestamp 1688980957
transform 1 0 23368 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _011_
timestamp 1688980957
transform 1 0 23368 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _012_
timestamp 1688980957
transform 1 0 23000 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _013_
timestamp 1688980957
transform 1 0 23644 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _014_
timestamp 1688980957
transform 1 0 23276 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _015_
timestamp 1688980957
transform 1 0 22172 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _016_
timestamp 1688980957
transform 1 0 23276 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _017_
timestamp 1688980957
transform 1 0 23644 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _018_
timestamp 1688980957
transform 1 0 23644 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _019_
timestamp 1688980957
transform 1 0 19780 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _020_
timestamp 1688980957
transform 1 0 20884 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _021_
timestamp 1688980957
transform 1 0 23460 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _022_
timestamp 1688980957
transform 1 0 23460 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _023_
timestamp 1688980957
transform 1 0 19228 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _024_
timestamp 1688980957
transform 1 0 20792 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _025_
timestamp 1688980957
transform 1 0 22816 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _026_
timestamp 1688980957
transform 1 0 21528 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _027_
timestamp 1688980957
transform 1 0 19504 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _028_
timestamp 1688980957
transform 1 0 22724 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _029_
timestamp 1688980957
transform 1 0 20424 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _030_
timestamp 1688980957
transform 1 0 22908 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp 1688980957
transform 1 0 20976 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp 1688980957
transform 1 0 20516 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp 1688980957
transform 1 0 20792 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _034_
timestamp 1688980957
transform 1 0 20700 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp 1688980957
transform 1 0 21252 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp 1688980957
transform 1 0 20240 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp 1688980957
transform 1 0 18860 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp 1688980957
transform 1 0 21804 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _039_
timestamp 1688980957
transform 1 0 22080 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp 1688980957
transform 1 0 21160 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp 1688980957
transform 1 0 22816 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp 1688980957
transform 1 0 21252 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp 1688980957
transform 1 0 21436 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp 1688980957
transform 1 0 23368 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp 1688980957
transform 1 0 20148 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp 1688980957
transform 1 0 22540 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp 1688980957
transform 1 0 23092 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _048_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1688980957
transform 1 0 19964 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp 1688980957
transform 1 0 23184 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _051_
timestamp 1688980957
transform 1 0 23276 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_
timestamp 1688980957
transform 1 0 10948 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp 1688980957
transform 1 0 3404 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp 1688980957
transform 1 0 12328 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _055_
timestamp 1688980957
transform 1 0 15088 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1688980957
transform 1 0 4968 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1688980957
transform 1 0 4692 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1688980957
transform 1 0 5244 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1688980957
transform 1 0 3404 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1688980957
transform 1 0 2760 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1688980957
transform 1 0 5796 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1688980957
transform 1 0 6624 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1688980957
transform 1 0 5520 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1688980957
transform 1 0 4048 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1688980957
transform 1 0 6900 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1688980957
transform 1 0 4692 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1688980957
transform 1 0 4968 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1688980957
transform 1 0 5428 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1688980957
transform 1 0 6164 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1688980957
transform 1 0 3772 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1688980957
transform 1 0 6808 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform 1 0 7268 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1688980957
transform 1 0 5796 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform 1 0 7728 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform 1 0 8096 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform 1 0 8372 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1688980957
transform 1 0 10028 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform 1 0 10672 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform 1 0 7728 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1688980957
transform 1 0 10304 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1688980957
transform 1 0 16928 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1688980957
transform 1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1688980957
transform 1 0 11960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1688980957
transform 1 0 15272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1688980957
transform 1 0 13064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1688980957
transform 1 0 11868 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1688980957
transform 1 0 13340 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1688980957
transform 1 0 14076 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1688980957
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1688980957
transform 1 0 11684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1688980957
transform 1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1688980957
transform 1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1688980957
transform 1 0 13616 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1688980957
transform 1 0 15824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1688980957
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1688980957
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1688980957
transform 1 0 17296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1688980957
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1688980957
transform 1 0 19412 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1688980957
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1688980957
transform 1 0 17480 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1688980957
transform 1 0 24104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1688980957
transform 1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1688980957
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1688980957
transform 1 0 1472 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1688980957
transform 1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1688980957
transform 1 0 4048 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1688980957
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1688980957
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1688980957
transform 1 0 3772 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1688980957
transform 1 0 3404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1688980957
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1688980957
transform 1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1688980957
transform 1 0 5152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1688980957
transform 1 0 4692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1688980957
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp 1688980957
transform 1 0 5704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1688980957
transform 1 0 1472 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1688980957
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _145_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _146_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _147_
timestamp 1688980957
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1688980957
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1688980957
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _152_
timestamp 1688980957
transform 1 0 16928 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1688980957
transform 1 0 3772 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1688980957
transform 1 0 1748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1688980957
transform 1 0 10396 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1688980957
transform 1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1688980957
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1688980957
transform 1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1688980957
transform 1 0 3772 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1688980957
transform 1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1688980957
transform 1 0 3404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _163_
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _167_
timestamp 1688980957
transform 1 0 9752 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1688980957
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _171_
timestamp 1688980957
transform 1 0 9200 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12972 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 12328 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 18492 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 18492 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 9384 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1688980957
transform 1 0 11776 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1688980957
transform 1 0 23000 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1688980957
transform 1 0 4968 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1688980957
transform 1 0 4508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1688980957
transform 1 0 12328 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1688980957
transform 1 0 5336 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1688980957
transform 1 0 7176 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1688980957
transform 1 0 23000 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1688980957
transform 1 0 5612 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1688980957
transform 1 0 13248 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1688980957
transform 1 0 13800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_0._0_
timestamp 1688980957
transform 1 0 22448 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_1._0_
timestamp 1688980957
transform 1 0 22448 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_2._0_
timestamp 1688980957
transform 1 0 23092 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_3._0_
timestamp 1688980957
transform 1 0 20332 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_4._0_
timestamp 1688980957
transform 1 0 23184 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_5._0_
timestamp 1688980957
transform 1 0 23092 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_6._0_
timestamp 1688980957
transform 1 0 23000 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_7._0_
timestamp 1688980957
transform 1 0 23460 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_8._0_
timestamp 1688980957
transform 1 0 23184 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_9._0_
timestamp 1688980957
transform 1 0 21804 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_10._0_
timestamp 1688980957
transform 1 0 22080 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_11._0_
timestamp 1688980957
transform 1 0 22172 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_12._0_
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_13._0_
timestamp 1688980957
transform 1 0 23000 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_14._0_
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_15._0_
timestamp 1688980957
transform 1 0 20608 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_16._0_
timestamp 1688980957
transform 1 0 22356 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_17._0_
timestamp 1688980957
transform 1 0 23552 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_18._0_
timestamp 1688980957
transform 1 0 21528 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_19._0_
timestamp 1688980957
transform 1 0 18584 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_20._0_
timestamp 1688980957
transform 1 0 19504 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_21._0_
timestamp 1688980957
transform 1 0 21712 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_22._0_
timestamp 1688980957
transform 1 0 21896 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_23._0_
timestamp 1688980957
transform 1 0 18124 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_24._0_
timestamp 1688980957
transform 1 0 19412 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_25._0_
timestamp 1688980957
transform 1 0 21344 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_26._0_
timestamp 1688980957
transform 1 0 21896 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_27._0_
timestamp 1688980957
transform 1 0 19596 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_28._0_
timestamp 1688980957
transform 1 0 22080 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_29._0_
timestamp 1688980957
transform 1 0 20884 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_30._0_
timestamp 1688980957
transform 1 0 23000 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_31._0_
timestamp 1688980957
transform 1 0 21804 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_0._0_
timestamp 1688980957
transform 1 0 23092 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_1._0_
timestamp 1688980957
transform 1 0 23184 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_2._0_
timestamp 1688980957
transform 1 0 23368 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_3._0_
timestamp 1688980957
transform 1 0 21160 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_4._0_
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_5._0_
timestamp 1688980957
transform 1 0 23552 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_6._0_
timestamp 1688980957
transform 1 0 22724 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_7._0_
timestamp 1688980957
transform 1 0 23736 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_8._0_
timestamp 1688980957
transform 1 0 23276 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_9._0_
timestamp 1688980957
transform 1 0 22632 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_10._0_
timestamp 1688980957
transform 1 0 23000 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_11._0_
timestamp 1688980957
transform 1 0 23000 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_12._0_
timestamp 1688980957
transform 1 0 22448 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_13._0_
timestamp 1688980957
transform 1 0 22724 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_14._0_
timestamp 1688980957
transform 1 0 22448 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_15._0_
timestamp 1688980957
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_16._0_
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_17._0_
timestamp 1688980957
transform 1 0 23644 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_18._0_
timestamp 1688980957
transform 1 0 22356 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_19._0_
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_20._0_
timestamp 1688980957
transform 1 0 20148 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_21._0_
timestamp 1688980957
transform 1 0 22448 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_22._0_
timestamp 1688980957
transform 1 0 22908 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_23._0_
timestamp 1688980957
transform 1 0 18676 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_24._0_
timestamp 1688980957
transform 1 0 20148 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_25._0_
timestamp 1688980957
transform 1 0 22080 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_26._0_
timestamp 1688980957
transform 1 0 21620 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_27._0_
timestamp 1688980957
transform 1 0 22448 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_28._0_
timestamp 1688980957
transform 1 0 18308 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_29._0_
timestamp 1688980957
transform 1 0 21804 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_30._0_
timestamp 1688980957
transform 1 0 22908 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_31._0_
timestamp 1688980957
transform 1 0 19872 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_76
timestamp 1688980957
transform 1 0 8096 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_120
timestamp 1688980957
transform 1 0 12144 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_130
timestamp 1688980957
transform 1 0 13064 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_151
timestamp 1688980957
transform 1 0 14996 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_187
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_191
timestamp 1688980957
transform 1 0 18676 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_222
timestamp 1688980957
transform 1 0 21528 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_231
timestamp 1688980957
transform 1 0 22356 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_17
timestamp 1688980957
transform 1 0 2668 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_101
timestamp 1688980957
transform 1 0 10396 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_127
timestamp 1688980957
transform 1 0 12788 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_131
timestamp 1688980957
transform 1 0 13156 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_139
timestamp 1688980957
transform 1 0 13892 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_156
timestamp 1688980957
transform 1 0 15456 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_245
timestamp 1688980957
transform 1 0 23644 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_253
timestamp 1688980957
transform 1 0 24380 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_14
timestamp 1688980957
transform 1 0 2392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 1688980957
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_35
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_114
timestamp 1688980957
transform 1 0 11592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_129
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_163
timestamp 1688980957
transform 1 0 16100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_167
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_194
timestamp 1688980957
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_200
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_23
timestamp 1688980957
transform 1 0 3220 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_91
timestamp 1688980957
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_136
timestamp 1688980957
transform 1 0 13616 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_148
timestamp 1688980957
transform 1 0 14720 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_160
timestamp 1688980957
transform 1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_164
timestamp 1688980957
transform 1 0 16192 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_21
timestamp 1688980957
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_44
timestamp 1688980957
transform 1 0 5152 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_52
timestamp 1688980957
transform 1 0 5888 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_88
timestamp 1688980957
transform 1 0 9200 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_116
timestamp 1688980957
transform 1 0 11776 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_124
timestamp 1688980957
transform 1 0 12512 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_134
timestamp 1688980957
transform 1 0 13432 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_184
timestamp 1688980957
transform 1 0 18032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_200
timestamp 1688980957
transform 1 0 19504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_232
timestamp 1688980957
transform 1 0 22448 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1688980957
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_49
timestamp 1688980957
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_91
timestamp 1688980957
transform 1 0 9476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_103
timestamp 1688980957
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_117
timestamp 1688980957
transform 1 0 11868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_136
timestamp 1688980957
transform 1 0 13616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_140
timestamp 1688980957
transform 1 0 13984 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_146
timestamp 1688980957
transform 1 0 14536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_177
timestamp 1688980957
transform 1 0 17388 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_185
timestamp 1688980957
transform 1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_191
timestamp 1688980957
transform 1 0 18676 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_219
timestamp 1688980957
transform 1 0 21252 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_37
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_42
timestamp 1688980957
transform 1 0 4968 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_54
timestamp 1688980957
transform 1 0 6072 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_66 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7176 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_113
timestamp 1688980957
transform 1 0 11500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_129
timestamp 1688980957
transform 1 0 12972 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 1688980957
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_156
timestamp 1688980957
transform 1 0 15456 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_168
timestamp 1688980957
transform 1 0 16560 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_174
timestamp 1688980957
transform 1 0 17112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_246
timestamp 1688980957
transform 1 0 23736 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_72
timestamp 1688980957
transform 1 0 7728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_84
timestamp 1688980957
transform 1 0 8832 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_90
timestamp 1688980957
transform 1 0 9384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_157
timestamp 1688980957
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1688980957
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_189
timestamp 1688980957
transform 1 0 18492 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_214
timestamp 1688980957
transform 1 0 20792 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 1688980957
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_250
timestamp 1688980957
transform 1 0 24104 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_47
timestamp 1688980957
transform 1 0 5428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_69
timestamp 1688980957
transform 1 0 7452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 1688980957
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_102
timestamp 1688980957
transform 1 0 10488 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_136
timestamp 1688980957
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_205
timestamp 1688980957
transform 1 0 19964 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_227
timestamp 1688980957
transform 1 0 21988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_52
timestamp 1688980957
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_94
timestamp 1688980957
transform 1 0 9752 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_106
timestamp 1688980957
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_134
timestamp 1688980957
transform 1 0 13432 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_146
timestamp 1688980957
transform 1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_163
timestamp 1688980957
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_175
timestamp 1688980957
transform 1 0 17204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_198
timestamp 1688980957
transform 1 0 19320 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_210
timestamp 1688980957
transform 1 0 20424 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_238
timestamp 1688980957
transform 1 0 23000 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1688980957
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1688980957
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_100
timestamp 1688980957
transform 1 0 10304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_123
timestamp 1688980957
transform 1 0 12420 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_173
timestamp 1688980957
transform 1 0 17020 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_212
timestamp 1688980957
transform 1 0 20608 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_218
timestamp 1688980957
transform 1 0 21160 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_238
timestamp 1688980957
transform 1 0 23000 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_38
timestamp 1688980957
transform 1 0 4600 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_50
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_73
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_85
timestamp 1688980957
transform 1 0 8924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_91
timestamp 1688980957
transform 1 0 9476 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_109
timestamp 1688980957
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_156
timestamp 1688980957
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_219
timestamp 1688980957
transform 1 0 21252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_232
timestamp 1688980957
transform 1 0 22448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_236
timestamp 1688980957
transform 1 0 22816 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_244
timestamp 1688980957
transform 1 0 23552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_254
timestamp 1688980957
transform 1 0 24472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_100
timestamp 1688980957
transform 1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_104
timestamp 1688980957
transform 1 0 10672 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_120
timestamp 1688980957
transform 1 0 12144 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_132
timestamp 1688980957
transform 1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_176
timestamp 1688980957
transform 1 0 17296 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_188
timestamp 1688980957
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_214
timestamp 1688980957
transform 1 0 20792 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_31
timestamp 1688980957
transform 1 0 3956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_47
timestamp 1688980957
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_80
timestamp 1688980957
transform 1 0 8464 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_88
timestamp 1688980957
transform 1 0 9200 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_106
timestamp 1688980957
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_117
timestamp 1688980957
transform 1 0 11868 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_154
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1688980957
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_184
timestamp 1688980957
transform 1 0 18032 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_196
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_204
timestamp 1688980957
transform 1 0 19872 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1688980957
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_233
timestamp 1688980957
transform 1 0 22540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_50
timestamp 1688980957
transform 1 0 5704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_58
timestamp 1688980957
transform 1 0 6440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1688980957
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_110
timestamp 1688980957
transform 1 0 11224 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_116
timestamp 1688980957
transform 1 0 11776 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_132
timestamp 1688980957
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_149
timestamp 1688980957
transform 1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_188
timestamp 1688980957
transform 1 0 18400 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_203
timestamp 1688980957
transform 1 0 19780 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_226
timestamp 1688980957
transform 1 0 21896 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_234
timestamp 1688980957
transform 1 0 22632 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_65
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_97
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1688980957
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_131
timestamp 1688980957
transform 1 0 13156 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_143
timestamp 1688980957
transform 1 0 14260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_155
timestamp 1688980957
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_215
timestamp 1688980957
transform 1 0 20884 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_241
timestamp 1688980957
transform 1 0 23276 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_35
timestamp 1688980957
transform 1 0 4324 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_67
timestamp 1688980957
transform 1 0 7268 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_79
timestamp 1688980957
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_106
timestamp 1688980957
transform 1 0 10856 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_122
timestamp 1688980957
transform 1 0 12328 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_156
timestamp 1688980957
transform 1 0 15456 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_168
timestamp 1688980957
transform 1 0 16560 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_180
timestamp 1688980957
transform 1 0 17664 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_188
timestamp 1688980957
transform 1 0 18400 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 1688980957
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_203
timestamp 1688980957
transform 1 0 19780 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_12
timestamp 1688980957
transform 1 0 2208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_32
timestamp 1688980957
transform 1 0 4048 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_52
timestamp 1688980957
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_78
timestamp 1688980957
transform 1 0 8280 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_90
timestamp 1688980957
transform 1 0 9384 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_96
timestamp 1688980957
transform 1 0 9936 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_131
timestamp 1688980957
transform 1 0 13156 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_189
timestamp 1688980957
transform 1 0 18492 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_216
timestamp 1688980957
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_241
timestamp 1688980957
transform 1 0 23276 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_6
timestamp 1688980957
transform 1 0 1656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_51
timestamp 1688980957
transform 1 0 5796 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_63
timestamp 1688980957
transform 1 0 6900 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_75
timestamp 1688980957
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_102
timestamp 1688980957
transform 1 0 10488 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_114
timestamp 1688980957
transform 1 0 11592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_130
timestamp 1688980957
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1688980957
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_212
timestamp 1688980957
transform 1 0 20608 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_224
timestamp 1688980957
transform 1 0 21712 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_228
timestamp 1688980957
transform 1 0 22080 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1688980957
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_9
timestamp 1688980957
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_43
timestamp 1688980957
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_61
timestamp 1688980957
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_92
timestamp 1688980957
transform 1 0 9568 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_108
timestamp 1688980957
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_148
timestamp 1688980957
transform 1 0 14720 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_160
timestamp 1688980957
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_199
timestamp 1688980957
transform 1 0 19412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_228
timestamp 1688980957
transform 1 0 22080 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_249
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_35
timestamp 1688980957
transform 1 0 4324 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_93
timestamp 1688980957
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_127
timestamp 1688980957
transform 1 0 12788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_159
timestamp 1688980957
transform 1 0 15732 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_187
timestamp 1688980957
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_230
timestamp 1688980957
transform 1 0 22264 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_37
timestamp 1688980957
transform 1 0 4508 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_72
timestamp 1688980957
transform 1 0 7728 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_84
timestamp 1688980957
transform 1 0 8832 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_116
timestamp 1688980957
transform 1 0 11776 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_124
timestamp 1688980957
transform 1 0 12512 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_177
timestamp 1688980957
transform 1 0 17388 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_202
timestamp 1688980957
transform 1 0 19688 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_214
timestamp 1688980957
transform 1 0 20792 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_11
timestamp 1688980957
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_56
timestamp 1688980957
transform 1 0 6256 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_68
timestamp 1688980957
transform 1 0 7360 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_136
timestamp 1688980957
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_157
timestamp 1688980957
transform 1 0 15548 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_179
timestamp 1688980957
transform 1 0 17572 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_201
timestamp 1688980957
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_233
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1688980957
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_47
timestamp 1688980957
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_77
timestamp 1688980957
transform 1 0 8188 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_97
timestamp 1688980957
transform 1 0 10028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 1688980957
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_141
timestamp 1688980957
transform 1 0 14076 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_214
timestamp 1688980957
transform 1 0 20792 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_218
timestamp 1688980957
transform 1 0 21160 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1688980957
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_253
timestamp 1688980957
transform 1 0 24380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_9
timestamp 1688980957
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_35
timestamp 1688980957
transform 1 0 4324 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_39
timestamp 1688980957
transform 1 0 4692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_47
timestamp 1688980957
transform 1 0 5428 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_63
timestamp 1688980957
transform 1 0 6900 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_79
timestamp 1688980957
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_120
timestamp 1688980957
transform 1 0 12144 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_132
timestamp 1688980957
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_171
timestamp 1688980957
transform 1 0 16836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_183
timestamp 1688980957
transform 1 0 17940 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_201
timestamp 1688980957
transform 1 0 19596 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_206
timestamp 1688980957
transform 1 0 20056 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_212
timestamp 1688980957
transform 1 0 20608 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_235
timestamp 1688980957
transform 1 0 22724 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_32
timestamp 1688980957
transform 1 0 4048 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_40
timestamp 1688980957
transform 1 0 4784 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_82
timestamp 1688980957
transform 1 0 8648 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_90
timestamp 1688980957
transform 1 0 9384 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_108
timestamp 1688980957
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_131
timestamp 1688980957
transform 1 0 13156 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_139
timestamp 1688980957
transform 1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_163
timestamp 1688980957
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_185
timestamp 1688980957
transform 1 0 18124 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_202
timestamp 1688980957
transform 1 0 19688 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_214
timestamp 1688980957
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_222
timestamp 1688980957
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_32
timestamp 1688980957
transform 1 0 4048 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_40
timestamp 1688980957
transform 1 0 4784 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_44
timestamp 1688980957
transform 1 0 5152 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_79
timestamp 1688980957
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_89
timestamp 1688980957
transform 1 0 9292 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_111
timestamp 1688980957
transform 1 0 11316 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_115
timestamp 1688980957
transform 1 0 11684 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_134
timestamp 1688980957
transform 1 0 13432 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1688980957
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_225
timestamp 1688980957
transform 1 0 21804 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_233
timestamp 1688980957
transform 1 0 22540 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_244
timestamp 1688980957
transform 1 0 23552 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_9
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_50
timestamp 1688980957
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_110
timestamp 1688980957
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_133
timestamp 1688980957
transform 1 0 13340 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_152
timestamp 1688980957
transform 1 0 15088 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_164
timestamp 1688980957
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_194
timestamp 1688980957
transform 1 0 18952 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_240
timestamp 1688980957
transform 1 0 23184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_254
timestamp 1688980957
transform 1 0 24472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_47
timestamp 1688980957
transform 1 0 5428 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_59
timestamp 1688980957
transform 1 0 6532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 1688980957
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_120
timestamp 1688980957
transform 1 0 12144 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_124
timestamp 1688980957
transform 1 0 12512 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_192
timestamp 1688980957
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_215
timestamp 1688980957
transform 1 0 20884 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1688980957
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_32
timestamp 1688980957
transform 1 0 4048 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_44
timestamp 1688980957
transform 1 0 5152 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_90
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_106
timestamp 1688980957
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_130
timestamp 1688980957
transform 1 0 13064 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_138
timestamp 1688980957
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_143
timestamp 1688980957
transform 1 0 14260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 1688980957
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_203
timestamp 1688980957
transform 1 0 19780 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_215
timestamp 1688980957
transform 1 0 20884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_228
timestamp 1688980957
transform 1 0 22080 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_35
timestamp 1688980957
transform 1 0 4324 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_66
timestamp 1688980957
transform 1 0 7176 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_78
timestamp 1688980957
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_107
timestamp 1688980957
transform 1 0 10948 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_129
timestamp 1688980957
transform 1 0 12972 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_137
timestamp 1688980957
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_171
timestamp 1688980957
transform 1 0 16836 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_175
timestamp 1688980957
transform 1 0 17204 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_183
timestamp 1688980957
transform 1 0 17940 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_187
timestamp 1688980957
transform 1 0 18308 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_191
timestamp 1688980957
transform 1 0 18676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_212
timestamp 1688980957
transform 1 0 20608 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_228
timestamp 1688980957
transform 1 0 22080 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 1688980957
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_52
timestamp 1688980957
transform 1 0 5888 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_75
timestamp 1688980957
transform 1 0 8004 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_97
timestamp 1688980957
transform 1 0 10028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_104
timestamp 1688980957
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_119
timestamp 1688980957
transform 1 0 12052 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_148
timestamp 1688980957
transform 1 0 14720 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_152
timestamp 1688980957
transform 1 0 15088 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_205
timestamp 1688980957
transform 1 0 19964 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_222
timestamp 1688980957
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_235
timestamp 1688980957
transform 1 0 22724 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_11
timestamp 1688980957
transform 1 0 2116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_33
timestamp 1688980957
transform 1 0 4140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_49
timestamp 1688980957
transform 1 0 5612 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1688980957
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_156
timestamp 1688980957
transform 1 0 15456 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_180
timestamp 1688980957
transform 1 0 17664 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_192
timestamp 1688980957
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_204
timestamp 1688980957
transform 1 0 19872 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_210
timestamp 1688980957
transform 1 0 20424 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_214
timestamp 1688980957
transform 1 0 20792 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_218
timestamp 1688980957
transform 1 0 21160 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_222
timestamp 1688980957
transform 1 0 21528 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_234
timestamp 1688980957
transform 1 0 22632 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_37
timestamp 1688980957
transform 1 0 4508 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_49
timestamp 1688980957
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_84
timestamp 1688980957
transform 1 0 8832 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_100
timestamp 1688980957
transform 1 0 10304 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_164
timestamp 1688980957
transform 1 0 16192 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_184
timestamp 1688980957
transform 1 0 18032 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_196
timestamp 1688980957
transform 1 0 19136 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_208
timestamp 1688980957
transform 1 0 20240 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_220
timestamp 1688980957
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_231
timestamp 1688980957
transform 1 0 22356 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_247
timestamp 1688980957
transform 1 0 23828 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_32
timestamp 1688980957
transform 1 0 4048 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_44
timestamp 1688980957
transform 1 0 5152 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_60
timestamp 1688980957
transform 1 0 6624 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_72
timestamp 1688980957
transform 1 0 7728 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_129
timestamp 1688980957
transform 1 0 12972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_160
timestamp 1688980957
transform 1 0 15824 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_172
timestamp 1688980957
transform 1 0 16928 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_200
timestamp 1688980957
transform 1 0 19504 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_228
timestamp 1688980957
transform 1 0 22080 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_16
timestamp 1688980957
transform 1 0 2576 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_35
timestamp 1688980957
transform 1 0 4324 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_85
timestamp 1688980957
transform 1 0 8924 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_106
timestamp 1688980957
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_121
timestamp 1688980957
transform 1 0 12236 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_127
timestamp 1688980957
transform 1 0 12788 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_139
timestamp 1688980957
transform 1 0 13892 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_151
timestamp 1688980957
transform 1 0 14996 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_163
timestamp 1688980957
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_188
timestamp 1688980957
transform 1 0 18400 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_193
timestamp 1688980957
transform 1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_218
timestamp 1688980957
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_233
timestamp 1688980957
transform 1 0 22540 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_254
timestamp 1688980957
transform 1 0 24472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_10
timestamp 1688980957
transform 1 0 2024 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_26
timestamp 1688980957
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_37
timestamp 1688980957
transform 1 0 4508 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_54
timestamp 1688980957
transform 1 0 6072 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_62
timestamp 1688980957
transform 1 0 6808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_89
timestamp 1688980957
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_105
timestamp 1688980957
transform 1 0 10764 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_134
timestamp 1688980957
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_149
timestamp 1688980957
transform 1 0 14812 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_201
timestamp 1688980957
transform 1 0 19596 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_205
timestamp 1688980957
transform 1 0 19964 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_217
timestamp 1688980957
transform 1 0 21068 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_233
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_250
timestamp 1688980957
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_42
timestamp 1688980957
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 1688980957
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_75
timestamp 1688980957
transform 1 0 8004 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_92
timestamp 1688980957
transform 1 0 9568 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_104
timestamp 1688980957
transform 1 0 10672 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_128
timestamp 1688980957
transform 1 0 12880 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_147
timestamp 1688980957
transform 1 0 14628 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_163
timestamp 1688980957
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_190
timestamp 1688980957
transform 1 0 18584 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_208
timestamp 1688980957
transform 1 0 20240 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_217
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_254
timestamp 1688980957
transform 1 0 24472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_21
timestamp 1688980957
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_45
timestamp 1688980957
transform 1 0 5244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_57
timestamp 1688980957
transform 1 0 6348 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_73
timestamp 1688980957
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_81
timestamp 1688980957
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_106
timestamp 1688980957
transform 1 0 10856 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_166
timestamp 1688980957
transform 1 0 16376 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_178
timestamp 1688980957
transform 1 0 17480 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_190
timestamp 1688980957
transform 1 0 18584 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1688980957
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_201
timestamp 1688980957
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_206
timestamp 1688980957
transform 1 0 20056 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_224
timestamp 1688980957
transform 1 0 21712 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_228
timestamp 1688980957
transform 1 0 22080 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_247
timestamp 1688980957
transform 1 0 23828 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_21
timestamp 1688980957
transform 1 0 3036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_32
timestamp 1688980957
transform 1 0 4048 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_90
timestamp 1688980957
transform 1 0 9384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_118
timestamp 1688980957
transform 1 0 11960 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_141
timestamp 1688980957
transform 1 0 14076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_160
timestamp 1688980957
transform 1 0 15824 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_210
timestamp 1688980957
transform 1 0 20424 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 1688980957
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_241
timestamp 1688980957
transform 1 0 23276 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_248
timestamp 1688980957
transform 1 0 23920 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_37
timestamp 1688980957
transform 1 0 4508 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_55
timestamp 1688980957
transform 1 0 6164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_61
timestamp 1688980957
transform 1 0 6716 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_88
timestamp 1688980957
transform 1 0 9200 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_111
timestamp 1688980957
transform 1 0 11316 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_123
timestamp 1688980957
transform 1 0 12420 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_135
timestamp 1688980957
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_176
timestamp 1688980957
transform 1 0 17296 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_183
timestamp 1688980957
transform 1 0 17940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_230
timestamp 1688980957
transform 1 0 22264 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_238
timestamp 1688980957
transform 1 0 23000 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_28
timestamp 1688980957
transform 1 0 3680 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_34
timestamp 1688980957
transform 1 0 4232 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_75
timestamp 1688980957
transform 1 0 8004 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_91
timestamp 1688980957
transform 1 0 9476 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_103
timestamp 1688980957
transform 1 0 10580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_128
timestamp 1688980957
transform 1 0 12880 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_140
timestamp 1688980957
transform 1 0 13984 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_148
timestamp 1688980957
transform 1 0 14720 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_166
timestamp 1688980957
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_191
timestamp 1688980957
transform 1 0 18676 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_203
timestamp 1688980957
transform 1 0 19780 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_211
timestamp 1688980957
transform 1 0 20516 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_217
timestamp 1688980957
transform 1 0 21068 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_247
timestamp 1688980957
transform 1 0 23828 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_23
timestamp 1688980957
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_44
timestamp 1688980957
transform 1 0 5152 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_56
timestamp 1688980957
transform 1 0 6256 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_68
timestamp 1688980957
transform 1 0 7360 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_80
timestamp 1688980957
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_103
timestamp 1688980957
transform 1 0 10580 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_111
timestamp 1688980957
transform 1 0 11316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_135
timestamp 1688980957
transform 1 0 13524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_162
timestamp 1688980957
transform 1 0 16008 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_169
timestamp 1688980957
transform 1 0 16652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_188
timestamp 1688980957
transform 1 0 18400 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_200
timestamp 1688980957
transform 1 0 19504 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_225
timestamp 1688980957
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_246
timestamp 1688980957
transform 1 0 23736 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_21
timestamp 1688980957
transform 1 0 3036 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_41
timestamp 1688980957
transform 1 0 4876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_53
timestamp 1688980957
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_72
timestamp 1688980957
transform 1 0 7728 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_119
timestamp 1688980957
transform 1 0 12052 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_135
timestamp 1688980957
transform 1 0 13524 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_147
timestamp 1688980957
transform 1 0 14628 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_159
timestamp 1688980957
transform 1 0 15732 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_163
timestamp 1688980957
transform 1 0 16100 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_175
timestamp 1688980957
transform 1 0 17204 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_179
timestamp 1688980957
transform 1 0 17572 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_187
timestamp 1688980957
transform 1 0 18308 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_220
timestamp 1688980957
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_229
timestamp 1688980957
transform 1 0 22172 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_236
timestamp 1688980957
transform 1 0 22816 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_247
timestamp 1688980957
transform 1 0 23828 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_12
timestamp 1688980957
transform 1 0 2208 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_37
timestamp 1688980957
transform 1 0 4508 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_72
timestamp 1688980957
transform 1 0 7728 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_114
timestamp 1688980957
transform 1 0 11592 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_138
timestamp 1688980957
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_162
timestamp 1688980957
transform 1 0 16008 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_174
timestamp 1688980957
transform 1 0 17112 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_178
timestamp 1688980957
transform 1 0 17480 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_194
timestamp 1688980957
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_205
timestamp 1688980957
transform 1 0 19964 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_212
timestamp 1688980957
transform 1 0 20608 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_224
timestamp 1688980957
transform 1 0 21712 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_236
timestamp 1688980957
transform 1 0 22816 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_242
timestamp 1688980957
transform 1 0 23368 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_18
timestamp 1688980957
transform 1 0 2760 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_30
timestamp 1688980957
transform 1 0 3864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_49
timestamp 1688980957
transform 1 0 5612 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_62
timestamp 1688980957
transform 1 0 6808 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_85
timestamp 1688980957
transform 1 0 8924 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_177
timestamp 1688980957
transform 1 0 17388 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_205
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_209
timestamp 1688980957
transform 1 0 20332 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_213
timestamp 1688980957
transform 1 0 20700 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_220
timestamp 1688980957
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_229
timestamp 1688980957
transform 1 0 22172 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_243
timestamp 1688980957
transform 1 0 23460 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_6
timestamp 1688980957
transform 1 0 1656 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_22
timestamp 1688980957
transform 1 0 3128 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_33
timestamp 1688980957
transform 1 0 4140 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_49
timestamp 1688980957
transform 1 0 5612 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_61
timestamp 1688980957
transform 1 0 6716 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_82
timestamp 1688980957
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_128
timestamp 1688980957
transform 1 0 12880 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_183
timestamp 1688980957
transform 1 0 17940 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_187
timestamp 1688980957
transform 1 0 18308 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_191
timestamp 1688980957
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_23
timestamp 1688980957
transform 1 0 3220 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_44
timestamp 1688980957
transform 1 0 5152 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_88
timestamp 1688980957
transform 1 0 9200 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_104
timestamp 1688980957
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_156
timestamp 1688980957
transform 1 0 15456 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_184
timestamp 1688980957
transform 1 0 18032 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_196
timestamp 1688980957
transform 1 0 19136 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_208
timestamp 1688980957
transform 1 0 20240 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_220
timestamp 1688980957
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_253
timestamp 1688980957
transform 1 0 24380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_32
timestamp 1688980957
transform 1 0 4048 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_71
timestamp 1688980957
transform 1 0 7636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_105
timestamp 1688980957
transform 1 0 10764 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_115
timestamp 1688980957
transform 1 0 11684 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_132
timestamp 1688980957
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_157
timestamp 1688980957
transform 1 0 15548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_169
timestamp 1688980957
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_181
timestamp 1688980957
transform 1 0 17756 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_189
timestamp 1688980957
transform 1 0 18492 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_193
timestamp 1688980957
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_201
timestamp 1688980957
transform 1 0 19596 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_207
timestamp 1688980957
transform 1 0 20148 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_219
timestamp 1688980957
transform 1 0 21252 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_231
timestamp 1688980957
transform 1 0 22356 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_235
timestamp 1688980957
transform 1 0 22724 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_54
timestamp 1688980957
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_65
timestamp 1688980957
transform 1 0 7084 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_117
timestamp 1688980957
transform 1 0 11868 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_129
timestamp 1688980957
transform 1 0 12972 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_141
timestamp 1688980957
transform 1 0 14076 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_164
timestamp 1688980957
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_215
timestamp 1688980957
transform 1 0 20884 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_221
timestamp 1688980957
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_229
timestamp 1688980957
transform 1 0 22172 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_235
timestamp 1688980957
transform 1 0 22724 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_239
timestamp 1688980957
transform 1 0 23092 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_243
timestamp 1688980957
transform 1 0 23460 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_248
timestamp 1688980957
transform 1 0 23920 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_11
timestamp 1688980957
transform 1 0 2116 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_47
timestamp 1688980957
transform 1 0 5428 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_55
timestamp 1688980957
transform 1 0 6164 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_71
timestamp 1688980957
transform 1 0 7636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_201
timestamp 1688980957
transform 1 0 19596 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_208
timestamp 1688980957
transform 1 0 20240 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_228
timestamp 1688980957
transform 1 0 22080 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_24
timestamp 1688980957
transform 1 0 3312 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_35
timestamp 1688980957
transform 1 0 4324 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_54
timestamp 1688980957
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_102
timestamp 1688980957
transform 1 0 10488 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_110
timestamp 1688980957
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_117
timestamp 1688980957
transform 1 0 11868 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_121
timestamp 1688980957
transform 1 0 12236 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_156
timestamp 1688980957
transform 1 0 15456 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_188
timestamp 1688980957
transform 1 0 18400 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_200
timestamp 1688980957
transform 1 0 19504 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_212
timestamp 1688980957
transform 1 0 20608 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_221
timestamp 1688980957
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_234
timestamp 1688980957
transform 1 0 22632 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_243
timestamp 1688980957
transform 1 0 23460 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_248
timestamp 1688980957
transform 1 0 23920 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_19
timestamp 1688980957
transform 1 0 2852 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_23
timestamp 1688980957
transform 1 0 3220 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_75
timestamp 1688980957
transform 1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_93
timestamp 1688980957
transform 1 0 9660 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_137
timestamp 1688980957
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_171
timestamp 1688980957
transform 1 0 16836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_183
timestamp 1688980957
transform 1 0 17940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_219
timestamp 1688980957
transform 1 0 21252 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_235
timestamp 1688980957
transform 1 0 22724 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_242
timestamp 1688980957
transform 1 0 23368 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_13
timestamp 1688980957
transform 1 0 2300 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_33
timestamp 1688980957
transform 1 0 4140 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_37
timestamp 1688980957
transform 1 0 4508 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_90
timestamp 1688980957
transform 1 0 9384 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_120
timestamp 1688980957
transform 1 0 12144 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_124
timestamp 1688980957
transform 1 0 12512 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_129
timestamp 1688980957
transform 1 0 12972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_141
timestamp 1688980957
transform 1 0 14076 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_145
timestamp 1688980957
transform 1 0 14444 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_231
timestamp 1688980957
transform 1 0 22356 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_247
timestamp 1688980957
transform 1 0 23828 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_32
timestamp 1688980957
transform 1 0 4048 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_56
timestamp 1688980957
transform 1 0 6256 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_68
timestamp 1688980957
transform 1 0 7360 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_116
timestamp 1688980957
transform 1 0 11776 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_120
timestamp 1688980957
transform 1 0 12144 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_123
timestamp 1688980957
transform 1 0 12420 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_175
timestamp 1688980957
transform 1 0 17204 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_194
timestamp 1688980957
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_206
timestamp 1688980957
transform 1 0 20056 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_214
timestamp 1688980957
transform 1 0 20792 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_218
timestamp 1688980957
transform 1 0 21160 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_230
timestamp 1688980957
transform 1 0 22264 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_244
timestamp 1688980957
transform 1 0 23552 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_7
timestamp 1688980957
transform 1 0 1748 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_32
timestamp 1688980957
transform 1 0 4048 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_40
timestamp 1688980957
transform 1 0 4784 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_75
timestamp 1688980957
transform 1 0 8004 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_91
timestamp 1688980957
transform 1 0 9476 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_103
timestamp 1688980957
transform 1 0 10580 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_143
timestamp 1688980957
transform 1 0 14260 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_151
timestamp 1688980957
transform 1 0 14996 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_186
timestamp 1688980957
transform 1 0 18216 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_198
timestamp 1688980957
transform 1 0 19320 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_210
timestamp 1688980957
transform 1 0 20424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_222
timestamp 1688980957
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_243
timestamp 1688980957
transform 1 0 23460 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_248
timestamp 1688980957
transform 1 0 23920 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_24
timestamp 1688980957
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_48
timestamp 1688980957
transform 1 0 5520 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_114
timestamp 1688980957
transform 1 0 11592 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_118
timestamp 1688980957
transform 1 0 11960 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_135
timestamp 1688980957
transform 1 0 13524 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_157
timestamp 1688980957
transform 1 0 15548 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_179
timestamp 1688980957
transform 1 0 17572 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_191
timestamp 1688980957
transform 1 0 18676 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_229
timestamp 1688980957
transform 1 0 22172 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_24
timestamp 1688980957
transform 1 0 3312 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_28
timestamp 1688980957
transform 1 0 3680 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_44
timestamp 1688980957
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_91
timestamp 1688980957
transform 1 0 9476 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_118
timestamp 1688980957
transform 1 0 11960 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_130
timestamp 1688980957
transform 1 0 13064 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_138
timestamp 1688980957
transform 1 0 13800 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_157
timestamp 1688980957
transform 1 0 15548 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_165
timestamp 1688980957
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_217
timestamp 1688980957
transform 1 0 21068 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_241
timestamp 1688980957
transform 1 0 23276 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_24
timestamp 1688980957
transform 1 0 3312 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_47
timestamp 1688980957
transform 1 0 5428 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_51
timestamp 1688980957
transform 1 0 5796 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_71
timestamp 1688980957
transform 1 0 7636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_92
timestamp 1688980957
transform 1 0 9568 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_179
timestamp 1688980957
transform 1 0 17572 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_223
timestamp 1688980957
transform 1 0 21620 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_228
timestamp 1688980957
transform 1 0 22080 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_237
timestamp 1688980957
transform 1 0 22908 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_247
timestamp 1688980957
transform 1 0 23828 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_21
timestamp 1688980957
transform 1 0 3036 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_40
timestamp 1688980957
transform 1 0 4784 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_52
timestamp 1688980957
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_106
timestamp 1688980957
transform 1 0 10856 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_135
timestamp 1688980957
transform 1 0 13524 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_160
timestamp 1688980957
transform 1 0 15824 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_173
timestamp 1688980957
transform 1 0 17020 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_177
timestamp 1688980957
transform 1 0 17388 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_188
timestamp 1688980957
transform 1 0 18400 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_194
timestamp 1688980957
transform 1 0 18952 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_210
timestamp 1688980957
transform 1 0 20424 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_222
timestamp 1688980957
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_231
timestamp 1688980957
transform 1 0 22356 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_241
timestamp 1688980957
transform 1 0 23276 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_245
timestamp 1688980957
transform 1 0 23644 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_24
timestamp 1688980957
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_47
timestamp 1688980957
transform 1 0 5428 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_63
timestamp 1688980957
transform 1 0 6900 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_79
timestamp 1688980957
transform 1 0 8372 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_95
timestamp 1688980957
transform 1 0 9844 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_102
timestamp 1688980957
transform 1 0 10488 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_114
timestamp 1688980957
transform 1 0 11592 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_135
timestamp 1688980957
transform 1 0 13524 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_171
timestamp 1688980957
transform 1 0 16836 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_180
timestamp 1688980957
transform 1 0 17664 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_192
timestamp 1688980957
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_224
timestamp 1688980957
transform 1 0 21712 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_228
timestamp 1688980957
transform 1 0 22080 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_235
timestamp 1688980957
transform 1 0 22724 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_241
timestamp 1688980957
transform 1 0 23276 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_19
timestamp 1688980957
transform 1 0 2852 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_72
timestamp 1688980957
transform 1 0 7728 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_90
timestamp 1688980957
transform 1 0 9384 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_102
timestamp 1688980957
transform 1 0 10488 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_110
timestamp 1688980957
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_156
timestamp 1688980957
transform 1 0 15456 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_184
timestamp 1688980957
transform 1 0 18032 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_196
timestamp 1688980957
transform 1 0 19136 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_208
timestamp 1688980957
transform 1 0 20240 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_215
timestamp 1688980957
transform 1 0 20884 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_228
timestamp 1688980957
transform 1 0 22080 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_244
timestamp 1688980957
transform 1 0 23552 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_248
timestamp 1688980957
transform 1 0 23920 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_26
timestamp 1688980957
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_47
timestamp 1688980957
transform 1 0 5428 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_82
timestamp 1688980957
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_134
timestamp 1688980957
transform 1 0 13432 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_200
timestamp 1688980957
transform 1 0 19504 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_223
timestamp 1688980957
transform 1 0 21620 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_232
timestamp 1688980957
transform 1 0 22448 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_9
timestamp 1688980957
transform 1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_13
timestamp 1688980957
transform 1 0 2300 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_132
timestamp 1688980957
transform 1 0 13248 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_140
timestamp 1688980957
transform 1 0 13984 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_156
timestamp 1688980957
transform 1 0 15456 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_177
timestamp 1688980957
transform 1 0 17388 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_200
timestamp 1688980957
transform 1 0 19504 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_240
timestamp 1688980957
transform 1 0 23184 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_247
timestamp 1688980957
transform 1 0 23828 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_9
timestamp 1688980957
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_66
timestamp 1688980957
transform 1 0 7176 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_78
timestamp 1688980957
transform 1 0 8280 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_89
timestamp 1688980957
transform 1 0 9292 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_120
timestamp 1688980957
transform 1 0 12144 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_136
timestamp 1688980957
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_177
timestamp 1688980957
transform 1 0 17388 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_188
timestamp 1688980957
transform 1 0 18400 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_194
timestamp 1688980957
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_200
timestamp 1688980957
transform 1 0 19504 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_225
timestamp 1688980957
transform 1 0 21804 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_239
timestamp 1688980957
transform 1 0 23092 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_18
timestamp 1688980957
transform 1 0 2760 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_53
timestamp 1688980957
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_65
timestamp 1688980957
transform 1 0 7084 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_72
timestamp 1688980957
transform 1 0 7728 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_84
timestamp 1688980957
transform 1 0 8832 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_92
timestamp 1688980957
transform 1 0 9568 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_110
timestamp 1688980957
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_161
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_189
timestamp 1688980957
transform 1 0 18492 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_193
timestamp 1688980957
transform 1 0 18860 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_199
timestamp 1688980957
transform 1 0 19412 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_203
timestamp 1688980957
transform 1 0 19780 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_215
timestamp 1688980957
transform 1 0 20884 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 1688980957
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_234
timestamp 1688980957
transform 1 0 22632 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_240
timestamp 1688980957
transform 1 0 23184 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_248
timestamp 1688980957
transform 1 0 23920 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_24
timestamp 1688980957
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_58
timestamp 1688980957
transform 1 0 6440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_78
timestamp 1688980957
transform 1 0 8280 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_100
timestamp 1688980957
transform 1 0 10304 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_112
timestamp 1688980957
transform 1 0 11408 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_124
timestamp 1688980957
transform 1 0 12512 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_136
timestamp 1688980957
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1688980957
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 1688980957
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1688980957
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_200
timestamp 1688980957
transform 1 0 19504 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_206
timestamp 1688980957
transform 1 0 20056 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_210
timestamp 1688980957
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_222
timestamp 1688980957
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_227
timestamp 1688980957
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_231
timestamp 1688980957
transform 1 0 22356 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_235
timestamp 1688980957
transform 1 0 22724 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_243
timestamp 1688980957
transform 1 0 23460 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_36
timestamp 1688980957
transform 1 0 4416 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_53
timestamp 1688980957
transform 1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_65
timestamp 1688980957
transform 1 0 7084 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_71
timestamp 1688980957
transform 1 0 7636 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_77
timestamp 1688980957
transform 1 0 8188 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_96
timestamp 1688980957
transform 1 0 9936 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_108
timestamp 1688980957
transform 1 0 11040 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_141
timestamp 1688980957
transform 1 0 14076 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_153
timestamp 1688980957
transform 1 0 15180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_165
timestamp 1688980957
transform 1 0 16284 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_181
timestamp 1688980957
transform 1 0 17756 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_188
timestamp 1688980957
transform 1 0 18400 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_200
timestamp 1688980957
transform 1 0 19504 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_212
timestamp 1688980957
transform 1 0 20608 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_218
timestamp 1688980957
transform 1 0 21160 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_229
timestamp 1688980957
transform 1 0 22172 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_240
timestamp 1688980957
transform 1 0 23184 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_248
timestamp 1688980957
transform 1 0 23920 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_26
timestamp 1688980957
transform 1 0 3496 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_44
timestamp 1688980957
transform 1 0 5152 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_56
timestamp 1688980957
transform 1 0 6256 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_68
timestamp 1688980957
transform 1 0 7360 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_114
timestamp 1688980957
transform 1 0 11592 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_118
timestamp 1688980957
transform 1 0 11960 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 1688980957
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_189
timestamp 1688980957
transform 1 0 18492 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_194
timestamp 1688980957
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_202
timestamp 1688980957
transform 1 0 19688 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_210
timestamp 1688980957
transform 1 0 20424 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_246
timestamp 1688980957
transform 1 0 23736 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_253
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_38
timestamp 1688980957
transform 1 0 4600 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_50
timestamp 1688980957
transform 1 0 5704 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_63
timestamp 1688980957
transform 1 0 6900 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_137
timestamp 1688980957
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_149
timestamp 1688980957
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_161
timestamp 1688980957
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_167
timestamp 1688980957
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 1688980957
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_193
timestamp 1688980957
transform 1 0 18860 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_200
timestamp 1688980957
transform 1 0 19504 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_206
timestamp 1688980957
transform 1 0 20056 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_213
timestamp 1688980957
transform 1 0 20700 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_220
timestamp 1688980957
transform 1 0 21344 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_228
timestamp 1688980957
transform 1 0 22080 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_236
timestamp 1688980957
transform 1 0 22816 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_9
timestamp 1688980957
transform 1 0 1932 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_32
timestamp 1688980957
transform 1 0 4048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_75
timestamp 1688980957
transform 1 0 8004 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_103
timestamp 1688980957
transform 1 0 10580 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_136
timestamp 1688980957
transform 1 0 13616 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_165
timestamp 1688980957
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_177
timestamp 1688980957
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_189
timestamp 1688980957
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_195
timestamp 1688980957
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_209
timestamp 1688980957
transform 1 0 20332 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_213
timestamp 1688980957
transform 1 0 20700 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_241
timestamp 1688980957
transform 1 0 23276 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_246
timestamp 1688980957
transform 1 0 23736 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_253
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_39
timestamp 1688980957
transform 1 0 4692 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_74
timestamp 1688980957
transform 1 0 7912 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_98
timestamp 1688980957
transform 1 0 10120 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_110
timestamp 1688980957
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1688980957
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 1688980957
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 1688980957
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 1688980957
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 1688980957
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1688980957
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_193
timestamp 1688980957
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_214
timestamp 1688980957
transform 1 0 20792 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_234
timestamp 1688980957
transform 1 0 22632 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_245
timestamp 1688980957
transform 1 0 23644 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_93
timestamp 1688980957
transform 1 0 9660 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_116
timestamp 1688980957
transform 1 0 11776 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_128
timestamp 1688980957
transform 1 0 12880 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 1688980957
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_177
timestamp 1688980957
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_189
timestamp 1688980957
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_195
timestamp 1688980957
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_231
timestamp 1688980957
transform 1 0 22356 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_236
timestamp 1688980957
transform 1 0 22816 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_253
timestamp 1688980957
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_54
timestamp 1688980957
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_66
timestamp 1688980957
transform 1 0 7176 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_78
timestamp 1688980957
transform 1 0 8280 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_90
timestamp 1688980957
transform 1 0 9384 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_94
timestamp 1688980957
transform 1 0 9752 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_116
timestamp 1688980957
transform 1 0 11776 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_128
timestamp 1688980957
transform 1 0 12880 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_140
timestamp 1688980957
transform 1 0 13984 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_152
timestamp 1688980957
transform 1 0 15088 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_164
timestamp 1688980957
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_181
timestamp 1688980957
transform 1 0 17756 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_189
timestamp 1688980957
transform 1 0 18492 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_197
timestamp 1688980957
transform 1 0 19228 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_202
timestamp 1688980957
transform 1 0 19688 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_213
timestamp 1688980957
transform 1 0 20700 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_217
timestamp 1688980957
transform 1 0 21068 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_231
timestamp 1688980957
transform 1 0 22356 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_253
timestamp 1688980957
transform 1 0 24380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_45
timestamp 1688980957
transform 1 0 5244 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_50
timestamp 1688980957
transform 1 0 5704 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_54
timestamp 1688980957
transform 1 0 6072 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_58
timestamp 1688980957
transform 1 0 6440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_70
timestamp 1688980957
transform 1 0 7544 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_75
timestamp 1688980957
transform 1 0 8004 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_82
timestamp 1688980957
transform 1 0 8648 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_88
timestamp 1688980957
transform 1 0 9200 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_92
timestamp 1688980957
transform 1 0 9568 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1688980957
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 1688980957
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 1688980957
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_153
timestamp 1688980957
transform 1 0 15180 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_161
timestamp 1688980957
transform 1 0 15916 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_170
timestamp 1688980957
transform 1 0 16744 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_182
timestamp 1688980957
transform 1 0 17848 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_186
timestamp 1688980957
transform 1 0 18216 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_212
timestamp 1688980957
transform 1 0 20608 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_253
timestamp 1688980957
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_44
timestamp 1688980957
transform 1 0 5152 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_48
timestamp 1688980957
transform 1 0 5520 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_64
timestamp 1688980957
transform 1 0 6992 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_84
timestamp 1688980957
transform 1 0 8832 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_101
timestamp 1688980957
transform 1 0 10396 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75_109
timestamp 1688980957
transform 1 0 11132 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 1688980957
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_161
timestamp 1688980957
transform 1 0 15916 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_204
timestamp 1688980957
transform 1 0 19872 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_217
timestamp 1688980957
transform 1 0 21068 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_14
timestamp 1688980957
transform 1 0 2392 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_77
timestamp 1688980957
transform 1 0 8188 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_88
timestamp 1688980957
transform 1 0 9200 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_96
timestamp 1688980957
transform 1 0 9936 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_103
timestamp 1688980957
transform 1 0 10580 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_110
timestamp 1688980957
transform 1 0 11224 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_120
timestamp 1688980957
transform 1 0 12144 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_125
timestamp 1688980957
transform 1 0 12604 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_132
timestamp 1688980957
transform 1 0 13248 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_150
timestamp 1688980957
transform 1 0 14904 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_158
timestamp 1688980957
transform 1 0 15640 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_166
timestamp 1688980957
transform 1 0 16376 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_217
timestamp 1688980957
transform 1 0 21068 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_251
timestamp 1688980957
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_253
timestamp 1688980957
transform 1 0 24380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_54
timestamp 1688980957
transform 1 0 6072 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_66
timestamp 1688980957
transform 1 0 7176 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_89
timestamp 1688980957
transform 1 0 9292 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_117
timestamp 1688980957
transform 1 0 11868 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_130
timestamp 1688980957
transform 1 0 13064 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_145
timestamp 1688980957
transform 1 0 14444 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_155
timestamp 1688980957
transform 1 0 15364 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_194
timestamp 1688980957
transform 1 0 18952 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_200
timestamp 1688980957
transform 1 0 19504 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_253
timestamp 1688980957
transform 1 0 24380 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1688980957
transform 1 0 2760 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 1932 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 2760 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1688980957
transform 1 0 2760 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform 1 0 3404 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 3128 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 3312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 2300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 1748 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 3496 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 3772 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 3312 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1688980957
transform 1 0 1748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1688980957
transform 1 0 1932 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1688980957
transform 1 0 5428 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1688980957
transform 1 0 3404 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 3220 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 2760 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 3496 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 3036 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 2760 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 3312 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 1656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 1932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 2760 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 1932 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 2208 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input50
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input51
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input52
timestamp 1688980957
transform 1 0 1932 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input53
timestamp 1688980957
transform 1 0 3772 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input54
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input55
timestamp 1688980957
transform 1 0 2760 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input56
timestamp 1688980957
transform 1 0 4324 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input57
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input58
timestamp 1688980957
transform 1 0 2392 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input59
timestamp 1688980957
transform 1 0 3312 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input60
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input61
timestamp 1688980957
transform 1 0 4324 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input62
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input63
timestamp 1688980957
transform 1 0 2392 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input64
timestamp 1688980957
transform 1 0 2944 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input65 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input66
timestamp 1688980957
transform 1 0 3864 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input67
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input68
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input69
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input70
timestamp 1688980957
transform 1 0 2300 0 -1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input71
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input72
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input73
timestamp 1688980957
transform 1 0 2392 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input74
timestamp 1688980957
transform 1 0 1932 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input75
timestamp 1688980957
transform 1 0 2760 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input76
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1688980957
transform 1 0 2760 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input78
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input80
timestamp 1688980957
transform 1 0 4324 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  input81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20424 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input82
timestamp 1688980957
transform 1 0 23736 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1688980957
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1688980957
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input85
timestamp 1688980957
transform 1 0 19688 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1688980957
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1688980957
transform 1 0 20884 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input88
timestamp 1688980957
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1688980957
transform 1 0 24196 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input90
timestamp 1688980957
transform 1 0 19688 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 1688980957
transform 1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  input92
timestamp 1688980957
transform 1 0 20608 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  input93 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20608 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  input94
timestamp 1688980957
transform 1 0 22448 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  input95
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  input96
timestamp 1688980957
transform 1 0 22632 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input97
timestamp 1688980957
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input98
timestamp 1688980957
transform 1 0 21988 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input99
timestamp 1688980957
transform 1 0 22632 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input100
timestamp 1688980957
transform 1 0 19320 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input102 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1748 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1688980957
transform 1 0 2300 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1688980957
transform 1 0 3312 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1688980957
transform 1 0 3864 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input107
timestamp 1688980957
transform 1 0 4140 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input108
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1688980957
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input110
timestamp 1688980957
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input111
timestamp 1688980957
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input112
timestamp 1688980957
transform 1 0 4232 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 1688980957
transform 1 0 1748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input114
timestamp 1688980957
transform 1 0 1472 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1688980957
transform 1 0 1840 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input116
timestamp 1688980957
transform 1 0 2208 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input117
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input118
timestamp 1688980957
transform 1 0 2760 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1688980957
transform 1 0 3128 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input120
timestamp 1688980957
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1688980957
transform 1 0 4508 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1688980957
transform 1 0 5060 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input128
timestamp 1688980957
transform 1 0 5336 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input129
timestamp 1688980957
transform 1 0 5888 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1688980957
transform 1 0 7360 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1688980957
transform 1 0 6440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1688980957
transform 1 0 6716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1688980957
transform 1 0 6992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1688980957
transform 1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1688980957
transform 1 0 3864 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input137
timestamp 1688980957
transform 1 0 24196 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input138
timestamp 1688980957
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1688980957
transform 1 0 22816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input141
timestamp 1688980957
transform 1 0 22080 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input142
timestamp 1688980957
transform 1 0 21160 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input143
timestamp 1688980957
transform 1 0 23000 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input144
timestamp 1688980957
transform 1 0 23276 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input145
timestamp 1688980957
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input146
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input147
timestamp 1688980957
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input148
timestamp 1688980957
transform 1 0 23736 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1688980957
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input150
timestamp 1688980957
transform 1 0 22264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input151
timestamp 1688980957
transform 1 0 18768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input152
timestamp 1688980957
transform 1 0 23828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input153
timestamp 1688980957
transform 1 0 9936 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input154
timestamp 1688980957
transform 1 0 10304 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input155
timestamp 1688980957
transform 1 0 10672 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1688980957
transform 1 0 11040 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input157
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input158
timestamp 1688980957
transform 1 0 11592 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input159
timestamp 1688980957
transform 1 0 11868 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input160
timestamp 1688980957
transform 1 0 12052 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input161
timestamp 1688980957
transform 1 0 12328 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input162
timestamp 1688980957
transform 1 0 12696 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input163
timestamp 1688980957
transform 1 0 12972 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input164
timestamp 1688980957
transform 1 0 14076 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input165
timestamp 1688980957
transform 1 0 13616 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input166
timestamp 1688980957
transform 1 0 14628 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input167
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input168
timestamp 1688980957
transform 1 0 14352 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input169
timestamp 1688980957
transform 1 0 14628 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input170
timestamp 1688980957
transform 1 0 14996 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input171
timestamp 1688980957
transform 1 0 15364 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input172
timestamp 1688980957
transform 1 0 15456 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input173
timestamp 1688980957
transform 1 0 15824 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input174
timestamp 1688980957
transform 1 0 17296 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input175
timestamp 1688980957
transform 1 0 17020 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input176
timestamp 1688980957
transform 1 0 19596 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input177
timestamp 1688980957
transform 1 0 18584 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input178
timestamp 1688980957
transform 1 0 18584 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input179
timestamp 1688980957
transform 1 0 20332 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input180
timestamp 1688980957
transform 1 0 16192 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input181
timestamp 1688980957
transform 1 0 16652 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input182
timestamp 1688980957
transform 1 0 16560 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input183
timestamp 1688980957
transform 1 0 17572 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input184
timestamp 1688980957
transform 1 0 17848 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input185
timestamp 1688980957
transform 1 0 18124 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input186
timestamp 1688980957
transform 1 0 18400 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input187
timestamp 1688980957
transform 1 0 18676 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input188
timestamp 1688980957
transform 1 0 24012 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  inst_clk_buf
timestamp 1688980957
transform 1 0 19228 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._0_
timestamp 1688980957
transform 1 0 23920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._1_
timestamp 1688980957
transform 1 0 22172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._2_
timestamp 1688980957
transform 1 0 22448 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._3_
timestamp 1688980957
transform 1 0 22356 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 20056 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 22632 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 22356 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._2_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19412 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._3_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19596 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19412 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18400 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19688 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 21252 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 22448 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20516 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22172 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 22816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 23276 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 24196 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 23092 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22356 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 23276 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 23368 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 24104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22448 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23092 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 20700 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 20976 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 22172 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 19136 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 22172 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 22908 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 22172 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21252 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22448 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 22448 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23000 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 23184 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22724 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 23368 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22632 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23092 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 20608 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 21528 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 21160 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19688 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 18216 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 20608 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 19044 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19320 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 20056 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 19688 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19780 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 22264 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23184 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23276 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 22540 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 22264 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21068 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22264 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 20516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 21528 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 21160 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19504 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20792 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 18492 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 20608 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 17664 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 18032 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19688 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 19964 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20056 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 22540 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 22356 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 22172 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21160 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22816 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18676 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 19136 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18124 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 19320 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 19964 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19780 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18584 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19688 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 19964 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 17664 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 19320 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 22080 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20424 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 23460 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23552 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22540 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23000 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18676 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 19412 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 19044 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18124 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19412 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 21160 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20884 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 20792 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19596 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 20240 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 22356 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19596 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 17480 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 22172 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20792 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21804 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23184 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 23644 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23460 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 21436 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 22080 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20056 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 19504 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17940 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19780 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 18124 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 17572 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19596 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 20148 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 19688 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18676 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19872 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 22172 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20792 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21896 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 20148 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 21068 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20700 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19688 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21344 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 18400 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 19412 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19044 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18032 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19688 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 19228 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 20056 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 23092 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18952 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 20516 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19320 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18676 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20976 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 19872 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 21344 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 20148 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20700 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21620 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 23092 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 23644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 22264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23000 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 18032 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 20792 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 23092 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 21528 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18676 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 19320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 18676 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 21160 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 20516 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 23092 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20240 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 22172 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21252 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 17572 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 19136 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 17940 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 20516 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18584 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 18032 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17296 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 19688 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 19964 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 20148 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20240 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18584 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 17940 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17664 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19412 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20976 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 20516 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 18032 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 22816 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 22448 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 23092 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 17480 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 22632 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 22908 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 23184 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22632 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22356 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 21712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 21252 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 18584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 23184 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22080 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23828 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit1
timestamp 1688980957
transform 1 0 11684 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit2
timestamp 1688980957
transform 1 0 2024 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit3
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit4
timestamp 1688980957
transform 1 0 6992 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit5
timestamp 1688980957
transform 1 0 9200 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit6
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit7
timestamp 1688980957
transform 1 0 12604 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit8
timestamp 1688980957
transform 1 0 9016 0 -1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit9
timestamp 1688980957
transform 1 0 9752 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit10
timestamp 1688980957
transform 1 0 4140 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit11
timestamp 1688980957
transform 1 0 4876 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit12
timestamp 1688980957
transform 1 0 5520 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit13
timestamp 1688980957
transform 1 0 6072 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit14
timestamp 1688980957
transform 1 0 9476 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit15
timestamp 1688980957
transform 1 0 9936 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit16
timestamp 1688980957
transform 1 0 4876 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit17
timestamp 1688980957
transform 1 0 4876 0 -1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit18
timestamp 1688980957
transform 1 0 4876 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit19
timestamp 1688980957
transform 1 0 5520 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit20
timestamp 1688980957
transform 1 0 4876 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit21
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit22
timestamp 1688980957
transform 1 0 11592 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit23
timestamp 1688980957
transform 1 0 12236 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit24
timestamp 1688980957
transform 1 0 10764 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit25
timestamp 1688980957
transform 1 0 11684 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit26
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit27
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit28
timestamp 1688980957
transform 1 0 9752 0 1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit29
timestamp 1688980957
transform 1 0 10028 0 -1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit30
timestamp 1688980957
transform 1 0 12604 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit31
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit0
timestamp 1688980957
transform 1 0 12420 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit1
timestamp 1688980957
transform 1 0 12880 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit2
timestamp 1688980957
transform 1 0 3128 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit3
timestamp 1688980957
transform 1 0 3772 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit4
timestamp 1688980957
transform 1 0 12236 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit5
timestamp 1688980957
transform 1 0 12696 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit6
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit7
timestamp 1688980957
transform 1 0 18032 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit8
timestamp 1688980957
transform 1 0 10948 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit9
timestamp 1688980957
transform 1 0 11868 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit10
timestamp 1688980957
transform 1 0 2392 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit11
timestamp 1688980957
transform 1 0 3220 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit12
timestamp 1688980957
transform 1 0 7452 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit13
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit14
timestamp 1688980957
transform 1 0 12696 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit15
timestamp 1688980957
transform 1 0 14076 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit16
timestamp 1688980957
transform 1 0 9752 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit17
timestamp 1688980957
transform 1 0 10856 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit18
timestamp 1688980957
transform 1 0 2300 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit19
timestamp 1688980957
transform 1 0 4600 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit20
timestamp 1688980957
transform 1 0 7268 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit21
timestamp 1688980957
transform 1 0 8004 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit22
timestamp 1688980957
transform 1 0 13340 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit23
timestamp 1688980957
transform 1 0 14536 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit24
timestamp 1688980957
transform 1 0 10764 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit25
timestamp 1688980957
transform 1 0 11776 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit26
timestamp 1688980957
transform 1 0 2300 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit27
timestamp 1688980957
transform 1 0 3312 0 -1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit28
timestamp 1688980957
transform 1 0 7452 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit29
timestamp 1688980957
transform 1 0 9016 0 -1 42432
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit30
timestamp 1688980957
transform 1 0 12604 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit31
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit0
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit1
timestamp 1688980957
transform 1 0 11868 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit2
timestamp 1688980957
transform 1 0 4048 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit3
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit4
timestamp 1688980957
transform 1 0 9384 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit5
timestamp 1688980957
transform 1 0 10212 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit6
timestamp 1688980957
transform 1 0 14536 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit7
timestamp 1688980957
transform 1 0 15180 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit8
timestamp 1688980957
transform 1 0 12604 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit9
timestamp 1688980957
transform 1 0 14168 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit10
timestamp 1688980957
transform 1 0 3772 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit11
timestamp 1688980957
transform 1 0 4232 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit12
timestamp 1688980957
transform 1 0 11224 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit13
timestamp 1688980957
transform 1 0 12144 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit14
timestamp 1688980957
transform 1 0 15180 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit15
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit16
timestamp 1688980957
transform 1 0 15180 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit17
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit18
timestamp 1688980957
transform 1 0 6624 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit19
timestamp 1688980957
transform 1 0 7544 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit20
timestamp 1688980957
transform 1 0 4416 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit21
timestamp 1688980957
transform 1 0 5796 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit22
timestamp 1688980957
transform 1 0 14168 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit23
timestamp 1688980957
transform 1 0 14720 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit24
timestamp 1688980957
transform 1 0 14996 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit25
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit26
timestamp 1688980957
transform 1 0 7360 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit27
timestamp 1688980957
transform 1 0 8188 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit28
timestamp 1688980957
transform 1 0 4692 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit29
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit30
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit31
timestamp 1688980957
transform 1 0 11224 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit0
timestamp 1688980957
transform 1 0 15180 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit1
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit2
timestamp 1688980957
transform 1 0 6808 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit3
timestamp 1688980957
transform 1 0 8188 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit4
timestamp 1688980957
transform 1 0 2392 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit5
timestamp 1688980957
transform 1 0 4048 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit6
timestamp 1688980957
transform 1 0 9568 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit7
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit8
timestamp 1688980957
transform 1 0 14996 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit9
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit10
timestamp 1688980957
transform 1 0 7176 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit11
timestamp 1688980957
transform 1 0 8004 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit12
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit13
timestamp 1688980957
transform 1 0 4232 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit14
timestamp 1688980957
transform 1 0 8648 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit15
timestamp 1688980957
transform 1 0 9476 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit16
timestamp 1688980957
transform 1 0 11500 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit17
timestamp 1688980957
transform 1 0 12144 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit18
timestamp 1688980957
transform 1 0 2300 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit19
timestamp 1688980957
transform 1 0 3036 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit20
timestamp 1688980957
transform 1 0 9844 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit21
timestamp 1688980957
transform 1 0 10764 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit22
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit23
timestamp 1688980957
transform 1 0 15456 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit24
timestamp 1688980957
transform 1 0 12144 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit25
timestamp 1688980957
transform 1 0 12696 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit26
timestamp 1688980957
transform 1 0 2300 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit27
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit28
timestamp 1688980957
transform 1 0 9752 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit29
timestamp 1688980957
transform 1 0 10028 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit30
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit31
timestamp 1688980957
transform 1 0 17020 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit0
timestamp 1688980957
transform 1 0 15180 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit1
timestamp 1688980957
transform 1 0 17112 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit2
timestamp 1688980957
transform 1 0 4876 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit3
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit4
timestamp 1688980957
transform 1 0 2668 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit5
timestamp 1688980957
transform 1 0 4048 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit6
timestamp 1688980957
transform 1 0 9108 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit7
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit8
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit9
timestamp 1688980957
transform 1 0 18032 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit10
timestamp 1688980957
transform 1 0 6440 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit11
timestamp 1688980957
transform 1 0 7084 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit12
timestamp 1688980957
transform 1 0 2300 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit13
timestamp 1688980957
transform 1 0 3128 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit14
timestamp 1688980957
transform 1 0 7452 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit15
timestamp 1688980957
transform 1 0 8372 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit16
timestamp 1688980957
transform 1 0 15088 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit17
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit18
timestamp 1688980957
transform 1 0 6992 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit19
timestamp 1688980957
transform 1 0 6992 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit20
timestamp 1688980957
transform 1 0 3496 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit21
timestamp 1688980957
transform 1 0 4048 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit22
timestamp 1688980957
transform 1 0 7176 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit23
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit24
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit25
timestamp 1688980957
transform 1 0 15456 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit26
timestamp 1688980957
transform 1 0 5704 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit27
timestamp 1688980957
transform 1 0 6532 0 -1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit28
timestamp 1688980957
transform 1 0 4324 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit29
timestamp 1688980957
transform 1 0 4876 0 -1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit30
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit31
timestamp 1688980957
transform 1 0 12696 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit0
timestamp 1688980957
transform 1 0 14720 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit1
timestamp 1688980957
transform 1 0 17112 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit2
timestamp 1688980957
transform 1 0 1656 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit3
timestamp 1688980957
transform 1 0 2208 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit4
timestamp 1688980957
transform 1 0 1656 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit5
timestamp 1688980957
transform 1 0 2024 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit6
timestamp 1688980957
transform 1 0 6072 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit7
timestamp 1688980957
transform 1 0 7452 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit8
timestamp 1688980957
transform 1 0 10120 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit9
timestamp 1688980957
transform 1 0 10856 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit10
timestamp 1688980957
transform 1 0 4048 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit11
timestamp 1688980957
transform 1 0 7360 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit12
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit13
timestamp 1688980957
transform 1 0 1656 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit14
timestamp 1688980957
transform 1 0 1932 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit15
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit16
timestamp 1688980957
transform 1 0 14628 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit17
timestamp 1688980957
transform 1 0 16008 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit18
timestamp 1688980957
transform 1 0 1656 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit19
timestamp 1688980957
transform 1 0 2116 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit20
timestamp 1688980957
transform 1 0 1748 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit21
timestamp 1688980957
transform 1 0 2208 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit22
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit23
timestamp 1688980957
transform 1 0 7452 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit24
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit25
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit26
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit27
timestamp 1688980957
transform 1 0 5888 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit28
timestamp 1688980957
transform 1 0 3680 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit29
timestamp 1688980957
transform 1 0 4232 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit30
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit31
timestamp 1688980957
transform 1 0 8648 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit0
timestamp 1688980957
transform 1 0 7268 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit1
timestamp 1688980957
transform 1 0 7268 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit2
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit3
timestamp 1688980957
transform 1 0 14444 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit4
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit5
timestamp 1688980957
transform 1 0 14076 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit6
timestamp 1688980957
transform 1 0 17020 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit7
timestamp 1688980957
transform 1 0 3864 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit8
timestamp 1688980957
transform 1 0 4784 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit9
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit10
timestamp 1688980957
transform 1 0 9108 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit11
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit12
timestamp 1688980957
transform 1 0 11684 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit13
timestamp 1688980957
transform 1 0 14996 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit14
timestamp 1688980957
transform 1 0 17020 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit15
timestamp 1688980957
transform 1 0 17664 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit16
timestamp 1688980957
transform 1 0 9108 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit17
timestamp 1688980957
transform 1 0 10212 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit18
timestamp 1688980957
transform 1 0 2116 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit19
timestamp 1688980957
transform 1 0 2208 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit20
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit21
timestamp 1688980957
transform 1 0 9476 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit22
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit23
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit24
timestamp 1688980957
transform 1 0 9752 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit25
timestamp 1688980957
transform 1 0 10764 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit26
timestamp 1688980957
transform 1 0 4876 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit27
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit28
timestamp 1688980957
transform 1 0 2024 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit29
timestamp 1688980957
transform 1 0 2392 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit30
timestamp 1688980957
transform 1 0 3312 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit31
timestamp 1688980957
transform 1 0 4048 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit0
timestamp 1688980957
transform 1 0 9200 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit1
timestamp 1688980957
transform 1 0 9936 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit2
timestamp 1688980957
transform 1 0 10028 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit3
timestamp 1688980957
transform 1 0 4600 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit4
timestamp 1688980957
transform 1 0 5060 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit5
timestamp 1688980957
transform 1 0 6532 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit6
timestamp 1688980957
transform 1 0 6992 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit7
timestamp 1688980957
transform 1 0 7452 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit8
timestamp 1688980957
transform 1 0 9476 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit9
timestamp 1688980957
transform 1 0 15456 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit10
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit11
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit12
timestamp 1688980957
transform 1 0 8924 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit13
timestamp 1688980957
transform 1 0 9384 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit14
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit15
timestamp 1688980957
transform 1 0 5704 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit16
timestamp 1688980957
transform 1 0 12052 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit17
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit18
timestamp 1688980957
transform 1 0 12604 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit19
timestamp 1688980957
transform 1 0 14076 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit20
timestamp 1688980957
transform 1 0 9660 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit21
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit22
timestamp 1688980957
transform 1 0 4600 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit23
timestamp 1688980957
transform 1 0 6256 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit24
timestamp 1688980957
transform 1 0 7452 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit25
timestamp 1688980957
transform 1 0 8096 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit26
timestamp 1688980957
transform 1 0 12144 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit27
timestamp 1688980957
transform 1 0 12604 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit28
timestamp 1688980957
transform 1 0 12696 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit29
timestamp 1688980957
transform 1 0 12604 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit30
timestamp 1688980957
transform 1 0 4692 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit31
timestamp 1688980957
transform 1 0 5244 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit0
timestamp 1688980957
transform 1 0 19412 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit1
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit2
timestamp 1688980957
transform 1 0 22080 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit3
timestamp 1688980957
transform 1 0 19780 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit4
timestamp 1688980957
transform 1 0 22816 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit5
timestamp 1688980957
transform 1 0 22724 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit6
timestamp 1688980957
transform 1 0 22632 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit7
timestamp 1688980957
transform 1 0 22816 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit8
timestamp 1688980957
transform 1 0 8648 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit9
timestamp 1688980957
transform 1 0 9292 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit10
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit11
timestamp 1688980957
transform 1 0 1472 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit12
timestamp 1688980957
transform 1 0 10028 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit13
timestamp 1688980957
transform 1 0 10856 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit14
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit15
timestamp 1688980957
transform 1 0 14076 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit16
timestamp 1688980957
transform 1 0 7544 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit17
timestamp 1688980957
transform 1 0 8096 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit18
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit19
timestamp 1688980957
transform 1 0 1472 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit20
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit21
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit22
timestamp 1688980957
transform 1 0 1840 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit23
timestamp 1688980957
transform 1 0 2300 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit24
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit25
timestamp 1688980957
transform 1 0 1748 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit26
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit27
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit28
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit29
timestamp 1688980957
transform 1 0 1748 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit30
timestamp 1688980957
transform 1 0 5796 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit31
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit0
timestamp 1688980957
transform 1 0 17204 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit1
timestamp 1688980957
transform 1 0 18768 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit2
timestamp 1688980957
transform 1 0 18032 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit3
timestamp 1688980957
transform 1 0 19596 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit4
timestamp 1688980957
transform 1 0 17204 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit5
timestamp 1688980957
transform 1 0 22632 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit6
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit7
timestamp 1688980957
transform 1 0 23184 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit8
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit9
timestamp 1688980957
transform 1 0 21344 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit10
timestamp 1688980957
transform 1 0 17756 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit11
timestamp 1688980957
transform 1 0 19504 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit12
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit13
timestamp 1688980957
transform 1 0 22448 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit14
timestamp 1688980957
transform 1 0 18032 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit15
timestamp 1688980957
transform 1 0 19872 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit16
timestamp 1688980957
transform 1 0 21160 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit17
timestamp 1688980957
transform 1 0 22816 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit18
timestamp 1688980957
transform 1 0 20240 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit19
timestamp 1688980957
transform 1 0 17940 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit20
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit21
timestamp 1688980957
transform 1 0 20884 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit22
timestamp 1688980957
transform 1 0 19688 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit23
timestamp 1688980957
transform 1 0 17572 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit24
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit25
timestamp 1688980957
transform 1 0 20700 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit26
timestamp 1688980957
transform 1 0 22816 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit27
timestamp 1688980957
transform 1 0 22724 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit28
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit29
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit30
timestamp 1688980957
transform 1 0 22448 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit31
timestamp 1688980957
transform 1 0 19780 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit24
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit25
timestamp 1688980957
transform 1 0 19504 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit26
timestamp 1688980957
transform 1 0 22264 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit27
timestamp 1688980957
transform 1 0 20884 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit28
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit29
timestamp 1688980957
transform 1 0 19412 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit30
timestamp 1688980957
transform 1 0 22356 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit31
timestamp 1688980957
transform 1 0 20884 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._32_
timestamp 1688980957
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._33_
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._34_
timestamp 1688980957
transform 1 0 3404 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._35_
timestamp 1688980957
transform 1 0 3772 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._36_
timestamp 1688980957
transform 1 0 4324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._37_
timestamp 1688980957
transform 1 0 4416 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._38_
timestamp 1688980957
transform 1 0 4600 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._39_
timestamp 1688980957
transform 1 0 5244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._40_
timestamp 1688980957
transform 1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._41_
timestamp 1688980957
transform 1 0 11408 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._42_
timestamp 1688980957
transform 1 0 11592 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._43_
timestamp 1688980957
transform 1 0 11684 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._44_
timestamp 1688980957
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._45_
timestamp 1688980957
transform 1 0 13156 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._46_
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._47_
timestamp 1688980957
transform 1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0_395 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15732 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7176 0 1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1_396
timestamp 1688980957
transform 1 0 6900 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2_397
timestamp 1688980957
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3_398
timestamp 1688980957
transform 1 0 15548 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3
timestamp 1688980957
transform 1 0 14444 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0_399
timestamp 1688980957
transform 1 0 16376 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0
timestamp 1688980957
transform 1 0 15364 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1_400
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1
timestamp 1688980957
transform 1 0 7728 0 -1 22848
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2_401
timestamp 1688980957
transform 1 0 6532 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2
timestamp 1688980957
transform 1 0 6072 0 1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3
timestamp 1688980957
transform 1 0 11500 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3_402
timestamp 1688980957
transform 1 0 12512 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0_403
timestamp 1688980957
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0
timestamp 1688980957
transform 1 0 12788 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1_404
timestamp 1688980957
transform 1 0 4508 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2_405
timestamp 1688980957
transform 1 0 13432 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2
timestamp 1688980957
transform 1 0 12052 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3_409
timestamp 1688980957
transform 1 0 18032 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3
timestamp 1688980957
transform 1 0 17020 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I0
timestamp 1688980957
transform 1 0 11868 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I1
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I2
timestamp 1688980957
transform 1 0 10120 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I3
timestamp 1688980957
transform 1 0 15272 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I0
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I1
timestamp 1688980957
transform 1 0 3220 0 -1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I2
timestamp 1688980957
transform 1 0 9660 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I3
timestamp 1688980957
transform 1 0 17204 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I0
timestamp 1688980957
transform 1 0 11592 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I1
timestamp 1688980957
transform 1 0 4416 0 -1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I2
timestamp 1688980957
transform 1 0 9476 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I3
timestamp 1688980957
transform 1 0 15272 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I0
timestamp 1688980957
transform 1 0 13524 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I1
timestamp 1688980957
transform 1 0 3956 0 -1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I2
timestamp 1688980957
transform 1 0 11592 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I3
timestamp 1688980957
transform 1 0 16008 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0_406
timestamp 1688980957
transform 1 0 11776 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0
timestamp 1688980957
transform 1 0 11316 0 1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1_407
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2_408
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2
timestamp 1688980957
transform 1 0 9844 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3_394
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3
timestamp 1688980957
transform 1 0 13432 0 -1 16320
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG0
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG1
timestamp 1688980957
transform 1 0 4600 0 1 30464
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG2
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG3
timestamp 1688980957
transform 1 0 9752 0 -1 22848
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG4
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG5
timestamp 1688980957
transform 1 0 5336 0 1 15232
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG6
timestamp 1688980957
transform 1 0 6348 0 1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG7
timestamp 1688980957
transform 1 0 11960 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG0
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG1
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG2
timestamp 1688980957
transform 1 0 8280 0 -1 38080
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG3
timestamp 1688980957
transform 1 0 13616 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG4
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG5
timestamp 1688980957
transform 1 0 2944 0 -1 36992
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG6
timestamp 1688980957
transform 1 0 7820 0 -1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG7
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG8
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG9
timestamp 1688980957
transform 1 0 3036 0 -1 40256
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG10
timestamp 1688980957
transform 1 0 8464 0 -1 40256
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG11
timestamp 1688980957
transform 1 0 13524 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG12
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG13
timestamp 1688980957
transform 1 0 2944 0 -1 39168
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG14
timestamp 1688980957
transform 1 0 8372 0 -1 39168
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG15
timestamp 1688980957
transform 1 0 11960 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG0
timestamp 1688980957
transform 1 0 9108 0 1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG1
timestamp 1688980957
transform 1 0 1564 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG2
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG3
timestamp 1688980957
transform 1 0 13892 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG0
timestamp 1688980957
transform 1 0 7820 0 -1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG1
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG2
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG3
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG4
timestamp 1688980957
transform 1 0 1564 0 1 23936
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG5
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG6
timestamp 1688980957
transform 1 0 1564 0 -1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG7
timestamp 1688980957
transform 1 0 7176 0 1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG0
timestamp 1688980957
transform 1 0 9200 0 -1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG1
timestamp 1688980957
transform 1 0 4600 0 -1 34816
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG2
timestamp 1688980957
transform 1 0 11592 0 -1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG3
timestamp 1688980957
transform 1 0 13892 0 -1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG0
timestamp 1688980957
transform 1 0 11040 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG1
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG2
timestamp 1688980957
transform 1 0 7728 0 -1 30464
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG3
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG4
timestamp 1688980957
transform 1 0 12972 0 -1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG5
timestamp 1688980957
transform 1 0 4600 0 -1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG6
timestamp 1688980957
transform 1 0 7544 0 -1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG7
timestamp 1688980957
transform 1 0 14260 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG0
timestamp 1688980957
transform 1 0 9476 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG1
timestamp 1688980957
transform 1 0 2668 0 -1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG2
timestamp 1688980957
transform 1 0 9292 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG3
timestamp 1688980957
transform 1 0 13616 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG0
timestamp 1688980957
transform 1 0 10488 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG1
timestamp 1688980957
transform 1 0 5520 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG2
timestamp 1688980957
transform 1 0 1748 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG3
timestamp 1688980957
transform 1 0 3680 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG4
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG5
timestamp 1688980957
transform 1 0 2024 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG6
timestamp 1688980957
transform 1 0 1748 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG7
timestamp 1688980957
transform 1 0 7544 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb0
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb1
timestamp 1688980957
transform 1 0 5428 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb2
timestamp 1688980957
transform 1 0 1656 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb3
timestamp 1688980957
transform 1 0 3312 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb4
timestamp 1688980957
transform 1 0 14628 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb5
timestamp 1688980957
transform 1 0 1748 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb6
timestamp 1688980957
transform 1 0 2024 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb7
timestamp 1688980957
transform 1 0 7544 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG0
timestamp 1688980957
transform 1 0 14168 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG1
timestamp 1688980957
transform 1 0 6072 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG2
timestamp 1688980957
transform 1 0 4140 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG3
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG4
timestamp 1688980957
transform 1 0 15640 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG5
timestamp 1688980957
transform 1 0 6900 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG6
timestamp 1688980957
transform 1 0 3772 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG7
timestamp 1688980957
transform 1 0 9384 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG8
timestamp 1688980957
transform 1 0 15456 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG9
timestamp 1688980957
transform 1 0 7636 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG10
timestamp 1688980957
transform 1 0 3956 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG11
timestamp 1688980957
transform 1 0 9016 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG0
timestamp 1688980957
transform 1 0 16468 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG1
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG2
timestamp 1688980957
transform 1 0 3864 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG3
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG4
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG5
timestamp 1688980957
transform 1 0 4968 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG6
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG7
timestamp 1688980957
transform 1 0 9384 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG8
timestamp 1688980957
transform 1 0 16376 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG9
timestamp 1688980957
transform 1 0 6716 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG10
timestamp 1688980957
transform 1 0 2024 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG11
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG12
timestamp 1688980957
transform 1 0 15364 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG13
timestamp 1688980957
transform 1 0 6716 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG14
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG15
timestamp 1688980957
transform 1 0 7820 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 11408 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 11868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 11592 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 9660 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 9476 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 7176 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 7360 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 7912 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 6900 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 4324 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 4968 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 10212 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 9936 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 9200 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 9568 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 9292 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 7544 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 7544 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 17112 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 17388 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17296 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17112 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 15364 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 15640 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 16744 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 17664 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 18032 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16192 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17296 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 6808 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 6900 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 6440 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 7544 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 4324 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 4324 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 12236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 12420 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 13064 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 11868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 11960 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 9752 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 9476 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 18492 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18308 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18584 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 16376 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_0._0_
timestamp 1688980957
transform 1 0 4692 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_1._0_
timestamp 1688980957
transform 1 0 5704 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_2._0_
timestamp 1688980957
transform 1 0 6532 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_3._0_
timestamp 1688980957
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_4._0_
timestamp 1688980957
transform 1 0 6440 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_5._0_
timestamp 1688980957
transform 1 0 6716 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_6._0_
timestamp 1688980957
transform 1 0 8004 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_7._0_
timestamp 1688980957
transform 1 0 7912 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_8._0_
timestamp 1688980957
transform 1 0 7728 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_9._0_
timestamp 1688980957
transform 1 0 8004 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_10._0_
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_11._0_
timestamp 1688980957
transform 1 0 9476 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_0._0_
timestamp 1688980957
transform 1 0 6992 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_1._0_
timestamp 1688980957
transform 1 0 6624 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_2._0_
timestamp 1688980957
transform 1 0 6440 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_3._0_
timestamp 1688980957
transform 1 0 6808 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_4._0_
timestamp 1688980957
transform 1 0 7176 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_5._0_
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_6._0_
timestamp 1688980957
transform 1 0 7544 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_7._0_
timestamp 1688980957
transform 1 0 7912 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_8._0_
timestamp 1688980957
transform 1 0 8280 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_9._0_
timestamp 1688980957
transform 1 0 8648 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_10._0_
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_11._0_
timestamp 1688980957
transform 1 0 9200 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output189
timestamp 1688980957
transform 1 0 23460 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output190
timestamp 1688980957
transform 1 0 23460 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output191
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output192
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output193
timestamp 1688980957
transform 1 0 23552 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output194
timestamp 1688980957
transform 1 0 23920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output195
timestamp 1688980957
transform 1 0 23644 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output196
timestamp 1688980957
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output197
timestamp 1688980957
transform 1 0 24012 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output198
timestamp 1688980957
transform 1 0 24012 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output199
timestamp 1688980957
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output200
timestamp 1688980957
transform 1 0 23368 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1688980957
transform 1 0 24196 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output202
timestamp 1688980957
transform 1 0 23460 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output203
timestamp 1688980957
transform 1 0 23552 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1688980957
transform 1 0 23184 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output205
timestamp 1688980957
transform 1 0 23736 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output206
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output207
timestamp 1688980957
transform 1 0 23736 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output208
timestamp 1688980957
transform 1 0 23828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1688980957
transform 1 0 23460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output210
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1688980957
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output212
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output213
timestamp 1688980957
transform 1 0 23552 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output214
timestamp 1688980957
transform 1 0 23920 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1688980957
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output216
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1688980957
transform 1 0 24196 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output218
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output219
timestamp 1688980957
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output220
timestamp 1688980957
transform 1 0 23368 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1688980957
transform 1 0 23368 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1688980957
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output223
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1688980957
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output225
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output226
timestamp 1688980957
transform 1 0 23736 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output227
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output228
timestamp 1688980957
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output229
timestamp 1688980957
transform 1 0 24012 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1688980957
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output231
timestamp 1688980957
transform 1 0 24012 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output232
timestamp 1688980957
transform 1 0 24012 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1688980957
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output234
timestamp 1688980957
transform 1 0 24012 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1688980957
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output236
timestamp 1688980957
transform 1 0 24012 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output237
timestamp 1688980957
transform 1 0 23736 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output238
timestamp 1688980957
transform 1 0 23276 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output239
timestamp 1688980957
transform 1 0 24012 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output240
timestamp 1688980957
transform 1 0 22724 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output241
timestamp 1688980957
transform 1 0 23460 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output242
timestamp 1688980957
transform 1 0 21988 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1688980957
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output244
timestamp 1688980957
transform 1 0 23184 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output245
timestamp 1688980957
transform 1 0 22356 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output246
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output247
timestamp 1688980957
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output248
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output249
timestamp 1688980957
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output250
timestamp 1688980957
transform 1 0 24012 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output251
timestamp 1688980957
transform 1 0 23736 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output252
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output253
timestamp 1688980957
transform 1 0 20240 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output254
timestamp 1688980957
transform 1 0 23460 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output255
timestamp 1688980957
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output256
timestamp 1688980957
transform 1 0 21804 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output257
timestamp 1688980957
transform 1 0 23736 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output258
timestamp 1688980957
transform 1 0 22908 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output259
timestamp 1688980957
transform 1 0 23828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output260
timestamp 1688980957
transform 1 0 22632 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output261
timestamp 1688980957
transform 1 0 21436 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output262
timestamp 1688980957
transform 1 0 23184 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output263
timestamp 1688980957
transform 1 0 21160 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output264
timestamp 1688980957
transform 1 0 20792 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1688980957
transform 1 0 21344 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output266
timestamp 1688980957
transform 1 0 21804 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output267
timestamp 1688980957
transform 1 0 22356 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output268
timestamp 1688980957
transform 1 0 22908 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output269
timestamp 1688980957
transform 1 0 22080 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output270
timestamp 1688980957
transform 1 0 22540 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output271
timestamp 1688980957
transform 1 0 19688 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output272
timestamp 1688980957
transform 1 0 23092 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output273
timestamp 1688980957
transform 1 0 4600 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output274
timestamp 1688980957
transform 1 0 4048 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output275
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output276
timestamp 1688980957
transform 1 0 2392 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output277
timestamp 1688980957
transform 1 0 3496 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output278
timestamp 1688980957
transform 1 0 2944 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output279
timestamp 1688980957
transform 1 0 1748 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output280
timestamp 1688980957
transform 1 0 1656 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output281
timestamp 1688980957
transform 1 0 2208 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output282
timestamp 1688980957
transform 1 0 2576 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output283
timestamp 1688980957
transform 1 0 2760 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output284
timestamp 1688980957
transform 1 0 3128 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output285
timestamp 1688980957
transform 1 0 4324 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output286
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output287
timestamp 1688980957
transform 1 0 4140 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output288
timestamp 1688980957
transform 1 0 4048 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output289
timestamp 1688980957
transform 1 0 3312 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output290
timestamp 1688980957
transform 1 0 4968 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output291
timestamp 1688980957
transform 1 0 4600 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output292
timestamp 1688980957
transform 1 0 4968 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output293
timestamp 1688980957
transform 1 0 5520 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output294
timestamp 1688980957
transform 1 0 7728 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output295
timestamp 1688980957
transform 1 0 8280 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output296
timestamp 1688980957
transform 1 0 8924 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output297
timestamp 1688980957
transform 1 0 9384 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output298
timestamp 1688980957
transform 1 0 8280 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output299
timestamp 1688980957
transform 1 0 9384 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output300
timestamp 1688980957
transform 1 0 5888 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output301
timestamp 1688980957
transform 1 0 5520 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output302
timestamp 1688980957
transform 1 0 6440 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output303
timestamp 1688980957
transform 1 0 6624 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output304
timestamp 1688980957
transform 1 0 6992 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output305
timestamp 1688980957
transform 1 0 7360 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output306
timestamp 1688980957
transform 1 0 7544 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output307
timestamp 1688980957
transform 1 0 7360 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output308
timestamp 1688980957
transform 1 0 8280 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output309
timestamp 1688980957
transform 1 0 9568 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output310
timestamp 1688980957
transform 1 0 10488 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output311
timestamp 1688980957
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output312
timestamp 1688980957
transform 1 0 10856 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output313
timestamp 1688980957
transform 1 0 13248 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output314
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output315
timestamp 1688980957
transform 1 0 14628 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output316
timestamp 1688980957
transform 1 0 14444 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output317
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output318
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output319
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output320
timestamp 1688980957
transform 1 0 16100 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output321
timestamp 1688980957
transform 1 0 9936 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output322
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output323
timestamp 1688980957
transform 1 0 11684 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output324
timestamp 1688980957
transform 1 0 10488 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output325
timestamp 1688980957
transform 1 0 12512 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output326
timestamp 1688980957
transform 1 0 12236 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output327
timestamp 1688980957
transform 1 0 11040 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output328
timestamp 1688980957
transform 1 0 13616 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output329
timestamp 1688980957
transform 1 0 15548 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output330
timestamp 1688980957
transform 1 0 20056 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output331
timestamp 1688980957
transform 1 0 17204 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output332
timestamp 1688980957
transform 1 0 19504 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output333
timestamp 1688980957
transform 1 0 19596 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output334
timestamp 1688980957
transform 1 0 20148 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output335
timestamp 1688980957
transform 1 0 20700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output336
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output337
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output338
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output339
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output340
timestamp 1688980957
transform 1 0 18860 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output341
timestamp 1688980957
transform 1 0 18124 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output342
timestamp 1688980957
transform 1 0 17572 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output343
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output344
timestamp 1688980957
transform 1 0 18308 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  output345
timestamp 1688980957
transform 1 0 21528 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output346
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output347
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output348
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output349
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output350
timestamp 1688980957
transform 1 0 2116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output351
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output352
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output353
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output354
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output355
timestamp 1688980957
transform 1 0 3036 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output356
timestamp 1688980957
transform 1 0 2668 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output357
timestamp 1688980957
transform 1 0 1564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output358
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output359
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output360
timestamp 1688980957
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output361
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output362
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output363
timestamp 1688980957
transform 1 0 1472 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output364
timestamp 1688980957
transform 1 0 2116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output365
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output366
timestamp 1688980957
transform 1 0 1564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output367
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output368
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output369
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output370
timestamp 1688980957
transform 1 0 1564 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output371
timestamp 1688980957
transform 1 0 3496 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output372
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output373
timestamp 1688980957
transform 1 0 1564 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output374
timestamp 1688980957
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output375
timestamp 1688980957
transform 1 0 2668 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output376
timestamp 1688980957
transform 1 0 2116 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output377
timestamp 1688980957
transform 1 0 1564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output378
timestamp 1688980957
transform 1 0 2668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output379
timestamp 1688980957
transform 1 0 2116 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output380
timestamp 1688980957
transform 1 0 5704 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output381
timestamp 1688980957
transform 1 0 2300 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output382
timestamp 1688980957
transform 1 0 1472 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output383
timestamp 1688980957
transform 1 0 2852 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output384
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output385
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output386
timestamp 1688980957
transform 1 0 1564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output387
timestamp 1688980957
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output388
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output389
timestamp 1688980957
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output390
timestamp 1688980957
transform 1 0 1932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output391
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output392
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output393
timestamp 1688980957
transform 1 0 3956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 24840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 24840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 24840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 24840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 24840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 24840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 24840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 24840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 24840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 24840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 24840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 24840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 24840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 24840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 24840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 24840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 24840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 24840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 24840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 24840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 24840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 24840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 24840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 24840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 24840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 24840 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 24840 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 24840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 24840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 24840 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 24840 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 24840 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 24840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 24840 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 24840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 24840 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 24840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 24840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 24840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 24840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 24840 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 24840 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 24840 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 24840 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 24840 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 24840 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 24840 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 24840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 24840 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 24840 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 24840 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 24840 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 24840 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 24840 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 24840 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 24840 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 24840 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 24840 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 24840 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 24840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 24840 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 24840 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 24840 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 24840 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 24840 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 24840 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 24840 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 24840 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 24840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 24840 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 24840 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_0._0_
timestamp 1688980957
transform 1 0 16008 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_1._0_
timestamp 1688980957
transform 1 0 16376 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_2._0_
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_3._0_
timestamp 1688980957
transform 1 0 17020 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_4._0_
timestamp 1688980957
transform 1 0 17388 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_5._0_
timestamp 1688980957
transform 1 0 17756 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_6._0_
timestamp 1688980957
transform 1 0 18124 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_7._0_
timestamp 1688980957
transform 1 0 18492 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_8._0_
timestamp 1688980957
transform 1 0 18860 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_9._0_
timestamp 1688980957
transform 1 0 19228 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_10._0_
timestamp 1688980957
transform 1 0 18860 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_11._0_
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_0._0_
timestamp 1688980957
transform 1 0 16284 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_1._0_
timestamp 1688980957
transform 1 0 16008 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_2._0_
timestamp 1688980957
transform 1 0 17204 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_3._0_
timestamp 1688980957
transform 1 0 17480 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_4._0_
timestamp 1688980957
transform 1 0 17756 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_5._0_
timestamp 1688980957
transform 1 0 18032 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_6._0_
timestamp 1688980957
transform 1 0 18308 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_7._0_
timestamp 1688980957
transform 1 0 18584 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_8._0_
timestamp 1688980957
transform 1 0 18860 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_9._0_
timestamp 1688980957
transform 1 0 19228 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_10._0_
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_11._0_
timestamp 1688980957
transform 1 0 19412 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0._0_
timestamp 1688980957
transform 1 0 19780 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1._0_
timestamp 1688980957
transform 1 0 20056 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2._0_
timestamp 1688980957
transform 1 0 20424 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3._0_
timestamp 1688980957
transform 1 0 20424 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4._0_
timestamp 1688980957
transform 1 0 20792 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_inbuf_5._0_
timestamp 1688980957
transform 1 0 21804 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6._0_
timestamp 1688980957
transform 1 0 21436 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7._0_
timestamp 1688980957
transform 1 0 21804 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8._0_
timestamp 1688980957
transform 1 0 22172 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9._0_
timestamp 1688980957
transform 1 0 22632 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_10._0_
timestamp 1688980957
transform 1 0 22448 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_11._0_
timestamp 1688980957
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12._0_
timestamp 1688980957
transform 1 0 23460 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13._0_
timestamp 1688980957
transform 1 0 23460 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14._0_
timestamp 1688980957
transform 1 0 23368 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15._0_
timestamp 1688980957
transform 1 0 23368 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16._0_
timestamp 1688980957
transform 1 0 23644 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17._0_
timestamp 1688980957
transform 1 0 23184 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18._0_
timestamp 1688980957
transform 1 0 22724 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19._0_
timestamp 1688980957
transform 1 0 23184 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0._0_
timestamp 1688980957
transform 1 0 19964 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1._0_
timestamp 1688980957
transform 1 0 20240 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_2._0_
timestamp 1688980957
transform 1 0 20516 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3._0_
timestamp 1688980957
transform 1 0 20700 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4._0_
timestamp 1688980957
transform 1 0 20976 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5._0_
timestamp 1688980957
transform 1 0 21160 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6._0_
timestamp 1688980957
transform 1 0 20148 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7._0_
timestamp 1688980957
transform 1 0 21160 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8._0_
timestamp 1688980957
transform 1 0 22356 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9._0_
timestamp 1688980957
transform 1 0 22540 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10._0_
timestamp 1688980957
transform 1 0 21068 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11._0_
timestamp 1688980957
transform 1 0 22448 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12._0_
timestamp 1688980957
transform 1 0 19872 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13._0_
timestamp 1688980957
transform 1 0 23184 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14._0_
timestamp 1688980957
transform 1 0 23184 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15._0_
timestamp 1688980957
transform 1 0 23736 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16._0_
timestamp 1688980957
transform 1 0 23736 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17._0_
timestamp 1688980957
transform 1 0 23736 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18._0_
timestamp 1688980957
transform 1 0 23460 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19._0_
timestamp 1688980957
transform 1 0 23644 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 3680 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 8832 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 13984 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 19136 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 24288 0 -1 43520
box -38 -48 130 592
<< labels >>
flabel metal3 s 25840 9528 26000 9648 0 FreeSans 480 0 0 0 Config_accessC_bit0
port 0 nsew signal tristate
flabel metal3 s 25840 10072 26000 10192 0 FreeSans 480 0 0 0 Config_accessC_bit1
port 1 nsew signal tristate
flabel metal3 s 25840 10616 26000 10736 0 FreeSans 480 0 0 0 Config_accessC_bit2
port 2 nsew signal tristate
flabel metal3 s 25840 11160 26000 11280 0 FreeSans 480 0 0 0 Config_accessC_bit3
port 3 nsew signal tristate
flabel metal3 s 0 18232 160 18352 0 FreeSans 480 0 0 0 E1END[0]
port 4 nsew signal input
flabel metal3 s 0 18504 160 18624 0 FreeSans 480 0 0 0 E1END[1]
port 5 nsew signal input
flabel metal3 s 0 18776 160 18896 0 FreeSans 480 0 0 0 E1END[2]
port 6 nsew signal input
flabel metal3 s 0 19048 160 19168 0 FreeSans 480 0 0 0 E1END[3]
port 7 nsew signal input
flabel metal3 s 0 21496 160 21616 0 FreeSans 480 0 0 0 E2END[0]
port 8 nsew signal input
flabel metal3 s 0 21768 160 21888 0 FreeSans 480 0 0 0 E2END[1]
port 9 nsew signal input
flabel metal3 s 0 22040 160 22160 0 FreeSans 480 0 0 0 E2END[2]
port 10 nsew signal input
flabel metal3 s 0 22312 160 22432 0 FreeSans 480 0 0 0 E2END[3]
port 11 nsew signal input
flabel metal3 s 0 22584 160 22704 0 FreeSans 480 0 0 0 E2END[4]
port 12 nsew signal input
flabel metal3 s 0 22856 160 22976 0 FreeSans 480 0 0 0 E2END[5]
port 13 nsew signal input
flabel metal3 s 0 23128 160 23248 0 FreeSans 480 0 0 0 E2END[6]
port 14 nsew signal input
flabel metal3 s 0 23400 160 23520 0 FreeSans 480 0 0 0 E2END[7]
port 15 nsew signal input
flabel metal3 s 0 19320 160 19440 0 FreeSans 480 0 0 0 E2MID[0]
port 16 nsew signal input
flabel metal3 s 0 19592 160 19712 0 FreeSans 480 0 0 0 E2MID[1]
port 17 nsew signal input
flabel metal3 s 0 19864 160 19984 0 FreeSans 480 0 0 0 E2MID[2]
port 18 nsew signal input
flabel metal3 s 0 20136 160 20256 0 FreeSans 480 0 0 0 E2MID[3]
port 19 nsew signal input
flabel metal3 s 0 20408 160 20528 0 FreeSans 480 0 0 0 E2MID[4]
port 20 nsew signal input
flabel metal3 s 0 20680 160 20800 0 FreeSans 480 0 0 0 E2MID[5]
port 21 nsew signal input
flabel metal3 s 0 20952 160 21072 0 FreeSans 480 0 0 0 E2MID[6]
port 22 nsew signal input
flabel metal3 s 0 21224 160 21344 0 FreeSans 480 0 0 0 E2MID[7]
port 23 nsew signal input
flabel metal3 s 0 28024 160 28144 0 FreeSans 480 0 0 0 E6END[0]
port 24 nsew signal input
flabel metal3 s 0 30744 160 30864 0 FreeSans 480 0 0 0 E6END[10]
port 25 nsew signal input
flabel metal3 s 0 31016 160 31136 0 FreeSans 480 0 0 0 E6END[11]
port 26 nsew signal input
flabel metal3 s 0 28296 160 28416 0 FreeSans 480 0 0 0 E6END[1]
port 27 nsew signal input
flabel metal3 s 0 28568 160 28688 0 FreeSans 480 0 0 0 E6END[2]
port 28 nsew signal input
flabel metal3 s 0 28840 160 28960 0 FreeSans 480 0 0 0 E6END[3]
port 29 nsew signal input
flabel metal3 s 0 29112 160 29232 0 FreeSans 480 0 0 0 E6END[4]
port 30 nsew signal input
flabel metal3 s 0 29384 160 29504 0 FreeSans 480 0 0 0 E6END[5]
port 31 nsew signal input
flabel metal3 s 0 29656 160 29776 0 FreeSans 480 0 0 0 E6END[6]
port 32 nsew signal input
flabel metal3 s 0 29928 160 30048 0 FreeSans 480 0 0 0 E6END[7]
port 33 nsew signal input
flabel metal3 s 0 30200 160 30320 0 FreeSans 480 0 0 0 E6END[8]
port 34 nsew signal input
flabel metal3 s 0 30472 160 30592 0 FreeSans 480 0 0 0 E6END[9]
port 35 nsew signal input
flabel metal3 s 0 23672 160 23792 0 FreeSans 480 0 0 0 EE4END[0]
port 36 nsew signal input
flabel metal3 s 0 26392 160 26512 0 FreeSans 480 0 0 0 EE4END[10]
port 37 nsew signal input
flabel metal3 s 0 26664 160 26784 0 FreeSans 480 0 0 0 EE4END[11]
port 38 nsew signal input
flabel metal3 s 0 26936 160 27056 0 FreeSans 480 0 0 0 EE4END[12]
port 39 nsew signal input
flabel metal3 s 0 27208 160 27328 0 FreeSans 480 0 0 0 EE4END[13]
port 40 nsew signal input
flabel metal3 s 0 27480 160 27600 0 FreeSans 480 0 0 0 EE4END[14]
port 41 nsew signal input
flabel metal3 s 0 27752 160 27872 0 FreeSans 480 0 0 0 EE4END[15]
port 42 nsew signal input
flabel metal3 s 0 23944 160 24064 0 FreeSans 480 0 0 0 EE4END[1]
port 43 nsew signal input
flabel metal3 s 0 24216 160 24336 0 FreeSans 480 0 0 0 EE4END[2]
port 44 nsew signal input
flabel metal3 s 0 24488 160 24608 0 FreeSans 480 0 0 0 EE4END[3]
port 45 nsew signal input
flabel metal3 s 0 24760 160 24880 0 FreeSans 480 0 0 0 EE4END[4]
port 46 nsew signal input
flabel metal3 s 0 25032 160 25152 0 FreeSans 480 0 0 0 EE4END[5]
port 47 nsew signal input
flabel metal3 s 0 25304 160 25424 0 FreeSans 480 0 0 0 EE4END[6]
port 48 nsew signal input
flabel metal3 s 0 25576 160 25696 0 FreeSans 480 0 0 0 EE4END[7]
port 49 nsew signal input
flabel metal3 s 0 25848 160 25968 0 FreeSans 480 0 0 0 EE4END[8]
port 50 nsew signal input
flabel metal3 s 0 26120 160 26240 0 FreeSans 480 0 0 0 EE4END[9]
port 51 nsew signal input
flabel metal3 s 25840 16056 26000 16176 0 FreeSans 480 0 0 0 FAB2RAM_A0_O0
port 52 nsew signal tristate
flabel metal3 s 25840 16600 26000 16720 0 FreeSans 480 0 0 0 FAB2RAM_A0_O1
port 53 nsew signal tristate
flabel metal3 s 25840 17144 26000 17264 0 FreeSans 480 0 0 0 FAB2RAM_A0_O2
port 54 nsew signal tristate
flabel metal3 s 25840 17688 26000 17808 0 FreeSans 480 0 0 0 FAB2RAM_A0_O3
port 55 nsew signal tristate
flabel metal3 s 25840 13880 26000 14000 0 FreeSans 480 0 0 0 FAB2RAM_A1_O0
port 56 nsew signal tristate
flabel metal3 s 25840 14424 26000 14544 0 FreeSans 480 0 0 0 FAB2RAM_A1_O1
port 57 nsew signal tristate
flabel metal3 s 25840 14968 26000 15088 0 FreeSans 480 0 0 0 FAB2RAM_A1_O2
port 58 nsew signal tristate
flabel metal3 s 25840 15512 26000 15632 0 FreeSans 480 0 0 0 FAB2RAM_A1_O3
port 59 nsew signal tristate
flabel metal3 s 25840 11704 26000 11824 0 FreeSans 480 0 0 0 FAB2RAM_C_O0
port 60 nsew signal tristate
flabel metal3 s 25840 12248 26000 12368 0 FreeSans 480 0 0 0 FAB2RAM_C_O1
port 61 nsew signal tristate
flabel metal3 s 25840 12792 26000 12912 0 FreeSans 480 0 0 0 FAB2RAM_C_O2
port 62 nsew signal tristate
flabel metal3 s 25840 13336 26000 13456 0 FreeSans 480 0 0 0 FAB2RAM_C_O3
port 63 nsew signal tristate
flabel metal3 s 25840 24760 26000 24880 0 FreeSans 480 0 0 0 FAB2RAM_D0_O0
port 64 nsew signal tristate
flabel metal3 s 25840 25304 26000 25424 0 FreeSans 480 0 0 0 FAB2RAM_D0_O1
port 65 nsew signal tristate
flabel metal3 s 25840 25848 26000 25968 0 FreeSans 480 0 0 0 FAB2RAM_D0_O2
port 66 nsew signal tristate
flabel metal3 s 25840 26392 26000 26512 0 FreeSans 480 0 0 0 FAB2RAM_D0_O3
port 67 nsew signal tristate
flabel metal3 s 25840 22584 26000 22704 0 FreeSans 480 0 0 0 FAB2RAM_D1_O0
port 68 nsew signal tristate
flabel metal3 s 25840 23128 26000 23248 0 FreeSans 480 0 0 0 FAB2RAM_D1_O1
port 69 nsew signal tristate
flabel metal3 s 25840 23672 26000 23792 0 FreeSans 480 0 0 0 FAB2RAM_D1_O2
port 70 nsew signal tristate
flabel metal3 s 25840 24216 26000 24336 0 FreeSans 480 0 0 0 FAB2RAM_D1_O3
port 71 nsew signal tristate
flabel metal3 s 25840 20408 26000 20528 0 FreeSans 480 0 0 0 FAB2RAM_D2_O0
port 72 nsew signal tristate
flabel metal3 s 25840 20952 26000 21072 0 FreeSans 480 0 0 0 FAB2RAM_D2_O1
port 73 nsew signal tristate
flabel metal3 s 25840 21496 26000 21616 0 FreeSans 480 0 0 0 FAB2RAM_D2_O2
port 74 nsew signal tristate
flabel metal3 s 25840 22040 26000 22160 0 FreeSans 480 0 0 0 FAB2RAM_D2_O3
port 75 nsew signal tristate
flabel metal3 s 25840 18232 26000 18352 0 FreeSans 480 0 0 0 FAB2RAM_D3_O0
port 76 nsew signal tristate
flabel metal3 s 25840 18776 26000 18896 0 FreeSans 480 0 0 0 FAB2RAM_D3_O1
port 77 nsew signal tristate
flabel metal3 s 25840 19320 26000 19440 0 FreeSans 480 0 0 0 FAB2RAM_D3_O2
port 78 nsew signal tristate
flabel metal3 s 25840 19864 26000 19984 0 FreeSans 480 0 0 0 FAB2RAM_D3_O3
port 79 nsew signal tristate
flabel metal3 s 0 31288 160 31408 0 FreeSans 480 0 0 0 FrameData[0]
port 80 nsew signal input
flabel metal3 s 0 34008 160 34128 0 FreeSans 480 0 0 0 FrameData[10]
port 81 nsew signal input
flabel metal3 s 0 34280 160 34400 0 FreeSans 480 0 0 0 FrameData[11]
port 82 nsew signal input
flabel metal3 s 0 34552 160 34672 0 FreeSans 480 0 0 0 FrameData[12]
port 83 nsew signal input
flabel metal3 s 0 34824 160 34944 0 FreeSans 480 0 0 0 FrameData[13]
port 84 nsew signal input
flabel metal3 s 0 35096 160 35216 0 FreeSans 480 0 0 0 FrameData[14]
port 85 nsew signal input
flabel metal3 s 0 35368 160 35488 0 FreeSans 480 0 0 0 FrameData[15]
port 86 nsew signal input
flabel metal3 s 0 35640 160 35760 0 FreeSans 480 0 0 0 FrameData[16]
port 87 nsew signal input
flabel metal3 s 0 35912 160 36032 0 FreeSans 480 0 0 0 FrameData[17]
port 88 nsew signal input
flabel metal3 s 0 36184 160 36304 0 FreeSans 480 0 0 0 FrameData[18]
port 89 nsew signal input
flabel metal3 s 0 36456 160 36576 0 FreeSans 480 0 0 0 FrameData[19]
port 90 nsew signal input
flabel metal3 s 0 31560 160 31680 0 FreeSans 480 0 0 0 FrameData[1]
port 91 nsew signal input
flabel metal3 s 0 36728 160 36848 0 FreeSans 480 0 0 0 FrameData[20]
port 92 nsew signal input
flabel metal3 s 0 37000 160 37120 0 FreeSans 480 0 0 0 FrameData[21]
port 93 nsew signal input
flabel metal3 s 0 37272 160 37392 0 FreeSans 480 0 0 0 FrameData[22]
port 94 nsew signal input
flabel metal3 s 0 37544 160 37664 0 FreeSans 480 0 0 0 FrameData[23]
port 95 nsew signal input
flabel metal3 s 0 37816 160 37936 0 FreeSans 480 0 0 0 FrameData[24]
port 96 nsew signal input
flabel metal3 s 0 38088 160 38208 0 FreeSans 480 0 0 0 FrameData[25]
port 97 nsew signal input
flabel metal3 s 0 38360 160 38480 0 FreeSans 480 0 0 0 FrameData[26]
port 98 nsew signal input
flabel metal3 s 0 38632 160 38752 0 FreeSans 480 0 0 0 FrameData[27]
port 99 nsew signal input
flabel metal3 s 0 38904 160 39024 0 FreeSans 480 0 0 0 FrameData[28]
port 100 nsew signal input
flabel metal3 s 0 39176 160 39296 0 FreeSans 480 0 0 0 FrameData[29]
port 101 nsew signal input
flabel metal3 s 0 31832 160 31952 0 FreeSans 480 0 0 0 FrameData[2]
port 102 nsew signal input
flabel metal3 s 0 39448 160 39568 0 FreeSans 480 0 0 0 FrameData[30]
port 103 nsew signal input
flabel metal3 s 0 39720 160 39840 0 FreeSans 480 0 0 0 FrameData[31]
port 104 nsew signal input
flabel metal3 s 0 32104 160 32224 0 FreeSans 480 0 0 0 FrameData[3]
port 105 nsew signal input
flabel metal3 s 0 32376 160 32496 0 FreeSans 480 0 0 0 FrameData[4]
port 106 nsew signal input
flabel metal3 s 0 32648 160 32768 0 FreeSans 480 0 0 0 FrameData[5]
port 107 nsew signal input
flabel metal3 s 0 32920 160 33040 0 FreeSans 480 0 0 0 FrameData[6]
port 108 nsew signal input
flabel metal3 s 0 33192 160 33312 0 FreeSans 480 0 0 0 FrameData[7]
port 109 nsew signal input
flabel metal3 s 0 33464 160 33584 0 FreeSans 480 0 0 0 FrameData[8]
port 110 nsew signal input
flabel metal3 s 0 33736 160 33856 0 FreeSans 480 0 0 0 FrameData[9]
port 111 nsew signal input
flabel metal3 s 25840 26936 26000 27056 0 FreeSans 480 0 0 0 FrameData_O[0]
port 112 nsew signal tristate
flabel metal3 s 25840 32376 26000 32496 0 FreeSans 480 0 0 0 FrameData_O[10]
port 113 nsew signal tristate
flabel metal3 s 25840 32920 26000 33040 0 FreeSans 480 0 0 0 FrameData_O[11]
port 114 nsew signal tristate
flabel metal3 s 25840 33464 26000 33584 0 FreeSans 480 0 0 0 FrameData_O[12]
port 115 nsew signal tristate
flabel metal3 s 25840 34008 26000 34128 0 FreeSans 480 0 0 0 FrameData_O[13]
port 116 nsew signal tristate
flabel metal3 s 25840 34552 26000 34672 0 FreeSans 480 0 0 0 FrameData_O[14]
port 117 nsew signal tristate
flabel metal3 s 25840 35096 26000 35216 0 FreeSans 480 0 0 0 FrameData_O[15]
port 118 nsew signal tristate
flabel metal3 s 25840 35640 26000 35760 0 FreeSans 480 0 0 0 FrameData_O[16]
port 119 nsew signal tristate
flabel metal3 s 25840 36184 26000 36304 0 FreeSans 480 0 0 0 FrameData_O[17]
port 120 nsew signal tristate
flabel metal3 s 25840 36728 26000 36848 0 FreeSans 480 0 0 0 FrameData_O[18]
port 121 nsew signal tristate
flabel metal3 s 25840 37272 26000 37392 0 FreeSans 480 0 0 0 FrameData_O[19]
port 122 nsew signal tristate
flabel metal3 s 25840 27480 26000 27600 0 FreeSans 480 0 0 0 FrameData_O[1]
port 123 nsew signal tristate
flabel metal3 s 25840 37816 26000 37936 0 FreeSans 480 0 0 0 FrameData_O[20]
port 124 nsew signal tristate
flabel metal3 s 25840 38360 26000 38480 0 FreeSans 480 0 0 0 FrameData_O[21]
port 125 nsew signal tristate
flabel metal3 s 25840 38904 26000 39024 0 FreeSans 480 0 0 0 FrameData_O[22]
port 126 nsew signal tristate
flabel metal3 s 25840 39448 26000 39568 0 FreeSans 480 0 0 0 FrameData_O[23]
port 127 nsew signal tristate
flabel metal3 s 25840 39992 26000 40112 0 FreeSans 480 0 0 0 FrameData_O[24]
port 128 nsew signal tristate
flabel metal3 s 25840 40536 26000 40656 0 FreeSans 480 0 0 0 FrameData_O[25]
port 129 nsew signal tristate
flabel metal3 s 25840 41080 26000 41200 0 FreeSans 480 0 0 0 FrameData_O[26]
port 130 nsew signal tristate
flabel metal3 s 25840 41624 26000 41744 0 FreeSans 480 0 0 0 FrameData_O[27]
port 131 nsew signal tristate
flabel metal3 s 25840 42168 26000 42288 0 FreeSans 480 0 0 0 FrameData_O[28]
port 132 nsew signal tristate
flabel metal3 s 25840 42712 26000 42832 0 FreeSans 480 0 0 0 FrameData_O[29]
port 133 nsew signal tristate
flabel metal3 s 25840 28024 26000 28144 0 FreeSans 480 0 0 0 FrameData_O[2]
port 134 nsew signal tristate
flabel metal3 s 25840 43256 26000 43376 0 FreeSans 480 0 0 0 FrameData_O[30]
port 135 nsew signal tristate
flabel metal3 s 25840 43800 26000 43920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 136 nsew signal tristate
flabel metal3 s 25840 28568 26000 28688 0 FreeSans 480 0 0 0 FrameData_O[3]
port 137 nsew signal tristate
flabel metal3 s 25840 29112 26000 29232 0 FreeSans 480 0 0 0 FrameData_O[4]
port 138 nsew signal tristate
flabel metal3 s 25840 29656 26000 29776 0 FreeSans 480 0 0 0 FrameData_O[5]
port 139 nsew signal tristate
flabel metal3 s 25840 30200 26000 30320 0 FreeSans 480 0 0 0 FrameData_O[6]
port 140 nsew signal tristate
flabel metal3 s 25840 30744 26000 30864 0 FreeSans 480 0 0 0 FrameData_O[7]
port 141 nsew signal tristate
flabel metal3 s 25840 31288 26000 31408 0 FreeSans 480 0 0 0 FrameData_O[8]
port 142 nsew signal tristate
flabel metal3 s 25840 31832 26000 31952 0 FreeSans 480 0 0 0 FrameData_O[9]
port 143 nsew signal tristate
flabel metal2 s 20350 0 20406 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 144 nsew signal input
flabel metal2 s 23110 0 23166 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 145 nsew signal input
flabel metal2 s 23386 0 23442 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 146 nsew signal input
flabel metal2 s 23662 0 23718 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 147 nsew signal input
flabel metal2 s 23938 0 23994 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 148 nsew signal input
flabel metal2 s 24214 0 24270 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 149 nsew signal input
flabel metal2 s 24490 0 24546 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 150 nsew signal input
flabel metal2 s 24766 0 24822 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 151 nsew signal input
flabel metal2 s 25042 0 25098 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 152 nsew signal input
flabel metal2 s 25318 0 25374 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 153 nsew signal input
flabel metal2 s 25594 0 25650 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 154 nsew signal input
flabel metal2 s 20626 0 20682 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 155 nsew signal input
flabel metal2 s 20902 0 20958 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 156 nsew signal input
flabel metal2 s 21178 0 21234 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 157 nsew signal input
flabel metal2 s 21454 0 21510 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 158 nsew signal input
flabel metal2 s 21730 0 21786 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 159 nsew signal input
flabel metal2 s 22006 0 22062 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 160 nsew signal input
flabel metal2 s 22282 0 22338 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 161 nsew signal input
flabel metal2 s 22558 0 22614 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 162 nsew signal input
flabel metal2 s 22834 0 22890 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 163 nsew signal input
flabel metal2 s 20350 44840 20406 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 164 nsew signal tristate
flabel metal2 s 23110 44840 23166 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 165 nsew signal tristate
flabel metal2 s 23386 44840 23442 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 166 nsew signal tristate
flabel metal2 s 23662 44840 23718 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 167 nsew signal tristate
flabel metal2 s 23938 44840 23994 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 168 nsew signal tristate
flabel metal2 s 24214 44840 24270 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 169 nsew signal tristate
flabel metal2 s 24490 44840 24546 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 170 nsew signal tristate
flabel metal2 s 24766 44840 24822 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 171 nsew signal tristate
flabel metal2 s 25042 44840 25098 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 172 nsew signal tristate
flabel metal2 s 25318 44840 25374 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 173 nsew signal tristate
flabel metal2 s 25594 44840 25650 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 174 nsew signal tristate
flabel metal2 s 20626 44840 20682 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 175 nsew signal tristate
flabel metal2 s 20902 44840 20958 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 176 nsew signal tristate
flabel metal2 s 21178 44840 21234 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 177 nsew signal tristate
flabel metal2 s 21454 44840 21510 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 178 nsew signal tristate
flabel metal2 s 21730 44840 21786 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 179 nsew signal tristate
flabel metal2 s 22006 44840 22062 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 180 nsew signal tristate
flabel metal2 s 22282 44840 22338 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 181 nsew signal tristate
flabel metal2 s 22558 44840 22614 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 182 nsew signal tristate
flabel metal2 s 22834 44840 22890 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 183 nsew signal tristate
flabel metal2 s 202 44840 258 45000 0 FreeSans 224 90 0 0 N1BEG[0]
port 184 nsew signal tristate
flabel metal2 s 478 44840 534 45000 0 FreeSans 224 90 0 0 N1BEG[1]
port 185 nsew signal tristate
flabel metal2 s 754 44840 810 45000 0 FreeSans 224 90 0 0 N1BEG[2]
port 186 nsew signal tristate
flabel metal2 s 1030 44840 1086 45000 0 FreeSans 224 90 0 0 N1BEG[3]
port 187 nsew signal tristate
flabel metal2 s 202 0 258 160 0 FreeSans 224 90 0 0 N1END[0]
port 188 nsew signal input
flabel metal2 s 478 0 534 160 0 FreeSans 224 90 0 0 N1END[1]
port 189 nsew signal input
flabel metal2 s 754 0 810 160 0 FreeSans 224 90 0 0 N1END[2]
port 190 nsew signal input
flabel metal2 s 1030 0 1086 160 0 FreeSans 224 90 0 0 N1END[3]
port 191 nsew signal input
flabel metal2 s 1306 44840 1362 45000 0 FreeSans 224 90 0 0 N2BEG[0]
port 192 nsew signal tristate
flabel metal2 s 1582 44840 1638 45000 0 FreeSans 224 90 0 0 N2BEG[1]
port 193 nsew signal tristate
flabel metal2 s 1858 44840 1914 45000 0 FreeSans 224 90 0 0 N2BEG[2]
port 194 nsew signal tristate
flabel metal2 s 2134 44840 2190 45000 0 FreeSans 224 90 0 0 N2BEG[3]
port 195 nsew signal tristate
flabel metal2 s 2410 44840 2466 45000 0 FreeSans 224 90 0 0 N2BEG[4]
port 196 nsew signal tristate
flabel metal2 s 2686 44840 2742 45000 0 FreeSans 224 90 0 0 N2BEG[5]
port 197 nsew signal tristate
flabel metal2 s 2962 44840 3018 45000 0 FreeSans 224 90 0 0 N2BEG[6]
port 198 nsew signal tristate
flabel metal2 s 3238 44840 3294 45000 0 FreeSans 224 90 0 0 N2BEG[7]
port 199 nsew signal tristate
flabel metal2 s 3514 44840 3570 45000 0 FreeSans 224 90 0 0 N2BEGb[0]
port 200 nsew signal tristate
flabel metal2 s 3790 44840 3846 45000 0 FreeSans 224 90 0 0 N2BEGb[1]
port 201 nsew signal tristate
flabel metal2 s 4066 44840 4122 45000 0 FreeSans 224 90 0 0 N2BEGb[2]
port 202 nsew signal tristate
flabel metal2 s 4342 44840 4398 45000 0 FreeSans 224 90 0 0 N2BEGb[3]
port 203 nsew signal tristate
flabel metal2 s 4618 44840 4674 45000 0 FreeSans 224 90 0 0 N2BEGb[4]
port 204 nsew signal tristate
flabel metal2 s 4894 44840 4950 45000 0 FreeSans 224 90 0 0 N2BEGb[5]
port 205 nsew signal tristate
flabel metal2 s 5170 44840 5226 45000 0 FreeSans 224 90 0 0 N2BEGb[6]
port 206 nsew signal tristate
flabel metal2 s 5446 44840 5502 45000 0 FreeSans 224 90 0 0 N2BEGb[7]
port 207 nsew signal tristate
flabel metal2 s 3514 0 3570 160 0 FreeSans 224 90 0 0 N2END[0]
port 208 nsew signal input
flabel metal2 s 3790 0 3846 160 0 FreeSans 224 90 0 0 N2END[1]
port 209 nsew signal input
flabel metal2 s 4066 0 4122 160 0 FreeSans 224 90 0 0 N2END[2]
port 210 nsew signal input
flabel metal2 s 4342 0 4398 160 0 FreeSans 224 90 0 0 N2END[3]
port 211 nsew signal input
flabel metal2 s 4618 0 4674 160 0 FreeSans 224 90 0 0 N2END[4]
port 212 nsew signal input
flabel metal2 s 4894 0 4950 160 0 FreeSans 224 90 0 0 N2END[5]
port 213 nsew signal input
flabel metal2 s 5170 0 5226 160 0 FreeSans 224 90 0 0 N2END[6]
port 214 nsew signal input
flabel metal2 s 5446 0 5502 160 0 FreeSans 224 90 0 0 N2END[7]
port 215 nsew signal input
flabel metal2 s 1306 0 1362 160 0 FreeSans 224 90 0 0 N2MID[0]
port 216 nsew signal input
flabel metal2 s 1582 0 1638 160 0 FreeSans 224 90 0 0 N2MID[1]
port 217 nsew signal input
flabel metal2 s 1858 0 1914 160 0 FreeSans 224 90 0 0 N2MID[2]
port 218 nsew signal input
flabel metal2 s 2134 0 2190 160 0 FreeSans 224 90 0 0 N2MID[3]
port 219 nsew signal input
flabel metal2 s 2410 0 2466 160 0 FreeSans 224 90 0 0 N2MID[4]
port 220 nsew signal input
flabel metal2 s 2686 0 2742 160 0 FreeSans 224 90 0 0 N2MID[5]
port 221 nsew signal input
flabel metal2 s 2962 0 3018 160 0 FreeSans 224 90 0 0 N2MID[6]
port 222 nsew signal input
flabel metal2 s 3238 0 3294 160 0 FreeSans 224 90 0 0 N2MID[7]
port 223 nsew signal input
flabel metal2 s 5722 44840 5778 45000 0 FreeSans 224 90 0 0 N4BEG[0]
port 224 nsew signal tristate
flabel metal2 s 8482 44840 8538 45000 0 FreeSans 224 90 0 0 N4BEG[10]
port 225 nsew signal tristate
flabel metal2 s 8758 44840 8814 45000 0 FreeSans 224 90 0 0 N4BEG[11]
port 226 nsew signal tristate
flabel metal2 s 9034 44840 9090 45000 0 FreeSans 224 90 0 0 N4BEG[12]
port 227 nsew signal tristate
flabel metal2 s 9310 44840 9366 45000 0 FreeSans 224 90 0 0 N4BEG[13]
port 228 nsew signal tristate
flabel metal2 s 9586 44840 9642 45000 0 FreeSans 224 90 0 0 N4BEG[14]
port 229 nsew signal tristate
flabel metal2 s 9862 44840 9918 45000 0 FreeSans 224 90 0 0 N4BEG[15]
port 230 nsew signal tristate
flabel metal2 s 5998 44840 6054 45000 0 FreeSans 224 90 0 0 N4BEG[1]
port 231 nsew signal tristate
flabel metal2 s 6274 44840 6330 45000 0 FreeSans 224 90 0 0 N4BEG[2]
port 232 nsew signal tristate
flabel metal2 s 6550 44840 6606 45000 0 FreeSans 224 90 0 0 N4BEG[3]
port 233 nsew signal tristate
flabel metal2 s 6826 44840 6882 45000 0 FreeSans 224 90 0 0 N4BEG[4]
port 234 nsew signal tristate
flabel metal2 s 7102 44840 7158 45000 0 FreeSans 224 90 0 0 N4BEG[5]
port 235 nsew signal tristate
flabel metal2 s 7378 44840 7434 45000 0 FreeSans 224 90 0 0 N4BEG[6]
port 236 nsew signal tristate
flabel metal2 s 7654 44840 7710 45000 0 FreeSans 224 90 0 0 N4BEG[7]
port 237 nsew signal tristate
flabel metal2 s 7930 44840 7986 45000 0 FreeSans 224 90 0 0 N4BEG[8]
port 238 nsew signal tristate
flabel metal2 s 8206 44840 8262 45000 0 FreeSans 224 90 0 0 N4BEG[9]
port 239 nsew signal tristate
flabel metal2 s 5722 0 5778 160 0 FreeSans 224 90 0 0 N4END[0]
port 240 nsew signal input
flabel metal2 s 8482 0 8538 160 0 FreeSans 224 90 0 0 N4END[10]
port 241 nsew signal input
flabel metal2 s 8758 0 8814 160 0 FreeSans 224 90 0 0 N4END[11]
port 242 nsew signal input
flabel metal2 s 9034 0 9090 160 0 FreeSans 224 90 0 0 N4END[12]
port 243 nsew signal input
flabel metal2 s 9310 0 9366 160 0 FreeSans 224 90 0 0 N4END[13]
port 244 nsew signal input
flabel metal2 s 9586 0 9642 160 0 FreeSans 224 90 0 0 N4END[14]
port 245 nsew signal input
flabel metal2 s 9862 0 9918 160 0 FreeSans 224 90 0 0 N4END[15]
port 246 nsew signal input
flabel metal2 s 5998 0 6054 160 0 FreeSans 224 90 0 0 N4END[1]
port 247 nsew signal input
flabel metal2 s 6274 0 6330 160 0 FreeSans 224 90 0 0 N4END[2]
port 248 nsew signal input
flabel metal2 s 6550 0 6606 160 0 FreeSans 224 90 0 0 N4END[3]
port 249 nsew signal input
flabel metal2 s 6826 0 6882 160 0 FreeSans 224 90 0 0 N4END[4]
port 250 nsew signal input
flabel metal2 s 7102 0 7158 160 0 FreeSans 224 90 0 0 N4END[5]
port 251 nsew signal input
flabel metal2 s 7378 0 7434 160 0 FreeSans 224 90 0 0 N4END[6]
port 252 nsew signal input
flabel metal2 s 7654 0 7710 160 0 FreeSans 224 90 0 0 N4END[7]
port 253 nsew signal input
flabel metal2 s 7930 0 7986 160 0 FreeSans 224 90 0 0 N4END[8]
port 254 nsew signal input
flabel metal2 s 8206 0 8262 160 0 FreeSans 224 90 0 0 N4END[9]
port 255 nsew signal input
flabel metal3 s 25840 7352 26000 7472 0 FreeSans 480 0 0 0 RAM2FAB_D0_I0
port 256 nsew signal input
flabel metal3 s 25840 7896 26000 8016 0 FreeSans 480 0 0 0 RAM2FAB_D0_I1
port 257 nsew signal input
flabel metal3 s 25840 8440 26000 8560 0 FreeSans 480 0 0 0 RAM2FAB_D0_I2
port 258 nsew signal input
flabel metal3 s 25840 8984 26000 9104 0 FreeSans 480 0 0 0 RAM2FAB_D0_I3
port 259 nsew signal input
flabel metal3 s 25840 5176 26000 5296 0 FreeSans 480 0 0 0 RAM2FAB_D1_I0
port 260 nsew signal input
flabel metal3 s 25840 5720 26000 5840 0 FreeSans 480 0 0 0 RAM2FAB_D1_I1
port 261 nsew signal input
flabel metal3 s 25840 6264 26000 6384 0 FreeSans 480 0 0 0 RAM2FAB_D1_I2
port 262 nsew signal input
flabel metal3 s 25840 6808 26000 6928 0 FreeSans 480 0 0 0 RAM2FAB_D1_I3
port 263 nsew signal input
flabel metal3 s 25840 3000 26000 3120 0 FreeSans 480 0 0 0 RAM2FAB_D2_I0
port 264 nsew signal input
flabel metal3 s 25840 3544 26000 3664 0 FreeSans 480 0 0 0 RAM2FAB_D2_I1
port 265 nsew signal input
flabel metal3 s 25840 4088 26000 4208 0 FreeSans 480 0 0 0 RAM2FAB_D2_I2
port 266 nsew signal input
flabel metal3 s 25840 4632 26000 4752 0 FreeSans 480 0 0 0 RAM2FAB_D2_I3
port 267 nsew signal input
flabel metal3 s 25840 824 26000 944 0 FreeSans 480 0 0 0 RAM2FAB_D3_I0
port 268 nsew signal input
flabel metal3 s 25840 1368 26000 1488 0 FreeSans 480 0 0 0 RAM2FAB_D3_I1
port 269 nsew signal input
flabel metal3 s 25840 1912 26000 2032 0 FreeSans 480 0 0 0 RAM2FAB_D3_I2
port 270 nsew signal input
flabel metal3 s 25840 2456 26000 2576 0 FreeSans 480 0 0 0 RAM2FAB_D3_I3
port 271 nsew signal input
flabel metal2 s 10138 0 10194 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 272 nsew signal tristate
flabel metal2 s 10414 0 10470 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 273 nsew signal tristate
flabel metal2 s 10690 0 10746 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 274 nsew signal tristate
flabel metal2 s 10966 0 11022 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 275 nsew signal tristate
flabel metal2 s 10138 44840 10194 45000 0 FreeSans 224 90 0 0 S1END[0]
port 276 nsew signal input
flabel metal2 s 10414 44840 10470 45000 0 FreeSans 224 90 0 0 S1END[1]
port 277 nsew signal input
flabel metal2 s 10690 44840 10746 45000 0 FreeSans 224 90 0 0 S1END[2]
port 278 nsew signal input
flabel metal2 s 10966 44840 11022 45000 0 FreeSans 224 90 0 0 S1END[3]
port 279 nsew signal input
flabel metal2 s 13450 0 13506 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 280 nsew signal tristate
flabel metal2 s 13726 0 13782 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 281 nsew signal tristate
flabel metal2 s 14002 0 14058 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 282 nsew signal tristate
flabel metal2 s 14278 0 14334 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 283 nsew signal tristate
flabel metal2 s 14554 0 14610 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 284 nsew signal tristate
flabel metal2 s 14830 0 14886 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 285 nsew signal tristate
flabel metal2 s 15106 0 15162 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 286 nsew signal tristate
flabel metal2 s 15382 0 15438 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 287 nsew signal tristate
flabel metal2 s 11242 0 11298 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 288 nsew signal tristate
flabel metal2 s 11518 0 11574 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 289 nsew signal tristate
flabel metal2 s 11794 0 11850 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 290 nsew signal tristate
flabel metal2 s 12070 0 12126 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 291 nsew signal tristate
flabel metal2 s 12346 0 12402 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 292 nsew signal tristate
flabel metal2 s 12622 0 12678 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 293 nsew signal tristate
flabel metal2 s 12898 0 12954 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 294 nsew signal tristate
flabel metal2 s 13174 0 13230 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 295 nsew signal tristate
flabel metal2 s 11242 44840 11298 45000 0 FreeSans 224 90 0 0 S2END[0]
port 296 nsew signal input
flabel metal2 s 11518 44840 11574 45000 0 FreeSans 224 90 0 0 S2END[1]
port 297 nsew signal input
flabel metal2 s 11794 44840 11850 45000 0 FreeSans 224 90 0 0 S2END[2]
port 298 nsew signal input
flabel metal2 s 12070 44840 12126 45000 0 FreeSans 224 90 0 0 S2END[3]
port 299 nsew signal input
flabel metal2 s 12346 44840 12402 45000 0 FreeSans 224 90 0 0 S2END[4]
port 300 nsew signal input
flabel metal2 s 12622 44840 12678 45000 0 FreeSans 224 90 0 0 S2END[5]
port 301 nsew signal input
flabel metal2 s 12898 44840 12954 45000 0 FreeSans 224 90 0 0 S2END[6]
port 302 nsew signal input
flabel metal2 s 13174 44840 13230 45000 0 FreeSans 224 90 0 0 S2END[7]
port 303 nsew signal input
flabel metal2 s 13450 44840 13506 45000 0 FreeSans 224 90 0 0 S2MID[0]
port 304 nsew signal input
flabel metal2 s 13726 44840 13782 45000 0 FreeSans 224 90 0 0 S2MID[1]
port 305 nsew signal input
flabel metal2 s 14002 44840 14058 45000 0 FreeSans 224 90 0 0 S2MID[2]
port 306 nsew signal input
flabel metal2 s 14278 44840 14334 45000 0 FreeSans 224 90 0 0 S2MID[3]
port 307 nsew signal input
flabel metal2 s 14554 44840 14610 45000 0 FreeSans 224 90 0 0 S2MID[4]
port 308 nsew signal input
flabel metal2 s 14830 44840 14886 45000 0 FreeSans 224 90 0 0 S2MID[5]
port 309 nsew signal input
flabel metal2 s 15106 44840 15162 45000 0 FreeSans 224 90 0 0 S2MID[6]
port 310 nsew signal input
flabel metal2 s 15382 44840 15438 45000 0 FreeSans 224 90 0 0 S2MID[7]
port 311 nsew signal input
flabel metal2 s 15658 0 15714 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 312 nsew signal tristate
flabel metal2 s 18418 0 18474 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 313 nsew signal tristate
flabel metal2 s 18694 0 18750 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 314 nsew signal tristate
flabel metal2 s 18970 0 19026 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 315 nsew signal tristate
flabel metal2 s 19246 0 19302 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 316 nsew signal tristate
flabel metal2 s 19522 0 19578 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 317 nsew signal tristate
flabel metal2 s 19798 0 19854 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 318 nsew signal tristate
flabel metal2 s 15934 0 15990 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 319 nsew signal tristate
flabel metal2 s 16210 0 16266 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 320 nsew signal tristate
flabel metal2 s 16486 0 16542 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 321 nsew signal tristate
flabel metal2 s 16762 0 16818 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 322 nsew signal tristate
flabel metal2 s 17038 0 17094 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 323 nsew signal tristate
flabel metal2 s 17314 0 17370 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 324 nsew signal tristate
flabel metal2 s 17590 0 17646 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 325 nsew signal tristate
flabel metal2 s 17866 0 17922 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 326 nsew signal tristate
flabel metal2 s 18142 0 18198 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 327 nsew signal tristate
flabel metal2 s 15658 44840 15714 45000 0 FreeSans 224 90 0 0 S4END[0]
port 328 nsew signal input
flabel metal2 s 18418 44840 18474 45000 0 FreeSans 224 90 0 0 S4END[10]
port 329 nsew signal input
flabel metal2 s 18694 44840 18750 45000 0 FreeSans 224 90 0 0 S4END[11]
port 330 nsew signal input
flabel metal2 s 18970 44840 19026 45000 0 FreeSans 224 90 0 0 S4END[12]
port 331 nsew signal input
flabel metal2 s 19246 44840 19302 45000 0 FreeSans 224 90 0 0 S4END[13]
port 332 nsew signal input
flabel metal2 s 19522 44840 19578 45000 0 FreeSans 224 90 0 0 S4END[14]
port 333 nsew signal input
flabel metal2 s 19798 44840 19854 45000 0 FreeSans 224 90 0 0 S4END[15]
port 334 nsew signal input
flabel metal2 s 15934 44840 15990 45000 0 FreeSans 224 90 0 0 S4END[1]
port 335 nsew signal input
flabel metal2 s 16210 44840 16266 45000 0 FreeSans 224 90 0 0 S4END[2]
port 336 nsew signal input
flabel metal2 s 16486 44840 16542 45000 0 FreeSans 224 90 0 0 S4END[3]
port 337 nsew signal input
flabel metal2 s 16762 44840 16818 45000 0 FreeSans 224 90 0 0 S4END[4]
port 338 nsew signal input
flabel metal2 s 17038 44840 17094 45000 0 FreeSans 224 90 0 0 S4END[5]
port 339 nsew signal input
flabel metal2 s 17314 44840 17370 45000 0 FreeSans 224 90 0 0 S4END[6]
port 340 nsew signal input
flabel metal2 s 17590 44840 17646 45000 0 FreeSans 224 90 0 0 S4END[7]
port 341 nsew signal input
flabel metal2 s 17866 44840 17922 45000 0 FreeSans 224 90 0 0 S4END[8]
port 342 nsew signal input
flabel metal2 s 18142 44840 18198 45000 0 FreeSans 224 90 0 0 S4END[9]
port 343 nsew signal input
flabel metal2 s 20074 0 20130 160 0 FreeSans 224 90 0 0 UserCLK
port 344 nsew signal input
flabel metal2 s 20074 44840 20130 45000 0 FreeSans 224 90 0 0 UserCLKo
port 345 nsew signal tristate
flabel metal4 s 6878 1040 7198 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 12812 1040 13132 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 18746 1040 19066 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 24680 1040 25000 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 3911 1040 4231 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 9845 1040 10165 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 15779 1040 16099 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 21713 1040 22033 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal3 s 0 5176 160 5296 0 FreeSans 480 0 0 0 W1BEG[0]
port 348 nsew signal tristate
flabel metal3 s 0 5448 160 5568 0 FreeSans 480 0 0 0 W1BEG[1]
port 349 nsew signal tristate
flabel metal3 s 0 5720 160 5840 0 FreeSans 480 0 0 0 W1BEG[2]
port 350 nsew signal tristate
flabel metal3 s 0 5992 160 6112 0 FreeSans 480 0 0 0 W1BEG[3]
port 351 nsew signal tristate
flabel metal3 s 0 6264 160 6384 0 FreeSans 480 0 0 0 W2BEG[0]
port 352 nsew signal tristate
flabel metal3 s 0 6536 160 6656 0 FreeSans 480 0 0 0 W2BEG[1]
port 353 nsew signal tristate
flabel metal3 s 0 6808 160 6928 0 FreeSans 480 0 0 0 W2BEG[2]
port 354 nsew signal tristate
flabel metal3 s 0 7080 160 7200 0 FreeSans 480 0 0 0 W2BEG[3]
port 355 nsew signal tristate
flabel metal3 s 0 7352 160 7472 0 FreeSans 480 0 0 0 W2BEG[4]
port 356 nsew signal tristate
flabel metal3 s 0 7624 160 7744 0 FreeSans 480 0 0 0 W2BEG[5]
port 357 nsew signal tristate
flabel metal3 s 0 7896 160 8016 0 FreeSans 480 0 0 0 W2BEG[6]
port 358 nsew signal tristate
flabel metal3 s 0 8168 160 8288 0 FreeSans 480 0 0 0 W2BEG[7]
port 359 nsew signal tristate
flabel metal3 s 0 8440 160 8560 0 FreeSans 480 0 0 0 W2BEGb[0]
port 360 nsew signal tristate
flabel metal3 s 0 8712 160 8832 0 FreeSans 480 0 0 0 W2BEGb[1]
port 361 nsew signal tristate
flabel metal3 s 0 8984 160 9104 0 FreeSans 480 0 0 0 W2BEGb[2]
port 362 nsew signal tristate
flabel metal3 s 0 9256 160 9376 0 FreeSans 480 0 0 0 W2BEGb[3]
port 363 nsew signal tristate
flabel metal3 s 0 9528 160 9648 0 FreeSans 480 0 0 0 W2BEGb[4]
port 364 nsew signal tristate
flabel metal3 s 0 9800 160 9920 0 FreeSans 480 0 0 0 W2BEGb[5]
port 365 nsew signal tristate
flabel metal3 s 0 10072 160 10192 0 FreeSans 480 0 0 0 W2BEGb[6]
port 366 nsew signal tristate
flabel metal3 s 0 10344 160 10464 0 FreeSans 480 0 0 0 W2BEGb[7]
port 367 nsew signal tristate
flabel metal3 s 0 14968 160 15088 0 FreeSans 480 0 0 0 W6BEG[0]
port 368 nsew signal tristate
flabel metal3 s 0 17688 160 17808 0 FreeSans 480 0 0 0 W6BEG[10]
port 369 nsew signal tristate
flabel metal3 s 0 17960 160 18080 0 FreeSans 480 0 0 0 W6BEG[11]
port 370 nsew signal tristate
flabel metal3 s 0 15240 160 15360 0 FreeSans 480 0 0 0 W6BEG[1]
port 371 nsew signal tristate
flabel metal3 s 0 15512 160 15632 0 FreeSans 480 0 0 0 W6BEG[2]
port 372 nsew signal tristate
flabel metal3 s 0 15784 160 15904 0 FreeSans 480 0 0 0 W6BEG[3]
port 373 nsew signal tristate
flabel metal3 s 0 16056 160 16176 0 FreeSans 480 0 0 0 W6BEG[4]
port 374 nsew signal tristate
flabel metal3 s 0 16328 160 16448 0 FreeSans 480 0 0 0 W6BEG[5]
port 375 nsew signal tristate
flabel metal3 s 0 16600 160 16720 0 FreeSans 480 0 0 0 W6BEG[6]
port 376 nsew signal tristate
flabel metal3 s 0 16872 160 16992 0 FreeSans 480 0 0 0 W6BEG[7]
port 377 nsew signal tristate
flabel metal3 s 0 17144 160 17264 0 FreeSans 480 0 0 0 W6BEG[8]
port 378 nsew signal tristate
flabel metal3 s 0 17416 160 17536 0 FreeSans 480 0 0 0 W6BEG[9]
port 379 nsew signal tristate
flabel metal3 s 0 10616 160 10736 0 FreeSans 480 0 0 0 WW4BEG[0]
port 380 nsew signal tristate
flabel metal3 s 0 13336 160 13456 0 FreeSans 480 0 0 0 WW4BEG[10]
port 381 nsew signal tristate
flabel metal3 s 0 13608 160 13728 0 FreeSans 480 0 0 0 WW4BEG[11]
port 382 nsew signal tristate
flabel metal3 s 0 13880 160 14000 0 FreeSans 480 0 0 0 WW4BEG[12]
port 383 nsew signal tristate
flabel metal3 s 0 14152 160 14272 0 FreeSans 480 0 0 0 WW4BEG[13]
port 384 nsew signal tristate
flabel metal3 s 0 14424 160 14544 0 FreeSans 480 0 0 0 WW4BEG[14]
port 385 nsew signal tristate
flabel metal3 s 0 14696 160 14816 0 FreeSans 480 0 0 0 WW4BEG[15]
port 386 nsew signal tristate
flabel metal3 s 0 10888 160 11008 0 FreeSans 480 0 0 0 WW4BEG[1]
port 387 nsew signal tristate
flabel metal3 s 0 11160 160 11280 0 FreeSans 480 0 0 0 WW4BEG[2]
port 388 nsew signal tristate
flabel metal3 s 0 11432 160 11552 0 FreeSans 480 0 0 0 WW4BEG[3]
port 389 nsew signal tristate
flabel metal3 s 0 11704 160 11824 0 FreeSans 480 0 0 0 WW4BEG[4]
port 390 nsew signal tristate
flabel metal3 s 0 11976 160 12096 0 FreeSans 480 0 0 0 WW4BEG[5]
port 391 nsew signal tristate
flabel metal3 s 0 12248 160 12368 0 FreeSans 480 0 0 0 WW4BEG[6]
port 392 nsew signal tristate
flabel metal3 s 0 12520 160 12640 0 FreeSans 480 0 0 0 WW4BEG[7]
port 393 nsew signal tristate
flabel metal3 s 0 12792 160 12912 0 FreeSans 480 0 0 0 WW4BEG[8]
port 394 nsew signal tristate
flabel metal3 s 0 13064 160 13184 0 FreeSans 480 0 0 0 WW4BEG[9]
port 395 nsew signal tristate
rlabel via1 13052 43520 13052 43520 0 VGND
rlabel metal1 12972 42976 12972 42976 0 VPWR
rlabel metal3 24928 9588 24928 9588 0 Config_accessC_bit0
rlabel metal3 24882 10132 24882 10132 0 Config_accessC_bit1
rlabel metal3 25204 10676 25204 10676 0 Config_accessC_bit2
rlabel metal1 24794 9622 24794 9622 0 Config_accessC_bit3
rlabel metal3 1441 18292 1441 18292 0 E1END[0]
rlabel metal3 452 18564 452 18564 0 E1END[1]
rlabel metal3 544 18836 544 18836 0 E1END[2]
rlabel metal3 452 19108 452 19108 0 E1END[3]
rlabel metal3 590 21556 590 21556 0 E2END[0]
rlabel metal3 498 21828 498 21828 0 E2END[1]
rlabel metal2 1380 21964 1380 21964 0 E2END[2]
rlabel metal3 774 22372 774 22372 0 E2END[3]
rlabel metal3 820 22644 820 22644 0 E2END[4]
rlabel metal3 728 22916 728 22916 0 E2END[5]
rlabel metal2 3450 23443 3450 23443 0 E2END[6]
rlabel metal3 728 23460 728 23460 0 E2END[7]
rlabel metal3 728 19380 728 19380 0 E2MID[0]
rlabel metal3 1740 19652 1740 19652 0 E2MID[1]
rlabel metal3 728 19924 728 19924 0 E2MID[2]
rlabel metal3 682 20196 682 20196 0 E2MID[3]
rlabel metal3 475 20468 475 20468 0 E2MID[4]
rlabel metal3 774 20740 774 20740 0 E2MID[5]
rlabel metal3 866 21012 866 21012 0 E2MID[6]
rlabel metal3 544 21284 544 21284 0 E2MID[7]
rlabel metal3 452 28084 452 28084 0 E6END[0]
rlabel metal3 636 30804 636 30804 0 E6END[10]
rlabel metal3 1763 31076 1763 31076 0 E6END[11]
rlabel metal2 3082 28985 3082 28985 0 E6END[1]
rlabel metal3 682 28628 682 28628 0 E6END[2]
rlabel metal3 912 28900 912 28900 0 E6END[3]
rlabel metal3 2016 29172 2016 29172 0 E6END[4]
rlabel metal3 728 29444 728 29444 0 E6END[5]
rlabel metal3 636 29716 636 29716 0 E6END[6]
rlabel metal3 843 29988 843 29988 0 E6END[7]
rlabel metal3 774 30260 774 30260 0 E6END[8]
rlabel metal3 728 30532 728 30532 0 E6END[9]
rlabel metal3 475 23732 475 23732 0 EE4END[0]
rlabel metal3 774 26452 774 26452 0 EE4END[10]
rlabel metal3 728 26724 728 26724 0 EE4END[11]
rlabel metal3 682 26996 682 26996 0 EE4END[12]
rlabel metal2 2806 27659 2806 27659 0 EE4END[13]
rlabel metal3 751 27540 751 27540 0 EE4END[14]
rlabel metal2 3818 27625 3818 27625 0 EE4END[15]
rlabel metal3 912 24004 912 24004 0 EE4END[1]
rlabel metal3 1050 24276 1050 24276 0 EE4END[2]
rlabel metal3 728 24548 728 24548 0 EE4END[3]
rlabel metal3 728 24820 728 24820 0 EE4END[4]
rlabel metal3 498 25092 498 25092 0 EE4END[5]
rlabel metal3 544 25364 544 25364 0 EE4END[6]
rlabel metal3 774 25636 774 25636 0 EE4END[7]
rlabel metal3 659 25908 659 25908 0 EE4END[8]
rlabel metal3 1326 26180 1326 26180 0 EE4END[9]
rlabel metal3 25503 16116 25503 16116 0 FAB2RAM_A0_O0
rlabel metal1 24380 16218 24380 16218 0 FAB2RAM_A0_O1
rlabel metal3 24974 17204 24974 17204 0 FAB2RAM_A0_O2
rlabel metal3 25411 17748 25411 17748 0 FAB2RAM_A0_O3
rlabel metal1 24472 12954 24472 12954 0 FAB2RAM_A1_O0
rlabel metal3 25158 14484 25158 14484 0 FAB2RAM_A1_O1
rlabel metal3 25227 15028 25227 15028 0 FAB2RAM_A1_O2
rlabel metal3 24836 15572 24836 15572 0 FAB2RAM_A1_O3
rlabel metal3 25158 11764 25158 11764 0 FAB2RAM_C_O0
rlabel metal3 24882 12308 24882 12308 0 FAB2RAM_C_O1
rlabel metal3 24974 12852 24974 12852 0 FAB2RAM_C_O2
rlabel metal3 25296 13396 25296 13396 0 FAB2RAM_C_O3
rlabel metal3 25020 24820 25020 24820 0 FAB2RAM_D0_O0
rlabel metal3 25158 25364 25158 25364 0 FAB2RAM_D0_O1
rlabel metal3 25526 25908 25526 25908 0 FAB2RAM_D0_O2
rlabel metal3 25066 26452 25066 26452 0 FAB2RAM_D0_O3
rlabel metal3 24790 22644 24790 22644 0 FAB2RAM_D1_O0
rlabel metal3 25158 23188 25158 23188 0 FAB2RAM_D1_O1
rlabel metal3 25020 23732 25020 23732 0 FAB2RAM_D1_O2
rlabel metal3 25158 24276 25158 24276 0 FAB2RAM_D1_O3
rlabel metal3 25227 20468 25227 20468 0 FAB2RAM_D2_O0
rlabel metal1 24380 20570 24380 20570 0 FAB2RAM_D2_O1
rlabel metal2 24150 21709 24150 21709 0 FAB2RAM_D2_O2
rlabel metal3 25158 22100 25158 22100 0 FAB2RAM_D2_O3
rlabel metal3 25158 18292 25158 18292 0 FAB2RAM_D3_O0
rlabel metal3 25158 18836 25158 18836 0 FAB2RAM_D3_O1
rlabel metal3 25066 19380 25066 19380 0 FAB2RAM_D3_O2
rlabel metal3 24836 19924 24836 19924 0 FAB2RAM_D3_O3
rlabel metal3 1464 31348 1464 31348 0 FrameData[0]
rlabel metal3 774 34068 774 34068 0 FrameData[10]
rlabel metal3 475 34340 475 34340 0 FrameData[11]
rlabel metal2 2898 35683 2898 35683 0 FrameData[12]
rlabel metal3 728 34884 728 34884 0 FrameData[13]
rlabel metal4 3220 35496 3220 35496 0 FrameData[14]
rlabel metal2 2806 36329 2806 36329 0 FrameData[15]
rlabel metal2 4370 35921 4370 35921 0 FrameData[16]
rlabel metal3 728 35972 728 35972 0 FrameData[17]
rlabel metal2 3082 37315 3082 37315 0 FrameData[18]
rlabel metal2 3266 37179 3266 37179 0 FrameData[19]
rlabel metal3 475 31620 475 31620 0 FrameData[1]
rlabel metal2 3910 37009 3910 37009 0 FrameData[20]
rlabel metal3 866 37060 866 37060 0 FrameData[21]
rlabel metal2 2806 38131 2806 38131 0 FrameData[22]
rlabel metal3 682 37604 682 37604 0 FrameData[23]
rlabel metal1 1426 41480 1426 41480 0 FrameData[24]
rlabel metal3 728 38148 728 38148 0 FrameData[25]
rlabel metal3 820 38420 820 38420 0 FrameData[26]
rlabel metal3 774 38692 774 38692 0 FrameData[27]
rlabel metal2 1472 42602 1472 42602 0 FrameData[28]
rlabel metal3 1234 39236 1234 39236 0 FrameData[29]
rlabel metal3 475 31892 475 31892 0 FrameData[2]
rlabel metal3 774 39508 774 39508 0 FrameData[30]
rlabel metal3 1280 39780 1280 39780 0 FrameData[31]
rlabel metal3 1050 32164 1050 32164 0 FrameData[3]
rlabel metal3 728 32436 728 32436 0 FrameData[4]
rlabel metal3 728 32708 728 32708 0 FrameData[5]
rlabel metal2 2806 33473 2806 33473 0 FrameData[6]
rlabel metal3 1027 33252 1027 33252 0 FrameData[7]
rlabel metal3 866 33524 866 33524 0 FrameData[8]
rlabel metal2 3910 33881 3910 33881 0 FrameData[9]
rlabel metal3 24744 26996 24744 26996 0 FrameData_O[0]
rlabel metal3 25020 32436 25020 32436 0 FrameData_O[10]
rlabel metal3 25503 32980 25503 32980 0 FrameData_O[11]
rlabel metal3 25020 33524 25020 33524 0 FrameData_O[12]
rlabel metal3 25503 34068 25503 34068 0 FrameData_O[13]
rlabel metal3 25066 34612 25066 34612 0 FrameData_O[14]
rlabel metal3 25158 35156 25158 35156 0 FrameData_O[15]
rlabel metal3 25227 35700 25227 35700 0 FrameData_O[16]
rlabel metal3 25158 36244 25158 36244 0 FrameData_O[17]
rlabel metal3 25020 36788 25020 36788 0 FrameData_O[18]
rlabel metal3 25158 37332 25158 37332 0 FrameData_O[19]
rlabel metal3 25158 27540 25158 27540 0 FrameData_O[1]
rlabel metal3 25020 37876 25020 37876 0 FrameData_O[20]
rlabel metal3 25503 38420 25503 38420 0 FrameData_O[21]
rlabel metal3 25020 38964 25020 38964 0 FrameData_O[22]
rlabel metal3 25158 39508 25158 39508 0 FrameData_O[23]
rlabel metal3 25066 40052 25066 40052 0 FrameData_O[24]
rlabel metal3 24790 40596 24790 40596 0 FrameData_O[25]
rlabel metal1 24794 42194 24794 42194 0 FrameData_O[26]
rlabel metal3 24560 41684 24560 41684 0 FrameData_O[27]
rlabel metal3 24974 42228 24974 42228 0 FrameData_O[28]
rlabel metal3 25020 42772 25020 42772 0 FrameData_O[29]
rlabel metal3 25020 28084 25020 28084 0 FrameData_O[2]
rlabel metal1 23644 41786 23644 41786 0 FrameData_O[30]
rlabel metal1 22908 42330 22908 42330 0 FrameData_O[31]
rlabel metal3 25158 28628 25158 28628 0 FrameData_O[3]
rlabel metal3 25066 29172 25066 29172 0 FrameData_O[4]
rlabel metal3 25158 29716 25158 29716 0 FrameData_O[5]
rlabel metal3 25066 30260 25066 30260 0 FrameData_O[6]
rlabel metal3 25158 30804 25158 30804 0 FrameData_O[7]
rlabel metal3 25227 31348 25227 31348 0 FrameData_O[8]
rlabel metal3 25158 31892 25158 31892 0 FrameData_O[9]
rlabel metal2 20431 68 20431 68 0 FrameStrobe[0]
rlabel metal1 23460 3502 23460 3502 0 FrameStrobe[10]
rlabel metal2 23414 2574 23414 2574 0 FrameStrobe[11]
rlabel metal1 23828 4522 23828 4522 0 FrameStrobe[12]
rlabel metal2 23966 670 23966 670 0 FrameStrobe[13]
rlabel metal2 21574 3468 21574 3468 0 FrameStrobe[14]
rlabel metal2 24465 68 24465 68 0 FrameStrobe[15]
rlabel metal2 24695 68 24695 68 0 FrameStrobe[16]
rlabel metal1 24702 5202 24702 5202 0 FrameStrobe[17]
rlabel metal2 25346 976 25346 976 0 FrameStrobe[18]
rlabel metal1 24058 3706 24058 3706 0 FrameStrobe[19]
rlabel metal2 20654 755 20654 755 0 FrameStrobe[1]
rlabel metal2 20877 68 20877 68 0 FrameStrobe[2]
rlabel metal2 22494 952 22494 952 0 FrameStrobe[3]
rlabel metal2 21429 68 21429 68 0 FrameStrobe[4]
rlabel metal2 21659 68 21659 68 0 FrameStrobe[5]
rlabel metal2 22034 755 22034 755 0 FrameStrobe[6]
rlabel metal1 22264 3026 22264 3026 0 FrameStrobe[7]
rlabel metal2 22639 68 22639 68 0 FrameStrobe[8]
rlabel metal2 22862 500 22862 500 0 FrameStrobe[9]
rlabel metal2 20431 44948 20431 44948 0 FrameStrobe_O[0]
rlabel metal2 23138 44176 23138 44176 0 FrameStrobe_O[10]
rlabel metal2 23414 44261 23414 44261 0 FrameStrobe_O[11]
rlabel metal1 23046 42262 23046 42262 0 FrameStrobe_O[12]
rlabel metal2 23966 43360 23966 43360 0 FrameStrobe_O[13]
rlabel metal1 23782 42330 23782 42330 0 FrameStrobe_O[14]
rlabel metal2 24419 44948 24419 44948 0 FrameStrobe_O[15]
rlabel metal1 23828 41718 23828 41718 0 FrameStrobe_O[16]
rlabel metal2 25070 43734 25070 43734 0 FrameStrobe_O[17]
rlabel metal1 24472 40698 24472 40698 0 FrameStrobe_O[18]
rlabel metal1 25622 42092 25622 42092 0 FrameStrobe_O[19]
rlabel metal2 20654 44176 20654 44176 0 FrameStrobe_O[1]
rlabel metal1 21298 43078 21298 43078 0 FrameStrobe_O[2]
rlabel metal2 21206 44533 21206 44533 0 FrameStrobe_O[3]
rlabel metal1 22586 43384 22586 43384 0 FrameStrobe_O[4]
rlabel metal2 21857 44948 21857 44948 0 FrameStrobe_O[5]
rlabel metal2 22126 42925 22126 42925 0 FrameStrobe_O[6]
rlabel metal2 22310 43836 22310 43836 0 FrameStrobe_O[7]
rlabel metal1 22586 43248 22586 43248 0 FrameStrobe_O[8]
rlabel metal2 22862 43853 22862 43853 0 FrameStrobe_O[9]
rlabel metal2 24150 8874 24150 8874 0 Inst_Config_accessConfig_access.ConfigBits\[0\]
rlabel metal1 22402 11084 22402 11084 0 Inst_Config_accessConfig_access.ConfigBits\[1\]
rlabel metal1 22678 11220 22678 11220 0 Inst_Config_accessConfig_access.ConfigBits\[2\]
rlabel metal1 22632 11730 22632 11730 0 Inst_Config_accessConfig_access.ConfigBits\[3\]
rlabel metal1 19964 17850 19964 17850 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 21758 18258 21758 18258 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 23598 16966 23598 16966 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 23736 21658 23736 21658 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18160 18258 18160 18258 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 9338 20434 9338 20434 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 19642 18088 19642 18088 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 20102 21896 20102 21896 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 19780 18258 19780 18258 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 22034 18224 22034 18224 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 22586 17612 22586 17612 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[2\]
rlabel metal2 23782 21182 23782 21182 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 18906 17850 18906 17850 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 19780 18394 19780 18394 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal2 19550 17612 19550 17612 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal2 19734 17850 19734 17850 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 21298 18768 21298 18768 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 22678 18190 22678 18190 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal2 21942 18428 21942 18428 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 22356 18190 22356 18190 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 23000 18258 23000 18258 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 23506 16592 23506 16592 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 24150 17102 24150 17102 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 24150 16762 24150 16762 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 22908 20910 22908 20910 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 23368 20570 23368 20570 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 23828 21114 23828 21114 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 23966 21454 23966 21454 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 22402 13294 22402 13294 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 23000 15878 23000 15878 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 23460 18734 23460 18734 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 21022 19822 21022 19822 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 21206 13906 21206 13906 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[0\]
rlabel via1 21293 16558 21293 16558 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[1\]
rlabel metal2 19366 24259 19366 24259 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[2\]
rlabel viali 19448 20502 19448 20502 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 22678 14348 22678 14348 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 22816 16558 22816 16558 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 23322 18700 23322 18700 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 21114 20400 21114 20400 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[3\]
rlabel metal2 22218 14212 22218 14212 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 23138 13328 23138 13328 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal2 22310 13872 22310 13872 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 22494 13430 22494 13430 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal2 22494 16762 22494 16762 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 23230 16524 23230 16524 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 22954 15674 22954 15674 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 23460 15538 23460 15538 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 22816 18734 22816 18734 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 23552 18258 23552 18258 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 23230 18870 23230 18870 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 23644 18394 23644 18394 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 20194 20434 20194 20434 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 21758 19890 21758 19890 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 21022 20026 21022 20026 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 21574 19890 21574 19890 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 20102 13345 20102 13345 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 22908 31654 22908 31654 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 22724 38182 22724 38182 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 21022 15470 21022 15470 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18431 14994 18431 14994 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 21666 32436 21666 32436 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 17418 38250 17418 38250 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 19131 16150 19131 16150 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 19826 14382 19826 14382 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 23368 32538 23368 32538 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[1\]
rlabel metal2 22494 38726 22494 38726 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 21022 16116 21022 16116 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 19366 14348 19366 14348 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 20286 13770 20286 13770 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19780 13498 19780 13498 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 20102 13362 20102 13362 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal2 21482 32096 21482 32096 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 23368 31790 23368 31790 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 22770 31824 22770 31824 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 23138 31824 23138 31824 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 21850 38964 21850 38964 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 22778 39001 22778 39001 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel via1 22402 38709 22402 38709 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 22770 37910 22770 37910 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 20056 15674 20056 15674 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 21758 15538 21758 15538 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 20976 15674 20976 15674 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 21574 15538 21574 15538 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 20516 24582 20516 24582 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 22218 28560 22218 28560 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 19228 35054 19228 35054 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 20194 27846 20194 27846 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18390 24786 18390 24786 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 7222 28424 7222 28424 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[1\]
rlabel via1 17981 35666 17981 35666 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 18384 28118 18384 28118 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 19964 24922 19964 24922 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 23046 28458 23046 28458 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 19274 35802 19274 35802 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 19688 28186 19688 28186 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 19734 24140 19734 24140 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 20562 25228 20562 25228 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19964 24242 19964 24242 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 20332 24242 20332 24242 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 22310 27982 22310 27982 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 22724 28730 22724 28730 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 22494 28458 22494 28458 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal2 22494 28764 22494 28764 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 18722 36108 18722 36108 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 19412 35054 19412 35054 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal2 19274 35904 19274 35904 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 19412 35258 19412 35258 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 19366 27404 19366 27404 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 20194 28492 20194 28492 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 19688 27506 19688 27506 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal2 20102 27948 20102 27948 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 22402 26554 22402 26554 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal2 23506 24310 23506 24310 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 19136 33490 19136 33490 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 20884 30226 20884 30226 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18982 26282 18982 26282 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[0\]
rlabel via2 4738 24667 4738 24667 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 17832 32810 17832 32810 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 19826 29580 19826 29580 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[3\]
rlabel metal2 21390 26758 21390 26758 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 23322 24378 23322 24378 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 19504 32402 19504 32402 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 21666 30260 21666 30260 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 21114 25840 21114 25840 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 21850 27064 21850 27064 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 21574 25670 21574 25670 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 22172 25806 22172 25806 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 23506 24242 23506 24242 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 23782 24752 23782 24752 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 23782 23290 23782 23290 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 24150 23188 24150 23188 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 18722 33456 18722 33456 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 19550 32538 19550 32538 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 18998 33286 18998 33286 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 19458 33422 19458 33422 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 20424 29478 20424 29478 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal2 21482 30532 21482 30532 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 21114 30090 21114 30090 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel viali 21112 30188 21112 30188 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 22172 21114 22172 21114 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 23782 25874 23782 25874 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 21620 35258 21620 35258 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 19136 30362 19136 30362 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 20792 21522 20792 21522 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[0\]
rlabel metal2 18262 27761 18262 27761 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 19810 35734 19810 35734 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 17981 30702 17981 30702 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 21850 21998 21850 21998 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 23736 25262 23736 25262 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 21984 35670 21984 35670 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 20010 30736 20010 30736 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 21482 21488 21482 21488 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 21896 22100 21896 22100 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 21758 21318 21758 21318 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 22218 21454 22218 21454 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 22908 25874 22908 25874 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 23460 25466 23460 25466 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 23414 25738 23414 25738 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 23644 25806 23644 25806 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel viali 21482 35665 21482 35665 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 22310 35598 22310 35598 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 21252 35530 21252 35530 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 21804 35598 21804 35598 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 18952 30702 18952 30702 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 19780 30702 19780 30702 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 19366 30192 19366 30192 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 19596 29682 19596 29682 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 19734 22032 19734 22032 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 21758 23698 21758 23698 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 20746 32810 20746 32810 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 18860 25874 18860 25874 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18584 21998 18584 21998 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 20270 24106 20270 24106 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 19826 33490 19826 33490 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 18078 26350 18078 26350 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 20102 22576 20102 22576 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 21712 24378 21712 24378 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 21528 32878 21528 32878 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 19918 25942 19918 25942 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 19182 21862 19182 21862 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 20378 22644 20378 22644 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19780 22202 19780 22202 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 20148 22134 20148 22134 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 21482 23732 21482 23732 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal2 22402 24140 22402 24140 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 21758 23494 21758 23494 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 22218 23630 22218 23630 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 20194 33558 20194 33558 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 21344 32878 21344 32878 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal2 20838 33184 20838 33184 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 21114 32946 21114 32946 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 18446 26384 18446 26384 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 19688 25874 19688 25874 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 19182 25908 19182 25908 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 19458 25806 19458 25806 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 20470 7854 20470 7854 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20378 8908 20378 8908 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal2 23322 8500 23322 8500 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 22586 10098 22586 10098 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal2 16192 13260 16192 13260 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[0\]
rlabel metal1 6946 15062 6946 15062 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[1\]
rlabel metal1 1840 17646 1840 17646 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[2\]
rlabel metal2 15318 10489 15318 10489 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[3\]
rlabel metal1 21206 7412 21206 7412 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 21666 8602 21666 8602 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[1\]
rlabel metal2 22034 7633 22034 7633 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[2\]
rlabel metal2 23230 10166 23230 10166 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 18998 7412 18998 7412 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 20884 7514 20884 7514 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19412 7514 19412 7514 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 20286 7888 20286 7888 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 20792 7174 20792 7174 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 21620 8942 21620 8942 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 20562 8976 20562 8976 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 21114 8976 21114 8976 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal2 23690 8024 23690 8024 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 22310 7344 22310 7344 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 23230 8602 23230 8602 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal2 24058 8228 24058 8228 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 21620 9690 21620 9690 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 22770 10064 22770 10064 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 22402 10438 22402 10438 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal2 22678 10438 22678 10438 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 19366 10812 19366 10812 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20838 12410 20838 12410 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal2 16330 3791 16330 3791 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal2 22126 7004 22126 7004 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 16146 13158 16146 13158 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[0\]
rlabel metal1 14214 11696 14214 11696 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[1\]
rlabel metal1 2300 18190 2300 18190 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[2\]
rlabel metal3 15548 6120 15548 6120 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[3\]
rlabel metal1 19596 9690 19596 9690 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 22218 11798 22218 11798 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 21114 6324 21114 6324 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 22862 6970 22862 6970 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 18998 10030 18998 10030 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 19550 10438 19550 10438 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 18860 10234 18860 10234 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 19366 10710 19366 10710 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 20930 12784 20930 12784 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 21620 11866 21620 11866 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal2 21022 12172 21022 12172 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal2 21344 11730 21344 11730 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 20470 5882 20470 5882 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 16514 3094 16514 3094 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 21068 6426 21068 6426 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 16514 2822 16514 2822 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal2 21298 7140 21298 7140 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 22494 7378 22494 7378 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 22218 6732 22218 6732 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 22494 6290 22494 6290 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 18308 6630 18308 6630 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel via1 20010 5066 20010 5066 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 18906 13328 18906 13328 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 20792 10438 20792 10438 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18262 7208 18262 7208 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[0\]
rlabel metal1 16974 4624 16974 4624 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[1\]
rlabel metal1 1702 17612 1702 17612 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[2\]
rlabel metal1 17526 5644 17526 5644 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[3\]
rlabel metal1 19136 6290 19136 6290 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 20102 4250 20102 4250 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 19504 12818 19504 12818 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 21758 4726 21758 4726 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 17986 6426 17986 6426 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 19136 6426 19136 6426 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 18492 6970 18492 6970 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 18722 7378 18722 7378 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 19734 4556 19734 4556 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal2 20194 4658 20194 4658 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal2 19826 4998 19826 4998 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 20424 4794 20424 4794 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 17710 12784 17710 12784 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal2 19458 13124 19458 13124 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 18170 13328 18170 13328 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 18768 13226 18768 13226 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 21298 5236 21298 5236 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 21206 5168 21206 5168 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 21344 5338 21344 5338 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 20976 5134 20976 5134 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 17940 4114 17940 4114 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 23506 15130 23506 15130 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 17802 3570 17802 3570 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 23092 5134 23092 5134 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 14766 4114 14766 4114 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[0\]
rlabel metal1 1932 15538 1932 15538 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[1\]
rlabel metal2 1794 4675 1794 4675 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[2\]
rlabel metal2 7866 6052 7866 6052 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[3\]
rlabel metal2 19504 3162 19504 3162 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 23414 14586 23414 14586 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 15778 2482 15778 2482 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 24058 1972 24058 1972 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 18170 3162 18170 3162 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 18446 3468 18446 3468 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 18400 3570 18400 3570 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 18216 4114 18216 4114 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 22678 13260 22678 13260 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 22770 15130 22770 15130 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal2 23690 14654 23690 14654 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 24150 13974 24150 13974 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal2 19734 5015 19734 5015 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 15594 2312 15594 2312 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal2 21666 4250 21666 4250 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel via2 17894 3451 17894 3451 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 18630 4556 18630 4556 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 23920 2074 23920 2074 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 18722 5032 18722 5032 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal2 23782 5678 23782 5678 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 13754 21930 13754 21930 0 Inst_RAM_IO_ConfigMem.ConfigBits\[100\]
rlabel metal1 13616 21862 13616 21862 0 Inst_RAM_IO_ConfigMem.ConfigBits\[101\]
rlabel metal2 5474 20570 5474 20570 0 Inst_RAM_IO_ConfigMem.ConfigBits\[102\]
rlabel metal1 5750 20026 5750 20026 0 Inst_RAM_IO_ConfigMem.ConfigBits\[103\]
rlabel metal2 8326 26724 8326 26724 0 Inst_RAM_IO_ConfigMem.ConfigBits\[104\]
rlabel metal1 8234 27030 8234 27030 0 Inst_RAM_IO_ConfigMem.ConfigBits\[105\]
rlabel metal1 15042 18938 15042 18938 0 Inst_RAM_IO_ConfigMem.ConfigBits\[106\]
rlabel metal2 15502 19516 15502 19516 0 Inst_RAM_IO_ConfigMem.ConfigBits\[107\]
rlabel metal1 14720 25330 14720 25330 0 Inst_RAM_IO_ConfigMem.ConfigBits\[108\]
rlabel metal2 15318 25755 15318 25755 0 Inst_RAM_IO_ConfigMem.ConfigBits\[109\]
rlabel metal2 18078 23868 18078 23868 0 Inst_RAM_IO_ConfigMem.ConfigBits\[110\]
rlabel metal2 5014 23052 5014 23052 0 Inst_RAM_IO_ConfigMem.ConfigBits\[111\]
rlabel metal1 5704 23290 5704 23290 0 Inst_RAM_IO_ConfigMem.ConfigBits\[112\]
rlabel metal1 7314 22406 7314 22406 0 Inst_RAM_IO_ConfigMem.ConfigBits\[113\]
rlabel metal1 10304 29682 10304 29682 0 Inst_RAM_IO_ConfigMem.ConfigBits\[114\]
rlabel metal1 10902 30158 10902 30158 0 Inst_RAM_IO_ConfigMem.ConfigBits\[115\]
rlabel metal1 12926 29750 12926 29750 0 Inst_RAM_IO_ConfigMem.ConfigBits\[116\]
rlabel metal1 16560 21046 16560 21046 0 Inst_RAM_IO_ConfigMem.ConfigBits\[117\]
rlabel metal2 17618 20740 17618 20740 0 Inst_RAM_IO_ConfigMem.ConfigBits\[118\]
rlabel metal1 18630 20026 18630 20026 0 Inst_RAM_IO_ConfigMem.ConfigBits\[119\]
rlabel metal2 10166 5338 10166 5338 0 Inst_RAM_IO_ConfigMem.ConfigBits\[120\]
rlabel metal1 10994 5134 10994 5134 0 Inst_RAM_IO_ConfigMem.ConfigBits\[121\]
rlabel metal1 3128 20774 3128 20774 0 Inst_RAM_IO_ConfigMem.ConfigBits\[122\]
rlabel metal2 3266 20876 3266 20876 0 Inst_RAM_IO_ConfigMem.ConfigBits\[123\]
rlabel metal1 9890 8058 9890 8058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[124\]
rlabel metal2 10534 8772 10534 8772 0 Inst_RAM_IO_ConfigMem.ConfigBits\[125\]
rlabel metal1 13800 5066 13800 5066 0 Inst_RAM_IO_ConfigMem.ConfigBits\[126\]
rlabel metal1 14996 4794 14996 4794 0 Inst_RAM_IO_ConfigMem.ConfigBits\[127\]
rlabel metal1 11132 6834 11132 6834 0 Inst_RAM_IO_ConfigMem.ConfigBits\[128\]
rlabel metal2 11730 7242 11730 7242 0 Inst_RAM_IO_ConfigMem.ConfigBits\[129\]
rlabel metal1 6072 5338 6072 5338 0 Inst_RAM_IO_ConfigMem.ConfigBits\[130\]
rlabel metal2 7406 5542 7406 5542 0 Inst_RAM_IO_ConfigMem.ConfigBits\[131\]
rlabel metal1 2438 11288 2438 11288 0 Inst_RAM_IO_ConfigMem.ConfigBits\[132\]
rlabel metal1 3220 10778 3220 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[133\]
rlabel metal2 4370 5746 4370 5746 0 Inst_RAM_IO_ConfigMem.ConfigBits\[134\]
rlabel metal1 5014 5882 5014 5882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[135\]
rlabel metal1 15778 5814 15778 5814 0 Inst_RAM_IO_ConfigMem.ConfigBits\[136\]
rlabel metal1 16744 5746 16744 5746 0 Inst_RAM_IO_ConfigMem.ConfigBits\[137\]
rlabel metal2 2714 12546 2714 12546 0 Inst_RAM_IO_ConfigMem.ConfigBits\[138\]
rlabel metal1 3634 12750 3634 12750 0 Inst_RAM_IO_ConfigMem.ConfigBits\[139\]
rlabel metal1 2576 3706 2576 3706 0 Inst_RAM_IO_ConfigMem.ConfigBits\[140\]
rlabel metal2 2990 5916 2990 5916 0 Inst_RAM_IO_ConfigMem.ConfigBits\[141\]
rlabel metal1 7682 3706 7682 3706 0 Inst_RAM_IO_ConfigMem.ConfigBits\[142\]
rlabel metal2 8786 4284 8786 4284 0 Inst_RAM_IO_ConfigMem.ConfigBits\[143\]
rlabel metal2 11178 5474 11178 5474 0 Inst_RAM_IO_ConfigMem.ConfigBits\[144\]
rlabel metal1 12328 5882 12328 5882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[145\]
rlabel metal1 5612 7990 5612 7990 0 Inst_RAM_IO_ConfigMem.ConfigBits\[146\]
rlabel metal1 7038 7922 7038 7922 0 Inst_RAM_IO_ConfigMem.ConfigBits\[147\]
rlabel metal1 2392 17782 2392 17782 0 Inst_RAM_IO_ConfigMem.ConfigBits\[148\]
rlabel metal2 2806 18020 2806 18020 0 Inst_RAM_IO_ConfigMem.ConfigBits\[149\]
rlabel metal1 3496 3978 3496 3978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[150\]
rlabel metal1 4692 3706 4692 3706 0 Inst_RAM_IO_ConfigMem.ConfigBits\[151\]
rlabel metal1 15548 3706 15548 3706 0 Inst_RAM_IO_ConfigMem.ConfigBits\[152\]
rlabel metal2 17066 3876 17066 3876 0 Inst_RAM_IO_ConfigMem.ConfigBits\[153\]
rlabel metal1 2484 15606 2484 15606 0 Inst_RAM_IO_ConfigMem.ConfigBits\[154\]
rlabel metal1 3082 15130 3082 15130 0 Inst_RAM_IO_ConfigMem.ConfigBits\[155\]
rlabel metal2 2806 8602 2806 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[156\]
rlabel metal2 3266 8262 3266 8262 0 Inst_RAM_IO_ConfigMem.ConfigBits\[157\]
rlabel metal1 8096 2618 8096 2618 0 Inst_RAM_IO_ConfigMem.ConfigBits\[158\]
rlabel metal2 8786 3196 8786 3196 0 Inst_RAM_IO_ConfigMem.ConfigBits\[159\]
rlabel metal1 17434 8602 17434 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[160\]
rlabel metal2 17664 8942 17664 8942 0 Inst_RAM_IO_ConfigMem.ConfigBits\[161\]
rlabel metal2 5566 10370 5566 10370 0 Inst_RAM_IO_ConfigMem.ConfigBits\[162\]
rlabel via2 6946 10251 6946 10251 0 Inst_RAM_IO_ConfigMem.ConfigBits\[163\]
rlabel metal1 4600 11254 4600 11254 0 Inst_RAM_IO_ConfigMem.ConfigBits\[164\]
rlabel metal1 5198 10778 5198 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[165\]
rlabel metal1 8970 9690 8970 9690 0 Inst_RAM_IO_ConfigMem.ConfigBits\[166\]
rlabel metal1 9936 9690 9936 9690 0 Inst_RAM_IO_ConfigMem.ConfigBits\[167\]
rlabel metal1 16054 10778 16054 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[168\]
rlabel metal1 17158 11254 17158 11254 0 Inst_RAM_IO_ConfigMem.ConfigBits\[169\]
rlabel metal1 5796 12410 5796 12410 0 Inst_RAM_IO_ConfigMem.ConfigBits\[170\]
rlabel metal1 7268 12614 7268 12614 0 Inst_RAM_IO_ConfigMem.ConfigBits\[171\]
rlabel metal1 4094 13430 4094 13430 0 Inst_RAM_IO_ConfigMem.ConfigBits\[172\]
rlabel metal2 5014 13532 5014 13532 0 Inst_RAM_IO_ConfigMem.ConfigBits\[173\]
rlabel metal2 10166 12682 10166 12682 0 Inst_RAM_IO_ConfigMem.ConfigBits\[174\]
rlabel metal1 10672 11866 10672 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[175\]
rlabel metal1 17526 11594 17526 11594 0 Inst_RAM_IO_ConfigMem.ConfigBits\[176\]
rlabel metal1 19090 11662 19090 11662 0 Inst_RAM_IO_ConfigMem.ConfigBits\[177\]
rlabel metal1 7452 7514 7452 7514 0 Inst_RAM_IO_ConfigMem.ConfigBits\[178\]
rlabel metal1 8050 8602 8050 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[179\]
rlabel metal2 2806 18360 2806 18360 0 Inst_RAM_IO_ConfigMem.ConfigBits\[180\]
rlabel metal2 3266 18700 3266 18700 0 Inst_RAM_IO_ConfigMem.ConfigBits\[181\]
rlabel metal1 9062 13430 9062 13430 0 Inst_RAM_IO_ConfigMem.ConfigBits\[182\]
rlabel metal2 9706 13770 9706 13770 0 Inst_RAM_IO_ConfigMem.ConfigBits\[183\]
rlabel metal1 16100 7990 16100 7990 0 Inst_RAM_IO_ConfigMem.ConfigBits\[184\]
rlabel metal1 17158 7514 17158 7514 0 Inst_RAM_IO_ConfigMem.ConfigBits\[185\]
rlabel metal2 7406 15130 7406 15130 0 Inst_RAM_IO_ConfigMem.ConfigBits\[186\]
rlabel metal1 8004 14586 8004 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[187\]
rlabel metal1 4462 9112 4462 9112 0 Inst_RAM_IO_ConfigMem.ConfigBits\[188\]
rlabel metal1 5060 8602 5060 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[189\]
rlabel metal1 8372 6222 8372 6222 0 Inst_RAM_IO_ConfigMem.ConfigBits\[190\]
rlabel metal2 9062 6460 9062 6460 0 Inst_RAM_IO_ConfigMem.ConfigBits\[191\]
rlabel metal1 14996 14586 14996 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[192\]
rlabel metal1 16376 14586 16376 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[193\]
rlabel metal2 6762 39950 6762 39950 0 Inst_RAM_IO_ConfigMem.ConfigBits\[194\]
rlabel metal1 7406 39474 7406 39474 0 Inst_RAM_IO_ConfigMem.ConfigBits\[195\]
rlabel metal1 4830 39576 4830 39576 0 Inst_RAM_IO_ConfigMem.ConfigBits\[196\]
rlabel metal1 5658 39474 5658 39474 0 Inst_RAM_IO_ConfigMem.ConfigBits\[197\]
rlabel metal2 13294 12954 13294 12954 0 Inst_RAM_IO_ConfigMem.ConfigBits\[198\]
rlabel via1 13846 12835 13846 12835 0 Inst_RAM_IO_ConfigMem.ConfigBits\[199\]
rlabel metal1 16284 13430 16284 13430 0 Inst_RAM_IO_ConfigMem.ConfigBits\[200\]
rlabel metal1 17296 13362 17296 13362 0 Inst_RAM_IO_ConfigMem.ConfigBits\[201\]
rlabel metal1 7728 11866 7728 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[202\]
rlabel metal1 8694 11866 8694 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[203\]
rlabel metal1 3956 15946 3956 15946 0 Inst_RAM_IO_ConfigMem.ConfigBits\[204\]
rlabel metal2 5014 16252 5014 16252 0 Inst_RAM_IO_ConfigMem.ConfigBits\[205\]
rlabel metal1 10074 15640 10074 15640 0 Inst_RAM_IO_ConfigMem.ConfigBits\[206\]
rlabel metal1 10672 15130 10672 15130 0 Inst_RAM_IO_ConfigMem.ConfigBits\[207\]
rlabel metal1 16146 16694 16146 16694 0 Inst_RAM_IO_ConfigMem.ConfigBits\[208\]
rlabel metal1 17066 16626 17066 16626 0 Inst_RAM_IO_ConfigMem.ConfigBits\[209\]
rlabel metal2 8326 16354 8326 16354 0 Inst_RAM_IO_ConfigMem.ConfigBits\[210\]
rlabel metal2 8878 16524 8878 16524 0 Inst_RAM_IO_ConfigMem.ConfigBits\[211\]
rlabel metal1 4600 18190 4600 18190 0 Inst_RAM_IO_ConfigMem.ConfigBits\[212\]
rlabel metal2 5198 18428 5198 18428 0 Inst_RAM_IO_ConfigMem.ConfigBits\[213\]
rlabel metal2 9706 18020 9706 18020 0 Inst_RAM_IO_ConfigMem.ConfigBits\[214\]
rlabel metal1 10396 17306 10396 17306 0 Inst_RAM_IO_ConfigMem.ConfigBits\[215\]
rlabel metal2 12558 25806 12558 25806 0 Inst_RAM_IO_ConfigMem.ConfigBits\[216\]
rlabel metal2 13202 25075 13202 25075 0 Inst_RAM_IO_ConfigMem.ConfigBits\[217\]
rlabel metal1 3588 28662 3588 28662 0 Inst_RAM_IO_ConfigMem.ConfigBits\[218\]
rlabel metal1 4232 28186 4232 28186 0 Inst_RAM_IO_ConfigMem.ConfigBits\[219\]
rlabel metal1 10856 35190 10856 35190 0 Inst_RAM_IO_ConfigMem.ConfigBits\[220\]
rlabel metal2 11362 35530 11362 35530 0 Inst_RAM_IO_ConfigMem.ConfigBits\[221\]
rlabel metal1 15916 27914 15916 27914 0 Inst_RAM_IO_ConfigMem.ConfigBits\[222\]
rlabel metal2 16514 29172 16514 29172 0 Inst_RAM_IO_ConfigMem.ConfigBits\[223\]
rlabel metal1 13984 26486 13984 26486 0 Inst_RAM_IO_ConfigMem.ConfigBits\[224\]
rlabel metal2 15318 26486 15318 26486 0 Inst_RAM_IO_ConfigMem.ConfigBits\[225\]
rlabel metal2 3358 24922 3358 24922 0 Inst_RAM_IO_ConfigMem.ConfigBits\[226\]
rlabel metal1 4324 24378 4324 24378 0 Inst_RAM_IO_ConfigMem.ConfigBits\[227\]
rlabel metal1 10350 31960 10350 31960 0 Inst_RAM_IO_ConfigMem.ConfigBits\[228\]
rlabel metal1 10994 31858 10994 31858 0 Inst_RAM_IO_ConfigMem.ConfigBits\[229\]
rlabel metal1 17802 28186 17802 28186 0 Inst_RAM_IO_ConfigMem.ConfigBits\[230\]
rlabel metal2 18446 28730 18446 28730 0 Inst_RAM_IO_ConfigMem.ConfigBits\[231\]
rlabel metal2 12282 24038 12282 24038 0 Inst_RAM_IO_ConfigMem.ConfigBits\[232\]
rlabel metal2 12880 24174 12880 24174 0 Inst_RAM_IO_ConfigMem.ConfigBits\[233\]
rlabel metal2 5106 28866 5106 28866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[234\]
rlabel metal1 5658 28934 5658 28934 0 Inst_RAM_IO_ConfigMem.ConfigBits\[235\]
rlabel metal1 10074 35530 10074 35530 0 Inst_RAM_IO_ConfigMem.ConfigBits\[236\]
rlabel metal1 10999 35598 10999 35598 0 Inst_RAM_IO_ConfigMem.ConfigBits\[237\]
rlabel metal1 15778 30362 15778 30362 0 Inst_RAM_IO_ConfigMem.ConfigBits\[238\]
rlabel metal2 16514 30940 16514 30940 0 Inst_RAM_IO_ConfigMem.ConfigBits\[239\]
rlabel metal1 14076 26894 14076 26894 0 Inst_RAM_IO_ConfigMem.ConfigBits\[240\]
rlabel metal2 14766 27132 14766 27132 0 Inst_RAM_IO_ConfigMem.ConfigBits\[241\]
rlabel metal2 4830 26282 4830 26282 0 Inst_RAM_IO_ConfigMem.ConfigBits\[242\]
rlabel metal2 4554 26078 4554 26078 0 Inst_RAM_IO_ConfigMem.ConfigBits\[243\]
rlabel metal2 12282 33218 12282 33218 0 Inst_RAM_IO_ConfigMem.ConfigBits\[244\]
rlabel metal1 13018 33422 13018 33422 0 Inst_RAM_IO_ConfigMem.ConfigBits\[245\]
rlabel metal1 16468 26010 16468 26010 0 Inst_RAM_IO_ConfigMem.ConfigBits\[246\]
rlabel metal1 17572 26418 17572 26418 0 Inst_RAM_IO_ConfigMem.ConfigBits\[247\]
rlabel metal1 16330 18394 16330 18394 0 Inst_RAM_IO_ConfigMem.ConfigBits\[248\]
rlabel metal1 17342 18802 17342 18802 0 Inst_RAM_IO_ConfigMem.ConfigBits\[249\]
rlabel metal2 7682 21148 7682 21148 0 Inst_RAM_IO_ConfigMem.ConfigBits\[250\]
rlabel metal1 8188 20570 8188 20570 0 Inst_RAM_IO_ConfigMem.ConfigBits\[251\]
rlabel metal1 6118 17850 6118 17850 0 Inst_RAM_IO_ConfigMem.ConfigBits\[252\]
rlabel metal1 6900 17850 6900 17850 0 Inst_RAM_IO_ConfigMem.ConfigBits\[253\]
rlabel metal2 15134 22270 15134 22270 0 Inst_RAM_IO_ConfigMem.ConfigBits\[254\]
rlabel metal1 15732 21658 15732 21658 0 Inst_RAM_IO_ConfigMem.ConfigBits\[255\]
rlabel metal1 16100 23222 16100 23222 0 Inst_RAM_IO_ConfigMem.ConfigBits\[256\]
rlabel metal2 16606 23290 16606 23290 0 Inst_RAM_IO_ConfigMem.ConfigBits\[257\]
rlabel metal2 8418 22746 8418 22746 0 Inst_RAM_IO_ConfigMem.ConfigBits\[258\]
rlabel metal1 8832 21658 8832 21658 0 Inst_RAM_IO_ConfigMem.ConfigBits\[259\]
rlabel metal1 5750 25364 5750 25364 0 Inst_RAM_IO_ConfigMem.ConfigBits\[260\]
rlabel metal1 7360 24922 7360 24922 0 Inst_RAM_IO_ConfigMem.ConfigBits\[261\]
rlabel metal2 12558 21216 12558 21216 0 Inst_RAM_IO_ConfigMem.ConfigBits\[262\]
rlabel metal1 12742 20944 12742 20944 0 Inst_RAM_IO_ConfigMem.ConfigBits\[263\]
rlabel metal2 13478 18394 13478 18394 0 Inst_RAM_IO_ConfigMem.ConfigBits\[264\]
rlabel metal2 14030 18700 14030 18700 0 Inst_RAM_IO_ConfigMem.ConfigBits\[265\]
rlabel metal1 4048 33286 4048 33286 0 Inst_RAM_IO_ConfigMem.ConfigBits\[266\]
rlabel metal1 4600 32538 4600 32538 0 Inst_RAM_IO_ConfigMem.ConfigBits\[267\]
rlabel metal1 12742 38488 12742 38488 0 Inst_RAM_IO_ConfigMem.ConfigBits\[268\]
rlabel metal1 13524 37978 13524 37978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[269\]
rlabel metal1 17710 15912 17710 15912 0 Inst_RAM_IO_ConfigMem.ConfigBits\[270\]
rlabel metal1 18354 16014 18354 16014 0 Inst_RAM_IO_ConfigMem.ConfigBits\[271\]
rlabel metal1 11960 9894 11960 9894 0 Inst_RAM_IO_ConfigMem.ConfigBits\[272\]
rlabel metal2 12282 9350 12282 9350 0 Inst_RAM_IO_ConfigMem.ConfigBits\[273\]
rlabel metal2 3450 35292 3450 35292 0 Inst_RAM_IO_ConfigMem.ConfigBits\[274\]
rlabel metal1 4232 34714 4232 34714 0 Inst_RAM_IO_ConfigMem.ConfigBits\[275\]
rlabel metal2 8510 37978 8510 37978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[276\]
rlabel metal1 9844 37434 9844 37434 0 Inst_RAM_IO_ConfigMem.ConfigBits\[277\]
rlabel metal1 13800 7514 13800 7514 0 Inst_RAM_IO_ConfigMem.ConfigBits\[278\]
rlabel metal1 14674 7514 14674 7514 0 Inst_RAM_IO_ConfigMem.ConfigBits\[279\]
rlabel metal1 10810 12308 10810 12308 0 Inst_RAM_IO_ConfigMem.ConfigBits\[280\]
rlabel metal2 11822 12206 11822 12206 0 Inst_RAM_IO_ConfigMem.ConfigBits\[281\]
rlabel metal2 3358 36516 3358 36516 0 Inst_RAM_IO_ConfigMem.ConfigBits\[282\]
rlabel metal1 3542 36856 3542 36856 0 Inst_RAM_IO_ConfigMem.ConfigBits\[283\]
rlabel metal1 8280 35258 8280 35258 0 Inst_RAM_IO_ConfigMem.ConfigBits\[284\]
rlabel metal1 8740 34714 8740 34714 0 Inst_RAM_IO_ConfigMem.ConfigBits\[285\]
rlabel metal1 14352 11866 14352 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[286\]
rlabel metal1 15134 12206 15134 12206 0 Inst_RAM_IO_ConfigMem.ConfigBits\[287\]
rlabel metal1 11776 14586 11776 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[288\]
rlabel metal2 12098 15198 12098 15198 0 Inst_RAM_IO_ConfigMem.ConfigBits\[289\]
rlabel metal1 3312 40358 3312 40358 0 Inst_RAM_IO_ConfigMem.ConfigBits\[290\]
rlabel metal1 3726 40086 3726 40086 0 Inst_RAM_IO_ConfigMem.ConfigBits\[291\]
rlabel metal2 8510 40154 8510 40154 0 Inst_RAM_IO_ConfigMem.ConfigBits\[292\]
rlabel metal1 9568 41990 9568 41990 0 Inst_RAM_IO_ConfigMem.ConfigBits\[293\]
rlabel metal2 13662 10404 13662 10404 0 Inst_RAM_IO_ConfigMem.ConfigBits\[294\]
rlabel metal1 14628 10234 14628 10234 0 Inst_RAM_IO_ConfigMem.ConfigBits\[295\]
rlabel metal1 11316 10506 11316 10506 0 Inst_RAM_IO_ConfigMem.ConfigBits\[296\]
rlabel metal2 12098 10846 12098 10846 0 Inst_RAM_IO_ConfigMem.ConfigBits\[297\]
rlabel metal2 3082 39066 3082 39066 0 Inst_RAM_IO_ConfigMem.ConfigBits\[298\]
rlabel metal2 4830 38726 4830 38726 0 Inst_RAM_IO_ConfigMem.ConfigBits\[299\]
rlabel metal1 8050 38828 8050 38828 0 Inst_RAM_IO_ConfigMem.ConfigBits\[300\]
rlabel metal2 10258 39168 10258 39168 0 Inst_RAM_IO_ConfigMem.ConfigBits\[301\]
rlabel metal1 13616 5882 13616 5882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[302\]
rlabel metal1 13064 6630 13064 6630 0 Inst_RAM_IO_ConfigMem.ConfigBits\[303\]
rlabel metal1 10166 2074 10166 2074 0 Inst_RAM_IO_ConfigMem.ConfigBits\[304\]
rlabel metal2 10258 3230 10258 3230 0 Inst_RAM_IO_ConfigMem.ConfigBits\[305\]
rlabel metal1 5152 31654 5152 31654 0 Inst_RAM_IO_ConfigMem.ConfigBits\[306\]
rlabel viali 5198 30700 5198 30700 0 Inst_RAM_IO_ConfigMem.ConfigBits\[307\]
rlabel metal2 6578 33388 6578 33388 0 Inst_RAM_IO_ConfigMem.ConfigBits\[308\]
rlabel metal1 6854 31994 6854 31994 0 Inst_RAM_IO_ConfigMem.ConfigBits\[309\]
rlabel metal2 10534 22372 10534 22372 0 Inst_RAM_IO_ConfigMem.ConfigBits\[310\]
rlabel metal1 10672 22678 10672 22678 0 Inst_RAM_IO_ConfigMem.ConfigBits\[311\]
rlabel metal1 5658 2822 5658 2822 0 Inst_RAM_IO_ConfigMem.ConfigBits\[312\]
rlabel metal1 5888 2074 5888 2074 0 Inst_RAM_IO_ConfigMem.ConfigBits\[313\]
rlabel metal1 5888 15130 5888 15130 0 Inst_RAM_IO_ConfigMem.ConfigBits\[314\]
rlabel metal1 6256 14586 6256 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[315\]
rlabel metal2 5934 29852 5934 29852 0 Inst_RAM_IO_ConfigMem.ConfigBits\[316\]
rlabel metal1 7176 29614 7176 29614 0 Inst_RAM_IO_ConfigMem.ConfigBits\[317\]
rlabel metal2 12374 4250 12374 4250 0 Inst_RAM_IO_ConfigMem.ConfigBits\[318\]
rlabel metal1 12926 3162 12926 3162 0 Inst_RAM_IO_ConfigMem.ConfigBits\[319\]
rlabel metal1 11776 16762 11776 16762 0 Inst_RAM_IO_ConfigMem.ConfigBits\[320\]
rlabel metal2 11914 17442 11914 17442 0 Inst_RAM_IO_ConfigMem.ConfigBits\[321\]
rlabel metal1 2300 37434 2300 37434 0 Inst_RAM_IO_ConfigMem.ConfigBits\[322\]
rlabel metal2 2622 38828 2622 38828 0 Inst_RAM_IO_ConfigMem.ConfigBits\[323\]
rlabel metal1 10672 40698 10672 40698 0 Inst_RAM_IO_ConfigMem.ConfigBits\[324\]
rlabel metal2 11086 40732 11086 40732 0 Inst_RAM_IO_ConfigMem.ConfigBits\[325\]
rlabel metal2 13662 16218 13662 16218 0 Inst_RAM_IO_ConfigMem.ConfigBits\[326\]
rlabel metal1 14168 16082 14168 16082 0 Inst_RAM_IO_ConfigMem.ConfigBits\[327\]
rlabel metal2 9706 27676 9706 27676 0 Inst_RAM_IO_ConfigMem.ConfigBits\[48\]
rlabel metal1 10028 27098 10028 27098 0 Inst_RAM_IO_ConfigMem.ConfigBits\[49\]
rlabel metal1 2346 34170 2346 34170 0 Inst_RAM_IO_ConfigMem.ConfigBits\[50\]
rlabel metal2 2806 34884 2806 34884 0 Inst_RAM_IO_ConfigMem.ConfigBits\[51\]
rlabel metal1 11638 38794 11638 38794 0 Inst_RAM_IO_ConfigMem.ConfigBits\[52\]
rlabel metal2 12742 39100 12742 39100 0 Inst_RAM_IO_ConfigMem.ConfigBits\[53\]
rlabel metal1 14628 33422 14628 33422 0 Inst_RAM_IO_ConfigMem.ConfigBits\[54\]
rlabel metal2 15134 33932 15134 33932 0 Inst_RAM_IO_ConfigMem.ConfigBits\[55\]
rlabel metal1 8326 25670 8326 25670 0 Inst_RAM_IO_ConfigMem.ConfigBits\[56\]
rlabel metal1 8786 23834 8786 23834 0 Inst_RAM_IO_ConfigMem.ConfigBits\[57\]
rlabel metal1 2254 28186 2254 28186 0 Inst_RAM_IO_ConfigMem.ConfigBits\[58\]
rlabel metal2 2622 29308 2622 29308 0 Inst_RAM_IO_ConfigMem.ConfigBits\[59\]
rlabel metal1 1932 32334 1932 32334 0 Inst_RAM_IO_ConfigMem.ConfigBits\[60\]
rlabel metal1 2530 31994 2530 31994 0 Inst_RAM_IO_ConfigMem.ConfigBits\[61\]
rlabel metal2 3082 30634 3082 30634 0 Inst_RAM_IO_ConfigMem.ConfigBits\[62\]
rlabel metal1 3174 30294 3174 30294 0 Inst_RAM_IO_ConfigMem.ConfigBits\[63\]
rlabel metal2 2438 24412 2438 24412 0 Inst_RAM_IO_ConfigMem.ConfigBits\[64\]
rlabel metal2 2162 23970 2162 23970 0 Inst_RAM_IO_ConfigMem.ConfigBits\[65\]
rlabel metal2 2392 22508 2392 22508 0 Inst_RAM_IO_ConfigMem.ConfigBits\[66\]
rlabel metal1 2208 21998 2208 21998 0 Inst_RAM_IO_ConfigMem.ConfigBits\[67\]
rlabel metal2 2438 27098 2438 27098 0 Inst_RAM_IO_ConfigMem.ConfigBits\[68\]
rlabel metal2 2162 26758 2162 26758 0 Inst_RAM_IO_ConfigMem.ConfigBits\[69\]
rlabel metal1 6854 18836 6854 18836 0 Inst_RAM_IO_ConfigMem.ConfigBits\[70\]
rlabel metal2 7774 19108 7774 19108 0 Inst_RAM_IO_ConfigMem.ConfigBits\[71\]
rlabel metal1 10120 24718 10120 24718 0 Inst_RAM_IO_ConfigMem.ConfigBits\[72\]
rlabel metal2 10902 25500 10902 25500 0 Inst_RAM_IO_ConfigMem.ConfigBits\[73\]
rlabel metal1 11316 28050 11316 28050 0 Inst_RAM_IO_ConfigMem.ConfigBits\[74\]
rlabel metal2 5658 36958 5658 36958 0 Inst_RAM_IO_ConfigMem.ConfigBits\[75\]
rlabel metal2 6210 36652 6210 36652 0 Inst_RAM_IO_ConfigMem.ConfigBits\[76\]
rlabel metal1 7636 37434 7636 37434 0 Inst_RAM_IO_ConfigMem.ConfigBits\[77\]
rlabel metal1 8188 33422 8188 33422 0 Inst_RAM_IO_ConfigMem.ConfigBits\[78\]
rlabel metal2 8786 32946 8786 32946 0 Inst_RAM_IO_ConfigMem.ConfigBits\[79\]
rlabel metal1 9200 33966 9200 33966 0 Inst_RAM_IO_ConfigMem.ConfigBits\[80\]
rlabel metal1 16054 33048 16054 33048 0 Inst_RAM_IO_ConfigMem.ConfigBits\[81\]
rlabel metal2 16882 32402 16882 32402 0 Inst_RAM_IO_ConfigMem.ConfigBits\[82\]
rlabel metal1 17296 34714 17296 34714 0 Inst_RAM_IO_ConfigMem.ConfigBits\[83\]
rlabel metal1 11086 19482 11086 19482 0 Inst_RAM_IO_ConfigMem.ConfigBits\[84\]
rlabel metal1 10120 20502 10120 20502 0 Inst_RAM_IO_ConfigMem.ConfigBits\[85\]
rlabel metal1 5842 34619 5842 34619 0 Inst_RAM_IO_ConfigMem.ConfigBits\[86\]
rlabel metal1 5474 34646 5474 34646 0 Inst_RAM_IO_ConfigMem.ConfigBits\[87\]
rlabel metal2 13110 35428 13110 35428 0 Inst_RAM_IO_ConfigMem.ConfigBits\[88\]
rlabel metal2 12190 35836 12190 35836 0 Inst_RAM_IO_ConfigMem.ConfigBits\[89\]
rlabel metal2 13662 32538 13662 32538 0 Inst_RAM_IO_ConfigMem.ConfigBits\[90\]
rlabel metal2 14490 33966 14490 33966 0 Inst_RAM_IO_ConfigMem.ConfigBits\[91\]
rlabel metal1 11224 19958 11224 19958 0 Inst_RAM_IO_ConfigMem.ConfigBits\[92\]
rlabel metal1 12420 19482 12420 19482 0 Inst_RAM_IO_ConfigMem.ConfigBits\[93\]
rlabel metal1 5842 27574 5842 27574 0 Inst_RAM_IO_ConfigMem.ConfigBits\[94\]
rlabel metal1 6946 27438 6946 27438 0 Inst_RAM_IO_ConfigMem.ConfigBits\[95\]
rlabel metal1 8326 30566 8326 30566 0 Inst_RAM_IO_ConfigMem.ConfigBits\[96\]
rlabel metal1 8464 30294 8464 30294 0 Inst_RAM_IO_ConfigMem.ConfigBits\[97\]
rlabel metal1 13248 31654 13248 31654 0 Inst_RAM_IO_ConfigMem.ConfigBits\[98\]
rlabel metal1 13570 30906 13570 30906 0 Inst_RAM_IO_ConfigMem.ConfigBits\[99\]
rlabel metal2 9706 21257 9706 21257 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG0
rlabel metal1 2438 35122 2438 35122 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG1
rlabel metal2 12512 38930 12512 38930 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG2
rlabel metal1 17722 16014 17722 16014 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG3
rlabel metal2 16606 13396 16606 13396 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG0
rlabel metal1 3289 8398 3289 8398 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG1
rlabel metal1 7130 26010 7130 26010 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG2
rlabel metal1 15801 22066 15801 22066 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG3
rlabel metal1 2162 24038 2162 24038 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG4
rlabel via1 4922 20434 4922 20434 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG5
rlabel metal1 2622 5746 2622 5746 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG6
rlabel metal2 7682 18224 7682 18224 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG7
rlabel metal1 13156 25330 13156 25330 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG0
rlabel metal1 5244 34918 5244 34918 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG1
rlabel metal3 6532 12716 6532 12716 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG10
rlabel metal1 16422 20876 16422 20876 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG11
rlabel via1 15146 24242 15146 24242 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG12
rlabel metal1 4508 38726 4508 38726 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG13
rlabel metal1 8786 19754 8786 19754 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG14
rlabel via1 17446 20910 17446 20910 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG15
rlabel metal1 7820 16082 7820 16082 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG2
rlabel metal1 16100 21318 16100 21318 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG3
rlabel metal1 14352 24242 14352 24242 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG4
rlabel via1 5026 18258 5026 18258 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG5
rlabel metal1 9085 16014 9085 16014 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG6
rlabel metal1 16330 31654 16330 31654 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG7
rlabel metal1 13294 15130 13294 15130 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG8
rlabel via1 4842 16082 4842 16082 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG9
rlabel metal1 12556 27608 12556 27608 0 Inst_RAM_IO_switch_matrix.N1BEG0
rlabel metal1 3588 35258 3588 35258 0 Inst_RAM_IO_switch_matrix.N1BEG1
rlabel metal1 12834 39066 12834 39066 0 Inst_RAM_IO_switch_matrix.N1BEG2
rlabel metal1 15318 33626 15318 33626 0 Inst_RAM_IO_switch_matrix.N1BEG3
rlabel metal3 7291 39916 7291 39916 0 Inst_RAM_IO_switch_matrix.N2BEG0
rlabel metal1 4968 41038 4968 41038 0 Inst_RAM_IO_switch_matrix.N2BEG1
rlabel metal2 3266 33303 3266 33303 0 Inst_RAM_IO_switch_matrix.N2BEG2
rlabel metal2 5014 41106 5014 41106 0 Inst_RAM_IO_switch_matrix.N2BEG3
rlabel metal2 690 35964 690 35964 0 Inst_RAM_IO_switch_matrix.N2BEG4
rlabel metal2 920 26996 920 26996 0 Inst_RAM_IO_switch_matrix.N2BEG5
rlabel metal2 3082 27319 3082 27319 0 Inst_RAM_IO_switch_matrix.N2BEG6
rlabel metal2 17342 37315 17342 37315 0 Inst_RAM_IO_switch_matrix.N2BEG7
rlabel metal1 1886 2958 1886 2958 0 Inst_RAM_IO_switch_matrix.N2BEGb0
rlabel metal1 6624 41038 6624 41038 0 Inst_RAM_IO_switch_matrix.N2BEGb1
rlabel metal1 3542 32742 3542 32742 0 Inst_RAM_IO_switch_matrix.N2BEGb2
rlabel metal1 1012 33490 1012 33490 0 Inst_RAM_IO_switch_matrix.N2BEGb3
rlabel metal4 644 23596 644 23596 0 Inst_RAM_IO_switch_matrix.N2BEGb4
rlabel metal2 1196 18972 1196 18972 0 Inst_RAM_IO_switch_matrix.N2BEGb5
rlabel metal2 4830 30175 4830 30175 0 Inst_RAM_IO_switch_matrix.N2BEGb6
rlabel metal1 1656 43282 1656 43282 0 Inst_RAM_IO_switch_matrix.N2BEGb7
rlabel metal2 11086 34476 11086 34476 0 Inst_RAM_IO_switch_matrix.N4BEG0
rlabel metal1 8188 37162 8188 37162 0 Inst_RAM_IO_switch_matrix.N4BEG1
rlabel metal1 9982 34102 9982 34102 0 Inst_RAM_IO_switch_matrix.N4BEG2
rlabel metal1 16422 34442 16422 34442 0 Inst_RAM_IO_switch_matrix.N4BEG3
rlabel metal3 9729 2516 9729 2516 0 Inst_RAM_IO_switch_matrix.S1BEG0
rlabel metal2 368 15844 368 15844 0 Inst_RAM_IO_switch_matrix.S1BEG1
rlabel metal1 15870 18088 15870 18088 0 Inst_RAM_IO_switch_matrix.S1BEG2
rlabel via3 15525 2652 15525 2652 0 Inst_RAM_IO_switch_matrix.S1BEG3
rlabel metal1 13064 19686 13064 19686 0 Inst_RAM_IO_switch_matrix.S2BEG0
rlabel metal1 506 17102 506 17102 0 Inst_RAM_IO_switch_matrix.S2BEG1
rlabel metal1 13662 1938 13662 1938 0 Inst_RAM_IO_switch_matrix.S2BEG2
rlabel metal1 23506 2040 23506 2040 0 Inst_RAM_IO_switch_matrix.S2BEG3
rlabel metal1 14812 21318 14812 21318 0 Inst_RAM_IO_switch_matrix.S2BEG4
rlabel metal1 276 16082 276 16082 0 Inst_RAM_IO_switch_matrix.S2BEG5
rlabel via3 14835 2652 14835 2652 0 Inst_RAM_IO_switch_matrix.S2BEG6
rlabel via3 16491 1292 16491 1292 0 Inst_RAM_IO_switch_matrix.S2BEG7
rlabel metal1 11730 3026 11730 3026 0 Inst_RAM_IO_switch_matrix.S2BEGb0
rlabel via3 12029 2652 12029 2652 0 Inst_RAM_IO_switch_matrix.S2BEGb1
rlabel metal3 17664 2380 17664 2380 0 Inst_RAM_IO_switch_matrix.S2BEGb2
rlabel via3 11891 22236 11891 22236 0 Inst_RAM_IO_switch_matrix.S2BEGb3
rlabel metal1 12282 2346 12282 2346 0 Inst_RAM_IO_switch_matrix.S2BEGb4
rlabel metal2 13432 15334 13432 15334 0 Inst_RAM_IO_switch_matrix.S2BEGb5
rlabel metal1 13340 3026 13340 3026 0 Inst_RAM_IO_switch_matrix.S2BEGb6
rlabel metal1 13754 3366 13754 3366 0 Inst_RAM_IO_switch_matrix.S2BEGb7
rlabel metal3 20493 1292 20493 1292 0 Inst_RAM_IO_switch_matrix.S4BEG0
rlabel via2 18538 1309 18538 1309 0 Inst_RAM_IO_switch_matrix.S4BEG1
rlabel metal2 18492 17238 18492 17238 0 Inst_RAM_IO_switch_matrix.S4BEG2
rlabel metal2 20332 16388 20332 16388 0 Inst_RAM_IO_switch_matrix.S4BEG3
rlabel metal1 3542 4624 3542 4624 0 Inst_RAM_IO_switch_matrix.W1BEG0
rlabel metal2 920 17204 920 17204 0 Inst_RAM_IO_switch_matrix.W1BEG1
rlabel metal2 2898 4845 2898 4845 0 Inst_RAM_IO_switch_matrix.W1BEG2
rlabel metal1 11454 5168 11454 5168 0 Inst_RAM_IO_switch_matrix.W1BEG3
rlabel via2 1702 5661 1702 5661 0 Inst_RAM_IO_switch_matrix.W2BEG0
rlabel metal2 7406 6256 7406 6256 0 Inst_RAM_IO_switch_matrix.W2BEG1
rlabel metal1 4278 7446 4278 7446 0 Inst_RAM_IO_switch_matrix.W2BEG2
rlabel metal1 5704 6290 5704 6290 0 Inst_RAM_IO_switch_matrix.W2BEG3
rlabel metal1 15916 5542 15916 5542 0 Inst_RAM_IO_switch_matrix.W2BEG4
rlabel metal1 3864 7378 3864 7378 0 Inst_RAM_IO_switch_matrix.W2BEG5
rlabel metal2 3634 6086 3634 6086 0 Inst_RAM_IO_switch_matrix.W2BEG6
rlabel metal2 9430 4403 9430 4403 0 Inst_RAM_IO_switch_matrix.W2BEG7
rlabel metal2 6670 6426 6670 6426 0 Inst_RAM_IO_switch_matrix.W2BEGb0
rlabel metal1 4554 7412 4554 7412 0 Inst_RAM_IO_switch_matrix.W2BEGb1
rlabel metal1 4508 12342 4508 12342 0 Inst_RAM_IO_switch_matrix.W2BEGb2
rlabel metal2 5198 4420 5198 4420 0 Inst_RAM_IO_switch_matrix.W2BEGb3
rlabel metal2 14490 3808 14490 3808 0 Inst_RAM_IO_switch_matrix.W2BEGb4
rlabel metal2 5612 15164 5612 15164 0 Inst_RAM_IO_switch_matrix.W2BEGb5
rlabel metal2 1702 8772 1702 8772 0 Inst_RAM_IO_switch_matrix.W2BEGb6
rlabel metal2 1610 3332 1610 3332 0 Inst_RAM_IO_switch_matrix.W2BEGb7
rlabel metal2 2254 14433 2254 14433 0 Inst_RAM_IO_switch_matrix.W6BEG0
rlabel metal1 1426 40630 1426 40630 0 Inst_RAM_IO_switch_matrix.W6BEG1
rlabel metal2 1978 18207 1978 18207 0 Inst_RAM_IO_switch_matrix.W6BEG10
rlabel metal1 10810 17850 10810 17850 0 Inst_RAM_IO_switch_matrix.W6BEG11
rlabel metal1 1518 41072 1518 41072 0 Inst_RAM_IO_switch_matrix.W6BEG2
rlabel metal2 14490 14178 14490 14178 0 Inst_RAM_IO_switch_matrix.W6BEG3
rlabel metal2 17526 14586 17526 14586 0 Inst_RAM_IO_switch_matrix.W6BEG4
rlabel metal2 2346 15011 2346 15011 0 Inst_RAM_IO_switch_matrix.W6BEG5
rlabel metal2 1610 16388 1610 16388 0 Inst_RAM_IO_switch_matrix.W6BEG6
rlabel metal1 11224 15674 11224 15674 0 Inst_RAM_IO_switch_matrix.W6BEG7
rlabel metal2 17342 17204 17342 17204 0 Inst_RAM_IO_switch_matrix.W6BEG8
rlabel metal1 8142 16218 8142 16218 0 Inst_RAM_IO_switch_matrix.W6BEG9
rlabel metal2 7222 9316 7222 9316 0 Inst_RAM_IO_switch_matrix.WW4BEG0
rlabel metal2 3450 10030 3450 10030 0 Inst_RAM_IO_switch_matrix.WW4BEG1
rlabel metal1 1610 17748 1610 17748 0 Inst_RAM_IO_switch_matrix.WW4BEG10
rlabel metal2 10810 13702 10810 13702 0 Inst_RAM_IO_switch_matrix.WW4BEG11
rlabel metal1 14835 7718 14835 7718 0 Inst_RAM_IO_switch_matrix.WW4BEG12
rlabel metal1 3634 14484 3634 14484 0 Inst_RAM_IO_switch_matrix.WW4BEG13
rlabel metal1 1610 12172 1610 12172 0 Inst_RAM_IO_switch_matrix.WW4BEG14
rlabel metal2 9706 6902 9706 6902 0 Inst_RAM_IO_switch_matrix.WW4BEG15
rlabel metal1 5704 11050 5704 11050 0 Inst_RAM_IO_switch_matrix.WW4BEG2
rlabel metal1 7038 10200 7038 10200 0 Inst_RAM_IO_switch_matrix.WW4BEG3
rlabel metal1 10350 11288 10350 11288 0 Inst_RAM_IO_switch_matrix.WW4BEG4
rlabel metal1 3634 11764 3634 11764 0 Inst_RAM_IO_switch_matrix.WW4BEG5
rlabel metal1 1610 11152 1610 11152 0 Inst_RAM_IO_switch_matrix.WW4BEG6
rlabel metal1 11408 12818 11408 12818 0 Inst_RAM_IO_switch_matrix.WW4BEG7
rlabel metal1 2162 10676 2162 10676 0 Inst_RAM_IO_switch_matrix.WW4BEG8
rlabel via2 2162 7837 2162 7837 0 Inst_RAM_IO_switch_matrix.WW4BEG9
rlabel metal1 11822 25466 11822 25466 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A0
rlabel metal1 11454 24786 11454 24786 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A1
rlabel metal1 11914 27064 11914 27064 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[0\]
rlabel metal2 11638 27268 11638 27268 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[1\]
rlabel metal2 11270 27744 11270 27744 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._0_
rlabel metal1 11684 27642 11684 27642 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._1_
rlabel metal1 6762 35802 6762 35802 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A0
rlabel metal1 7268 36278 7268 36278 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A1
rlabel metal1 7084 36346 7084 36346 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[0\]
rlabel metal1 7544 36890 7544 36890 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[1\]
rlabel metal1 7682 36822 7682 36822 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._0_
rlabel metal2 8234 37468 8234 37468 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._1_
rlabel metal1 9522 33626 9522 33626 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A0
rlabel metal1 9476 32538 9476 32538 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A1
rlabel metal1 10258 33932 10258 33932 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[0\]
rlabel metal1 9384 33082 9384 33082 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[1\]
rlabel metal1 9246 34034 9246 34034 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._0_
rlabel metal1 9798 34034 9798 34034 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._1_
rlabel metal1 17388 32878 17388 32878 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A0
rlabel metal1 17434 31994 17434 31994 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A1
rlabel metal1 17250 33082 17250 33082 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[0\]
rlabel metal1 17388 33626 17388 33626 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[1\]
rlabel metal1 16790 34170 16790 34170 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._0_
rlabel metal1 16560 34510 16560 34510 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._1_
rlabel metal1 16192 24786 16192 24786 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A0
rlabel metal1 16054 24378 16054 24378 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A1
rlabel metal1 16790 24208 16790 24208 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[0\]
rlabel metal1 17848 23086 17848 23086 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[1\]
rlabel metal1 18216 23698 18216 23698 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._0_
rlabel metal1 18216 23290 18216 23290 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._1_
rlabel metal1 6440 23086 6440 23086 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A0
rlabel metal1 6992 21930 6992 21930 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A1
rlabel metal1 6854 23052 6854 23052 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[0\]
rlabel metal2 7590 22576 7590 22576 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[1\]
rlabel metal1 7222 21998 7222 21998 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._0_
rlabel metal1 7406 22950 7406 22950 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._1_
rlabel metal1 11868 29818 11868 29818 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A0
rlabel metal1 11776 29138 11776 29138 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A1
rlabel metal1 12282 30192 12282 30192 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[0\]
rlabel viali 12650 29140 12650 29140 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[1\]
rlabel metal2 12742 29818 12742 29818 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._0_
rlabel metal1 13156 29274 13156 29274 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._1_
rlabel via1 18542 20906 18542 20906 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A0
rlabel metal1 18814 20944 18814 20944 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A1
rlabel metal1 18906 20978 18906 20978 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[0\]
rlabel metal2 19458 20298 19458 20298 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[1\]
rlabel metal2 18630 20774 18630 20774 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._0_
rlabel metal1 18814 20332 18814 20332 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._1_
rlabel metal2 230 43088 230 43088 0 N1BEG[0]
rlabel metal2 506 43496 506 43496 0 N1BEG[1]
rlabel metal2 782 43258 782 43258 0 N1BEG[2]
rlabel metal2 1058 43632 1058 43632 0 N1BEG[3]
rlabel metal2 230 1010 230 1010 0 N1END[0]
rlabel metal2 605 68 605 68 0 N1END[1]
rlabel metal2 881 68 881 68 0 N1END[2]
rlabel metal2 1058 942 1058 942 0 N1END[3]
rlabel metal2 1334 43462 1334 43462 0 N2BEG[0]
rlabel metal2 1610 43598 1610 43598 0 N2BEG[1]
rlabel metal2 1985 44948 1985 44948 0 N2BEG[2]
rlabel metal1 2116 43418 2116 43418 0 N2BEG[3]
rlabel metal2 2438 44176 2438 44176 0 N2BEG[4]
rlabel metal2 2714 43836 2714 43836 0 N2BEG[5]
rlabel metal2 2990 44176 2990 44176 0 N2BEG[6]
rlabel metal2 3319 44948 3319 44948 0 N2BEG[7]
rlabel metal1 4232 41786 4232 41786 0 N2BEGb[0]
rlabel metal1 3910 42534 3910 42534 0 N2BEGb[1]
rlabel metal2 4094 44057 4094 44057 0 N2BEGb[2]
rlabel metal2 4370 44465 4370 44465 0 N2BEGb[3]
rlabel metal2 3542 43724 3542 43724 0 N2BEGb[4]
rlabel metal2 4922 43836 4922 43836 0 N2BEGb[5]
rlabel metal1 5014 43418 5014 43418 0 N2BEGb[6]
rlabel metal1 5428 43418 5428 43418 0 N2BEGb[7]
rlabel metal2 3542 1010 3542 1010 0 N2END[0]
rlabel metal2 3765 68 3765 68 0 N2END[1]
rlabel metal2 4094 636 4094 636 0 N2END[2]
rlabel metal2 4317 68 4317 68 0 N2END[3]
rlabel metal2 4646 1248 4646 1248 0 N2END[4]
rlabel metal2 4922 1248 4922 1248 0 N2END[5]
rlabel metal2 5251 68 5251 68 0 N2END[6]
rlabel metal2 5474 908 5474 908 0 N2END[7]
rlabel metal2 1334 755 1334 755 0 N2MID[0]
rlabel metal2 1610 670 1610 670 0 N2MID[1]
rlabel metal2 1939 68 1939 68 0 N2MID[2]
rlabel metal2 2215 68 2215 68 0 N2MID[3]
rlabel metal2 2438 687 2438 687 0 N2MID[4]
rlabel metal2 2714 1010 2714 1010 0 N2MID[5]
rlabel metal2 2990 670 2990 670 0 N2MID[6]
rlabel metal2 3266 1010 3266 1010 0 N2MID[7]
rlabel metal2 5750 44176 5750 44176 0 N4BEG[0]
rlabel metal1 8188 43418 8188 43418 0 N4BEG[10]
rlabel metal1 8740 42738 8740 42738 0 N4BEG[11]
rlabel metal1 9108 43418 9108 43418 0 N4BEG[12]
rlabel metal2 9437 44948 9437 44948 0 N4BEG[13]
rlabel metal1 8832 43418 8832 43418 0 N4BEG[14]
rlabel metal1 9844 43418 9844 43418 0 N4BEG[15]
rlabel metal2 6026 44329 6026 44329 0 N4BEG[1]
rlabel metal1 6026 42534 6026 42534 0 N4BEG[2]
rlabel metal2 6578 44329 6578 44329 0 N4BEG[3]
rlabel metal2 6801 44948 6801 44948 0 N4BEG[4]
rlabel metal2 7229 44948 7229 44948 0 N4BEG[5]
rlabel metal1 7498 42330 7498 42330 0 N4BEG[6]
rlabel metal1 7728 42534 7728 42534 0 N4BEG[7]
rlabel metal1 7774 43418 7774 43418 0 N4BEG[8]
rlabel metal2 8234 44261 8234 44261 0 N4BEG[9]
rlabel metal4 1012 19584 1012 19584 0 N4BEG_outbuf_0.A
rlabel metal1 5658 41650 5658 41650 0 N4BEG_outbuf_0.X
rlabel metal2 16652 22916 16652 22916 0 N4BEG_outbuf_1.A
rlabel metal1 6394 41616 6394 41616 0 N4BEG_outbuf_1.X
rlabel via2 9430 2635 9430 2635 0 N4BEG_outbuf_10.A
rlabel metal1 9062 41786 9062 41786 0 N4BEG_outbuf_10.X
rlabel via3 10741 16524 10741 16524 0 N4BEG_outbuf_11.A
rlabel metal1 10258 42704 10258 42704 0 N4BEG_outbuf_11.X
rlabel metal4 1196 21760 1196 21760 0 N4BEG_outbuf_2.A
rlabel metal1 6486 41786 6486 41786 0 N4BEG_outbuf_2.X
rlabel metal3 6693 1972 6693 1972 0 N4BEG_outbuf_3.A
rlabel metal1 7038 41548 7038 41548 0 N4BEG_outbuf_3.X
rlabel metal1 7728 1802 7728 1802 0 N4BEG_outbuf_4.A
rlabel metal1 6532 42330 6532 42330 0 N4BEG_outbuf_4.X
rlabel metal3 18699 14892 18699 14892 0 N4BEG_outbuf_5.A
rlabel metal1 7498 41616 7498 41616 0 N4BEG_outbuf_5.X
rlabel metal2 7774 2159 7774 2159 0 N4BEG_outbuf_6.A
rlabel metal1 7038 40902 7038 40902 0 N4BEG_outbuf_6.X
rlabel metal2 8142 2159 8142 2159 0 N4BEG_outbuf_7.A
rlabel metal1 7958 41684 7958 41684 0 N4BEG_outbuf_7.X
rlabel metal2 8510 2159 8510 2159 0 N4BEG_outbuf_8.A
rlabel metal1 8280 41582 8280 41582 0 N4BEG_outbuf_8.X
rlabel metal2 8878 2159 8878 2159 0 N4BEG_outbuf_9.A
rlabel metal1 8552 41582 8552 41582 0 N4BEG_outbuf_9.X
rlabel metal2 5750 551 5750 551 0 N4END[0]
rlabel metal2 8510 687 8510 687 0 N4END[10]
rlabel metal2 8786 1248 8786 1248 0 N4END[11]
rlabel metal2 9062 296 9062 296 0 N4END[12]
rlabel metal2 9338 1421 9338 1421 0 N4END[13]
rlabel metal2 9614 330 9614 330 0 N4END[14]
rlabel metal2 9890 211 9890 211 0 N4END[15]
rlabel metal2 6026 670 6026 670 0 N4END[1]
rlabel metal2 6302 704 6302 704 0 N4END[2]
rlabel metal2 6578 636 6578 636 0 N4END[3]
rlabel metal2 6755 68 6755 68 0 N4END[4]
rlabel metal2 7130 398 7130 398 0 N4END[5]
rlabel metal2 7314 3026 7314 3026 0 N4END[6]
rlabel metal1 7590 2958 7590 2958 0 N4END[7]
rlabel metal2 7859 68 7859 68 0 N4END[8]
rlabel metal2 8234 704 8234 704 0 N4END[9]
rlabel metal3 25066 7412 25066 7412 0 RAM2FAB_D0_I0
rlabel metal3 25618 7956 25618 7956 0 RAM2FAB_D0_I1
rlabel metal3 24928 8500 24928 8500 0 RAM2FAB_D0_I2
rlabel metal3 24882 9044 24882 9044 0 RAM2FAB_D0_I3
rlabel metal3 24008 5236 24008 5236 0 RAM2FAB_D1_I0
rlabel metal3 24744 5780 24744 5780 0 RAM2FAB_D1_I1
rlabel metal3 24560 6324 24560 6324 0 RAM2FAB_D1_I2
rlabel metal3 24698 6868 24698 6868 0 RAM2FAB_D1_I3
rlabel metal3 24146 3060 24146 3060 0 RAM2FAB_D2_I0
rlabel metal3 24514 3604 24514 3604 0 RAM2FAB_D2_I1
rlabel metal2 21390 5355 21390 5355 0 RAM2FAB_D2_I2
rlabel metal3 25411 4692 25411 4692 0 RAM2FAB_D2_I3
rlabel metal3 23502 884 23502 884 0 RAM2FAB_D3_I0
rlabel metal3 24238 1428 24238 1428 0 RAM2FAB_D3_I1
rlabel metal2 19274 3621 19274 3621 0 RAM2FAB_D3_I2
rlabel metal3 24974 2516 24974 2516 0 RAM2FAB_D3_I3
rlabel metal2 10067 68 10067 68 0 S1BEG[0]
rlabel metal2 10442 806 10442 806 0 S1BEG[1]
rlabel metal2 10718 1095 10718 1095 0 S1BEG[2]
rlabel metal2 10994 755 10994 755 0 S1BEG[3]
rlabel metal2 10067 44948 10067 44948 0 S1END[0]
rlabel metal2 10389 44948 10389 44948 0 S1END[1]
rlabel metal2 10718 44108 10718 44108 0 S1END[2]
rlabel metal2 10994 44533 10994 44533 0 S1END[3]
rlabel metal2 13478 636 13478 636 0 S2BEG[0]
rlabel metal2 13754 806 13754 806 0 S2BEG[1]
rlabel metal2 14030 636 14030 636 0 S2BEG[2]
rlabel metal2 14306 908 14306 908 0 S2BEG[3]
rlabel metal2 14681 68 14681 68 0 S2BEG[4]
rlabel metal2 14858 347 14858 347 0 S2BEG[5]
rlabel metal2 15134 755 15134 755 0 S2BEG[6]
rlabel metal2 15410 942 15410 942 0 S2BEG[7]
rlabel metal2 11217 68 11217 68 0 S2BEGb[0]
rlabel metal2 11546 347 11546 347 0 S2BEGb[1]
rlabel metal2 11875 68 11875 68 0 S2BEGb[2]
rlabel metal2 12098 483 12098 483 0 S2BEGb[3]
rlabel metal2 12558 1479 12558 1479 0 S2BEGb[4]
rlabel metal2 12650 908 12650 908 0 S2BEGb[5]
rlabel metal2 12926 534 12926 534 0 S2BEGb[6]
rlabel metal2 13301 68 13301 68 0 S2BEGb[7]
rlabel metal2 11270 44142 11270 44142 0 S2END[0]
rlabel metal2 11599 44948 11599 44948 0 S2END[1]
rlabel metal2 11875 44948 11875 44948 0 S2END[2]
rlabel metal2 12098 44108 12098 44108 0 S2END[3]
rlabel metal2 12466 43741 12466 43741 0 S2END[4]
rlabel metal2 12650 44142 12650 44142 0 S2END[5]
rlabel metal2 12827 44948 12827 44948 0 S2END[6]
rlabel metal2 13202 44176 13202 44176 0 S2END[7]
rlabel metal2 13478 44142 13478 44142 0 S2MID[0]
rlabel metal2 13754 43836 13754 43836 0 S2MID[1]
rlabel metal2 14083 44948 14083 44948 0 S2MID[2]
rlabel metal2 14359 44948 14359 44948 0 S2MID[3]
rlabel metal2 14681 44948 14681 44948 0 S2MID[4]
rlabel metal2 14858 44142 14858 44142 0 S2MID[5]
rlabel metal2 15134 43853 15134 43853 0 S2MID[6]
rlabel metal2 15410 44533 15410 44533 0 S2MID[7]
rlabel metal2 15686 908 15686 908 0 S4BEG[0]
rlabel metal2 18446 1452 18446 1452 0 S4BEG[10]
rlabel metal2 18669 68 18669 68 0 S4BEG[11]
rlabel metal2 19097 68 19097 68 0 S4BEG[12]
rlabel metal2 19274 1299 19274 1299 0 S4BEG[13]
rlabel metal2 19550 908 19550 908 0 S4BEG[14]
rlabel metal2 19879 68 19879 68 0 S4BEG[15]
rlabel metal2 16015 68 16015 68 0 S4BEG[1]
rlabel metal2 16238 738 16238 738 0 S4BEG[2]
rlabel metal2 16514 636 16514 636 0 S4BEG[3]
rlabel metal2 16843 68 16843 68 0 S4BEG[4]
rlabel metal2 17066 942 17066 942 0 S4BEG[5]
rlabel metal2 17395 68 17395 68 0 S4BEG[6]
rlabel metal2 17717 68 17717 68 0 S4BEG[7]
rlabel metal2 17894 908 17894 908 0 S4BEG[8]
rlabel metal2 18170 908 18170 908 0 S4BEG[9]
rlabel metal1 16238 41582 16238 41582 0 S4BEG_outbuf_0.A
rlabel metal3 16169 2516 16169 2516 0 S4BEG_outbuf_0.X
rlabel metal1 16468 41582 16468 41582 0 S4BEG_outbuf_1.A
rlabel metal1 16928 2414 16928 2414 0 S4BEG_outbuf_1.X
rlabel metal1 19090 41174 19090 41174 0 S4BEG_outbuf_10.A
rlabel metal2 19182 39168 19182 39168 0 S4BEG_outbuf_10.X
rlabel metal1 19412 40494 19412 40494 0 S4BEG_outbuf_11.A
rlabel metal3 19527 40052 19527 40052 0 S4BEG_outbuf_11.X
rlabel metal1 16790 42296 16790 42296 0 S4BEG_outbuf_2.A
rlabel metal1 16928 17510 16928 17510 0 S4BEG_outbuf_2.X
rlabel metal1 17250 42262 17250 42262 0 S4BEG_outbuf_3.A
rlabel via3 17733 4012 17733 4012 0 S4BEG_outbuf_3.X
rlabel metal1 17664 42262 17664 42262 0 S4BEG_outbuf_4.A
rlabel via3 17549 2652 17549 2652 0 S4BEG_outbuf_4.X
rlabel metal1 17986 42262 17986 42262 0 S4BEG_outbuf_5.A
rlabel metal3 18699 2652 18699 2652 0 S4BEG_outbuf_5.X
rlabel metal1 18262 42296 18262 42296 0 S4BEG_outbuf_6.A
rlabel metal2 19228 14348 19228 14348 0 S4BEG_outbuf_6.X
rlabel metal2 18630 42500 18630 42500 0 S4BEG_outbuf_7.A
rlabel metal2 18124 18700 18124 18700 0 S4BEG_outbuf_7.X
rlabel metal1 18722 42262 18722 42262 0 S4BEG_outbuf_8.A
rlabel metal2 17986 12614 17986 12614 0 S4BEG_outbuf_8.X
rlabel metal2 19366 42670 19366 42670 0 S4BEG_outbuf_9.A
rlabel metal3 15640 41684 15640 41684 0 S4BEG_outbuf_9.X
rlabel metal2 15686 44142 15686 44142 0 S4END[0]
rlabel metal2 18393 44948 18393 44948 0 S4END[10]
rlabel metal2 18623 44948 18623 44948 0 S4END[11]
rlabel metal2 18998 44329 18998 44329 0 S4END[12]
rlabel metal1 18676 41106 18676 41106 0 S4END[13]
rlabel metal2 19550 43258 19550 43258 0 S4END[14]
rlabel metal2 19826 43292 19826 43292 0 S4END[15]
rlabel metal2 15962 44125 15962 44125 0 S4END[1]
rlabel metal2 16238 44533 16238 44533 0 S4END[2]
rlabel metal2 16514 43802 16514 43802 0 S4END[3]
rlabel metal2 16790 44074 16790 44074 0 S4END[4]
rlabel metal2 17066 44346 17066 44346 0 S4END[5]
rlabel metal2 17342 44278 17342 44278 0 S4END[6]
rlabel metal2 17618 44312 17618 44312 0 S4END[7]
rlabel metal2 17894 44856 17894 44856 0 S4END[8]
rlabel metal2 23138 42993 23138 42993 0 S4END[9]
rlabel metal1 20240 22066 20240 22066 0 UserCLK
rlabel metal2 21712 41786 21712 41786 0 UserCLKo
rlabel metal3 199 5236 199 5236 0 W1BEG[0]
rlabel metal3 636 5508 636 5508 0 W1BEG[1]
rlabel metal1 2852 5338 2852 5338 0 W1BEG[2]
rlabel metal3 866 6052 866 6052 0 W1BEG[3]
rlabel metal3 682 6324 682 6324 0 W2BEG[0]
rlabel metal3 1142 6596 1142 6596 0 W2BEG[1]
rlabel via2 3358 6851 3358 6851 0 W2BEG[2]
rlabel metal3 728 7140 728 7140 0 W2BEG[3]
rlabel metal3 475 7412 475 7412 0 W2BEG[4]
rlabel metal3 728 7684 728 7684 0 W2BEG[5]
rlabel metal2 3082 7395 3082 7395 0 W2BEG[6]
rlabel metal3 567 8228 567 8228 0 W2BEG[7]
rlabel metal3 866 8500 866 8500 0 W2BEGb[0]
rlabel metal2 2898 8109 2898 8109 0 W2BEGb[1]
rlabel metal3 728 9044 728 9044 0 W2BEGb[2]
rlabel metal3 843 9316 843 9316 0 W2BEGb[3]
rlabel metal2 2898 9741 2898 9741 0 W2BEGb[4]
rlabel metal3 774 9860 774 9860 0 W2BEGb[5]
rlabel metal3 1234 10132 1234 10132 0 W2BEGb[6]
rlabel metal3 820 10404 820 10404 0 W2BEGb[7]
rlabel metal3 958 15028 958 15028 0 W6BEG[0]
rlabel metal3 728 17748 728 17748 0 W6BEG[10]
rlabel metal3 774 18020 774 18020 0 W6BEG[11]
rlabel metal2 4186 15300 4186 15300 0 W6BEG[1]
rlabel metal3 567 15572 567 15572 0 W6BEG[2]
rlabel metal2 3726 15487 3726 15487 0 W6BEG[3]
rlabel metal3 866 16116 866 16116 0 W6BEG[4]
rlabel metal3 958 16388 958 16388 0 W6BEG[5]
rlabel metal3 728 16660 728 16660 0 W6BEG[6]
rlabel metal3 728 16932 728 16932 0 W6BEG[7]
rlabel metal3 1004 17204 1004 17204 0 W6BEG[8]
rlabel metal3 544 17476 544 17476 0 W6BEG[9]
rlabel metal2 3174 10149 3174 10149 0 WW4BEG[0]
rlabel metal3 659 13396 659 13396 0 WW4BEG[10]
rlabel metal2 3542 13583 3542 13583 0 WW4BEG[11]
rlabel metal3 728 13940 728 13940 0 WW4BEG[12]
rlabel metal3 912 14212 912 14212 0 WW4BEG[13]
rlabel metal3 728 14484 728 14484 0 WW4BEG[14]
rlabel metal3 820 14756 820 14756 0 WW4BEG[15]
rlabel metal2 3358 10421 3358 10421 0 WW4BEG[1]
rlabel metal3 958 11220 958 11220 0 WW4BEG[2]
rlabel metal2 3266 10863 3266 10863 0 WW4BEG[3]
rlabel metal2 4002 11917 4002 11917 0 WW4BEG[4]
rlabel metal3 728 12036 728 12036 0 WW4BEG[5]
rlabel metal3 751 12308 751 12308 0 WW4BEG[6]
rlabel metal3 912 12580 912 12580 0 WW4BEG[7]
rlabel metal3 866 12852 866 12852 0 WW4BEG[8]
rlabel metal2 3542 13039 3542 13039 0 WW4BEG[9]
rlabel metal1 23322 27404 23322 27404 0 data_inbuf_0.X
rlabel metal1 23414 28016 23414 28016 0 data_inbuf_1.X
rlabel metal1 23230 32912 23230 32912 0 data_inbuf_10.X
rlabel metal1 23230 33524 23230 33524 0 data_inbuf_11.X
rlabel metal1 21482 34068 21482 34068 0 data_inbuf_12.X
rlabel metal1 23000 34578 23000 34578 0 data_inbuf_13.X
rlabel metal1 22678 34646 22678 34646 0 data_inbuf_14.X
rlabel metal1 21666 34612 21666 34612 0 data_inbuf_15.X
rlabel metal1 23138 35632 23138 35632 0 data_inbuf_16.X
rlabel metal1 23736 35802 23736 35802 0 data_inbuf_17.X
rlabel metal2 22310 36550 22310 36550 0 data_inbuf_18.X
rlabel metal1 19044 36890 19044 36890 0 data_inbuf_19.X
rlabel metal1 23598 28492 23598 28492 0 data_inbuf_2.X
rlabel metal1 19964 36890 19964 36890 0 data_inbuf_20.X
rlabel metal1 21919 37094 21919 37094 0 data_inbuf_21.X
rlabel metal1 23092 37842 23092 37842 0 data_inbuf_22.X
rlabel metal2 18170 38148 18170 38148 0 data_inbuf_23.X
rlabel metal1 19918 38182 19918 38182 0 data_inbuf_24.X
rlabel metal1 21390 39508 21390 39508 0 data_inbuf_25.X
rlabel metal1 21942 39406 21942 39406 0 data_inbuf_26.X
rlabel metal1 20286 40630 20286 40630 0 data_inbuf_27.X
rlabel metal3 19044 41616 19044 41616 0 data_inbuf_28.X
rlabel metal1 22034 40052 22034 40052 0 data_inbuf_29.X
rlabel metal1 20884 28730 20884 28730 0 data_inbuf_3.X
rlabel metal1 23092 38930 23092 38930 0 data_inbuf_30.X
rlabel metal1 20194 41106 20194 41106 0 data_inbuf_31.X
rlabel metal1 23184 29138 23184 29138 0 data_inbuf_4.X
rlabel metal1 23368 29818 23368 29818 0 data_inbuf_5.X
rlabel viali 22958 30226 22958 30226 0 data_inbuf_6.X
rlabel metal1 23552 31790 23552 31790 0 data_inbuf_7.X
rlabel metal1 23506 30736 23506 30736 0 data_inbuf_8.X
rlabel metal1 21965 32742 21965 32742 0 data_inbuf_9.X
rlabel metal1 23506 27574 23506 27574 0 data_outbuf_0.X
rlabel metal1 23414 28186 23414 28186 0 data_outbuf_1.X
rlabel metal1 23184 33082 23184 33082 0 data_outbuf_10.X
rlabel metal1 23184 33626 23184 33626 0 data_outbuf_11.X
rlabel metal1 23230 34034 23230 34034 0 data_outbuf_12.X
rlabel metal1 23736 34578 23736 34578 0 data_outbuf_13.X
rlabel metal1 23506 34544 23506 34544 0 data_outbuf_14.X
rlabel metal2 21482 34884 21482 34884 0 data_outbuf_15.X
rlabel metal1 23506 35700 23506 35700 0 data_outbuf_16.X
rlabel metal1 23782 37434 23782 37434 0 data_outbuf_17.X
rlabel metal1 23874 36788 23874 36788 0 data_outbuf_18.X
rlabel metal1 20010 37196 20010 37196 0 data_outbuf_19.X
rlabel metal2 23414 28866 23414 28866 0 data_outbuf_2.X
rlabel metal1 20654 37094 20654 37094 0 data_outbuf_20.X
rlabel metal2 22494 37876 22494 37876 0 data_outbuf_21.X
rlabel metal1 22770 37706 22770 37706 0 data_outbuf_22.X
rlabel metal1 19090 38522 19090 38522 0 data_outbuf_23.X
rlabel metal2 20194 39236 20194 39236 0 data_outbuf_24.X
rlabel metal1 23046 40052 23046 40052 0 data_outbuf_25.X
rlabel metal2 21666 40052 21666 40052 0 data_outbuf_26.X
rlabel metal1 21114 41480 21114 41480 0 data_outbuf_27.X
rlabel metal2 18354 40222 18354 40222 0 data_outbuf_28.X
rlabel metal1 21758 39814 21758 39814 0 data_outbuf_29.X
rlabel metal2 22126 28526 22126 28526 0 data_outbuf_3.X
rlabel metal2 22954 39780 22954 39780 0 data_outbuf_30.X
rlabel metal1 21298 40494 21298 40494 0 data_outbuf_31.X
rlabel metal2 22954 29274 22954 29274 0 data_outbuf_4.X
rlabel metal1 22770 30226 22770 30226 0 data_outbuf_5.X
rlabel metal1 23506 30192 23506 30192 0 data_outbuf_6.X
rlabel metal1 23460 32266 23460 32266 0 data_outbuf_7.X
rlabel metal1 23552 32402 23552 32402 0 data_outbuf_8.X
rlabel metal1 23690 32878 23690 32878 0 data_outbuf_9.X
rlabel metal1 3174 19346 3174 19346 0 net1
rlabel metal1 1656 32266 1656 32266 0 net10
rlabel metal2 20424 1972 20424 1972 0 net100
rlabel metal1 2300 2006 2300 2006 0 net101
rlabel metal1 2070 37400 2070 37400 0 net102
rlabel metal1 4554 2448 4554 2448 0 net103
rlabel metal1 2691 1802 2691 1802 0 net104
rlabel metal2 3358 1632 3358 1632 0 net105
rlabel metal2 736 17204 736 17204 0 net106
rlabel via3 4485 1292 4485 1292 0 net107
rlabel metal1 3910 2074 3910 2074 0 net108
rlabel metal1 6210 2312 6210 2312 0 net109
rlabel metal2 6946 27727 6946 27727 0 net11
rlabel metal1 4968 2618 4968 2618 0 net110
rlabel metal2 5198 3162 5198 3162 0 net111
rlabel metal2 4462 2227 4462 2227 0 net112
rlabel metal1 10994 3060 10994 3060 0 net113
rlabel metal1 1748 1326 1748 1326 0 net114
rlabel metal1 2116 1326 2116 1326 0 net115
rlabel metal1 2576 1326 2576 1326 0 net116
rlabel metal1 6256 2414 6256 2414 0 net117
rlabel metal1 2990 1904 2990 1904 0 net118
rlabel metal1 3634 1326 3634 1326 0 net119
rlabel metal1 11362 20978 11362 20978 0 net12
rlabel metal1 3450 2074 3450 2074 0 net120
rlabel metal1 12512 9554 12512 9554 0 net121
rlabel metal1 7820 2006 7820 2006 0 net122
rlabel metal1 8326 2006 8326 2006 0 net123
rlabel metal2 5106 1088 5106 1088 0 net124
rlabel metal1 8878 2006 8878 2006 0 net125
rlabel metal1 6440 1190 6440 1190 0 net126
rlabel metal1 8970 1258 8970 1258 0 net127
rlabel via3 5589 1972 5589 1972 0 net128
rlabel metal2 6118 969 6118 969 0 net129
rlabel metal1 14352 19346 14352 19346 0 net13
rlabel metal2 12742 1462 12742 1462 0 net130
rlabel metal1 6670 1394 6670 1394 0 net131
rlabel metal2 6762 2074 6762 2074 0 net132
rlabel metal1 6808 2890 6808 2890 0 net133
rlabel metal1 7130 2006 7130 2006 0 net134
rlabel metal2 3910 1054 3910 1054 0 net135
rlabel metal1 8096 1258 8096 1258 0 net136
rlabel metal1 20051 7446 20051 7446 0 net137
rlabel metal1 21022 7378 21022 7378 0 net138
rlabel metal1 23312 8466 23312 8466 0 net139
rlabel metal1 7774 20774 7774 20774 0 net14
rlabel metal1 22862 9520 22862 9520 0 net140
rlabel metal1 19458 9996 19458 9996 0 net141
rlabel metal1 21574 12818 21574 12818 0 net142
rlabel metal1 23220 6290 23220 6290 0 net143
rlabel metal1 21482 6868 21482 6868 0 net144
rlabel metal1 18395 6290 18395 6290 0 net145
rlabel metal1 21022 4590 21022 4590 0 net146
rlabel metal1 18579 12818 18579 12818 0 net147
rlabel metal1 21390 5712 21390 5712 0 net148
rlabel via1 19366 3025 19366 3025 0 net149
rlabel metal1 7590 18326 7590 18326 0 net15
rlabel metal1 22448 4794 22448 4794 0 net150
rlabel metal1 19642 2414 19642 2414 0 net151
rlabel metal1 22586 1326 22586 1326 0 net152
rlabel via2 11546 17595 11546 17595 0 net153
rlabel metal1 3358 40086 3358 40086 0 net154
rlabel metal1 8142 35734 8142 35734 0 net155
rlabel metal1 13892 16218 13892 16218 0 net156
rlabel metal3 16652 15980 16652 15980 0 net157
rlabel metal1 8050 41242 8050 41242 0 net158
rlabel metal2 7544 38012 7544 38012 0 net159
rlabel metal1 2530 20536 2530 20536 0 net16
rlabel metal3 11247 23460 11247 23460 0 net160
rlabel metal4 13524 10064 13524 10064 0 net161
rlabel via2 12926 43061 12926 43061 0 net162
rlabel metal1 13202 42568 13202 42568 0 net163
rlabel metal3 13961 13668 13961 13668 0 net164
rlabel metal3 13593 42908 13593 42908 0 net165
rlabel metal2 14812 42534 14812 42534 0 net166
rlabel metal2 13294 33201 13294 33201 0 net167
rlabel metal1 13984 42602 13984 42602 0 net168
rlabel via3 14973 42908 14973 42908 0 net169
rlabel metal1 1656 21114 1656 21114 0 net17
rlabel metal2 13386 16337 13386 16337 0 net170
rlabel metal1 13064 30294 13064 30294 0 net171
rlabel metal1 20102 8296 20102 8296 0 net172
rlabel metal1 15226 38726 15226 38726 0 net173
rlabel metal1 18538 42704 18538 42704 0 net174
rlabel metal1 18814 42772 18814 42772 0 net175
rlabel metal2 19642 42500 19642 42500 0 net176
rlabel metal1 19136 41242 19136 41242 0 net177
rlabel metal1 19458 41616 19458 41616 0 net178
rlabel metal1 19826 41106 19826 41106 0 net179
rlabel metal1 1449 20570 1449 20570 0 net18
rlabel metal1 3542 36754 3542 36754 0 net180
rlabel metal2 16882 43520 16882 43520 0 net181
rlabel metal1 12880 12682 12880 12682 0 net182
rlabel metal1 16974 42194 16974 42194 0 net183
rlabel via1 16238 42211 16238 42211 0 net184
rlabel metal1 17480 42670 17480 42670 0 net185
rlabel metal1 17802 42670 17802 42670 0 net186
rlabel metal1 18032 42670 18032 42670 0 net187
rlabel metal2 20102 42942 20102 42942 0 net188
rlabel metal1 23782 8058 23782 8058 0 net189
rlabel metal1 1748 29002 1748 29002 0 net19
rlabel metal1 23552 10710 23552 10710 0 net190
rlabel metal1 23920 10710 23920 10710 0 net191
rlabel metal1 23966 9622 23966 9622 0 net192
rlabel metal1 23690 16626 23690 16626 0 net193
rlabel metal1 24058 16184 24058 16184 0 net194
rlabel metal1 24150 17306 24150 17306 0 net195
rlabel metal1 24012 18734 24012 18734 0 net196
rlabel metal1 23322 12886 23322 12886 0 net197
rlabel metal1 23828 15062 23828 15062 0 net198
rlabel metal1 23736 15470 23736 15470 0 net199
rlabel metal1 5658 20502 5658 20502 0 net2
rlabel metal1 8694 21318 8694 21318 0 net20
rlabel metal1 21482 19720 21482 19720 0 net200
rlabel metal1 20010 13192 20010 13192 0 net201
rlabel metal1 24932 21522 24932 21522 0 net202
rlabel metal2 25668 17612 25668 17612 0 net203
rlabel metal1 23276 13294 23276 13294 0 net204
rlabel metal1 20746 24038 20746 24038 0 net205
rlabel metal1 24058 25942 24058 25942 0 net206
rlabel metal1 23828 27438 23828 27438 0 net207
rlabel metal2 21942 27200 21942 27200 0 net208
rlabel metal2 22586 24344 22586 24344 0 net209
rlabel viali 12834 18260 12834 18260 0 net21
rlabel metal2 24058 23494 24058 23494 0 net210
rlabel metal1 18952 33354 18952 33354 0 net211
rlabel metal1 21574 24820 21574 24820 0 net212
rlabel metal1 23690 20944 23690 20944 0 net213
rlabel metal1 23966 20502 23966 20502 0 net214
rlabel metal1 24840 21998 24840 21998 0 net215
rlabel metal2 20654 22746 20654 22746 0 net216
rlabel metal2 21022 20298 21022 20298 0 net217
rlabel metal1 24104 19414 24104 19414 0 net218
rlabel metal2 21022 31501 21022 31501 0 net219
rlabel metal1 7958 30328 7958 30328 0 net22
rlabel metal2 19274 25568 19274 25568 0 net220
rlabel metal1 23552 27438 23552 27438 0 net221
rlabel metal1 23920 32878 23920 32878 0 net222
rlabel metal1 23782 33558 23782 33558 0 net223
rlabel metal1 23966 33932 23966 33932 0 net224
rlabel metal1 23920 34646 23920 34646 0 net225
rlabel metal1 23460 34714 23460 34714 0 net226
rlabel metal1 23184 35190 23184 35190 0 net227
rlabel metal2 23322 36006 23322 36006 0 net228
rlabel metal1 24104 36822 24104 36822 0 net229
rlabel via2 5566 31467 5566 31467 0 net23
rlabel metal1 23828 36890 23828 36890 0 net230
rlabel metal1 19964 37094 19964 37094 0 net231
rlabel metal1 24150 28152 24150 28152 0 net232
rlabel metal1 21206 37978 21206 37978 0 net233
rlabel metal1 23782 38522 23782 38522 0 net234
rlabel metal1 23966 39440 23966 39440 0 net235
rlabel metal1 20930 38760 20930 38760 0 net236
rlabel metal2 20838 39389 20838 39389 0 net237
rlabel metal1 23000 40154 23000 40154 0 net238
rlabel metal1 21620 40630 21620 40630 0 net239
rlabel metal2 2622 28152 2622 28152 0 net24
rlabel metal1 19918 41446 19918 41446 0 net240
rlabel metal1 23184 39610 23184 39610 0 net241
rlabel metal1 20332 40698 20332 40698 0 net242
rlabel metal2 23966 28730 23966 28730 0 net243
rlabel metal1 23138 40698 23138 40698 0 net244
rlabel metal2 21022 41021 21022 41021 0 net245
rlabel metal1 21804 28186 21804 28186 0 net246
rlabel metal1 23690 29546 23690 29546 0 net247
rlabel metal1 23782 30294 23782 30294 0 net248
rlabel metal1 23598 30022 23598 30022 0 net249
rlabel metal1 1840 21862 1840 21862 0 net25
rlabel metal2 23046 31144 23046 31144 0 net250
rlabel metal1 23874 31824 23874 31824 0 net251
rlabel metal1 24150 32504 24150 32504 0 net252
rlabel metal1 20470 42330 20470 42330 0 net253
rlabel metal2 23460 42670 23460 42670 0 net254
rlabel metal1 21758 40154 21758 40154 0 net255
rlabel metal1 22931 42126 22931 42126 0 net256
rlabel metal1 20378 40902 20378 40902 0 net257
rlabel metal1 22816 42194 22816 42194 0 net258
rlabel metal1 23276 39882 23276 39882 0 net259
rlabel metal1 16652 16082 16652 16082 0 net26
rlabel metal1 23644 41446 23644 41446 0 net260
rlabel metal1 20010 40120 20010 40120 0 net261
rlabel metal2 23230 37842 23230 37842 0 net262
rlabel metal1 21298 42092 21298 42092 0 net263
rlabel metal1 20884 42330 20884 42330 0 net264
rlabel metal1 20930 40698 20930 40698 0 net265
rlabel metal1 21390 41786 21390 41786 0 net266
rlabel metal2 22126 43231 22126 43231 0 net267
rlabel metal2 22678 43520 22678 43520 0 net268
rlabel metal1 21896 40358 21896 40358 0 net269
rlabel metal1 10258 29070 10258 29070 0 net27
rlabel metal1 22540 42602 22540 42602 0 net270
rlabel metal1 21252 41242 21252 41242 0 net271
rlabel metal1 23046 42602 23046 42602 0 net272
rlabel metal1 11178 42296 11178 42296 0 net273
rlabel metal1 3634 41786 3634 41786 0 net274
rlabel metal2 12558 42432 12558 42432 0 net275
rlabel via2 2530 42211 2530 42211 0 net276
rlabel metal1 3726 40698 3726 40698 0 net277
rlabel metal1 4738 40970 4738 40970 0 net278
rlabel metal1 3027 41174 3027 41174 0 net279
rlabel metal2 3450 24344 3450 24344 0 net28
rlabel metal1 1794 43690 1794 43690 0 net280
rlabel metal1 3634 43384 3634 43384 0 net281
rlabel metal1 3266 39542 3266 39542 0 net282
rlabel metal1 2852 40154 2852 40154 0 net283
rlabel metal2 5842 41321 5842 41321 0 net284
rlabel metal1 4094 39610 4094 39610 0 net285
rlabel metal1 6486 40970 6486 40970 0 net286
rlabel metal1 4922 42534 4922 42534 0 net287
rlabel metal1 4186 40698 4186 40698 0 net288
rlabel metal1 6762 41242 6762 41242 0 net289
rlabel metal1 6394 29172 6394 29172 0 net29
rlabel metal1 4875 42602 4875 42602 0 net290
rlabel metal1 4830 41786 4830 41786 0 net291
rlabel metal1 5106 43214 5106 43214 0 net292
rlabel metal2 5474 42534 5474 42534 0 net293
rlabel metal1 8648 42874 8648 42874 0 net294
rlabel metal1 8832 42602 8832 42602 0 net295
rlabel metal1 10534 42534 10534 42534 0 net296
rlabel metal1 8694 40970 8694 40970 0 net297
rlabel metal1 10074 42806 10074 42806 0 net298
rlabel metal1 16974 42806 16974 42806 0 net299
rlabel metal2 12558 35088 12558 35088 0 net3
rlabel metal1 8096 24854 8096 24854 0 net30
rlabel metal1 6118 41786 6118 41786 0 net300
rlabel metal2 5566 42874 5566 42874 0 net301
rlabel metal2 6854 41939 6854 41939 0 net302
rlabel metal1 6762 43384 6762 43384 0 net303
rlabel metal2 7314 42194 7314 42194 0 net304
rlabel metal2 5842 42024 5842 42024 0 net305
rlabel metal1 7682 41786 7682 41786 0 net306
rlabel metal1 7820 41446 7820 41446 0 net307
rlabel metal2 8418 41990 8418 41990 0 net308
rlabel metal2 9614 1802 9614 1802 0 net309
rlabel metal1 1702 30668 1702 30668 0 net31
rlabel metal1 10166 1326 10166 1326 0 net310
rlabel metal1 10718 2346 10718 2346 0 net311
rlabel metal1 15318 2516 15318 2516 0 net312
rlabel metal1 13248 1326 13248 1326 0 net313
rlabel metal1 13662 1258 13662 1258 0 net314
rlabel metal1 14214 1326 14214 1326 0 net315
rlabel metal1 14490 1904 14490 1904 0 net316
rlabel metal1 14904 1938 14904 1938 0 net317
rlabel metal1 15042 1326 15042 1326 0 net318
rlabel metal1 15226 1258 15226 1258 0 net319
rlabel metal1 5060 34578 5060 34578 0 net32
rlabel metal1 16238 1530 16238 1530 0 net320
rlabel metal2 10902 1972 10902 1972 0 net321
rlabel metal1 11684 1326 11684 1326 0 net322
rlabel metal1 13662 2040 13662 2040 0 net323
rlabel metal2 13386 2176 13386 2176 0 net324
rlabel metal1 12650 1394 12650 1394 0 net325
rlabel metal2 8970 1054 8970 1054 0 net326
rlabel metal2 12466 1904 12466 1904 0 net327
rlabel metal2 13662 1530 13662 1530 0 net328
rlabel metal1 15778 2006 15778 2006 0 net329
rlabel metal1 12098 25194 12098 25194 0 net33
rlabel metal1 23460 1802 23460 1802 0 net330
rlabel metal1 17112 1938 17112 1938 0 net331
rlabel metal1 21390 1190 21390 1190 0 net332
rlabel metal1 18906 1224 18906 1224 0 net333
rlabel metal2 18906 3740 18906 3740 0 net334
rlabel metal1 20930 3434 20930 3434 0 net335
rlabel metal1 16744 1326 16744 1326 0 net336
rlabel metal1 17296 1326 17296 1326 0 net337
rlabel metal1 17802 1326 17802 1326 0 net338
rlabel metal1 17066 2006 17066 2006 0 net339
rlabel metal1 9522 35530 9522 35530 0 net34
rlabel metal1 18814 2006 18814 2006 0 net340
rlabel metal1 19412 2074 19412 2074 0 net341
rlabel metal1 17526 2346 17526 2346 0 net342
rlabel metal1 17756 2006 17756 2006 0 net343
rlabel via2 19251 2652 19251 2652 0 net344
rlabel metal1 21574 41616 21574 41616 0 net345
rlabel metal1 2139 4182 2139 4182 0 net346
rlabel metal2 2346 5066 2346 5066 0 net347
rlabel metal1 2576 4794 2576 4794 0 net348
rlabel metal1 1518 4658 1518 4658 0 net349
rlabel metal1 6394 27098 6394 27098 0 net35
rlabel metal1 1886 5882 1886 5882 0 net350
rlabel metal2 2070 5950 2070 5950 0 net351
rlabel metal1 3818 6766 3818 6766 0 net352
rlabel metal1 4922 6086 4922 6086 0 net353
rlabel metal1 2024 5202 2024 5202 0 net354
rlabel metal1 3496 7446 3496 7446 0 net355
rlabel metal1 3128 6426 3128 6426 0 net356
rlabel metal1 2254 4488 2254 4488 0 net357
rlabel metal1 2530 6358 2530 6358 0 net358
rlabel metal1 2070 7344 2070 7344 0 net359
rlabel metal1 9522 27404 9522 27404 0 net36
rlabel metal1 3266 8976 3266 8976 0 net360
rlabel metal2 1978 7174 1978 7174 0 net361
rlabel metal2 2714 7378 2714 7378 0 net362
rlabel metal1 1610 8398 1610 8398 0 net363
rlabel metal1 1886 9146 1886 9146 0 net364
rlabel metal1 1472 3706 1472 3706 0 net365
rlabel metal1 1886 13294 1886 13294 0 net366
rlabel metal1 3220 17238 3220 17238 0 net367
rlabel metal2 1518 17544 1518 17544 0 net368
rlabel metal2 1702 39389 1702 39389 0 net369
rlabel metal1 4232 25942 4232 25942 0 net37
rlabel metal3 1932 20944 1932 20944 0 net370
rlabel metal1 13754 15368 13754 15368 0 net371
rlabel metal1 1518 14416 1518 14416 0 net372
rlabel metal1 1932 15062 1932 15062 0 net373
rlabel metal1 1426 16456 1426 16456 0 net374
rlabel metal1 10304 16218 10304 16218 0 net375
rlabel via2 2254 17187 2254 17187 0 net376
rlabel metal1 2231 17238 2231 17238 0 net377
rlabel metal1 2944 9622 2944 9622 0 net378
rlabel metal1 2070 13974 2070 13974 0 net379
rlabel metal1 8602 29580 8602 29580 0 net38
rlabel metal1 6624 13294 6624 13294 0 net380
rlabel metal1 2484 14382 2484 14382 0 net381
rlabel metal1 2346 12784 2346 12784 0 net382
rlabel metal2 1426 13056 1426 13056 0 net383
rlabel metal2 2162 10625 2162 10625 0 net384
rlabel metal1 3588 9690 3588 9690 0 net385
rlabel metal1 1702 9520 1702 9520 0 net386
rlabel metal1 3174 9996 3174 9996 0 net387
rlabel metal1 5612 10778 5612 10778 0 net388
rlabel metal1 3312 11866 3312 11866 0 net389
rlabel via1 17078 26350 17078 26350 0 net39
rlabel metal1 1748 9962 1748 9962 0 net390
rlabel metal1 3082 10064 3082 10064 0 net391
rlabel metal1 1518 10744 1518 10744 0 net392
rlabel metal2 1978 10336 1978 10336 0 net393
rlabel metal1 14076 16150 14076 16150 0 net394
rlabel metal1 16606 18802 16606 18802 0 net395
rlabel metal1 7590 20842 7590 20842 0 net396
rlabel metal1 6210 18292 6210 18292 0 net397
rlabel metal1 15594 22406 15594 22406 0 net398
rlabel metal2 16330 23630 16330 23630 0 net399
rlabel metal2 16882 20417 16882 20417 0 net4
rlabel metal1 5014 28390 5014 28390 0 net40
rlabel metal1 8694 22678 8694 22678 0 net400
rlabel metal1 6348 25194 6348 25194 0 net401
rlabel metal1 12742 20468 12742 20468 0 net402
rlabel metal2 13800 18258 13800 18258 0 net403
rlabel metal2 4278 33082 4278 33082 0 net404
rlabel metal1 13340 38386 13340 38386 0 net405
rlabel metal1 11914 17646 11914 17646 0 net406
rlabel metal1 2530 36618 2530 36618 0 net407
rlabel via1 10810 40579 10810 40579 0 net408
rlabel metal2 17986 16864 17986 16864 0 net409
rlabel metal2 2162 25653 2162 25653 0 net41
rlabel metal2 15456 32878 15456 32878 0 net42
rlabel metal2 1610 25568 1610 25568 0 net43
rlabel metal1 3404 24922 3404 24922 0 net44
rlabel metal2 2162 26231 2162 26231 0 net45
rlabel metal2 1610 26401 1610 26401 0 net46
rlabel metal1 11592 25330 11592 25330 0 net47
rlabel metal1 4738 28424 4738 28424 0 net48
rlabel metal1 19533 13906 19533 13906 0 net49
rlabel metal2 2162 21097 2162 21097 0 net5
rlabel metal1 19366 33320 19366 33320 0 net50
rlabel metal1 21298 33932 21298 33932 0 net51
rlabel metal1 21528 33966 21528 33966 0 net52
rlabel metal1 21850 21080 21850 21080 0 net53
rlabel viali 18345 32432 18345 32432 0 net54
rlabel metal2 13478 7684 13478 7684 0 net55
rlabel metal1 20010 20910 20010 20910 0 net56
rlabel metal1 13155 36142 13155 36142 0 net57
rlabel metal1 2023 16558 2023 16558 0 net58
rlabel metal1 2989 21522 2989 21522 0 net59
rlabel metal1 7682 27030 7682 27030 0 net6
rlabel metal1 22155 31314 22155 31314 0 net60
rlabel metal1 19734 36788 19734 36788 0 net61
rlabel metal1 1978 38930 1978 38930 0 net62
rlabel metal1 2346 38794 2346 38794 0 net63
rlabel metal1 18354 37876 18354 37876 0 net64
rlabel metal2 19872 19890 19872 19890 0 net65
rlabel metal2 21022 17476 21022 17476 0 net66
rlabel metal2 2254 39729 2254 39729 0 net67
rlabel metal1 2392 38386 2392 38386 0 net68
rlabel metal1 2116 42602 2116 42602 0 net69
rlabel metal2 7360 18258 7360 18258 0 net7
rlabel metal1 21206 16048 21206 16048 0 net70
rlabel via3 1955 38692 1955 38692 0 net71
rlabel via2 2254 42109 2254 42109 0 net72
rlabel viali 20093 19792 20093 19792 0 net73
rlabel metal2 2714 33065 2714 33065 0 net74
rlabel via2 2714 16099 2714 16099 0 net75
rlabel metal2 1978 6868 1978 6868 0 net76
rlabel metal1 15869 30226 15869 30226 0 net77
rlabel metal1 21482 11628 21482 11628 0 net78
rlabel via2 1702 35581 1702 35581 0 net79
rlabel metal1 14490 21964 14490 21964 0 net8
rlabel metal3 16376 20740 16376 20740 0 net80
rlabel metal1 2070 39508 2070 39508 0 net81
rlabel via2 20746 6715 20746 6715 0 net82
rlabel metal1 23966 2414 23966 2414 0 net83
rlabel metal1 24472 38998 24472 38998 0 net84
rlabel metal2 20148 10778 20148 10778 0 net85
rlabel metal2 21436 18020 21436 18020 0 net86
rlabel metal1 21160 3910 21160 3910 0 net87
rlabel metal2 16974 9724 16974 9724 0 net88
rlabel metal2 24472 14348 24472 14348 0 net89
rlabel metal1 1702 23528 1702 23528 0 net9
rlabel metal1 20148 1938 20148 1938 0 net90
rlabel metal2 22586 5423 22586 5423 0 net91
rlabel metal1 2346 40460 2346 40460 0 net92
rlabel metal2 21574 15317 21574 15317 0 net93
rlabel metal1 18262 40562 18262 40562 0 net94
rlabel metal1 21620 2346 21620 2346 0 net95
rlabel metal1 1426 19380 1426 19380 0 net96
rlabel metal2 21252 40732 21252 40732 0 net97
rlabel metal1 17710 20366 17710 20366 0 net98
rlabel metal1 17940 19686 17940 19686 0 net99
rlabel metal1 19918 41786 19918 41786 0 strobe_inbuf_0.X
rlabel metal1 20286 41786 20286 41786 0 strobe_inbuf_1.X
rlabel metal3 21367 38692 21367 38692 0 strobe_inbuf_10.X
rlabel metal1 24380 2618 24380 2618 0 strobe_inbuf_11.X
rlabel metal2 23506 39151 23506 39151 0 strobe_inbuf_12.X
rlabel metal1 23460 36142 23460 36142 0 strobe_inbuf_13.X
rlabel metal2 23414 38454 23414 38454 0 strobe_inbuf_14.X
rlabel metal1 23506 36890 23506 36890 0 strobe_inbuf_15.X
rlabel metal1 23828 31450 23828 31450 0 strobe_inbuf_16.X
rlabel metal1 23460 37094 23460 37094 0 strobe_inbuf_17.X
rlabel metal2 22770 34374 22770 34374 0 strobe_inbuf_18.X
rlabel metal1 23874 22644 23874 22644 0 strobe_inbuf_19.X
rlabel metal1 20608 39066 20608 39066 0 strobe_inbuf_2.X
rlabel metal1 20562 41242 20562 41242 0 strobe_inbuf_3.X
rlabel metal1 21022 40902 21022 40902 0 strobe_inbuf_4.X
rlabel metal1 21804 20026 21804 20026 0 strobe_inbuf_5.X
rlabel metal1 20470 40494 20470 40494 0 strobe_inbuf_6.X
rlabel viali 21390 40030 21390 40030 0 strobe_inbuf_7.X
rlabel metal1 22402 39542 22402 39542 0 strobe_inbuf_8.X
rlabel metal1 22724 35802 22724 35802 0 strobe_inbuf_9.X
rlabel metal1 20746 42160 20746 42160 0 strobe_outbuf_0.X
rlabel metal1 21022 42126 21022 42126 0 strobe_outbuf_1.X
rlabel metal1 21298 39610 21298 39610 0 strobe_outbuf_10.X
rlabel metal1 21942 39984 21942 39984 0 strobe_outbuf_11.X
rlabel metal2 19918 40273 19918 40273 0 strobe_outbuf_12.X
rlabel metal1 22494 36312 22494 36312 0 strobe_outbuf_13.X
rlabel metal1 23184 39066 23184 39066 0 strobe_outbuf_14.X
rlabel metal1 23552 39066 23552 39066 0 strobe_outbuf_15.X
rlabel metal1 23736 33626 23736 33626 0 strobe_outbuf_16.X
rlabel metal2 20194 39967 20194 39967 0 strobe_outbuf_17.X
rlabel metal1 23460 35054 23460 35054 0 strobe_outbuf_18.X
rlabel metal1 23736 22746 23736 22746 0 strobe_outbuf_19.X
rlabel metal1 20746 40154 20746 40154 0 strobe_outbuf_2.X
rlabel metal1 21390 41582 21390 41582 0 strobe_outbuf_3.X
rlabel metal1 20746 41446 20746 41446 0 strobe_outbuf_4.X
rlabel metal2 19366 41684 19366 41684 0 strobe_outbuf_5.X
rlabel metal1 21942 40494 21942 40494 0 strobe_outbuf_6.X
rlabel metal1 21252 39882 21252 39882 0 strobe_outbuf_7.X
rlabel metal1 21390 41072 21390 41072 0 strobe_outbuf_8.X
rlabel metal1 23046 36176 23046 36176 0 strobe_outbuf_9.X
<< properties >>
string FIXED_BBOX 0 0 26000 45000
<< end >>
