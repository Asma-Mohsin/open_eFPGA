magic
tech sky130A
magscale 1 2
timestamp 1733308305
<< obsli1 >>
rect 1104 1071 46828 43537
<< obsm1 >>
rect 14 620 47918 44124
<< metal2 >>
rect 1122 44840 1178 45000
rect 1490 44840 1546 45000
rect 1858 44840 1914 45000
rect 2226 44840 2282 45000
rect 2594 44840 2650 45000
rect 2962 44840 3018 45000
rect 3330 44840 3386 45000
rect 3698 44840 3754 45000
rect 4066 44840 4122 45000
rect 4434 44840 4490 45000
rect 4802 44840 4858 45000
rect 5170 44840 5226 45000
rect 5538 44840 5594 45000
rect 5906 44840 5962 45000
rect 6274 44840 6330 45000
rect 6642 44840 6698 45000
rect 7010 44840 7066 45000
rect 7378 44840 7434 45000
rect 7746 44840 7802 45000
rect 8114 44840 8170 45000
rect 8482 44840 8538 45000
rect 8850 44840 8906 45000
rect 9218 44840 9274 45000
rect 9586 44840 9642 45000
rect 9954 44840 10010 45000
rect 10322 44840 10378 45000
rect 10690 44840 10746 45000
rect 11058 44840 11114 45000
rect 11426 44840 11482 45000
rect 11794 44840 11850 45000
rect 12162 44840 12218 45000
rect 12530 44840 12586 45000
rect 12898 44840 12954 45000
rect 13266 44840 13322 45000
rect 13634 44840 13690 45000
rect 14002 44840 14058 45000
rect 14370 44840 14426 45000
rect 14738 44840 14794 45000
rect 15106 44840 15162 45000
rect 15474 44840 15530 45000
rect 15842 44840 15898 45000
rect 16210 44840 16266 45000
rect 16578 44840 16634 45000
rect 16946 44840 17002 45000
rect 17314 44840 17370 45000
rect 17682 44840 17738 45000
rect 18050 44840 18106 45000
rect 18418 44840 18474 45000
rect 18786 44840 18842 45000
rect 19154 44840 19210 45000
rect 19522 44840 19578 45000
rect 19890 44840 19946 45000
rect 20258 44840 20314 45000
rect 20626 44840 20682 45000
rect 20994 44840 21050 45000
rect 21362 44840 21418 45000
rect 21730 44840 21786 45000
rect 22098 44840 22154 45000
rect 22466 44840 22522 45000
rect 22834 44840 22890 45000
rect 23202 44840 23258 45000
rect 23570 44840 23626 45000
rect 23938 44840 23994 45000
rect 24306 44840 24362 45000
rect 24674 44840 24730 45000
rect 25042 44840 25098 45000
rect 25410 44840 25466 45000
rect 25778 44840 25834 45000
rect 26146 44840 26202 45000
rect 26514 44840 26570 45000
rect 26882 44840 26938 45000
rect 27250 44840 27306 45000
rect 27618 44840 27674 45000
rect 27986 44840 28042 45000
rect 28354 44840 28410 45000
rect 28722 44840 28778 45000
rect 29090 44840 29146 45000
rect 29458 44840 29514 45000
rect 29826 44840 29882 45000
rect 30194 44840 30250 45000
rect 30562 44840 30618 45000
rect 30930 44840 30986 45000
rect 31298 44840 31354 45000
rect 31666 44840 31722 45000
rect 32034 44840 32090 45000
rect 32402 44840 32458 45000
rect 32770 44840 32826 45000
rect 33138 44840 33194 45000
rect 33506 44840 33562 45000
rect 33874 44840 33930 45000
rect 34242 44840 34298 45000
rect 34610 44840 34666 45000
rect 34978 44840 35034 45000
rect 35346 44840 35402 45000
rect 35714 44840 35770 45000
rect 36082 44840 36138 45000
rect 36450 44840 36506 45000
rect 36818 44840 36874 45000
rect 37186 44840 37242 45000
rect 37554 44840 37610 45000
rect 37922 44840 37978 45000
rect 38290 44840 38346 45000
rect 38658 44840 38714 45000
rect 39026 44840 39082 45000
rect 39394 44840 39450 45000
rect 39762 44840 39818 45000
rect 40130 44840 40186 45000
rect 40498 44840 40554 45000
rect 40866 44840 40922 45000
rect 41234 44840 41290 45000
rect 41602 44840 41658 45000
rect 41970 44840 42026 45000
rect 42338 44840 42394 45000
rect 42706 44840 42762 45000
rect 43074 44840 43130 45000
rect 43442 44840 43498 45000
rect 43810 44840 43866 45000
rect 44178 44840 44234 45000
rect 44546 44840 44602 45000
rect 44914 44840 44970 45000
rect 45282 44840 45338 45000
rect 45650 44840 45706 45000
rect 46018 44840 46074 45000
rect 46386 44840 46442 45000
rect 46754 44840 46810 45000
rect 1122 0 1178 160
rect 1490 0 1546 160
rect 1858 0 1914 160
rect 2226 0 2282 160
rect 2594 0 2650 160
rect 2962 0 3018 160
rect 3330 0 3386 160
rect 3698 0 3754 160
rect 4066 0 4122 160
rect 4434 0 4490 160
rect 4802 0 4858 160
rect 5170 0 5226 160
rect 5538 0 5594 160
rect 5906 0 5962 160
rect 6274 0 6330 160
rect 6642 0 6698 160
rect 7010 0 7066 160
rect 7378 0 7434 160
rect 7746 0 7802 160
rect 8114 0 8170 160
rect 8482 0 8538 160
rect 8850 0 8906 160
rect 9218 0 9274 160
rect 9586 0 9642 160
rect 9954 0 10010 160
rect 10322 0 10378 160
rect 10690 0 10746 160
rect 11058 0 11114 160
rect 11426 0 11482 160
rect 11794 0 11850 160
rect 12162 0 12218 160
rect 12530 0 12586 160
rect 12898 0 12954 160
rect 13266 0 13322 160
rect 13634 0 13690 160
rect 14002 0 14058 160
rect 14370 0 14426 160
rect 14738 0 14794 160
rect 15106 0 15162 160
rect 15474 0 15530 160
rect 15842 0 15898 160
rect 16210 0 16266 160
rect 16578 0 16634 160
rect 16946 0 17002 160
rect 17314 0 17370 160
rect 17682 0 17738 160
rect 18050 0 18106 160
rect 18418 0 18474 160
rect 18786 0 18842 160
rect 19154 0 19210 160
rect 19522 0 19578 160
rect 19890 0 19946 160
rect 20258 0 20314 160
rect 20626 0 20682 160
rect 20994 0 21050 160
rect 21362 0 21418 160
rect 21730 0 21786 160
rect 22098 0 22154 160
rect 22466 0 22522 160
rect 22834 0 22890 160
rect 23202 0 23258 160
rect 23570 0 23626 160
rect 23938 0 23994 160
rect 24306 0 24362 160
rect 24674 0 24730 160
rect 25042 0 25098 160
rect 25410 0 25466 160
rect 25778 0 25834 160
rect 26146 0 26202 160
rect 26514 0 26570 160
rect 26882 0 26938 160
rect 27250 0 27306 160
rect 27618 0 27674 160
rect 27986 0 28042 160
rect 28354 0 28410 160
rect 28722 0 28778 160
rect 29090 0 29146 160
rect 29458 0 29514 160
rect 29826 0 29882 160
rect 30194 0 30250 160
rect 30562 0 30618 160
rect 30930 0 30986 160
rect 31298 0 31354 160
rect 31666 0 31722 160
rect 32034 0 32090 160
rect 32402 0 32458 160
rect 32770 0 32826 160
rect 33138 0 33194 160
rect 33506 0 33562 160
rect 33874 0 33930 160
rect 34242 0 34298 160
rect 34610 0 34666 160
rect 34978 0 35034 160
rect 35346 0 35402 160
rect 35714 0 35770 160
rect 36082 0 36138 160
rect 36450 0 36506 160
rect 36818 0 36874 160
rect 37186 0 37242 160
rect 37554 0 37610 160
rect 37922 0 37978 160
rect 38290 0 38346 160
rect 38658 0 38714 160
rect 39026 0 39082 160
rect 39394 0 39450 160
rect 39762 0 39818 160
rect 40130 0 40186 160
rect 40498 0 40554 160
rect 40866 0 40922 160
rect 41234 0 41290 160
rect 41602 0 41658 160
rect 41970 0 42026 160
rect 42338 0 42394 160
rect 42706 0 42762 160
rect 43074 0 43130 160
rect 43442 0 43498 160
rect 43810 0 43866 160
rect 44178 0 44234 160
rect 44546 0 44602 160
rect 44914 0 44970 160
rect 45282 0 45338 160
rect 45650 0 45706 160
rect 46018 0 46074 160
rect 46386 0 46442 160
rect 46754 0 46810 160
<< obsm2 >>
rect 20 44784 1066 44962
rect 1234 44784 1434 44962
rect 1602 44784 1802 44962
rect 1970 44784 2170 44962
rect 2338 44784 2538 44962
rect 2706 44784 2906 44962
rect 3074 44784 3274 44962
rect 3442 44784 3642 44962
rect 3810 44784 4010 44962
rect 4178 44784 4378 44962
rect 4546 44784 4746 44962
rect 4914 44784 5114 44962
rect 5282 44784 5482 44962
rect 5650 44784 5850 44962
rect 6018 44784 6218 44962
rect 6386 44784 6586 44962
rect 6754 44784 6954 44962
rect 7122 44784 7322 44962
rect 7490 44784 7690 44962
rect 7858 44784 8058 44962
rect 8226 44784 8426 44962
rect 8594 44784 8794 44962
rect 8962 44784 9162 44962
rect 9330 44784 9530 44962
rect 9698 44784 9898 44962
rect 10066 44784 10266 44962
rect 10434 44784 10634 44962
rect 10802 44784 11002 44962
rect 11170 44784 11370 44962
rect 11538 44784 11738 44962
rect 11906 44784 12106 44962
rect 12274 44784 12474 44962
rect 12642 44784 12842 44962
rect 13010 44784 13210 44962
rect 13378 44784 13578 44962
rect 13746 44784 13946 44962
rect 14114 44784 14314 44962
rect 14482 44784 14682 44962
rect 14850 44784 15050 44962
rect 15218 44784 15418 44962
rect 15586 44784 15786 44962
rect 15954 44784 16154 44962
rect 16322 44784 16522 44962
rect 16690 44784 16890 44962
rect 17058 44784 17258 44962
rect 17426 44784 17626 44962
rect 17794 44784 17994 44962
rect 18162 44784 18362 44962
rect 18530 44784 18730 44962
rect 18898 44784 19098 44962
rect 19266 44784 19466 44962
rect 19634 44784 19834 44962
rect 20002 44784 20202 44962
rect 20370 44784 20570 44962
rect 20738 44784 20938 44962
rect 21106 44784 21306 44962
rect 21474 44784 21674 44962
rect 21842 44784 22042 44962
rect 22210 44784 22410 44962
rect 22578 44784 22778 44962
rect 22946 44784 23146 44962
rect 23314 44784 23514 44962
rect 23682 44784 23882 44962
rect 24050 44784 24250 44962
rect 24418 44784 24618 44962
rect 24786 44784 24986 44962
rect 25154 44784 25354 44962
rect 25522 44784 25722 44962
rect 25890 44784 26090 44962
rect 26258 44784 26458 44962
rect 26626 44784 26826 44962
rect 26994 44784 27194 44962
rect 27362 44784 27562 44962
rect 27730 44784 27930 44962
rect 28098 44784 28298 44962
rect 28466 44784 28666 44962
rect 28834 44784 29034 44962
rect 29202 44784 29402 44962
rect 29570 44784 29770 44962
rect 29938 44784 30138 44962
rect 30306 44784 30506 44962
rect 30674 44784 30874 44962
rect 31042 44784 31242 44962
rect 31410 44784 31610 44962
rect 31778 44784 31978 44962
rect 32146 44784 32346 44962
rect 32514 44784 32714 44962
rect 32882 44784 33082 44962
rect 33250 44784 33450 44962
rect 33618 44784 33818 44962
rect 33986 44784 34186 44962
rect 34354 44784 34554 44962
rect 34722 44784 34922 44962
rect 35090 44784 35290 44962
rect 35458 44784 35658 44962
rect 35826 44784 36026 44962
rect 36194 44784 36394 44962
rect 36562 44784 36762 44962
rect 36930 44784 37130 44962
rect 37298 44784 37498 44962
rect 37666 44784 37866 44962
rect 38034 44784 38234 44962
rect 38402 44784 38602 44962
rect 38770 44784 38970 44962
rect 39138 44784 39338 44962
rect 39506 44784 39706 44962
rect 39874 44784 40074 44962
rect 40242 44784 40442 44962
rect 40610 44784 40810 44962
rect 40978 44784 41178 44962
rect 41346 44784 41546 44962
rect 41714 44784 41914 44962
rect 42082 44784 42282 44962
rect 42450 44784 42650 44962
rect 42818 44784 43018 44962
rect 43186 44784 43386 44962
rect 43554 44784 43754 44962
rect 43922 44784 44122 44962
rect 44290 44784 44490 44962
rect 44658 44784 44858 44962
rect 45026 44784 45226 44962
rect 45394 44784 45594 44962
rect 45762 44784 45962 44962
rect 46130 44784 46330 44962
rect 46498 44784 46698 44962
rect 46866 44784 47992 44962
rect 20 216 47992 44784
rect 20 54 1066 216
rect 1234 54 1434 216
rect 1602 54 1802 216
rect 1970 54 2170 216
rect 2338 54 2538 216
rect 2706 54 2906 216
rect 3074 54 3274 216
rect 3442 54 3642 216
rect 3810 54 4010 216
rect 4178 54 4378 216
rect 4546 54 4746 216
rect 4914 54 5114 216
rect 5282 54 5482 216
rect 5650 54 5850 216
rect 6018 54 6218 216
rect 6386 54 6586 216
rect 6754 54 6954 216
rect 7122 54 7322 216
rect 7490 54 7690 216
rect 7858 54 8058 216
rect 8226 54 8426 216
rect 8594 54 8794 216
rect 8962 54 9162 216
rect 9330 54 9530 216
rect 9698 54 9898 216
rect 10066 54 10266 216
rect 10434 54 10634 216
rect 10802 54 11002 216
rect 11170 54 11370 216
rect 11538 54 11738 216
rect 11906 54 12106 216
rect 12274 54 12474 216
rect 12642 54 12842 216
rect 13010 54 13210 216
rect 13378 54 13578 216
rect 13746 54 13946 216
rect 14114 54 14314 216
rect 14482 54 14682 216
rect 14850 54 15050 216
rect 15218 54 15418 216
rect 15586 54 15786 216
rect 15954 54 16154 216
rect 16322 54 16522 216
rect 16690 54 16890 216
rect 17058 54 17258 216
rect 17426 54 17626 216
rect 17794 54 17994 216
rect 18162 54 18362 216
rect 18530 54 18730 216
rect 18898 54 19098 216
rect 19266 54 19466 216
rect 19634 54 19834 216
rect 20002 54 20202 216
rect 20370 54 20570 216
rect 20738 54 20938 216
rect 21106 54 21306 216
rect 21474 54 21674 216
rect 21842 54 22042 216
rect 22210 54 22410 216
rect 22578 54 22778 216
rect 22946 54 23146 216
rect 23314 54 23514 216
rect 23682 54 23882 216
rect 24050 54 24250 216
rect 24418 54 24618 216
rect 24786 54 24986 216
rect 25154 54 25354 216
rect 25522 54 25722 216
rect 25890 54 26090 216
rect 26258 54 26458 216
rect 26626 54 26826 216
rect 26994 54 27194 216
rect 27362 54 27562 216
rect 27730 54 27930 216
rect 28098 54 28298 216
rect 28466 54 28666 216
rect 28834 54 29034 216
rect 29202 54 29402 216
rect 29570 54 29770 216
rect 29938 54 30138 216
rect 30306 54 30506 216
rect 30674 54 30874 216
rect 31042 54 31242 216
rect 31410 54 31610 216
rect 31778 54 31978 216
rect 32146 54 32346 216
rect 32514 54 32714 216
rect 32882 54 33082 216
rect 33250 54 33450 216
rect 33618 54 33818 216
rect 33986 54 34186 216
rect 34354 54 34554 216
rect 34722 54 34922 216
rect 35090 54 35290 216
rect 35458 54 35658 216
rect 35826 54 36026 216
rect 36194 54 36394 216
rect 36562 54 36762 216
rect 36930 54 37130 216
rect 37298 54 37498 216
rect 37666 54 37866 216
rect 38034 54 38234 216
rect 38402 54 38602 216
rect 38770 54 38970 216
rect 39138 54 39338 216
rect 39506 54 39706 216
rect 39874 54 40074 216
rect 40242 54 40442 216
rect 40610 54 40810 216
rect 40978 54 41178 216
rect 41346 54 41546 216
rect 41714 54 41914 216
rect 42082 54 42282 216
rect 42450 54 42650 216
rect 42818 54 43018 216
rect 43186 54 43386 216
rect 43554 54 43754 216
rect 43922 54 44122 216
rect 44290 54 44490 216
rect 44658 54 44858 216
rect 45026 54 45226 216
rect 45394 54 45594 216
rect 45762 54 45962 216
rect 46130 54 46330 216
rect 46498 54 46698 216
rect 46866 54 47992 216
<< metal3 >>
rect 0 39720 160 39840
rect 0 39448 160 39568
rect 0 39176 160 39296
rect 0 38904 160 39024
rect 0 38632 160 38752
rect 0 38360 160 38480
rect 0 38088 160 38208
rect 0 37816 160 37936
rect 0 37544 160 37664
rect 0 37272 160 37392
rect 0 37000 160 37120
rect 0 36728 160 36848
rect 0 36456 160 36576
rect 0 36184 160 36304
rect 0 35912 160 36032
rect 0 35640 160 35760
rect 0 35368 160 35488
rect 0 35096 160 35216
rect 0 34824 160 34944
rect 0 34552 160 34672
rect 0 34280 160 34400
rect 0 34008 160 34128
rect 0 33736 160 33856
rect 0 33464 160 33584
rect 0 33192 160 33312
rect 0 32920 160 33040
rect 0 32648 160 32768
rect 0 32376 160 32496
rect 0 32104 160 32224
rect 0 31832 160 31952
rect 0 31560 160 31680
rect 0 31288 160 31408
rect 0 31016 160 31136
rect 0 30744 160 30864
rect 0 30472 160 30592
rect 0 30200 160 30320
rect 0 29928 160 30048
rect 0 29656 160 29776
rect 0 29384 160 29504
rect 0 29112 160 29232
rect 0 28840 160 28960
rect 0 28568 160 28688
rect 0 28296 160 28416
rect 0 28024 160 28144
rect 0 27752 160 27872
rect 0 27480 160 27600
rect 0 27208 160 27328
rect 0 26936 160 27056
rect 0 26664 160 26784
rect 0 26392 160 26512
rect 0 26120 160 26240
rect 0 25848 160 25968
rect 0 25576 160 25696
rect 0 25304 160 25424
rect 0 25032 160 25152
rect 0 24760 160 24880
rect 0 24488 160 24608
rect 0 24216 160 24336
rect 0 23944 160 24064
rect 0 23672 160 23792
rect 0 23400 160 23520
rect 0 23128 160 23248
rect 0 22856 160 22976
rect 0 22584 160 22704
rect 0 22312 160 22432
rect 0 22040 160 22160
rect 0 21768 160 21888
rect 0 21496 160 21616
rect 0 21224 160 21344
rect 0 20952 160 21072
rect 0 20680 160 20800
rect 0 20408 160 20528
rect 0 20136 160 20256
rect 0 19864 160 19984
rect 0 19592 160 19712
rect 0 19320 160 19440
rect 0 19048 160 19168
rect 0 18776 160 18896
rect 0 18504 160 18624
rect 0 18232 160 18352
rect 0 17960 160 18080
rect 0 17688 160 17808
rect 0 17416 160 17536
rect 0 17144 160 17264
rect 0 16872 160 16992
rect 0 16600 160 16720
rect 0 16328 160 16448
rect 0 16056 160 16176
rect 0 15784 160 15904
rect 0 15512 160 15632
rect 0 15240 160 15360
rect 0 14968 160 15088
rect 0 14696 160 14816
rect 0 14424 160 14544
rect 0 14152 160 14272
rect 0 13880 160 14000
rect 0 13608 160 13728
rect 0 13336 160 13456
rect 0 13064 160 13184
rect 0 12792 160 12912
rect 0 12520 160 12640
rect 0 12248 160 12368
rect 0 11976 160 12096
rect 0 11704 160 11824
rect 0 11432 160 11552
rect 0 11160 160 11280
rect 0 10888 160 11008
rect 0 10616 160 10736
rect 0 10344 160 10464
rect 0 10072 160 10192
rect 0 9800 160 9920
rect 0 9528 160 9648
rect 0 9256 160 9376
rect 0 8984 160 9104
rect 0 8712 160 8832
rect 0 8440 160 8560
rect 0 8168 160 8288
rect 0 7896 160 8016
rect 0 7624 160 7744
rect 0 7352 160 7472
rect 0 7080 160 7200
rect 0 6808 160 6928
rect 0 6536 160 6656
rect 0 6264 160 6384
rect 0 5992 160 6112
rect 0 5720 160 5840
rect 0 5448 160 5568
rect 0 5176 160 5296
rect 47840 39720 48000 39840
rect 47840 39448 48000 39568
rect 47840 39176 48000 39296
rect 47840 38904 48000 39024
rect 47840 38632 48000 38752
rect 47840 38360 48000 38480
rect 47840 38088 48000 38208
rect 47840 37816 48000 37936
rect 47840 37544 48000 37664
rect 47840 37272 48000 37392
rect 47840 37000 48000 37120
rect 47840 36728 48000 36848
rect 47840 36456 48000 36576
rect 47840 36184 48000 36304
rect 47840 35912 48000 36032
rect 47840 35640 48000 35760
rect 47840 35368 48000 35488
rect 47840 35096 48000 35216
rect 47840 34824 48000 34944
rect 47840 34552 48000 34672
rect 47840 34280 48000 34400
rect 47840 34008 48000 34128
rect 47840 33736 48000 33856
rect 47840 33464 48000 33584
rect 47840 33192 48000 33312
rect 47840 32920 48000 33040
rect 47840 32648 48000 32768
rect 47840 32376 48000 32496
rect 47840 32104 48000 32224
rect 47840 31832 48000 31952
rect 47840 31560 48000 31680
rect 47840 31288 48000 31408
rect 47840 31016 48000 31136
rect 47840 30744 48000 30864
rect 47840 30472 48000 30592
rect 47840 30200 48000 30320
rect 47840 29928 48000 30048
rect 47840 29656 48000 29776
rect 47840 29384 48000 29504
rect 47840 29112 48000 29232
rect 47840 28840 48000 28960
rect 47840 28568 48000 28688
rect 47840 28296 48000 28416
rect 47840 28024 48000 28144
rect 47840 27752 48000 27872
rect 47840 27480 48000 27600
rect 47840 27208 48000 27328
rect 47840 26936 48000 27056
rect 47840 26664 48000 26784
rect 47840 26392 48000 26512
rect 47840 26120 48000 26240
rect 47840 25848 48000 25968
rect 47840 25576 48000 25696
rect 47840 25304 48000 25424
rect 47840 25032 48000 25152
rect 47840 24760 48000 24880
rect 47840 24488 48000 24608
rect 47840 24216 48000 24336
rect 47840 23944 48000 24064
rect 47840 23672 48000 23792
rect 47840 23400 48000 23520
rect 47840 23128 48000 23248
rect 47840 22856 48000 22976
rect 47840 22584 48000 22704
rect 47840 22312 48000 22432
rect 47840 22040 48000 22160
rect 47840 21768 48000 21888
rect 47840 21496 48000 21616
rect 47840 21224 48000 21344
rect 47840 20952 48000 21072
rect 47840 20680 48000 20800
rect 47840 20408 48000 20528
rect 47840 20136 48000 20256
rect 47840 19864 48000 19984
rect 47840 19592 48000 19712
rect 47840 19320 48000 19440
rect 47840 19048 48000 19168
rect 47840 18776 48000 18896
rect 47840 18504 48000 18624
rect 47840 18232 48000 18352
rect 47840 17960 48000 18080
rect 47840 17688 48000 17808
rect 47840 17416 48000 17536
rect 47840 17144 48000 17264
rect 47840 16872 48000 16992
rect 47840 16600 48000 16720
rect 47840 16328 48000 16448
rect 47840 16056 48000 16176
rect 47840 15784 48000 15904
rect 47840 15512 48000 15632
rect 47840 15240 48000 15360
rect 47840 14968 48000 15088
rect 47840 14696 48000 14816
rect 47840 14424 48000 14544
rect 47840 14152 48000 14272
rect 47840 13880 48000 14000
rect 47840 13608 48000 13728
rect 47840 13336 48000 13456
rect 47840 13064 48000 13184
rect 47840 12792 48000 12912
rect 47840 12520 48000 12640
rect 47840 12248 48000 12368
rect 47840 11976 48000 12096
rect 47840 11704 48000 11824
rect 47840 11432 48000 11552
rect 47840 11160 48000 11280
rect 47840 10888 48000 11008
rect 47840 10616 48000 10736
rect 47840 10344 48000 10464
rect 47840 10072 48000 10192
rect 47840 9800 48000 9920
rect 47840 9528 48000 9648
rect 47840 9256 48000 9376
rect 47840 8984 48000 9104
rect 47840 8712 48000 8832
rect 47840 8440 48000 8560
rect 47840 8168 48000 8288
rect 47840 7896 48000 8016
rect 47840 7624 48000 7744
rect 47840 7352 48000 7472
rect 47840 7080 48000 7200
rect 47840 6808 48000 6928
rect 47840 6536 48000 6656
rect 47840 6264 48000 6384
rect 47840 5992 48000 6112
rect 47840 5720 48000 5840
rect 47840 5448 48000 5568
rect 47840 5176 48000 5296
<< obsm3 >>
rect 160 39920 47840 43553
rect 240 5096 47760 39920
rect 160 851 47840 5096
<< metal4 >>
rect 4208 1040 4528 43568
rect 19568 1040 19888 43568
rect 34928 1040 35248 43568
<< obsm4 >>
rect 427 960 4128 43349
rect 4608 960 19488 43349
rect 19968 960 34848 43349
rect 35328 960 45389 43349
rect 427 851 45389 960
<< labels >>
rlabel metal3 s 47840 18232 48000 18352 6 E1BEG[0]
port 1 nsew signal output
rlabel metal3 s 47840 18504 48000 18624 6 E1BEG[1]
port 2 nsew signal output
rlabel metal3 s 47840 18776 48000 18896 6 E1BEG[2]
port 3 nsew signal output
rlabel metal3 s 47840 19048 48000 19168 6 E1BEG[3]
port 4 nsew signal output
rlabel metal3 s 0 18232 160 18352 6 E1END[0]
port 5 nsew signal input
rlabel metal3 s 0 18504 160 18624 6 E1END[1]
port 6 nsew signal input
rlabel metal3 s 0 18776 160 18896 6 E1END[2]
port 7 nsew signal input
rlabel metal3 s 0 19048 160 19168 6 E1END[3]
port 8 nsew signal input
rlabel metal3 s 47840 19320 48000 19440 6 E2BEG[0]
port 9 nsew signal output
rlabel metal3 s 47840 19592 48000 19712 6 E2BEG[1]
port 10 nsew signal output
rlabel metal3 s 47840 19864 48000 19984 6 E2BEG[2]
port 11 nsew signal output
rlabel metal3 s 47840 20136 48000 20256 6 E2BEG[3]
port 12 nsew signal output
rlabel metal3 s 47840 20408 48000 20528 6 E2BEG[4]
port 13 nsew signal output
rlabel metal3 s 47840 20680 48000 20800 6 E2BEG[5]
port 14 nsew signal output
rlabel metal3 s 47840 20952 48000 21072 6 E2BEG[6]
port 15 nsew signal output
rlabel metal3 s 47840 21224 48000 21344 6 E2BEG[7]
port 16 nsew signal output
rlabel metal3 s 47840 21496 48000 21616 6 E2BEGb[0]
port 17 nsew signal output
rlabel metal3 s 47840 21768 48000 21888 6 E2BEGb[1]
port 18 nsew signal output
rlabel metal3 s 47840 22040 48000 22160 6 E2BEGb[2]
port 19 nsew signal output
rlabel metal3 s 47840 22312 48000 22432 6 E2BEGb[3]
port 20 nsew signal output
rlabel metal3 s 47840 22584 48000 22704 6 E2BEGb[4]
port 21 nsew signal output
rlabel metal3 s 47840 22856 48000 22976 6 E2BEGb[5]
port 22 nsew signal output
rlabel metal3 s 47840 23128 48000 23248 6 E2BEGb[6]
port 23 nsew signal output
rlabel metal3 s 47840 23400 48000 23520 6 E2BEGb[7]
port 24 nsew signal output
rlabel metal3 s 0 21496 160 21616 6 E2END[0]
port 25 nsew signal input
rlabel metal3 s 0 21768 160 21888 6 E2END[1]
port 26 nsew signal input
rlabel metal3 s 0 22040 160 22160 6 E2END[2]
port 27 nsew signal input
rlabel metal3 s 0 22312 160 22432 6 E2END[3]
port 28 nsew signal input
rlabel metal3 s 0 22584 160 22704 6 E2END[4]
port 29 nsew signal input
rlabel metal3 s 0 22856 160 22976 6 E2END[5]
port 30 nsew signal input
rlabel metal3 s 0 23128 160 23248 6 E2END[6]
port 31 nsew signal input
rlabel metal3 s 0 23400 160 23520 6 E2END[7]
port 32 nsew signal input
rlabel metal3 s 0 19320 160 19440 6 E2MID[0]
port 33 nsew signal input
rlabel metal3 s 0 19592 160 19712 6 E2MID[1]
port 34 nsew signal input
rlabel metal3 s 0 19864 160 19984 6 E2MID[2]
port 35 nsew signal input
rlabel metal3 s 0 20136 160 20256 6 E2MID[3]
port 36 nsew signal input
rlabel metal3 s 0 20408 160 20528 6 E2MID[4]
port 37 nsew signal input
rlabel metal3 s 0 20680 160 20800 6 E2MID[5]
port 38 nsew signal input
rlabel metal3 s 0 20952 160 21072 6 E2MID[6]
port 39 nsew signal input
rlabel metal3 s 0 21224 160 21344 6 E2MID[7]
port 40 nsew signal input
rlabel metal3 s 47840 28024 48000 28144 6 E6BEG[0]
port 41 nsew signal output
rlabel metal3 s 47840 30744 48000 30864 6 E6BEG[10]
port 42 nsew signal output
rlabel metal3 s 47840 31016 48000 31136 6 E6BEG[11]
port 43 nsew signal output
rlabel metal3 s 47840 28296 48000 28416 6 E6BEG[1]
port 44 nsew signal output
rlabel metal3 s 47840 28568 48000 28688 6 E6BEG[2]
port 45 nsew signal output
rlabel metal3 s 47840 28840 48000 28960 6 E6BEG[3]
port 46 nsew signal output
rlabel metal3 s 47840 29112 48000 29232 6 E6BEG[4]
port 47 nsew signal output
rlabel metal3 s 47840 29384 48000 29504 6 E6BEG[5]
port 48 nsew signal output
rlabel metal3 s 47840 29656 48000 29776 6 E6BEG[6]
port 49 nsew signal output
rlabel metal3 s 47840 29928 48000 30048 6 E6BEG[7]
port 50 nsew signal output
rlabel metal3 s 47840 30200 48000 30320 6 E6BEG[8]
port 51 nsew signal output
rlabel metal3 s 47840 30472 48000 30592 6 E6BEG[9]
port 52 nsew signal output
rlabel metal3 s 0 28024 160 28144 6 E6END[0]
port 53 nsew signal input
rlabel metal3 s 0 30744 160 30864 6 E6END[10]
port 54 nsew signal input
rlabel metal3 s 0 31016 160 31136 6 E6END[11]
port 55 nsew signal input
rlabel metal3 s 0 28296 160 28416 6 E6END[1]
port 56 nsew signal input
rlabel metal3 s 0 28568 160 28688 6 E6END[2]
port 57 nsew signal input
rlabel metal3 s 0 28840 160 28960 6 E6END[3]
port 58 nsew signal input
rlabel metal3 s 0 29112 160 29232 6 E6END[4]
port 59 nsew signal input
rlabel metal3 s 0 29384 160 29504 6 E6END[5]
port 60 nsew signal input
rlabel metal3 s 0 29656 160 29776 6 E6END[6]
port 61 nsew signal input
rlabel metal3 s 0 29928 160 30048 6 E6END[7]
port 62 nsew signal input
rlabel metal3 s 0 30200 160 30320 6 E6END[8]
port 63 nsew signal input
rlabel metal3 s 0 30472 160 30592 6 E6END[9]
port 64 nsew signal input
rlabel metal3 s 47840 23672 48000 23792 6 EE4BEG[0]
port 65 nsew signal output
rlabel metal3 s 47840 26392 48000 26512 6 EE4BEG[10]
port 66 nsew signal output
rlabel metal3 s 47840 26664 48000 26784 6 EE4BEG[11]
port 67 nsew signal output
rlabel metal3 s 47840 26936 48000 27056 6 EE4BEG[12]
port 68 nsew signal output
rlabel metal3 s 47840 27208 48000 27328 6 EE4BEG[13]
port 69 nsew signal output
rlabel metal3 s 47840 27480 48000 27600 6 EE4BEG[14]
port 70 nsew signal output
rlabel metal3 s 47840 27752 48000 27872 6 EE4BEG[15]
port 71 nsew signal output
rlabel metal3 s 47840 23944 48000 24064 6 EE4BEG[1]
port 72 nsew signal output
rlabel metal3 s 47840 24216 48000 24336 6 EE4BEG[2]
port 73 nsew signal output
rlabel metal3 s 47840 24488 48000 24608 6 EE4BEG[3]
port 74 nsew signal output
rlabel metal3 s 47840 24760 48000 24880 6 EE4BEG[4]
port 75 nsew signal output
rlabel metal3 s 47840 25032 48000 25152 6 EE4BEG[5]
port 76 nsew signal output
rlabel metal3 s 47840 25304 48000 25424 6 EE4BEG[6]
port 77 nsew signal output
rlabel metal3 s 47840 25576 48000 25696 6 EE4BEG[7]
port 78 nsew signal output
rlabel metal3 s 47840 25848 48000 25968 6 EE4BEG[8]
port 79 nsew signal output
rlabel metal3 s 47840 26120 48000 26240 6 EE4BEG[9]
port 80 nsew signal output
rlabel metal3 s 0 23672 160 23792 6 EE4END[0]
port 81 nsew signal input
rlabel metal3 s 0 26392 160 26512 6 EE4END[10]
port 82 nsew signal input
rlabel metal3 s 0 26664 160 26784 6 EE4END[11]
port 83 nsew signal input
rlabel metal3 s 0 26936 160 27056 6 EE4END[12]
port 84 nsew signal input
rlabel metal3 s 0 27208 160 27328 6 EE4END[13]
port 85 nsew signal input
rlabel metal3 s 0 27480 160 27600 6 EE4END[14]
port 86 nsew signal input
rlabel metal3 s 0 27752 160 27872 6 EE4END[15]
port 87 nsew signal input
rlabel metal3 s 0 23944 160 24064 6 EE4END[1]
port 88 nsew signal input
rlabel metal3 s 0 24216 160 24336 6 EE4END[2]
port 89 nsew signal input
rlabel metal3 s 0 24488 160 24608 6 EE4END[3]
port 90 nsew signal input
rlabel metal3 s 0 24760 160 24880 6 EE4END[4]
port 91 nsew signal input
rlabel metal3 s 0 25032 160 25152 6 EE4END[5]
port 92 nsew signal input
rlabel metal3 s 0 25304 160 25424 6 EE4END[6]
port 93 nsew signal input
rlabel metal3 s 0 25576 160 25696 6 EE4END[7]
port 94 nsew signal input
rlabel metal3 s 0 25848 160 25968 6 EE4END[8]
port 95 nsew signal input
rlabel metal3 s 0 26120 160 26240 6 EE4END[9]
port 96 nsew signal input
rlabel metal3 s 0 31288 160 31408 6 FrameData[0]
port 97 nsew signal input
rlabel metal3 s 0 34008 160 34128 6 FrameData[10]
port 98 nsew signal input
rlabel metal3 s 0 34280 160 34400 6 FrameData[11]
port 99 nsew signal input
rlabel metal3 s 0 34552 160 34672 6 FrameData[12]
port 100 nsew signal input
rlabel metal3 s 0 34824 160 34944 6 FrameData[13]
port 101 nsew signal input
rlabel metal3 s 0 35096 160 35216 6 FrameData[14]
port 102 nsew signal input
rlabel metal3 s 0 35368 160 35488 6 FrameData[15]
port 103 nsew signal input
rlabel metal3 s 0 35640 160 35760 6 FrameData[16]
port 104 nsew signal input
rlabel metal3 s 0 35912 160 36032 6 FrameData[17]
port 105 nsew signal input
rlabel metal3 s 0 36184 160 36304 6 FrameData[18]
port 106 nsew signal input
rlabel metal3 s 0 36456 160 36576 6 FrameData[19]
port 107 nsew signal input
rlabel metal3 s 0 31560 160 31680 6 FrameData[1]
port 108 nsew signal input
rlabel metal3 s 0 36728 160 36848 6 FrameData[20]
port 109 nsew signal input
rlabel metal3 s 0 37000 160 37120 6 FrameData[21]
port 110 nsew signal input
rlabel metal3 s 0 37272 160 37392 6 FrameData[22]
port 111 nsew signal input
rlabel metal3 s 0 37544 160 37664 6 FrameData[23]
port 112 nsew signal input
rlabel metal3 s 0 37816 160 37936 6 FrameData[24]
port 113 nsew signal input
rlabel metal3 s 0 38088 160 38208 6 FrameData[25]
port 114 nsew signal input
rlabel metal3 s 0 38360 160 38480 6 FrameData[26]
port 115 nsew signal input
rlabel metal3 s 0 38632 160 38752 6 FrameData[27]
port 116 nsew signal input
rlabel metal3 s 0 38904 160 39024 6 FrameData[28]
port 117 nsew signal input
rlabel metal3 s 0 39176 160 39296 6 FrameData[29]
port 118 nsew signal input
rlabel metal3 s 0 31832 160 31952 6 FrameData[2]
port 119 nsew signal input
rlabel metal3 s 0 39448 160 39568 6 FrameData[30]
port 120 nsew signal input
rlabel metal3 s 0 39720 160 39840 6 FrameData[31]
port 121 nsew signal input
rlabel metal3 s 0 32104 160 32224 6 FrameData[3]
port 122 nsew signal input
rlabel metal3 s 0 32376 160 32496 6 FrameData[4]
port 123 nsew signal input
rlabel metal3 s 0 32648 160 32768 6 FrameData[5]
port 124 nsew signal input
rlabel metal3 s 0 32920 160 33040 6 FrameData[6]
port 125 nsew signal input
rlabel metal3 s 0 33192 160 33312 6 FrameData[7]
port 126 nsew signal input
rlabel metal3 s 0 33464 160 33584 6 FrameData[8]
port 127 nsew signal input
rlabel metal3 s 0 33736 160 33856 6 FrameData[9]
port 128 nsew signal input
rlabel metal3 s 47840 31288 48000 31408 6 FrameData_O[0]
port 129 nsew signal output
rlabel metal3 s 47840 34008 48000 34128 6 FrameData_O[10]
port 130 nsew signal output
rlabel metal3 s 47840 34280 48000 34400 6 FrameData_O[11]
port 131 nsew signal output
rlabel metal3 s 47840 34552 48000 34672 6 FrameData_O[12]
port 132 nsew signal output
rlabel metal3 s 47840 34824 48000 34944 6 FrameData_O[13]
port 133 nsew signal output
rlabel metal3 s 47840 35096 48000 35216 6 FrameData_O[14]
port 134 nsew signal output
rlabel metal3 s 47840 35368 48000 35488 6 FrameData_O[15]
port 135 nsew signal output
rlabel metal3 s 47840 35640 48000 35760 6 FrameData_O[16]
port 136 nsew signal output
rlabel metal3 s 47840 35912 48000 36032 6 FrameData_O[17]
port 137 nsew signal output
rlabel metal3 s 47840 36184 48000 36304 6 FrameData_O[18]
port 138 nsew signal output
rlabel metal3 s 47840 36456 48000 36576 6 FrameData_O[19]
port 139 nsew signal output
rlabel metal3 s 47840 31560 48000 31680 6 FrameData_O[1]
port 140 nsew signal output
rlabel metal3 s 47840 36728 48000 36848 6 FrameData_O[20]
port 141 nsew signal output
rlabel metal3 s 47840 37000 48000 37120 6 FrameData_O[21]
port 142 nsew signal output
rlabel metal3 s 47840 37272 48000 37392 6 FrameData_O[22]
port 143 nsew signal output
rlabel metal3 s 47840 37544 48000 37664 6 FrameData_O[23]
port 144 nsew signal output
rlabel metal3 s 47840 37816 48000 37936 6 FrameData_O[24]
port 145 nsew signal output
rlabel metal3 s 47840 38088 48000 38208 6 FrameData_O[25]
port 146 nsew signal output
rlabel metal3 s 47840 38360 48000 38480 6 FrameData_O[26]
port 147 nsew signal output
rlabel metal3 s 47840 38632 48000 38752 6 FrameData_O[27]
port 148 nsew signal output
rlabel metal3 s 47840 38904 48000 39024 6 FrameData_O[28]
port 149 nsew signal output
rlabel metal3 s 47840 39176 48000 39296 6 FrameData_O[29]
port 150 nsew signal output
rlabel metal3 s 47840 31832 48000 31952 6 FrameData_O[2]
port 151 nsew signal output
rlabel metal3 s 47840 39448 48000 39568 6 FrameData_O[30]
port 152 nsew signal output
rlabel metal3 s 47840 39720 48000 39840 6 FrameData_O[31]
port 153 nsew signal output
rlabel metal3 s 47840 32104 48000 32224 6 FrameData_O[3]
port 154 nsew signal output
rlabel metal3 s 47840 32376 48000 32496 6 FrameData_O[4]
port 155 nsew signal output
rlabel metal3 s 47840 32648 48000 32768 6 FrameData_O[5]
port 156 nsew signal output
rlabel metal3 s 47840 32920 48000 33040 6 FrameData_O[6]
port 157 nsew signal output
rlabel metal3 s 47840 33192 48000 33312 6 FrameData_O[7]
port 158 nsew signal output
rlabel metal3 s 47840 33464 48000 33584 6 FrameData_O[8]
port 159 nsew signal output
rlabel metal3 s 47840 33736 48000 33856 6 FrameData_O[9]
port 160 nsew signal output
rlabel metal2 s 39762 0 39818 160 6 FrameStrobe[0]
port 161 nsew signal input
rlabel metal2 s 43442 0 43498 160 6 FrameStrobe[10]
port 162 nsew signal input
rlabel metal2 s 43810 0 43866 160 6 FrameStrobe[11]
port 163 nsew signal input
rlabel metal2 s 44178 0 44234 160 6 FrameStrobe[12]
port 164 nsew signal input
rlabel metal2 s 44546 0 44602 160 6 FrameStrobe[13]
port 165 nsew signal input
rlabel metal2 s 44914 0 44970 160 6 FrameStrobe[14]
port 166 nsew signal input
rlabel metal2 s 45282 0 45338 160 6 FrameStrobe[15]
port 167 nsew signal input
rlabel metal2 s 45650 0 45706 160 6 FrameStrobe[16]
port 168 nsew signal input
rlabel metal2 s 46018 0 46074 160 6 FrameStrobe[17]
port 169 nsew signal input
rlabel metal2 s 46386 0 46442 160 6 FrameStrobe[18]
port 170 nsew signal input
rlabel metal2 s 46754 0 46810 160 6 FrameStrobe[19]
port 171 nsew signal input
rlabel metal2 s 40130 0 40186 160 6 FrameStrobe[1]
port 172 nsew signal input
rlabel metal2 s 40498 0 40554 160 6 FrameStrobe[2]
port 173 nsew signal input
rlabel metal2 s 40866 0 40922 160 6 FrameStrobe[3]
port 174 nsew signal input
rlabel metal2 s 41234 0 41290 160 6 FrameStrobe[4]
port 175 nsew signal input
rlabel metal2 s 41602 0 41658 160 6 FrameStrobe[5]
port 176 nsew signal input
rlabel metal2 s 41970 0 42026 160 6 FrameStrobe[6]
port 177 nsew signal input
rlabel metal2 s 42338 0 42394 160 6 FrameStrobe[7]
port 178 nsew signal input
rlabel metal2 s 42706 0 42762 160 6 FrameStrobe[8]
port 179 nsew signal input
rlabel metal2 s 43074 0 43130 160 6 FrameStrobe[9]
port 180 nsew signal input
rlabel metal2 s 39762 44840 39818 45000 6 FrameStrobe_O[0]
port 181 nsew signal output
rlabel metal2 s 43442 44840 43498 45000 6 FrameStrobe_O[10]
port 182 nsew signal output
rlabel metal2 s 43810 44840 43866 45000 6 FrameStrobe_O[11]
port 183 nsew signal output
rlabel metal2 s 44178 44840 44234 45000 6 FrameStrobe_O[12]
port 184 nsew signal output
rlabel metal2 s 44546 44840 44602 45000 6 FrameStrobe_O[13]
port 185 nsew signal output
rlabel metal2 s 44914 44840 44970 45000 6 FrameStrobe_O[14]
port 186 nsew signal output
rlabel metal2 s 45282 44840 45338 45000 6 FrameStrobe_O[15]
port 187 nsew signal output
rlabel metal2 s 45650 44840 45706 45000 6 FrameStrobe_O[16]
port 188 nsew signal output
rlabel metal2 s 46018 44840 46074 45000 6 FrameStrobe_O[17]
port 189 nsew signal output
rlabel metal2 s 46386 44840 46442 45000 6 FrameStrobe_O[18]
port 190 nsew signal output
rlabel metal2 s 46754 44840 46810 45000 6 FrameStrobe_O[19]
port 191 nsew signal output
rlabel metal2 s 40130 44840 40186 45000 6 FrameStrobe_O[1]
port 192 nsew signal output
rlabel metal2 s 40498 44840 40554 45000 6 FrameStrobe_O[2]
port 193 nsew signal output
rlabel metal2 s 40866 44840 40922 45000 6 FrameStrobe_O[3]
port 194 nsew signal output
rlabel metal2 s 41234 44840 41290 45000 6 FrameStrobe_O[4]
port 195 nsew signal output
rlabel metal2 s 41602 44840 41658 45000 6 FrameStrobe_O[5]
port 196 nsew signal output
rlabel metal2 s 41970 44840 42026 45000 6 FrameStrobe_O[6]
port 197 nsew signal output
rlabel metal2 s 42338 44840 42394 45000 6 FrameStrobe_O[7]
port 198 nsew signal output
rlabel metal2 s 42706 44840 42762 45000 6 FrameStrobe_O[8]
port 199 nsew signal output
rlabel metal2 s 43074 44840 43130 45000 6 FrameStrobe_O[9]
port 200 nsew signal output
rlabel metal2 s 1122 44840 1178 45000 6 N1BEG[0]
port 201 nsew signal output
rlabel metal2 s 1490 44840 1546 45000 6 N1BEG[1]
port 202 nsew signal output
rlabel metal2 s 1858 44840 1914 45000 6 N1BEG[2]
port 203 nsew signal output
rlabel metal2 s 2226 44840 2282 45000 6 N1BEG[3]
port 204 nsew signal output
rlabel metal2 s 1122 0 1178 160 6 N1END[0]
port 205 nsew signal input
rlabel metal2 s 1490 0 1546 160 6 N1END[1]
port 206 nsew signal input
rlabel metal2 s 1858 0 1914 160 6 N1END[2]
port 207 nsew signal input
rlabel metal2 s 2226 0 2282 160 6 N1END[3]
port 208 nsew signal input
rlabel metal2 s 2594 44840 2650 45000 6 N2BEG[0]
port 209 nsew signal output
rlabel metal2 s 2962 44840 3018 45000 6 N2BEG[1]
port 210 nsew signal output
rlabel metal2 s 3330 44840 3386 45000 6 N2BEG[2]
port 211 nsew signal output
rlabel metal2 s 3698 44840 3754 45000 6 N2BEG[3]
port 212 nsew signal output
rlabel metal2 s 4066 44840 4122 45000 6 N2BEG[4]
port 213 nsew signal output
rlabel metal2 s 4434 44840 4490 45000 6 N2BEG[5]
port 214 nsew signal output
rlabel metal2 s 4802 44840 4858 45000 6 N2BEG[6]
port 215 nsew signal output
rlabel metal2 s 5170 44840 5226 45000 6 N2BEG[7]
port 216 nsew signal output
rlabel metal2 s 5538 44840 5594 45000 6 N2BEGb[0]
port 217 nsew signal output
rlabel metal2 s 5906 44840 5962 45000 6 N2BEGb[1]
port 218 nsew signal output
rlabel metal2 s 6274 44840 6330 45000 6 N2BEGb[2]
port 219 nsew signal output
rlabel metal2 s 6642 44840 6698 45000 6 N2BEGb[3]
port 220 nsew signal output
rlabel metal2 s 7010 44840 7066 45000 6 N2BEGb[4]
port 221 nsew signal output
rlabel metal2 s 7378 44840 7434 45000 6 N2BEGb[5]
port 222 nsew signal output
rlabel metal2 s 7746 44840 7802 45000 6 N2BEGb[6]
port 223 nsew signal output
rlabel metal2 s 8114 44840 8170 45000 6 N2BEGb[7]
port 224 nsew signal output
rlabel metal2 s 5538 0 5594 160 6 N2END[0]
port 225 nsew signal input
rlabel metal2 s 5906 0 5962 160 6 N2END[1]
port 226 nsew signal input
rlabel metal2 s 6274 0 6330 160 6 N2END[2]
port 227 nsew signal input
rlabel metal2 s 6642 0 6698 160 6 N2END[3]
port 228 nsew signal input
rlabel metal2 s 7010 0 7066 160 6 N2END[4]
port 229 nsew signal input
rlabel metal2 s 7378 0 7434 160 6 N2END[5]
port 230 nsew signal input
rlabel metal2 s 7746 0 7802 160 6 N2END[6]
port 231 nsew signal input
rlabel metal2 s 8114 0 8170 160 6 N2END[7]
port 232 nsew signal input
rlabel metal2 s 2594 0 2650 160 6 N2MID[0]
port 233 nsew signal input
rlabel metal2 s 2962 0 3018 160 6 N2MID[1]
port 234 nsew signal input
rlabel metal2 s 3330 0 3386 160 6 N2MID[2]
port 235 nsew signal input
rlabel metal2 s 3698 0 3754 160 6 N2MID[3]
port 236 nsew signal input
rlabel metal2 s 4066 0 4122 160 6 N2MID[4]
port 237 nsew signal input
rlabel metal2 s 4434 0 4490 160 6 N2MID[5]
port 238 nsew signal input
rlabel metal2 s 4802 0 4858 160 6 N2MID[6]
port 239 nsew signal input
rlabel metal2 s 5170 0 5226 160 6 N2MID[7]
port 240 nsew signal input
rlabel metal2 s 8482 44840 8538 45000 6 N4BEG[0]
port 241 nsew signal output
rlabel metal2 s 12162 44840 12218 45000 6 N4BEG[10]
port 242 nsew signal output
rlabel metal2 s 12530 44840 12586 45000 6 N4BEG[11]
port 243 nsew signal output
rlabel metal2 s 12898 44840 12954 45000 6 N4BEG[12]
port 244 nsew signal output
rlabel metal2 s 13266 44840 13322 45000 6 N4BEG[13]
port 245 nsew signal output
rlabel metal2 s 13634 44840 13690 45000 6 N4BEG[14]
port 246 nsew signal output
rlabel metal2 s 14002 44840 14058 45000 6 N4BEG[15]
port 247 nsew signal output
rlabel metal2 s 8850 44840 8906 45000 6 N4BEG[1]
port 248 nsew signal output
rlabel metal2 s 9218 44840 9274 45000 6 N4BEG[2]
port 249 nsew signal output
rlabel metal2 s 9586 44840 9642 45000 6 N4BEG[3]
port 250 nsew signal output
rlabel metal2 s 9954 44840 10010 45000 6 N4BEG[4]
port 251 nsew signal output
rlabel metal2 s 10322 44840 10378 45000 6 N4BEG[5]
port 252 nsew signal output
rlabel metal2 s 10690 44840 10746 45000 6 N4BEG[6]
port 253 nsew signal output
rlabel metal2 s 11058 44840 11114 45000 6 N4BEG[7]
port 254 nsew signal output
rlabel metal2 s 11426 44840 11482 45000 6 N4BEG[8]
port 255 nsew signal output
rlabel metal2 s 11794 44840 11850 45000 6 N4BEG[9]
port 256 nsew signal output
rlabel metal2 s 8482 0 8538 160 6 N4END[0]
port 257 nsew signal input
rlabel metal2 s 12162 0 12218 160 6 N4END[10]
port 258 nsew signal input
rlabel metal2 s 12530 0 12586 160 6 N4END[11]
port 259 nsew signal input
rlabel metal2 s 12898 0 12954 160 6 N4END[12]
port 260 nsew signal input
rlabel metal2 s 13266 0 13322 160 6 N4END[13]
port 261 nsew signal input
rlabel metal2 s 13634 0 13690 160 6 N4END[14]
port 262 nsew signal input
rlabel metal2 s 14002 0 14058 160 6 N4END[15]
port 263 nsew signal input
rlabel metal2 s 8850 0 8906 160 6 N4END[1]
port 264 nsew signal input
rlabel metal2 s 9218 0 9274 160 6 N4END[2]
port 265 nsew signal input
rlabel metal2 s 9586 0 9642 160 6 N4END[3]
port 266 nsew signal input
rlabel metal2 s 9954 0 10010 160 6 N4END[4]
port 267 nsew signal input
rlabel metal2 s 10322 0 10378 160 6 N4END[5]
port 268 nsew signal input
rlabel metal2 s 10690 0 10746 160 6 N4END[6]
port 269 nsew signal input
rlabel metal2 s 11058 0 11114 160 6 N4END[7]
port 270 nsew signal input
rlabel metal2 s 11426 0 11482 160 6 N4END[8]
port 271 nsew signal input
rlabel metal2 s 11794 0 11850 160 6 N4END[9]
port 272 nsew signal input
rlabel metal2 s 14370 44840 14426 45000 6 NN4BEG[0]
port 273 nsew signal output
rlabel metal2 s 18050 44840 18106 45000 6 NN4BEG[10]
port 274 nsew signal output
rlabel metal2 s 18418 44840 18474 45000 6 NN4BEG[11]
port 275 nsew signal output
rlabel metal2 s 18786 44840 18842 45000 6 NN4BEG[12]
port 276 nsew signal output
rlabel metal2 s 19154 44840 19210 45000 6 NN4BEG[13]
port 277 nsew signal output
rlabel metal2 s 19522 44840 19578 45000 6 NN4BEG[14]
port 278 nsew signal output
rlabel metal2 s 19890 44840 19946 45000 6 NN4BEG[15]
port 279 nsew signal output
rlabel metal2 s 14738 44840 14794 45000 6 NN4BEG[1]
port 280 nsew signal output
rlabel metal2 s 15106 44840 15162 45000 6 NN4BEG[2]
port 281 nsew signal output
rlabel metal2 s 15474 44840 15530 45000 6 NN4BEG[3]
port 282 nsew signal output
rlabel metal2 s 15842 44840 15898 45000 6 NN4BEG[4]
port 283 nsew signal output
rlabel metal2 s 16210 44840 16266 45000 6 NN4BEG[5]
port 284 nsew signal output
rlabel metal2 s 16578 44840 16634 45000 6 NN4BEG[6]
port 285 nsew signal output
rlabel metal2 s 16946 44840 17002 45000 6 NN4BEG[7]
port 286 nsew signal output
rlabel metal2 s 17314 44840 17370 45000 6 NN4BEG[8]
port 287 nsew signal output
rlabel metal2 s 17682 44840 17738 45000 6 NN4BEG[9]
port 288 nsew signal output
rlabel metal2 s 14370 0 14426 160 6 NN4END[0]
port 289 nsew signal input
rlabel metal2 s 18050 0 18106 160 6 NN4END[10]
port 290 nsew signal input
rlabel metal2 s 18418 0 18474 160 6 NN4END[11]
port 291 nsew signal input
rlabel metal2 s 18786 0 18842 160 6 NN4END[12]
port 292 nsew signal input
rlabel metal2 s 19154 0 19210 160 6 NN4END[13]
port 293 nsew signal input
rlabel metal2 s 19522 0 19578 160 6 NN4END[14]
port 294 nsew signal input
rlabel metal2 s 19890 0 19946 160 6 NN4END[15]
port 295 nsew signal input
rlabel metal2 s 14738 0 14794 160 6 NN4END[1]
port 296 nsew signal input
rlabel metal2 s 15106 0 15162 160 6 NN4END[2]
port 297 nsew signal input
rlabel metal2 s 15474 0 15530 160 6 NN4END[3]
port 298 nsew signal input
rlabel metal2 s 15842 0 15898 160 6 NN4END[4]
port 299 nsew signal input
rlabel metal2 s 16210 0 16266 160 6 NN4END[5]
port 300 nsew signal input
rlabel metal2 s 16578 0 16634 160 6 NN4END[6]
port 301 nsew signal input
rlabel metal2 s 16946 0 17002 160 6 NN4END[7]
port 302 nsew signal input
rlabel metal2 s 17314 0 17370 160 6 NN4END[8]
port 303 nsew signal input
rlabel metal2 s 17682 0 17738 160 6 NN4END[9]
port 304 nsew signal input
rlabel metal2 s 20258 0 20314 160 6 S1BEG[0]
port 305 nsew signal output
rlabel metal2 s 20626 0 20682 160 6 S1BEG[1]
port 306 nsew signal output
rlabel metal2 s 20994 0 21050 160 6 S1BEG[2]
port 307 nsew signal output
rlabel metal2 s 21362 0 21418 160 6 S1BEG[3]
port 308 nsew signal output
rlabel metal2 s 20258 44840 20314 45000 6 S1END[0]
port 309 nsew signal input
rlabel metal2 s 20626 44840 20682 45000 6 S1END[1]
port 310 nsew signal input
rlabel metal2 s 20994 44840 21050 45000 6 S1END[2]
port 311 nsew signal input
rlabel metal2 s 21362 44840 21418 45000 6 S1END[3]
port 312 nsew signal input
rlabel metal2 s 24674 0 24730 160 6 S2BEG[0]
port 313 nsew signal output
rlabel metal2 s 25042 0 25098 160 6 S2BEG[1]
port 314 nsew signal output
rlabel metal2 s 25410 0 25466 160 6 S2BEG[2]
port 315 nsew signal output
rlabel metal2 s 25778 0 25834 160 6 S2BEG[3]
port 316 nsew signal output
rlabel metal2 s 26146 0 26202 160 6 S2BEG[4]
port 317 nsew signal output
rlabel metal2 s 26514 0 26570 160 6 S2BEG[5]
port 318 nsew signal output
rlabel metal2 s 26882 0 26938 160 6 S2BEG[6]
port 319 nsew signal output
rlabel metal2 s 27250 0 27306 160 6 S2BEG[7]
port 320 nsew signal output
rlabel metal2 s 21730 0 21786 160 6 S2BEGb[0]
port 321 nsew signal output
rlabel metal2 s 22098 0 22154 160 6 S2BEGb[1]
port 322 nsew signal output
rlabel metal2 s 22466 0 22522 160 6 S2BEGb[2]
port 323 nsew signal output
rlabel metal2 s 22834 0 22890 160 6 S2BEGb[3]
port 324 nsew signal output
rlabel metal2 s 23202 0 23258 160 6 S2BEGb[4]
port 325 nsew signal output
rlabel metal2 s 23570 0 23626 160 6 S2BEGb[5]
port 326 nsew signal output
rlabel metal2 s 23938 0 23994 160 6 S2BEGb[6]
port 327 nsew signal output
rlabel metal2 s 24306 0 24362 160 6 S2BEGb[7]
port 328 nsew signal output
rlabel metal2 s 21730 44840 21786 45000 6 S2END[0]
port 329 nsew signal input
rlabel metal2 s 22098 44840 22154 45000 6 S2END[1]
port 330 nsew signal input
rlabel metal2 s 22466 44840 22522 45000 6 S2END[2]
port 331 nsew signal input
rlabel metal2 s 22834 44840 22890 45000 6 S2END[3]
port 332 nsew signal input
rlabel metal2 s 23202 44840 23258 45000 6 S2END[4]
port 333 nsew signal input
rlabel metal2 s 23570 44840 23626 45000 6 S2END[5]
port 334 nsew signal input
rlabel metal2 s 23938 44840 23994 45000 6 S2END[6]
port 335 nsew signal input
rlabel metal2 s 24306 44840 24362 45000 6 S2END[7]
port 336 nsew signal input
rlabel metal2 s 24674 44840 24730 45000 6 S2MID[0]
port 337 nsew signal input
rlabel metal2 s 25042 44840 25098 45000 6 S2MID[1]
port 338 nsew signal input
rlabel metal2 s 25410 44840 25466 45000 6 S2MID[2]
port 339 nsew signal input
rlabel metal2 s 25778 44840 25834 45000 6 S2MID[3]
port 340 nsew signal input
rlabel metal2 s 26146 44840 26202 45000 6 S2MID[4]
port 341 nsew signal input
rlabel metal2 s 26514 44840 26570 45000 6 S2MID[5]
port 342 nsew signal input
rlabel metal2 s 26882 44840 26938 45000 6 S2MID[6]
port 343 nsew signal input
rlabel metal2 s 27250 44840 27306 45000 6 S2MID[7]
port 344 nsew signal input
rlabel metal2 s 27618 0 27674 160 6 S4BEG[0]
port 345 nsew signal output
rlabel metal2 s 31298 0 31354 160 6 S4BEG[10]
port 346 nsew signal output
rlabel metal2 s 31666 0 31722 160 6 S4BEG[11]
port 347 nsew signal output
rlabel metal2 s 32034 0 32090 160 6 S4BEG[12]
port 348 nsew signal output
rlabel metal2 s 32402 0 32458 160 6 S4BEG[13]
port 349 nsew signal output
rlabel metal2 s 32770 0 32826 160 6 S4BEG[14]
port 350 nsew signal output
rlabel metal2 s 33138 0 33194 160 6 S4BEG[15]
port 351 nsew signal output
rlabel metal2 s 27986 0 28042 160 6 S4BEG[1]
port 352 nsew signal output
rlabel metal2 s 28354 0 28410 160 6 S4BEG[2]
port 353 nsew signal output
rlabel metal2 s 28722 0 28778 160 6 S4BEG[3]
port 354 nsew signal output
rlabel metal2 s 29090 0 29146 160 6 S4BEG[4]
port 355 nsew signal output
rlabel metal2 s 29458 0 29514 160 6 S4BEG[5]
port 356 nsew signal output
rlabel metal2 s 29826 0 29882 160 6 S4BEG[6]
port 357 nsew signal output
rlabel metal2 s 30194 0 30250 160 6 S4BEG[7]
port 358 nsew signal output
rlabel metal2 s 30562 0 30618 160 6 S4BEG[8]
port 359 nsew signal output
rlabel metal2 s 30930 0 30986 160 6 S4BEG[9]
port 360 nsew signal output
rlabel metal2 s 27618 44840 27674 45000 6 S4END[0]
port 361 nsew signal input
rlabel metal2 s 31298 44840 31354 45000 6 S4END[10]
port 362 nsew signal input
rlabel metal2 s 31666 44840 31722 45000 6 S4END[11]
port 363 nsew signal input
rlabel metal2 s 32034 44840 32090 45000 6 S4END[12]
port 364 nsew signal input
rlabel metal2 s 32402 44840 32458 45000 6 S4END[13]
port 365 nsew signal input
rlabel metal2 s 32770 44840 32826 45000 6 S4END[14]
port 366 nsew signal input
rlabel metal2 s 33138 44840 33194 45000 6 S4END[15]
port 367 nsew signal input
rlabel metal2 s 27986 44840 28042 45000 6 S4END[1]
port 368 nsew signal input
rlabel metal2 s 28354 44840 28410 45000 6 S4END[2]
port 369 nsew signal input
rlabel metal2 s 28722 44840 28778 45000 6 S4END[3]
port 370 nsew signal input
rlabel metal2 s 29090 44840 29146 45000 6 S4END[4]
port 371 nsew signal input
rlabel metal2 s 29458 44840 29514 45000 6 S4END[5]
port 372 nsew signal input
rlabel metal2 s 29826 44840 29882 45000 6 S4END[6]
port 373 nsew signal input
rlabel metal2 s 30194 44840 30250 45000 6 S4END[7]
port 374 nsew signal input
rlabel metal2 s 30562 44840 30618 45000 6 S4END[8]
port 375 nsew signal input
rlabel metal2 s 30930 44840 30986 45000 6 S4END[9]
port 376 nsew signal input
rlabel metal2 s 33506 0 33562 160 6 SS4BEG[0]
port 377 nsew signal output
rlabel metal2 s 37186 0 37242 160 6 SS4BEG[10]
port 378 nsew signal output
rlabel metal2 s 37554 0 37610 160 6 SS4BEG[11]
port 379 nsew signal output
rlabel metal2 s 37922 0 37978 160 6 SS4BEG[12]
port 380 nsew signal output
rlabel metal2 s 38290 0 38346 160 6 SS4BEG[13]
port 381 nsew signal output
rlabel metal2 s 38658 0 38714 160 6 SS4BEG[14]
port 382 nsew signal output
rlabel metal2 s 39026 0 39082 160 6 SS4BEG[15]
port 383 nsew signal output
rlabel metal2 s 33874 0 33930 160 6 SS4BEG[1]
port 384 nsew signal output
rlabel metal2 s 34242 0 34298 160 6 SS4BEG[2]
port 385 nsew signal output
rlabel metal2 s 34610 0 34666 160 6 SS4BEG[3]
port 386 nsew signal output
rlabel metal2 s 34978 0 35034 160 6 SS4BEG[4]
port 387 nsew signal output
rlabel metal2 s 35346 0 35402 160 6 SS4BEG[5]
port 388 nsew signal output
rlabel metal2 s 35714 0 35770 160 6 SS4BEG[6]
port 389 nsew signal output
rlabel metal2 s 36082 0 36138 160 6 SS4BEG[7]
port 390 nsew signal output
rlabel metal2 s 36450 0 36506 160 6 SS4BEG[8]
port 391 nsew signal output
rlabel metal2 s 36818 0 36874 160 6 SS4BEG[9]
port 392 nsew signal output
rlabel metal2 s 33506 44840 33562 45000 6 SS4END[0]
port 393 nsew signal input
rlabel metal2 s 37186 44840 37242 45000 6 SS4END[10]
port 394 nsew signal input
rlabel metal2 s 37554 44840 37610 45000 6 SS4END[11]
port 395 nsew signal input
rlabel metal2 s 37922 44840 37978 45000 6 SS4END[12]
port 396 nsew signal input
rlabel metal2 s 38290 44840 38346 45000 6 SS4END[13]
port 397 nsew signal input
rlabel metal2 s 38658 44840 38714 45000 6 SS4END[14]
port 398 nsew signal input
rlabel metal2 s 39026 44840 39082 45000 6 SS4END[15]
port 399 nsew signal input
rlabel metal2 s 33874 44840 33930 45000 6 SS4END[1]
port 400 nsew signal input
rlabel metal2 s 34242 44840 34298 45000 6 SS4END[2]
port 401 nsew signal input
rlabel metal2 s 34610 44840 34666 45000 6 SS4END[3]
port 402 nsew signal input
rlabel metal2 s 34978 44840 35034 45000 6 SS4END[4]
port 403 nsew signal input
rlabel metal2 s 35346 44840 35402 45000 6 SS4END[5]
port 404 nsew signal input
rlabel metal2 s 35714 44840 35770 45000 6 SS4END[6]
port 405 nsew signal input
rlabel metal2 s 36082 44840 36138 45000 6 SS4END[7]
port 406 nsew signal input
rlabel metal2 s 36450 44840 36506 45000 6 SS4END[8]
port 407 nsew signal input
rlabel metal2 s 36818 44840 36874 45000 6 SS4END[9]
port 408 nsew signal input
rlabel metal2 s 39394 0 39450 160 6 UserCLK
port 409 nsew signal input
rlabel metal2 s 39394 44840 39450 45000 6 UserCLKo
port 410 nsew signal output
rlabel metal4 s 19568 1040 19888 43568 6 VGND
port 411 nsew ground bidirectional
rlabel metal4 s 4208 1040 4528 43568 6 VPWR
port 412 nsew power bidirectional
rlabel metal4 s 34928 1040 35248 43568 6 VPWR
port 412 nsew power bidirectional
rlabel metal3 s 0 5176 160 5296 6 W1BEG[0]
port 413 nsew signal output
rlabel metal3 s 0 5448 160 5568 6 W1BEG[1]
port 414 nsew signal output
rlabel metal3 s 0 5720 160 5840 6 W1BEG[2]
port 415 nsew signal output
rlabel metal3 s 0 5992 160 6112 6 W1BEG[3]
port 416 nsew signal output
rlabel metal3 s 47840 5176 48000 5296 6 W1END[0]
port 417 nsew signal input
rlabel metal3 s 47840 5448 48000 5568 6 W1END[1]
port 418 nsew signal input
rlabel metal3 s 47840 5720 48000 5840 6 W1END[2]
port 419 nsew signal input
rlabel metal3 s 47840 5992 48000 6112 6 W1END[3]
port 420 nsew signal input
rlabel metal3 s 0 6264 160 6384 6 W2BEG[0]
port 421 nsew signal output
rlabel metal3 s 0 6536 160 6656 6 W2BEG[1]
port 422 nsew signal output
rlabel metal3 s 0 6808 160 6928 6 W2BEG[2]
port 423 nsew signal output
rlabel metal3 s 0 7080 160 7200 6 W2BEG[3]
port 424 nsew signal output
rlabel metal3 s 0 7352 160 7472 6 W2BEG[4]
port 425 nsew signal output
rlabel metal3 s 0 7624 160 7744 6 W2BEG[5]
port 426 nsew signal output
rlabel metal3 s 0 7896 160 8016 6 W2BEG[6]
port 427 nsew signal output
rlabel metal3 s 0 8168 160 8288 6 W2BEG[7]
port 428 nsew signal output
rlabel metal3 s 0 8440 160 8560 6 W2BEGb[0]
port 429 nsew signal output
rlabel metal3 s 0 8712 160 8832 6 W2BEGb[1]
port 430 nsew signal output
rlabel metal3 s 0 8984 160 9104 6 W2BEGb[2]
port 431 nsew signal output
rlabel metal3 s 0 9256 160 9376 6 W2BEGb[3]
port 432 nsew signal output
rlabel metal3 s 0 9528 160 9648 6 W2BEGb[4]
port 433 nsew signal output
rlabel metal3 s 0 9800 160 9920 6 W2BEGb[5]
port 434 nsew signal output
rlabel metal3 s 0 10072 160 10192 6 W2BEGb[6]
port 435 nsew signal output
rlabel metal3 s 0 10344 160 10464 6 W2BEGb[7]
port 436 nsew signal output
rlabel metal3 s 47840 8440 48000 8560 6 W2END[0]
port 437 nsew signal input
rlabel metal3 s 47840 8712 48000 8832 6 W2END[1]
port 438 nsew signal input
rlabel metal3 s 47840 8984 48000 9104 6 W2END[2]
port 439 nsew signal input
rlabel metal3 s 47840 9256 48000 9376 6 W2END[3]
port 440 nsew signal input
rlabel metal3 s 47840 9528 48000 9648 6 W2END[4]
port 441 nsew signal input
rlabel metal3 s 47840 9800 48000 9920 6 W2END[5]
port 442 nsew signal input
rlabel metal3 s 47840 10072 48000 10192 6 W2END[6]
port 443 nsew signal input
rlabel metal3 s 47840 10344 48000 10464 6 W2END[7]
port 444 nsew signal input
rlabel metal3 s 47840 6264 48000 6384 6 W2MID[0]
port 445 nsew signal input
rlabel metal3 s 47840 6536 48000 6656 6 W2MID[1]
port 446 nsew signal input
rlabel metal3 s 47840 6808 48000 6928 6 W2MID[2]
port 447 nsew signal input
rlabel metal3 s 47840 7080 48000 7200 6 W2MID[3]
port 448 nsew signal input
rlabel metal3 s 47840 7352 48000 7472 6 W2MID[4]
port 449 nsew signal input
rlabel metal3 s 47840 7624 48000 7744 6 W2MID[5]
port 450 nsew signal input
rlabel metal3 s 47840 7896 48000 8016 6 W2MID[6]
port 451 nsew signal input
rlabel metal3 s 47840 8168 48000 8288 6 W2MID[7]
port 452 nsew signal input
rlabel metal3 s 0 14968 160 15088 6 W6BEG[0]
port 453 nsew signal output
rlabel metal3 s 0 17688 160 17808 6 W6BEG[10]
port 454 nsew signal output
rlabel metal3 s 0 17960 160 18080 6 W6BEG[11]
port 455 nsew signal output
rlabel metal3 s 0 15240 160 15360 6 W6BEG[1]
port 456 nsew signal output
rlabel metal3 s 0 15512 160 15632 6 W6BEG[2]
port 457 nsew signal output
rlabel metal3 s 0 15784 160 15904 6 W6BEG[3]
port 458 nsew signal output
rlabel metal3 s 0 16056 160 16176 6 W6BEG[4]
port 459 nsew signal output
rlabel metal3 s 0 16328 160 16448 6 W6BEG[5]
port 460 nsew signal output
rlabel metal3 s 0 16600 160 16720 6 W6BEG[6]
port 461 nsew signal output
rlabel metal3 s 0 16872 160 16992 6 W6BEG[7]
port 462 nsew signal output
rlabel metal3 s 0 17144 160 17264 6 W6BEG[8]
port 463 nsew signal output
rlabel metal3 s 0 17416 160 17536 6 W6BEG[9]
port 464 nsew signal output
rlabel metal3 s 47840 14968 48000 15088 6 W6END[0]
port 465 nsew signal input
rlabel metal3 s 47840 17688 48000 17808 6 W6END[10]
port 466 nsew signal input
rlabel metal3 s 47840 17960 48000 18080 6 W6END[11]
port 467 nsew signal input
rlabel metal3 s 47840 15240 48000 15360 6 W6END[1]
port 468 nsew signal input
rlabel metal3 s 47840 15512 48000 15632 6 W6END[2]
port 469 nsew signal input
rlabel metal3 s 47840 15784 48000 15904 6 W6END[3]
port 470 nsew signal input
rlabel metal3 s 47840 16056 48000 16176 6 W6END[4]
port 471 nsew signal input
rlabel metal3 s 47840 16328 48000 16448 6 W6END[5]
port 472 nsew signal input
rlabel metal3 s 47840 16600 48000 16720 6 W6END[6]
port 473 nsew signal input
rlabel metal3 s 47840 16872 48000 16992 6 W6END[7]
port 474 nsew signal input
rlabel metal3 s 47840 17144 48000 17264 6 W6END[8]
port 475 nsew signal input
rlabel metal3 s 47840 17416 48000 17536 6 W6END[9]
port 476 nsew signal input
rlabel metal3 s 0 10616 160 10736 6 WW4BEG[0]
port 477 nsew signal output
rlabel metal3 s 0 13336 160 13456 6 WW4BEG[10]
port 478 nsew signal output
rlabel metal3 s 0 13608 160 13728 6 WW4BEG[11]
port 479 nsew signal output
rlabel metal3 s 0 13880 160 14000 6 WW4BEG[12]
port 480 nsew signal output
rlabel metal3 s 0 14152 160 14272 6 WW4BEG[13]
port 481 nsew signal output
rlabel metal3 s 0 14424 160 14544 6 WW4BEG[14]
port 482 nsew signal output
rlabel metal3 s 0 14696 160 14816 6 WW4BEG[15]
port 483 nsew signal output
rlabel metal3 s 0 10888 160 11008 6 WW4BEG[1]
port 484 nsew signal output
rlabel metal3 s 0 11160 160 11280 6 WW4BEG[2]
port 485 nsew signal output
rlabel metal3 s 0 11432 160 11552 6 WW4BEG[3]
port 486 nsew signal output
rlabel metal3 s 0 11704 160 11824 6 WW4BEG[4]
port 487 nsew signal output
rlabel metal3 s 0 11976 160 12096 6 WW4BEG[5]
port 488 nsew signal output
rlabel metal3 s 0 12248 160 12368 6 WW4BEG[6]
port 489 nsew signal output
rlabel metal3 s 0 12520 160 12640 6 WW4BEG[7]
port 490 nsew signal output
rlabel metal3 s 0 12792 160 12912 6 WW4BEG[8]
port 491 nsew signal output
rlabel metal3 s 0 13064 160 13184 6 WW4BEG[9]
port 492 nsew signal output
rlabel metal3 s 47840 10616 48000 10736 6 WW4END[0]
port 493 nsew signal input
rlabel metal3 s 47840 13336 48000 13456 6 WW4END[10]
port 494 nsew signal input
rlabel metal3 s 47840 13608 48000 13728 6 WW4END[11]
port 495 nsew signal input
rlabel metal3 s 47840 13880 48000 14000 6 WW4END[12]
port 496 nsew signal input
rlabel metal3 s 47840 14152 48000 14272 6 WW4END[13]
port 497 nsew signal input
rlabel metal3 s 47840 14424 48000 14544 6 WW4END[14]
port 498 nsew signal input
rlabel metal3 s 47840 14696 48000 14816 6 WW4END[15]
port 499 nsew signal input
rlabel metal3 s 47840 10888 48000 11008 6 WW4END[1]
port 500 nsew signal input
rlabel metal3 s 47840 11160 48000 11280 6 WW4END[2]
port 501 nsew signal input
rlabel metal3 s 47840 11432 48000 11552 6 WW4END[3]
port 502 nsew signal input
rlabel metal3 s 47840 11704 48000 11824 6 WW4END[4]
port 503 nsew signal input
rlabel metal3 s 47840 11976 48000 12096 6 WW4END[5]
port 504 nsew signal input
rlabel metal3 s 47840 12248 48000 12368 6 WW4END[6]
port 505 nsew signal input
rlabel metal3 s 47840 12520 48000 12640 6 WW4END[7]
port 506 nsew signal input
rlabel metal3 s 47840 12792 48000 12912 6 WW4END[8]
port 507 nsew signal input
rlabel metal3 s 47840 13064 48000 13184 6 WW4END[9]
port 508 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 48000 45000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7626878
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/RegFile/runs/24_12_04_10_28/results/signoff/RegFile.magic.gds
string GDS_START 292334
<< end >>

