* NGSPICE file created from DSP.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxbp_1 abstract view
.subckt sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

.subckt DSP Tile_X0Y0_E1BEG[0] Tile_X0Y0_E1BEG[1] Tile_X0Y0_E1BEG[2] Tile_X0Y0_E1BEG[3]
+ Tile_X0Y0_E1END[0] Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2] Tile_X0Y0_E1END[3] Tile_X0Y0_E2BEG[0]
+ Tile_X0Y0_E2BEG[1] Tile_X0Y0_E2BEG[2] Tile_X0Y0_E2BEG[3] Tile_X0Y0_E2BEG[4] Tile_X0Y0_E2BEG[5]
+ Tile_X0Y0_E2BEG[6] Tile_X0Y0_E2BEG[7] Tile_X0Y0_E2BEGb[0] Tile_X0Y0_E2BEGb[1] Tile_X0Y0_E2BEGb[2]
+ Tile_X0Y0_E2BEGb[3] Tile_X0Y0_E2BEGb[4] Tile_X0Y0_E2BEGb[5] Tile_X0Y0_E2BEGb[6]
+ Tile_X0Y0_E2BEGb[7] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1] Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6] Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3] Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6BEG[0] Tile_X0Y0_E6BEG[10] Tile_X0Y0_E6BEG[11]
+ Tile_X0Y0_E6BEG[1] Tile_X0Y0_E6BEG[2] Tile_X0Y0_E6BEG[3] Tile_X0Y0_E6BEG[4] Tile_X0Y0_E6BEG[5]
+ Tile_X0Y0_E6BEG[6] Tile_X0Y0_E6BEG[7] Tile_X0Y0_E6BEG[8] Tile_X0Y0_E6BEG[9] Tile_X0Y0_E6END[0]
+ Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11] Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3]
+ Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5] Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8]
+ Tile_X0Y0_E6END[9] Tile_X0Y0_EE4BEG[0] Tile_X0Y0_EE4BEG[10] Tile_X0Y0_EE4BEG[11]
+ Tile_X0Y0_EE4BEG[12] Tile_X0Y0_EE4BEG[13] Tile_X0Y0_EE4BEG[14] Tile_X0Y0_EE4BEG[15]
+ Tile_X0Y0_EE4BEG[1] Tile_X0Y0_EE4BEG[2] Tile_X0Y0_EE4BEG[3] Tile_X0Y0_EE4BEG[4]
+ Tile_X0Y0_EE4BEG[5] Tile_X0Y0_EE4BEG[6] Tile_X0Y0_EE4BEG[7] Tile_X0Y0_EE4BEG[8]
+ Tile_X0Y0_EE4BEG[9] Tile_X0Y0_EE4END[0] Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13] Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15]
+ Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2] Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4]
+ Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11]
+ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15]
+ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19]
+ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22]
+ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26]
+ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2]
+ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4]
+ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8]
+ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0] Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11]
+ Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13] Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15]
+ Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17] Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19]
+ Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20] Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22]
+ Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24] Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26]
+ Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28] Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2]
+ Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31] Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4]
+ Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6] Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8]
+ Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0] Tile_X0Y0_FrameStrobe_O[10]
+ Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12] Tile_X0Y0_FrameStrobe_O[13]
+ Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15] Tile_X0Y0_FrameStrobe_O[16]
+ Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18] Tile_X0Y0_FrameStrobe_O[19]
+ Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2] Tile_X0Y0_FrameStrobe_O[3]
+ Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5] Tile_X0Y0_FrameStrobe_O[6]
+ Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8] Tile_X0Y0_FrameStrobe_O[9]
+ Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2] Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0]
+ Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3] Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5]
+ Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0] Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2]
+ Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4] Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6]
+ Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10] Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12]
+ Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14] Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2]
+ Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4] Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7]
+ Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9] Tile_X0Y0_NN4BEG[0] Tile_X0Y0_NN4BEG[10] Tile_X0Y0_NN4BEG[11]
+ Tile_X0Y0_NN4BEG[12] Tile_X0Y0_NN4BEG[13] Tile_X0Y0_NN4BEG[14] Tile_X0Y0_NN4BEG[15]
+ Tile_X0Y0_NN4BEG[1] Tile_X0Y0_NN4BEG[2] Tile_X0Y0_NN4BEG[3] Tile_X0Y0_NN4BEG[4]
+ Tile_X0Y0_NN4BEG[5] Tile_X0Y0_NN4BEG[6] Tile_X0Y0_NN4BEG[7] Tile_X0Y0_NN4BEG[8]
+ Tile_X0Y0_NN4BEG[9] Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2] Tile_X0Y0_S1END[3]
+ Tile_X0Y0_S2END[0] Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3] Tile_X0Y0_S2END[4]
+ Tile_X0Y0_S2END[5] Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0] Tile_X0Y0_S2MID[1]
+ Tile_X0Y0_S2MID[2] Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5] Tile_X0Y0_S2MID[6]
+ Tile_X0Y0_S2MID[7] Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11] Tile_X0Y0_S4END[12]
+ Tile_X0Y0_S4END[13] Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15] Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2]
+ Tile_X0Y0_S4END[3] Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5] Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7]
+ Tile_X0Y0_S4END[8] Tile_X0Y0_S4END[9] Tile_X0Y0_SS4END[0] Tile_X0Y0_SS4END[10] Tile_X0Y0_SS4END[11]
+ Tile_X0Y0_SS4END[12] Tile_X0Y0_SS4END[13] Tile_X0Y0_SS4END[14] Tile_X0Y0_SS4END[15]
+ Tile_X0Y0_SS4END[1] Tile_X0Y0_SS4END[2] Tile_X0Y0_SS4END[3] Tile_X0Y0_SS4END[4]
+ Tile_X0Y0_SS4END[5] Tile_X0Y0_SS4END[6] Tile_X0Y0_SS4END[7] Tile_X0Y0_SS4END[8]
+ Tile_X0Y0_SS4END[9] Tile_X0Y0_UserCLKo Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2]
+ Tile_X0Y0_W1BEG[3] Tile_X0Y0_W1END[0] Tile_X0Y0_W1END[1] Tile_X0Y0_W1END[2] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_W2BEG[0] Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3] Tile_X0Y0_W2BEG[4]
+ Tile_X0Y0_W2BEG[5] Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0] Tile_X0Y0_W2BEGb[1]
+ Tile_X0Y0_W2BEGb[2] Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4] Tile_X0Y0_W2BEGb[5]
+ Tile_X0Y0_W2BEGb[6] Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W2END[0] Tile_X0Y0_W2END[1] Tile_X0Y0_W2END[2]
+ Tile_X0Y0_W2END[3] Tile_X0Y0_W2END[4] Tile_X0Y0_W2END[5] Tile_X0Y0_W2END[6] Tile_X0Y0_W2END[7]
+ Tile_X0Y0_W2MID[0] Tile_X0Y0_W2MID[1] Tile_X0Y0_W2MID[2] Tile_X0Y0_W2MID[3] Tile_X0Y0_W2MID[4]
+ Tile_X0Y0_W2MID[5] Tile_X0Y0_W2MID[6] Tile_X0Y0_W2MID[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10]
+ Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1] Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4]
+ Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6] Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9]
+ Tile_X0Y0_W6END[0] Tile_X0Y0_W6END[10] Tile_X0Y0_W6END[11] Tile_X0Y0_W6END[1] Tile_X0Y0_W6END[2]
+ Tile_X0Y0_W6END[3] Tile_X0Y0_W6END[4] Tile_X0Y0_W6END[5] Tile_X0Y0_W6END[6] Tile_X0Y0_W6END[7]
+ Tile_X0Y0_W6END[8] Tile_X0Y0_W6END[9] Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10] Tile_X0Y0_WW4BEG[11]
+ Tile_X0Y0_WW4BEG[12] Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14] Tile_X0Y0_WW4BEG[15]
+ Tile_X0Y0_WW4BEG[1] Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3] Tile_X0Y0_WW4BEG[4]
+ Tile_X0Y0_WW4BEG[5] Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7] Tile_X0Y0_WW4BEG[8]
+ Tile_X0Y0_WW4BEG[9] Tile_X0Y0_WW4END[0] Tile_X0Y0_WW4END[10] Tile_X0Y0_WW4END[11]
+ Tile_X0Y0_WW4END[12] Tile_X0Y0_WW4END[13] Tile_X0Y0_WW4END[14] Tile_X0Y0_WW4END[15]
+ Tile_X0Y0_WW4END[1] Tile_X0Y0_WW4END[2] Tile_X0Y0_WW4END[3] Tile_X0Y0_WW4END[4]
+ Tile_X0Y0_WW4END[5] Tile_X0Y0_WW4END[6] Tile_X0Y0_WW4END[7] Tile_X0Y0_WW4END[8]
+ Tile_X0Y0_WW4END[9] Tile_X0Y1_E1BEG[0] Tile_X0Y1_E1BEG[1] Tile_X0Y1_E1BEG[2] Tile_X0Y1_E1BEG[3]
+ Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2] Tile_X0Y1_E1END[3] Tile_X0Y1_E2BEG[0]
+ Tile_X0Y1_E2BEG[1] Tile_X0Y1_E2BEG[2] Tile_X0Y1_E2BEG[3] Tile_X0Y1_E2BEG[4] Tile_X0Y1_E2BEG[5]
+ Tile_X0Y1_E2BEG[6] Tile_X0Y1_E2BEG[7] Tile_X0Y1_E2BEGb[0] Tile_X0Y1_E2BEGb[1] Tile_X0Y1_E2BEGb[2]
+ Tile_X0Y1_E2BEGb[3] Tile_X0Y1_E2BEGb[4] Tile_X0Y1_E2BEGb[5] Tile_X0Y1_E2BEGb[6]
+ Tile_X0Y1_E2BEGb[7] Tile_X0Y1_E2END[0] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3]
+ Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5] Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0]
+ Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2] Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7] Tile_X0Y1_E6BEG[0] Tile_X0Y1_E6BEG[10] Tile_X0Y1_E6BEG[11]
+ Tile_X0Y1_E6BEG[1] Tile_X0Y1_E6BEG[2] Tile_X0Y1_E6BEG[3] Tile_X0Y1_E6BEG[4] Tile_X0Y1_E6BEG[5]
+ Tile_X0Y1_E6BEG[6] Tile_X0Y1_E6BEG[7] Tile_X0Y1_E6BEG[8] Tile_X0Y1_E6BEG[9] Tile_X0Y1_E6END[0]
+ Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11] Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2] Tile_X0Y1_E6END[3]
+ Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5] Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7] Tile_X0Y1_E6END[8]
+ Tile_X0Y1_E6END[9] Tile_X0Y1_EE4BEG[0] Tile_X0Y1_EE4BEG[10] Tile_X0Y1_EE4BEG[11]
+ Tile_X0Y1_EE4BEG[12] Tile_X0Y1_EE4BEG[13] Tile_X0Y1_EE4BEG[14] Tile_X0Y1_EE4BEG[15]
+ Tile_X0Y1_EE4BEG[1] Tile_X0Y1_EE4BEG[2] Tile_X0Y1_EE4BEG[3] Tile_X0Y1_EE4BEG[4]
+ Tile_X0Y1_EE4BEG[5] Tile_X0Y1_EE4BEG[6] Tile_X0Y1_EE4BEG[7] Tile_X0Y1_EE4BEG[8]
+ Tile_X0Y1_EE4BEG[9] Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13] Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11]
+ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15]
+ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19]
+ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22]
+ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26]
+ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2]
+ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4]
+ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8]
+ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0] Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11]
+ Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13] Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15]
+ Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17] Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19]
+ Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20] Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22]
+ Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24] Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26]
+ Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28] Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2]
+ Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31] Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4]
+ Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6] Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8]
+ Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11]
+ Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13] Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15]
+ Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17] Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19]
+ Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4]
+ Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8]
+ Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0] Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1] Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3]
+ Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6] Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0]
+ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3] Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0] Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11]
+ Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13] Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15]
+ Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3] Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5]
+ Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8] Tile_X0Y1_N4END[9] Tile_X0Y1_NN4END[0]
+ Tile_X0Y1_NN4END[10] Tile_X0Y1_NN4END[11] Tile_X0Y1_NN4END[12] Tile_X0Y1_NN4END[13]
+ Tile_X0Y1_NN4END[14] Tile_X0Y1_NN4END[15] Tile_X0Y1_NN4END[1] Tile_X0Y1_NN4END[2]
+ Tile_X0Y1_NN4END[3] Tile_X0Y1_NN4END[4] Tile_X0Y1_NN4END[5] Tile_X0Y1_NN4END[6]
+ Tile_X0Y1_NN4END[7] Tile_X0Y1_NN4END[8] Tile_X0Y1_NN4END[9] Tile_X0Y1_S1BEG[0] Tile_X0Y1_S1BEG[1]
+ Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3] Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1] Tile_X0Y1_S2BEG[2]
+ Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4] Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6] Tile_X0Y1_S2BEG[7]
+ Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1] Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3]
+ Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5] Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7]
+ Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11] Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13]
+ Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15] Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3]
+ Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5] Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8]
+ Tile_X0Y1_S4BEG[9] Tile_X0Y1_SS4BEG[0] Tile_X0Y1_SS4BEG[10] Tile_X0Y1_SS4BEG[11]
+ Tile_X0Y1_SS4BEG[12] Tile_X0Y1_SS4BEG[13] Tile_X0Y1_SS4BEG[14] Tile_X0Y1_SS4BEG[15]
+ Tile_X0Y1_SS4BEG[1] Tile_X0Y1_SS4BEG[2] Tile_X0Y1_SS4BEG[3] Tile_X0Y1_SS4BEG[4]
+ Tile_X0Y1_SS4BEG[5] Tile_X0Y1_SS4BEG[6] Tile_X0Y1_SS4BEG[7] Tile_X0Y1_SS4BEG[8]
+ Tile_X0Y1_SS4BEG[9] Tile_X0Y1_UserCLK Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2]
+ Tile_X0Y1_W1BEG[3] Tile_X0Y1_W1END[0] Tile_X0Y1_W1END[1] Tile_X0Y1_W1END[2] Tile_X0Y1_W1END[3]
+ Tile_X0Y1_W2BEG[0] Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3] Tile_X0Y1_W2BEG[4]
+ Tile_X0Y1_W2BEG[5] Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0] Tile_X0Y1_W2BEGb[1]
+ Tile_X0Y1_W2BEGb[2] Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4] Tile_X0Y1_W2BEGb[5]
+ Tile_X0Y1_W2BEGb[6] Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W2END[0] Tile_X0Y1_W2END[1] Tile_X0Y1_W2END[2]
+ Tile_X0Y1_W2END[3] Tile_X0Y1_W2END[4] Tile_X0Y1_W2END[5] Tile_X0Y1_W2END[6] Tile_X0Y1_W2END[7]
+ Tile_X0Y1_W2MID[0] Tile_X0Y1_W2MID[1] Tile_X0Y1_W2MID[2] Tile_X0Y1_W2MID[3] Tile_X0Y1_W2MID[4]
+ Tile_X0Y1_W2MID[5] Tile_X0Y1_W2MID[6] Tile_X0Y1_W2MID[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10]
+ Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1] Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4]
+ Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6] Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9]
+ Tile_X0Y1_W6END[0] Tile_X0Y1_W6END[10] Tile_X0Y1_W6END[11] Tile_X0Y1_W6END[1] Tile_X0Y1_W6END[2]
+ Tile_X0Y1_W6END[3] Tile_X0Y1_W6END[4] Tile_X0Y1_W6END[5] Tile_X0Y1_W6END[6] Tile_X0Y1_W6END[7]
+ Tile_X0Y1_W6END[8] Tile_X0Y1_W6END[9] Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10] Tile_X0Y1_WW4BEG[11]
+ Tile_X0Y1_WW4BEG[12] Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14] Tile_X0Y1_WW4BEG[15]
+ Tile_X0Y1_WW4BEG[1] Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3] Tile_X0Y1_WW4BEG[4]
+ Tile_X0Y1_WW4BEG[5] Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7] Tile_X0Y1_WW4BEG[8]
+ Tile_X0Y1_WW4BEG[9] Tile_X0Y1_WW4END[0] Tile_X0Y1_WW4END[10] Tile_X0Y1_WW4END[11]
+ Tile_X0Y1_WW4END[12] Tile_X0Y1_WW4END[13] Tile_X0Y1_WW4END[14] Tile_X0Y1_WW4END[15]
+ Tile_X0Y1_WW4END[1] Tile_X0Y1_WW4END[2] Tile_X0Y1_WW4END[3] Tile_X0Y1_WW4END[4]
+ Tile_X0Y1_WW4END[5] Tile_X0Y1_WW4END[6] Tile_X0Y1_WW4END[7] Tile_X0Y1_WW4END[8]
+ Tile_X0Y1_WW4END[9] VGND VPWR
XTile_X0Y1_DSP_bot_Inst_MULADD__1555_ Tile_X0Y1_DSP_bot_Inst_MULADD__1554_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1554_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1554_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1556_/B
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1486_ Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/X sky130_fd_sc_hd__and4_1
XFILLER_0_89_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_NN4END_inbuf_0__0_ net327 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/NN4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__58_ Tile_X0Y1_DSP_bot/JS2BEG\[4\] VGND
+ VGND VPWR VPWR net671 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_N4BEG_outbuf_3__0_ ANTENNA_75/DIODE VGND VGND VPWR VPWR net511
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[21\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_213 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_202 Tile_X0Y0_SS4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_data_outbuf_5__0_ Tile_X0Y1_DSP_bot_data_inbuf_5__0_/X VGND VGND
+ VPWR VPWR net658 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit28 net249 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[316\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit17 net237 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[305\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1
+ net88 net110 net140 net156 Tile_X0Y0_DSP_top/ConfigBits\[350\] Tile_X0Y0_DSP_top/ConfigBits\[351\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_data_outbuf_27__0_ Tile_X0Y1_DSP_bot_data_inbuf_27__0_/X VGND VGND
+ VPWR VPWR net650 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1340_ Tile_X0Y1_DSP_bot_Inst_MULADD__1255_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1338_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1339_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1342_/A
+ sky130_fd_sc_hd__o21a_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1271_ Tile_X0Y1_DSP_bot_Inst_MULADD__1093_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1095_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/B
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit9 net260 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[393\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_86_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG0 Tile_X0Y1_N2BEG\[7\]
+ net20 net100 net152 Tile_X0Y0_DSP_top/ConfigBits\[190\] Tile_X0Y0_DSP_top/ConfigBits\[191\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[0\] sky130_fd_sc_hd__mux4_1
Xoutput401 net401 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0986_ Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/B Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0973_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0986_/Y sky130_fd_sc_hd__a221oi_2
Xoutput434 net434 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[13] sky130_fd_sc_hd__buf_2
Xoutput412 net412 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput423 net423 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_data_inbuf_29__0_ net250 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_29__0_/X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput467 net467 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[14] sky130_fd_sc_hd__clkbuf_4
Xoutput478 net478 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[6] sky130_fd_sc_hd__clkbuf_4
Xoutput445 net445 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput456 net456 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[4] sky130_fd_sc_hd__buf_2
Xoutput489 net489 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit1 net240 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[97\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit0 net49 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[278\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_data_outbuf_18__0_ Tile_X0Y1_DSP_bot_data_inbuf_18__0_/X VGND VGND
+ VPWR VPWR net640 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1607_ Tile_X0Y1_DSP_bot_Inst_MULADD__1629_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1629_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1606_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1620_/B
+ sky130_fd_sc_hd__a21boi_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1538_ Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1479_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1488_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1484_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1538_/X sky130_fd_sc_hd__o311a_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1469_ Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1716_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1469_/X sky130_fd_sc_hd__and2_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_S4BEG_outbuf_7__0_ Tile_X0Y1_DSP_bot/S4BEG_i\[7\] VGND VGND VPWR
+ VPWR net696 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_W6BEG_outbuf_3__0_ Tile_X0Y0_DSP_top/W6BEG_i\[3\] VGND VGND VPWR
+ VPWR net560 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[146\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit10 net50 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[160\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit21 net62 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[171\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[1\] Tile_X0Y1_N2BEGb\[5\] net2 net10 Tile_X0Y0_DSP_top/ConfigBits\[262\]
+ Tile_X0Y0_DSP_top/ConfigBits\[263\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_141_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1323_ Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/C
+ sky130_fd_sc_hd__nand3_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_S1BEG2 Tile_X0Y1_bot2top\[6\]
+ Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[1\] Tile_X0Y0_DSP_top/JE2BEG\[1\] Tile_X0Y0_DSP_top/J_l_GH_BEG\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[60\] Tile_X0Y0_DSP_top/ConfigBits\[61\] VGND VGND
+ VPWR VPWR Tile_X0Y0_S1BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_91_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1254_ Tile_X0Y1_DSP_bot_Inst_MULADD__1339_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1339_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1255_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1185_ Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1733_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_115_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0969_ Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1736_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0969_/X sky130_fd_sc_hd__and2_2
XTile_X0Y0_DSP_top_E6END_inbuf_1__0_ net26 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/E6BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[8\] Tile_X0Y0_DSP_top/J2MID_EFb_BEG\[1\] Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2END_CD_BEG\[2\] Tile_X0Y0_DSP_top/ConfigBits\[98\] Tile_X0Y0_DSP_top/ConfigBits\[99\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[0\] Tile_X0Y0_S1BEG\[2\] Tile_X0Y0_S2BEGb\[6\] net336 Tile_X0Y1_DSP_bot/ConfigBits\[372\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[373\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit16 net236 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[336\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit27 net248 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[347\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[27\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_NN4BEG\[13\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_data_outbuf_23__0_ Tile_X0Y0_DSP_top_data_inbuf_23__0_/X VGND VGND
+ VPWR VPWR net445 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1
+ net109 net125 net139 net153 Tile_X0Y0_DSP_top/ConfigBits\[314\] Tile_X0Y0_DSP_top/ConfigBits\[315\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[38\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit4 net255 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[196\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_W1BEG0 Tile_X0Y1_DSP_bot/Q5
+ Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[3\] Tile_X0Y1_DSP_bot/JS2BEG\[3\] Tile_X0Y1_DSP_bot/J_l_CD_BEG\[1\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[90\] Tile_X0Y1_DSP_bot/ConfigBits\[91\] VGND VGND
+ VPWR VPWR net715 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_data_outbuf_14__0_ Tile_X0Y0_DSP_top_data_inbuf_14__0_/X VGND VGND
+ VPWR VPWR net435 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit3 net74 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[377\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1306_ Tile_X0Y1_DSP_bot_Inst_MULADD__1306_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1306_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1306_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_66_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1237_ Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_S4BEG_outbuf_3__0_ Tile_X0Y0_DSP_top/S4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_S4BEG\[3\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1168_ Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1712_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1099_ Tile_X0Y1_DSP_bot_Inst_MULADD__1097_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0895_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1099_/Y
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit20 net61 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[202\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0
+ net281 net285 net181 net213 Tile_X0Y1_DSP_bot/ConfigBits\[284\] Tile_X0Y1_DSP_bot/ConfigBits\[285\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit31 net73 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[213\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_E6END_inbuf_1__0_ net206 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/E6BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1022_ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1054_/C sky130_fd_sc_hd__nand4_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__91_ Tile_X0Y1_DSP_bot/Q15 VGND VGND
+ VPWR VPWR Tile_X0Y1_bot2top\[5\] sky130_fd_sc_hd__buf_12
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[100\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_strobe_outbuf_7__0_ Tile_X0Y0_DSP_top_strobe_inbuf_7__0_/X VGND
+ VGND VPWR VPWR net479 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit15 net235 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[367\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit26 net247 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[378\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit24 net65 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[110\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit13 net53 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[99\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[278\] Tile_X0Y0_DSP_top/ConfigBits\[279\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_153_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[1\] Tile_X0Y0_S2BEGb\[5\] net335 net337 Tile_X0Y1_DSP_bot/ConfigBits\[336\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[337\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_data_inbuf_4__0_ net255 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_4__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__12_ net17 VGND VGND VPWR VPWR net398
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit9 net80 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[159\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_NN4END_inbuf_9__0_ Tile_X0Y1_NN4BEG\[13\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/NN4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[6\] Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[1\] Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2END_GH_BEG\[3\] Tile_X0Y0_DSP_top/ConfigBits\[72\] Tile_X0Y0_DSP_top/ConfigBits\[73\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
Xinput301 Tile_X0Y1_N4END[0] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_2
Xinput312 Tile_X0Y1_N4END[5] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_1
Xinput345 Tile_X0Y1_W2END[7] VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkbuf_4
Xinput334 Tile_X0Y1_W1END[0] VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkbuf_4
Xinput323 Tile_X0Y1_NN4END[15] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_1
Xinput378 Tile_X0Y1_WW4END[6] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_1
Xinput367 Tile_X0Y1_WW4END[10] VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput356 Tile_X0Y1_W6END[11] VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_strobe_outbuf_0__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_0__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[0\] sky130_fd_sc_hd__buf_8
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[104\] Tile_X0Y0_DSP_top/ConfigBits\[105\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_5 Tile_X0Y0_S2BEG\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1640_ Tile_X0Y1_DSP_bot_Inst_MULADD__1664_/S Tile_X0Y1_DSP_bot_Inst_MULADD__1640_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1640_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_67_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_WW4BEG_outbuf_5__0_ Tile_X0Y0_DSP_top/WW4BEG_i\[5\] VGND VGND VPWR
+ VPWR net578 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1571_ Tile_X0Y1_DSP_bot_Inst_MULADD__1588_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1560_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1570_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1578_/A
+ sky130_fd_sc_hd__o21ai_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[260\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[261\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit7 net258 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[295\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[44\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit30 net72 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[244\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit19 net239 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[275\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__74_ net342 VGND VGND VPWR VPWR net723
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1005_ Tile_X0Y1_DSP_bot_Inst_MULADD__1006_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1006_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1006_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1007_/A
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_inbuf_15__0_ net267 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_15__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput120 Tile_X0Y0_SS4END[12] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
Xinput131 Tile_X0Y0_SS4END[8] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
Xinput153 Tile_X0Y0_W6END[0] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_4
Xinput142 Tile_X0Y0_W2END[5] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
Xinput164 Tile_X0Y0_W6END[9] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_1
Xinput175 Tile_X0Y0_WW4END[4] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
Xinput186 Tile_X0Y1_E2END[1] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
Xinput197 Tile_X0Y1_E2MID[4] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__buf_2
XFILLER_0_128_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit14 net234 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[398\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit25 net246 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[409\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_N4END_inbuf_5__0_ Tile_X0Y1_N4BEG\[9\] VGND VGND VPWR VPWR ANTENNA_76/DIODE
+ sky130_fd_sc_hd__buf_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit12 net52 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[130\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 net764 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[300\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[301\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit23 net64 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[141\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput627 net627 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput616 net616 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput605 net605 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[11] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG0 Tile_X0Y1_N2BEG\[6\]
+ net99 net151 Tile_X0Y0_DSP_top/JN2BEG\[3\] Tile_X0Y0_DSP_top/ConfigBits\[150\] Tile_X0Y0_DSP_top/ConfigBits\[151\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_111_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput638 net638 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[16] sky130_fd_sc_hd__buf_2
Xoutput649 net649 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[26] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1623_ Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1721_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1554_ Tile_X0Y1_DSP_bot_Inst_MULADD__1554_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1554_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1554_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1556_/A
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1485_ Tile_X0Y1_DSP_bot_Inst_MULADD__1019_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1484_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1485_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_134_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__57_ Tile_X0Y1_DSP_bot/JS2BEG\[3\] VGND
+ VGND VPWR VPWR net670 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[106\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[21\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_203 Tile_X0Y0_SS4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_WW4END_inbuf_1__0_ net377 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/WW4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit29 net250 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[317\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit18 net238 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[306\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[350\] Tile_X0Y0_DSP_top/ConfigBits\[351\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1270_ Tile_X0Y1_DSP_bot_Inst_MULADD__0895_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1268_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1270_/Y sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y1_DSP_bot_strobe_inbuf_8__0_ net279 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_8__0_/X
+ sky130_fd_sc_hd__buf_1
XFILLER_0_148_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG1 Tile_X0Y1_N2BEG\[3\]
+ net16 net96 net148 Tile_X0Y0_DSP_top/ConfigBits\[192\] Tile_X0Y0_DSP_top/ConfigBits\[193\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_N4END_inbuf_5__0_ net316 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/N4BEG_i\[5\]
+ sky130_fd_sc_hd__buf_2
Xoutput402 net402 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_0_124_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__0985_ Tile_X0Y1_DSP_bot_Inst_MULADD__0974_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/B Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0984_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/B sky130_fd_sc_hd__o2111ai_4
Xoutput435 net435 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[14] sky130_fd_sc_hd__buf_2
Xoutput413 net413 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput424 net424 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput468 net468 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[15] sky130_fd_sc_hd__clkbuf_4
Xoutput446 net446 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput457 net457 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput479 net479 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[7] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit2 net251 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[98\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1606_ Tile_X0Y1_DSP_bot_Inst_MULADD__1604_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1518_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1605_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1581_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1606_/Y sky130_fd_sc_hd__o211ai_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_S4BEG0 net24 net87
+ net108 Tile_X0Y1_bot2top\[0\] Tile_X0Y0_DSP_top/ConfigBits\[64\] Tile_X0Y0_DSP_top/ConfigBits\[65\]
+ VGND VGND VPWR VPWR Tile_X0Y0_S4BEG\[12\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit1 net60 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[279\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1537_ Tile_X0Y1_DSP_bot_Inst_MULADD__1536_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1536_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1541_/C
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1468_ Tile_X0Y1_DSP_bot_Inst_MULADD__1465_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1604_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1465_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1690_/C sky130_fd_sc_hd__a22o_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1399_ Tile_X0Y1_DSP_bot_Inst_MULADD__1398_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1297_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1311_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1294_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1399_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit11 net51 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[161\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit22 net63 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[172\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1
+ net82 net90 net134 net136 Tile_X0Y0_DSP_top/ConfigBits\[262\] Tile_X0Y0_DSP_top/ConfigBits\[263\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG0 net310
+ net213 Tile_X0Y0_S4BEG\[3\] Tile_X0Y1_DSP_bot/JN2BEG\[4\] Tile_X0Y1_DSP_bot/ConfigBits\[408\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[409\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_GH_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1322_ Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/B
+ sky130_fd_sc_hd__a21o_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_S1BEG3 Tile_X0Y1_bot2top\[7\]
+ Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[2\] Tile_X0Y0_DSP_top/JE2BEG\[2\] ANTENNA_65/DIODE
+ Tile_X0Y0_DSP_top/ConfigBits\[62\] Tile_X0Y0_DSP_top/ConfigBits\[63\] VGND VGND
+ VPWR VPWR Tile_X0Y0_S1BEG\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_78_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1253_ Tile_X0Y1_DSP_bot_Inst_MULADD__1251_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1713_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1614_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1339_/B
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1184_ Tile_X0Y1_DSP_bot/A7 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1184_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_86_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__0968_ Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/A ANTENNA_97/DIODE
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0968_/Y sky130_fd_sc_hd__nor2b_4
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0899_ Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1378_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[372\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[373\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit17 net237 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[337\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit28 net249 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[348\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[27\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[3\] Tile_X0Y1_N2BEGb\[7\] net4 net12 Tile_X0Y0_DSP_top/ConfigBits\[302\]
+ Tile_X0Y0_DSP_top/ConfigBits\[303\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[314\] Tile_X0Y0_DSP_top/ConfigBits\[315\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top_strobe_inbuf_4__0_ Tile_X0Y1_FrameStrobe_O\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_4__0_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_W1BEG1 net763 Tile_X0Y1_DSP_bot/J2MID_EFb_BEG\[0\]
+ Tile_X0Y1_DSP_bot/JS2BEG\[0\] Tile_X0Y1_DSP_bot/J_l_EF_BEG\[2\] Tile_X0Y1_DSP_bot/ConfigBits\[92\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[93\] VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit5 net256 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[197\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit4 net75 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[378\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1305_ Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1306_/B sky130_fd_sc_hd__nand4_1
XFILLER_0_149_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1236_ Tile_X0Y1_DSP_bot_Inst_MULADD__1233_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1234_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1235_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1236_/Y
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1167_ Tile_X0Y1_DSP_bot_Inst_MULADD__1167_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1167_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1683_/B sky130_fd_sc_hd__xor2_2
XTile_X0Y0_DSP_top_NN4BEG_outbuf_8__0_ ANTENNA_79/DIODE VGND VGND VPWR VPWR net532
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1098_ Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/A Tile_X0Y1_DSP_bot/A4
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/Y sky130_fd_sc_hd__nor2b_4
XFILLER_0_117_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit10 net50 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[192\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[0\] Tile_X0Y0_S2BEGb\[0\] net334 net336 Tile_X0Y1_DSP_bot/ConfigBits\[284\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[285\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit21 net62 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[203\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_NN4BEG_outbuf_1__0_ Tile_X0Y1_DSP_bot/NN4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y1_NN4BEG\[1\] sky130_fd_sc_hd__buf_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_SS4END_inbuf_3__0_ Tile_X0Y0_SS4BEG\[7\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/SS4BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG0 net300
+ net200 Tile_X0Y0_S2BEG\[7\] net353 Tile_X0Y1_DSP_bot/ConfigBits\[208\] Tile_X0Y1_DSP_bot/ConfigBits\[209\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_EFb_BEG\[0\] sky130_fd_sc_hd__mux4_2
XFILLER_0_88_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__90_ Tile_X0Y1_DSP_bot/Q14 VGND VGND
+ VPWR VPWR Tile_X0Y1_bot2top\[4\] sky130_fd_sc_hd__buf_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1021_ Tile_X0Y1_DSP_bot_Inst_MULADD__0968_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0969_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/B sky130_fd_sc_hd__o211ai_4
XFILLER_0_146_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[100\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_SS4BEG_outbuf_4__0_ Tile_X0Y1_DSP_bot/SS4BEG_i\[4\] VGND VGND VPWR
+ VPWR net709 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit16 net236 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[368\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit27 net248 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[379\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit25 net66 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[111\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit14 net54 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[100\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[278\] Tile_X0Y0_DSP_top/ConfigBits\[279\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[336\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[337\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1219_ Tile_X0Y1_DSP_bot_Inst_MULADD__1196_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1197_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1289_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1289_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1219_/X sky130_fd_sc_hd__o211a_2
XFILLER_0_137_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__11_ net16 VGND VGND VPWR VPWR net397
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput302 Tile_X0Y1_N4END[10] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkbuf_1
Xinput335 Tile_X0Y1_W1END[1] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__buf_4
Xinput324 Tile_X0Y1_NN4END[1] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkbuf_2
Xinput313 Tile_X0Y1_N4END[6] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_1
Xinput379 Tile_X0Y1_WW4END[7] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_1
Xinput346 Tile_X0Y1_W2MID[0] VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__clkbuf_4
Xinput368 Tile_X0Y1_WW4END[11] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_1
Xinput357 Tile_X0Y1_W6END[1] VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[1\] Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[1\] Tile_X0Y0_DSP_top/J2MID_EFb_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[1\] Tile_X0Y0_DSP_top/ConfigBits\[104\] Tile_X0Y0_DSP_top/ConfigBits\[105\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_6 Tile_X0Y0_S2BEG\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_EE4END_inbuf_2__0_ net225 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/EE4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_NN4BEG_outbuf_10__0_ Tile_X0Y1_DSP_bot/NN4BEG_i\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y1_NN4BEG\[10\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1570_ Tile_X0Y1_DSP_bot_Inst_MULADD__1593_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1593_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1570_/Y sky130_fd_sc_hd__nor2_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[262\] Tile_X0Y1_DSP_bot/ConfigBits\[263\] VGND VGND
+ VPWR VPWR ANTENNA_106/DIODE sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_83_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit31 net73 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[245\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit20 net61 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[234\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_88_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit8 net259 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[296\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_107_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__73_ net341 VGND VGND VPWR VPWR net722
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1004_ Tile_X0Y1_DSP_bot_Inst_MULADD__0953_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1003_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0953_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1006_/B
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_127_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[74\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR Tile_X0Y0_SS4BEG\[12\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1699_ Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1699_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1721_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_94_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput110 Tile_X0Y0_S4END[3] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xinput132 Tile_X0Y0_SS4END[9] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
Xinput121 Tile_X0Y0_SS4END[13] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
Xinput154 Tile_X0Y0_W6END[10] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_1
Xinput143 Tile_X0Y0_W2END[6] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput176 Tile_X0Y0_WW4END[5] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
Xinput165 Tile_X0Y0_WW4END[0] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
Xinput187 Tile_X0Y1_E2END[2] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_4
Xinput198 Tile_X0Y1_E2MID[5] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_strobe_outbuf_10__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_10__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[10\] sky130_fd_sc_hd__buf_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit15 net235 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[399\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit26 net247 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[410\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_160_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit13 net53 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[131\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit24 net65 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[142\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[300\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[301\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput617 net617 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput606 net606 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[1] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG1 net15
+ net95 net147 Tile_X0Y0_DSP_top/JE2BEG\[3\] Tile_X0Y0_DSP_top/ConfigBits\[152\] Tile_X0Y0_DSP_top/ConfigBits\[153\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[1\] sky130_fd_sc_hd__mux4_1
Xoutput628 net628 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput639 net639 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[17] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_WW4END_inbuf_11__0_ net171 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/WW4BEG_i\[11\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1622_ Tile_X0Y1_DSP_bot_Inst_MULADD__1622_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1622_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1699_/B sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1553_ Tile_X0Y1_DSP_bot_Inst_MULADD__1553_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1553_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1554_/C sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1484_ Tile_X0Y1_DSP_bot_Inst_MULADD__1479_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1482_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1483_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1484_/X
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot_E6BEG_outbuf_6__0_ ANTENNA_98/DIODE VGND VGND VPWR VPWR net611
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__56_ Tile_X0Y1_DSP_bot/JS2BEG\[2\] VGND
+ VGND VPWR VPWR net669 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[106\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit0 net229 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[64\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_204 Tile_X0Y0_SS4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_S4END_inbuf_8__0_ net104 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/S4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit30 net72 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[276\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit19 net239 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[307\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[350\] Tile_X0Y0_DSP_top/ConfigBits\[351\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG2 Tile_X0Y1_N2BEG\[5\]
+ net18 net98 net150 Tile_X0Y0_DSP_top/ConfigBits\[194\] Tile_X0Y0_DSP_top/ConfigBits\[195\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[2\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[0\] Tile_X0Y1_N2BEGb\[0\] net1 net5 Tile_X0Y0_DSP_top/ConfigBits\[338\]
+ Tile_X0Y0_DSP_top/ConfigBits\[339\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0984_ Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/B Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0973_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0984_/X sky130_fd_sc_hd__a221o_2
Xoutput403 net403 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput425 net425 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput414 net414 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput469 net469 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[16] sky130_fd_sc_hd__clkbuf_4
Xoutput447 net447 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[25] sky130_fd_sc_hd__buf_2
Xoutput436 net436 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput458 net458 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG0 Tile_X0Y1_N4BEG\[3\]
+ net8 net140 Tile_X0Y0_DSP_top/JN2BEG\[3\] Tile_X0Y0_DSP_top/ConfigBits\[390\] Tile_X0Y0_DSP_top/ConfigBits\[391\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_EF_BEG\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_129_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1605_ Tile_X0Y1_DSP_bot_Inst_MULADD__1605_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1605_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1605_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_129_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit3 net254 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[99\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_EE4BEG_outbuf_11__0_ Tile_X0Y0_DSP_top/EE4BEG_i\[11\] VGND VGND
+ VPWR VPWR net416 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_S4BEG1 net21 net88
+ net109 Tile_X0Y1_bot2top\[1\] Tile_X0Y0_DSP_top/ConfigBits\[66\] Tile_X0Y0_DSP_top/ConfigBits\[67\]
+ VGND VGND VPWR VPWR Tile_X0Y0_S4BEG\[13\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit2 net71 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[280\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1536_ Tile_X0Y1_DSP_bot_Inst_MULADD__1536_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1536_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1541_/B
+ sky130_fd_sc_hd__and3_2
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1467_ Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/Y sky130_fd_sc_hd__nand2_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1398_ Tile_X0Y1_DSP_bot_Inst_MULADD__1398_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1398_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1398_/Y sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[80\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__39_ ANTENNA_106/DIODE VGND VGND VPWR
+ VPWR Tile_X0Y1_N2BEG\[1\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit23 net64 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[173\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit12 net52 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[162\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[262\] Tile_X0Y0_DSP_top/ConfigBits\[263\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_138_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG1 net309
+ Tile_X0Y0_SS4BEG\[2\] net340 Tile_X0Y1_DSP_bot/JE2BEG\[4\] Tile_X0Y1_DSP_bot/ConfigBits\[410\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[411\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_GH_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_S4END_inbuf_8__0_ Tile_X0Y0_S4BEG\[12\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/S4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1321_ Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/C sky130_fd_sc_hd__a31o_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1252_ Tile_X0Y1_DSP_bot_Inst_MULADD__1252_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1614_/S sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_E6BEG_outbuf_2__0_ Tile_X0Y0_DSP_top/E6BEG_i\[2\] VGND VGND VPWR
+ VPWR net406 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1183_ Tile_X0Y1_DSP_bot_Inst_MULADD__1183_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1183_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_129_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_EE4BEG_outbuf_4__0_ Tile_X0Y1_DSP_bot/EE4BEG_i\[4\] VGND VGND VPWR
+ VPWR net625 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__0967_ Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0965_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0966_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/C
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0898_ Tile_X0Y1_DSP_bot_Inst_MULADD__1032_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/A sky130_fd_sc_hd__clkbuf_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1519_ Tile_X0Y1_DSP_bot_Inst_MULADD__1518_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1518_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1605_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1518_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1520_/B sky130_fd_sc_hd__o22a_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit30 net252 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[30\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q4 wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[372\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[373\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit18 net238 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[338\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit29 net250 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[349\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_92_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1
+ net82 net84 net92 net136 Tile_X0Y0_DSP_top/ConfigBits\[302\] Tile_X0Y0_DSP_top/ConfigBits\[303\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[314\] Tile_X0Y0_DSP_top/ConfigBits\[315\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG0 net199
+ Tile_X0Y0_S2BEG\[6\] net352 Tile_X0Y1_DSP_bot/JN2BEG\[4\] Tile_X0Y1_DSP_bot/ConfigBits\[168\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[169\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG0 Tile_X0Y1_NN4BEG\[3\]
+ net11 net91 net143 Tile_X0Y0_DSP_top/ConfigBits\[222\] Tile_X0Y0_DSP_top/ConfigBits\[223\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_CD_BEG\[0\] sky130_fd_sc_hd__mux4_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_W1BEG2 Tile_X0Y1_DSP_bot/Q7
+ Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[1\] Tile_X0Y1_DSP_bot/JS2BEG\[1\] Tile_X0Y1_DSP_bot/J_l_GH_BEG\[3\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[94\] Tile_X0Y1_DSP_bot/ConfigBits\[95\] VGND VGND
+ VPWR VPWR net717 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit6 net257 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[198\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_data_inbuf_10__0_ net50 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_10__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit5 net76 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[379\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1304_ Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1306_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_149_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1235_ Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1183_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1235_/Y
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1166_ Tile_X0Y1_DSP_bot_Inst_MULADD__1166_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1166_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1167_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1097_ Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1730_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1097_/X sky130_fd_sc_hd__and2_2
XFILLER_0_62_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit11 net51 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[193\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 net764 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[284\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[285\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit22 net63 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[204\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG1 net296
+ net196 Tile_X0Y0_S2BEG\[3\] net349 Tile_X0Y1_DSP_bot/ConfigBits\[210\] Tile_X0Y1_DSP_bot/ConfigBits\[211\]
+ VGND VGND VPWR VPWR ANTENNA_105/DIODE sky130_fd_sc_hd__mux4_2
XFILLER_0_88_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1020_ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1019_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0875_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/A sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_139_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_21_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_inbuf_1__0_ net60 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_1__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit28 net249 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[380\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit17 net237 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[369\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit15 net55 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[101\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit26 net67 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[112\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_inst_clk_buf net333 VGND VGND VPWR VPWR Tile_X0Y1_UserCLKo sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_data_inbuf_10__0_ net230 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_10__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[280\] Tile_X0Y0_DSP_top/ConfigBits\[281\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JE2BEG\[0\] sky130_fd_sc_hd__mux4_2
XFILLER_0_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1218_ Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1218_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1218_/Y sky130_fd_sc_hd__nand2_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1149_ Tile_X0Y1_DSP_bot_Inst_MULADD__1026_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1062_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1149_/Y sky130_fd_sc_hd__o211ai_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[336\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[337\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__10_ net15 VGND VGND VPWR VPWR net396
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_strobe_outbuf_18__0_ Tile_X0Y0_DSP_top_strobe_inbuf_18__0_/X VGND
+ VGND VPWR VPWR net471 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput303 Tile_X0Y1_N4END[11] VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkbuf_1
Xinput336 Tile_X0Y1_W1END[2] VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__buf_4
Xinput325 Tile_X0Y1_NN4END[2] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_2
Xinput314 Tile_X0Y1_N4END[7] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__buf_2
Xinput347 Tile_X0Y1_W2MID[1] VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__buf_2
Xinput369 Tile_X0Y1_WW4END[12] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkbuf_1
Xinput358 Tile_X0Y1_W6END[2] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_data_outbuf_8__0_ Tile_X0Y0_DSP_top_data_inbuf_8__0_/X VGND VGND
+ VPWR VPWR net460 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[106\] Tile_X0Y0_DSP_top/ConfigBits\[107\] VGND VGND
+ VPWR VPWR net556 sky130_fd_sc_hd__mux4_1
XFILLER_0_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_7 Tile_X0Y0_SS4BEG\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit10 net50 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[224\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit21 net62 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[235\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit9 net260 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[297\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__72_ Tile_X0Y1_DSP_bot/JW2BEG\[2\] VGND
+ VGND VPWR VPWR net721 sky130_fd_sc_hd__buf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1003_ Tile_X0Y1_DSP_bot_Inst_MULADD__1252_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0922_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0950_/B Tile_X0Y1_DSP_bot_Inst_MULADD__0950_/C Tile_X0Y1_DSP_bot_Inst_MULADD__0923_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1003_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[74\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_SS4END_inbuf_10__0_ Tile_X0Y0_SS4BEG\[14\] VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot/SS4BEG_i\[10\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit0 net49 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[182\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1698_ Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1698_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1698_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1720_/D
+ sky130_fd_sc_hd__nor3_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_NN4END_inbuf_3__0_ net330 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/NN4BEG_i\[3\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_N4BEG_outbuf_6__0_ Tile_X0Y0_DSP_top/N4BEG_i\[6\] VGND VGND VPWR
+ VPWR net514 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput111 Tile_X0Y0_S4END[4] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_1
Xinput100 Tile_X0Y0_S2MID[7] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_4
Xinput122 Tile_X0Y0_SS4END[14] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
Xinput144 Tile_X0Y0_W2END[7] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_4
Xinput133 Tile_X0Y0_W1END[0] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__buf_4
Xinput155 Tile_X0Y0_W6END[11] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_1
Xinput166 Tile_X0Y0_WW4END[10] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_1
Xinput177 Tile_X0Y0_WW4END[6] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
Xinput199 Tile_X0Y1_E2MID[6] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_4
Xinput188 Tile_X0Y1_E2END[3] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit16 net236 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[400\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit27 net248 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[411\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_data_outbuf_8__0_ Tile_X0Y1_DSP_bot_data_inbuf_8__0_/X VGND VGND
+ VPWR VPWR net661 sky130_fd_sc_hd__clkbuf_1
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit25 net66 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[143\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit14 net54 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[132\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[302\] Tile_X0Y1_DSP_bot/ConfigBits\[303\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JE2BEG\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_81_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput618 net618 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput607 net607 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[2] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG2 Tile_X0Y1_N2BEG\[4\]
+ net17 net149 Tile_X0Y0_DSP_top/JS2BEG\[3\] Tile_X0Y0_DSP_top/ConfigBits\[154\] Tile_X0Y0_DSP_top/ConfigBits\[155\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[2\] sky130_fd_sc_hd__mux4_2
Xoutput629 net629 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[8] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1621_ Tile_X0Y1_DSP_bot_Inst_MULADD__1619_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1698_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1622_/B sky130_fd_sc_hd__a2bb2oi_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1552_ Tile_X0Y1_DSP_bot_Inst_MULADD__1718_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1614_/S
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1553_/B sky130_fd_sc_hd__and2b_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1483_ Tile_X0Y1_DSP_bot_Inst_MULADD__1089_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1091_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1483_/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__55_ Tile_X0Y1_DSP_bot/JS2BEG\[1\] VGND
+ VGND VPWR VPWR net668 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit1 net240 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[65\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_216 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_W6BEG_outbuf_6__0_ ANTENNA_96/DIODE VGND VGND VPWR VPWR net563
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit20 net61 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[266\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit31 net73 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[277\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[352\] Tile_X0Y0_DSP_top/ConfigBits\[353\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JW2BEG\[2\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0
+ net284 net286 net186 net204 Tile_X0Y1_DSP_bot/ConfigBits\[352\] Tile_X0Y1_DSP_bot/ConfigBits\[353\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG3 Tile_X0Y1_N2BEG\[1\]
+ net14 net94 net146 Tile_X0Y0_DSP_top/ConfigBits\[196\] Tile_X0Y0_DSP_top/ConfigBits\[197\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[3\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1
+ net81 net85 net133 net135 Tile_X0Y0_DSP_top/ConfigBits\[338\] Tile_X0Y0_DSP_top/ConfigBits\[339\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0983_ Tile_X0Y1_DSP_bot_Inst_MULADD__0983_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/A sky130_fd_sc_hd__clkbuf_4
Xoutput404 net404 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[11] sky130_fd_sc_hd__buf_2
Xoutput415 net415 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput426 net426 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput448 net448 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[26] sky130_fd_sc_hd__clkbuf_4
Xoutput437 net437 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[16] sky130_fd_sc_hd__clkbuf_4
Xoutput459 net459 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_10_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG1 Tile_X0Y1_NN4BEG\[2\]
+ net7 net109 Tile_X0Y0_DSP_top/JE2BEG\[3\] Tile_X0Y0_DSP_top/ConfigBits\[392\] Tile_X0Y0_DSP_top/ConfigBits\[393\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_EF_BEG\[1\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1604_ Tile_X0Y1_DSP_bot_Inst_MULADD__1604_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1604_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1604_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit4 net255 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[100\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_S4BEG2 net85 net110
+ net156 Tile_X0Y1_bot2top\[2\] Tile_X0Y0_DSP_top/ConfigBits\[68\] Tile_X0Y0_DSP_top/ConfigBits\[69\]
+ VGND VGND VPWR VPWR Tile_X0Y0_S4BEG\[14\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit3 net74 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[281\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1535_ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/A sky130_fd_sc_hd__nand4_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1466_ Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1465_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1690_/B
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit0 net49 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[22\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1397_ Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1396_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1397_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[80\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__38_ Tile_X0Y1_DSP_bot/JN2BEG\[0\] VGND
+ VGND VPWR VPWR Tile_X0Y1_N2BEG\[0\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_E6END_inbuf_4__0_ net29 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/E6BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit24 net65 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[174\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit13 net53 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[163\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[262\] Tile_X0Y0_DSP_top/ConfigBits\[263\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG2 net204
+ Tile_X0Y0_S4BEG\[1\] net375 Tile_X0Y1_DSP_bot/JS2BEG\[4\] Tile_X0Y1_DSP_bot/ConfigBits\[412\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[413\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_GH_BEG\[2\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_strobe_inbuf_12__0_ Tile_X0Y1_FrameStrobe_O\[12\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_12__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_outbuf_26__0_ Tile_X0Y0_DSP_top_data_inbuf_26__0_/X VGND VGND
+ VPWR VPWR net448 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1320_ Tile_X0Y1_DSP_bot_Inst_MULADD__1314_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1318_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1220_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1236_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1319_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/B sky130_fd_sc_hd__o221ai_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1251_ Tile_X0Y1_DSP_bot/C7 Tile_X0Y1_DSP_bot_Inst_MULADD__1749_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1459_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1251_/X
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1182_ Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1180_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1181_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1183_/A sky130_fd_sc_hd__o22ai_4
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0966_ Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1730_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0966_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0897_ Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0885_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0886_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1032_/B
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y0_DSP_top_data_outbuf_17__0_ Tile_X0Y0_DSP_top_data_inbuf_17__0_/X VGND VGND
+ VPWR VPWR net438 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1518_ Tile_X0Y1_DSP_bot_Inst_MULADD__1518_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1518_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1605_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1518_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1520_/A sky130_fd_sc_hd__nor4_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit20 net241 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[20\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit31 net253 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[31\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1449_ Tile_X0Y1_DSP_bot_Inst_MULADD__1452_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/Y
+ sky130_fd_sc_hd__nand3b_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[374\] Tile_X0Y1_DSP_bot/ConfigBits\[375\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JW2BEG\[5\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit30 net72 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[308\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_S4BEG_outbuf_6__0_ ANTENNA_91/DIODE VGND VGND VPWR VPWR Tile_X0Y0_S4BEG\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit19 net239 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[339\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_81_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[302\] Tile_X0Y0_DSP_top/ConfigBits\[303\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_E6END_inbuf_4__0_ net209 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/E6BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[316\] Tile_X0Y0_DSP_top/ConfigBits\[317\] VGND VGND
+ VPWR VPWR ANTENNA_63/DIODE sky130_fd_sc_hd__mux4_2
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG1 net295
+ net195 net348 Tile_X0Y1_DSP_bot/JE2BEG\[4\] Tile_X0Y1_DSP_bot/ConfigBits\[170\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[171\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG1 Tile_X0Y1_N2BEGb\[2\]
+ net7 net87 net173 Tile_X0Y0_DSP_top/ConfigBits\[224\] Tile_X0Y0_DSP_top/ConfigBits\[225\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_CD_BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_W1BEG3 Tile_X0Y1_DSP_bot/Q0
+ Tile_X0Y1_DSP_bot/J2MID_ABb_BEG\[2\] Tile_X0Y1_DSP_bot/JS2BEG\[2\] Tile_X0Y1_DSP_bot/J_l_AB_BEG\[0\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[96\] Tile_X0Y1_DSP_bot/ConfigBits\[97\] VGND VGND
+ VPWR VPWR net718 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit7 net258 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[199\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit6 net77 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[380\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_126_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1303_ Tile_X0Y1_DSP_bot_Inst_MULADD__0887_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1128_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1211_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1201_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/C sky130_fd_sc_hd__o221ai_4
XFILLER_0_149_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1234_ Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1215_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1117_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1234_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_59_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1165_ Tile_X0Y1_DSP_bot_Inst_MULADD__1165_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1165_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1165_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1166_/B
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_157_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_EE4END_inbuf_10__0_ net218 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/EE4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1096_ Tile_X0Y1_DSP_bot_Inst_MULADD__0854_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0854_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1093_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1095_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1096_/Y sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit23 net64 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[205\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[284\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[285\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit12 net52 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[194\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0949_ Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0950_/C
+ sky130_fd_sc_hd__and3_1
XFILLER_0_65_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_data_inbuf_7__0_ net258 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_7__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG0 net326
+ Tile_X0Y0_S4BEG\[3\] net366 ANTENNA_106/DIODE Tile_X0Y1_DSP_bot/ConfigBits\[384\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[385\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_AB_BEG\[0\]
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_strobe_outbuf_3__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_3__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[3\] sky130_fd_sc_hd__buf_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG2 net298
+ net198 Tile_X0Y0_S2BEG\[5\] net351 Tile_X0Y1_DSP_bot/ConfigBits\[212\] Tile_X0Y1_DSP_bot/ConfigBits\[213\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_EFb_BEG\[2\] sky130_fd_sc_hd__mux4_1
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit30 net252 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[62\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_141_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_WW4BEG_outbuf_8__0_ Tile_X0Y0_DSP_top/WW4BEG_i\[8\] VGND VGND VPWR
+ VPWR net581 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit29 net250 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[381\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit18 net238 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[370\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit16 net56 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[102\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit27 net68 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[113\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_79_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1217_ Tile_X0Y1_DSP_bot_Inst_MULADD__1207_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1213_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1216_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1217_/Y
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1148_ Tile_X0Y1_DSP_bot_Inst_MULADD__1140_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1140_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1131_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1135_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1148_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[338\] Tile_X0Y1_DSP_bot/ConfigBits\[339\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JS2BEG\[4\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1079_ Tile_X0Y1_DSP_bot_Inst_MULADD__1026_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1044_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1048_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1049_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1079_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_0_132_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst0
+ net284 Tile_X0Y0_S1BEG\[3\] net337 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[101\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[102\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
Xinput326 Tile_X0Y1_NN4END[3] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_2
Xinput315 Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_1
Xinput304 Tile_X0Y1_N4END[12] VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_WW4BEG_outbuf_1__0_ Tile_X0Y1_DSP_bot/WW4BEG_i\[1\] VGND VGND VPWR
+ VPWR net754 sky130_fd_sc_hd__clkbuf_1
Xinput348 Tile_X0Y1_W2MID[2] VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__clkbuf_4
Xinput337 Tile_X0Y1_W1END[3] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__buf_4
Xinput359 Tile_X0Y1_W6END[3] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_strobe_inbuf_18__0_ net270 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_18__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_8 Tile_X0Y0_SS4BEG\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit11 net51 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[225\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit22 net63 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[236\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_107_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_N4END_inbuf_8__0_ Tile_X0Y1_N4BEG\[12\] VGND VGND VPWR VPWR ANTENNA_180/DIODE
+ sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__71_ Tile_X0Y1_DSP_bot/JW2BEG\[1\] VGND
+ VGND VPWR VPWR net720 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1002_ Tile_X0Y1_DSP_bot_Inst_MULADD__1002_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1002_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1002_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1006_/A
+ sky130_fd_sc_hd__and3_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit1 net60 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[183\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1697_ Tile_X0Y1_DSP_bot_Inst_MULADD__1697_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1719_/D sky130_fd_sc_hd__clkbuf_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput101 Tile_X0Y0_S4END[0] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_2
XFILLER_0_101_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput112 Tile_X0Y0_S4END[5] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
Xinput123 Tile_X0Y0_SS4END[15] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xinput145 Tile_X0Y0_W2MID[0] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_2
Xinput134 Tile_X0Y0_W1END[1] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_4
Xinput156 Tile_X0Y0_W6END[1] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_4
Xinput167 Tile_X0Y0_WW4END[11] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_1
Xinput178 Tile_X0Y0_WW4END[7] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput189 Tile_X0Y1_E2END[4] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit17 net237 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[401\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit28 net249 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[412\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit26 net67 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[144\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit15 net55 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[133\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_WW4END_inbuf_4__0_ net380 VGND VGND VPWR VPWR ANTENNA_113/DIODE
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput608 net608 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput619 net619 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[13] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG3 Tile_X0Y1_N2BEG\[0\]
+ net13 net93 Tile_X0Y0_DSP_top/JW2BEG\[3\] Tile_X0Y0_DSP_top/ConfigBits\[156\] Tile_X0Y0_DSP_top/ConfigBits\[157\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[3\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1620_ Tile_X0Y1_DSP_bot_Inst_MULADD__1620_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1620_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1698_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1551_ Tile_X0Y1_DSP_bot_Inst_MULADD__1614_/S Tile_X0Y1_DSP_bot_Inst_MULADD__1551_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1553_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1482_ Tile_X0Y1_DSP_bot_Inst_MULADD__0926_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0958_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1480_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1482_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_89_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__54_ Tile_X0Y1_DSP_bot/JS2BEG\[0\] VGND
+ VGND VPWR VPWR net667 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_N4END_inbuf_8__0_ net304 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/N4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_cus_mux41_buf_inst0
+ Tile_X0Y1_DSP_bot/JN2BEG\[5\] ANTENNA_183/DIODE Tile_X0Y1_DSP_bot/JE2BEG\[5\] Tile_X0Y1_DSP_bot/JE2BEG\[7\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[153\] Tile_X0Y1_DSP_bot/ConfigBits\[154\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_SS4BEG_outbuf_1__0_ ANTENNA_94/DIODE VGND VGND VPWR VPWR Tile_X0Y0_SS4BEG\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit2 net251 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[66\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_110_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1749_ net333 Tile_X0Y1_DSP_bot/C7 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1749_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_206 ANTENNA_206/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_217 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit10 net50 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[256\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit21 net62 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[267\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1
+ Tile_X0Y0_S2BEGb\[1\] Tile_X0Y0_S4BEG\[1\] net339 net357 Tile_X0Y1_DSP_bot/ConfigBits\[352\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[353\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[338\] Tile_X0Y0_DSP_top/ConfigBits\[339\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__0982_ Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/C Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0983_/A sky130_fd_sc_hd__or4_1
Xoutput405 net405 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput416 net416 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput449 net449 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[27] sky130_fd_sc_hd__clkbuf_4
Xoutput438 net438 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[17] sky130_fd_sc_hd__clkbuf_4
Xoutput427 net427 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[7] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG2 Tile_X0Y1_N4BEG\[1\]
+ net124 net141 Tile_X0Y0_DSP_top/JS2BEG\[3\] Tile_X0Y0_DSP_top/ConfigBits\[394\]
+ Tile_X0Y0_DSP_top/ConfigBits\[395\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_EF_BEG\[2\]
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1603_ Tile_X0Y1_DSP_bot_Inst_MULADD__1560_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1553_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1553_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1579_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1629_/D sky130_fd_sc_hd__o41ai_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit5 net256 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[101\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit4 net75 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[282\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_S4BEG3 net86 net101
+ net153 Tile_X0Y1_bot2top\[3\] Tile_X0Y0_DSP_top/ConfigBits\[70\] Tile_X0Y0_DSP_top/ConfigBits\[71\]
+ VGND VGND VPWR VPWR Tile_X0Y0_S4BEG\[15\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1534_ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1536_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1465_ Tile_X0Y1_DSP_bot_Inst_MULADD__1465_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1465_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1604_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1465_/Y
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_145_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit1 net60 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[23\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1396_ Tile_X0Y1_DSP_bot_Inst_MULADD__1421_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1421_/C
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1396_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_159_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_147_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__37_ net200 VGND VGND VPWR VPWR net602
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit14 net54 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[164\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit25 net66 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[175\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[264\] Tile_X0Y0_DSP_top/ConfigBits\[265\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JN2BEG\[4\] sky130_fd_sc_hd__mux4_2
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG3 net317
+ net201 net338 Tile_X0Y1_DSP_bot/JW2BEG\[4\] Tile_X0Y1_DSP_bot/ConfigBits\[414\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[415\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_GH_BEG\[3\]
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0
+ net288 net310 net182 net188 Tile_X0Y1_DSP_bot/ConfigBits\[264\] Tile_X0Y1_DSP_bot/ConfigBits\[265\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_WW4END_inbuf_0__0_ net175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/WW4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1250_ Tile_X0Y1_DSP_bot_Inst_MULADD__1171_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1246_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1249_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1339_/A
+ sky130_fd_sc_hd__o21a_1
XTile_X0Y0_DSP_top_strobe_inbuf_7__0_ Tile_X0Y1_FrameStrobe_O\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_7__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1181_ Tile_X0Y1_DSP_bot_Inst_MULADD__1128_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1113_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1172_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1181_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_115_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0965_ Tile_X0Y1_DSP_bot/A4 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0965_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_112_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0896_ Tile_X0Y1_DSP_bot/A0 Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0849_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0896_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1517_ Tile_X0Y1_DSP_bot_Inst_MULADD__1523_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1523_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1523_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1518_/D
+ sky130_fd_sc_hd__and3_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit10 net230 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[10\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit21 net242 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[21\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_156_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst0
+ net282 net182 Tile_X0Y0_S1BEG\[1\] Tile_X0Y1_DSP_bot/Q5 Tile_X0Y1_DSP_bot/ConfigBits\[51\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[52\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1448_ Tile_X0Y1_DSP_bot_Inst_MULADD__1291_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1318_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1387_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1447_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1448_/Y sky130_fd_sc_hd__a41oi_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit20 net61 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[298\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit31 net73 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[309\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1379_ Tile_X0Y1_DSP_bot_Inst_MULADD__1379_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1379_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1379_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[302\] Tile_X0Y0_DSP_top/ConfigBits\[303\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG2 Tile_X0Y1_N2BEGb\[4\]
+ net9 net125 net141 Tile_X0Y0_DSP_top/ConfigBits\[226\] Tile_X0Y0_DSP_top/ConfigBits\[227\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_CD_BEG\[2\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG2 net297
+ net197 Tile_X0Y0_S2BEG\[4\] Tile_X0Y1_DSP_bot/JS2BEG\[4\] Tile_X0Y1_DSP_bot/ConfigBits\[172\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[173\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[2\]
+ sky130_fd_sc_hd__mux4_2
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_NN4BEG_outbuf_4__0_ Tile_X0Y1_DSP_bot/NN4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y1_NN4BEG\[4\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_SS4END_inbuf_6__0_ Tile_X0Y0_SS4BEG\[10\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/SS4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit8 net259 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[200\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1302_ Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1300_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1301_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/A
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_126_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit7 net78 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[381\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1233_ Tile_X0Y1_DSP_bot_Inst_MULADD__1231_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1219_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1218_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1233_/Y sky130_fd_sc_hd__o2bb2ai_2
XFILLER_0_149_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1164_ Tile_X0Y1_DSP_bot_Inst_MULADD__1164_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1164_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1165_/C sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot_SS4BEG_outbuf_7__0_ Tile_X0Y1_DSP_bot/SS4BEG_i\[7\] VGND VGND VPWR
+ VPWR net712 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1095_ Tile_X0Y1_DSP_bot_Inst_MULADD__1095_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1095_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit24 net65 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[206\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[286\] Tile_X0Y1_DSP_bot/ConfigBits\[287\] VGND VGND
+ VPWR VPWR ANTENNA_183/DIODE sky130_fd_sc_hd__mux4_2
XFILLER_0_70_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit13 net53 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[195\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0948_ Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/D VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0950_/B
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_140_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0879_ Tile_X0Y1_DSP_bot_Inst_MULADD__0878_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0906_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0878_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0880_/B
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot_S4BEG_outbuf_11__0_ Tile_X0Y1_DSP_bot/S4BEG_i\[11\] VGND VGND VPWR
+ VPWR net685 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG1 net221
+ Tile_X0Y0_S4BEG\[2\] net345 Tile_X0Y1_DSP_bot/JE2BEG\[1\] Tile_X0Y1_DSP_bot/ConfigBits\[386\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[387\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_AB_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG3 net294
+ net194 Tile_X0Y0_S2BEG\[1\] net347 Tile_X0Y1_DSP_bot/ConfigBits\[214\] Tile_X0Y1_DSP_bot/ConfigBits\[215\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_EFb_BEG\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit20 net241 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[52\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_W6END_inbuf_2__0_ net159 VGND VGND VPWR VPWR ANTENNA_95/DIODE sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit31 net253 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[63\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_122_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_EE4END_inbuf_5__0_ net228 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/EE4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit30 net72 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[340\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_122_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit19 net239 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[371\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit28 net69 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[114\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit17 net57 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[103\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1216_ Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1215_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1117_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1216_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1147_ Tile_X0Y1_DSP_bot_Inst_MULADD__1050_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1078_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1135_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1146_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1141_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1147_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_0_157_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1078_ Tile_X0Y1_DSP_bot_Inst_MULADD__1051_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1052_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1078_/Y
+ sky130_fd_sc_hd__a21oi_4
XTile_X0Y0_DSP_top_EE4BEG_outbuf_1__0_ Tile_X0Y0_DSP_top/EE4BEG_i\[1\] VGND VGND VPWR
+ VPWR net421 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[2\] Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2END_EF_BEG\[2\] Tile_X0Y1_DSP_bot/ConfigBits\[101\] Tile_X0Y1_DSP_bot/ConfigBits\[102\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_87_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput327 Tile_X0Y1_NN4END[4] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_1
Xinput316 Tile_X0Y1_N4END[9] VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_1
Xinput305 Tile_X0Y1_N4END[13] VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_1
Xinput338 Tile_X0Y1_W2END[0] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__buf_2
Xinput349 Tile_X0Y1_W2MID[3] VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkbuf_4
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_9 Tile_X0Y0_SS4BEG\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[3\] net4 net136 Tile_X0Y1_bot2top\[3\] Tile_X0Y0_DSP_top/ConfigBits\[19\]
+ Tile_X0Y0_DSP_top/ConfigBits\[20\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_SS4END_inbuf_2__0_ net129 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/SS4BEG_i\[2\]
+ sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit12 net52 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[226\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_107_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit23 net64 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[237\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_strobe_outbuf_13__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_13__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[13\] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__70_ net338 VGND VGND VPWR VPWR net719
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1001_ Tile_X0Y1_DSP_bot_Inst_MULADD__1001_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1006_/C sky130_fd_sc_hd__inv_2
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_W6END_inbuf_2__0_ net360 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/W6BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit2 net71 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[184\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1696_ Tile_X0Y1_DSP_bot_Inst_MULADD__1674_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1696_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1697_/A sky130_fd_sc_hd__and2b_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_E6BEG_outbuf_9__0_ Tile_X0Y1_DSP_bot/E6BEG_i\[9\] VGND VGND VPWR
+ VPWR net614 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput102 Tile_X0Y0_S4END[10] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput124 Tile_X0Y0_SS4END[1] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__buf_2
Xinput113 Tile_X0Y0_S4END[6] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
Xinput135 Tile_X0Y0_W1END[2] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_4
Xinput157 Tile_X0Y0_W6END[2] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
Xinput168 Tile_X0Y0_WW4END[12] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
Xinput146 Tile_X0Y0_W2MID[1] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_2
Xinput179 Tile_X0Y0_WW4END[8] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit30 net252 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[94\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit0 net229 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[320\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit29 net250 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[413\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit18 net238 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[402\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit27 net68 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[145\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit16 net56 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[134\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput609 net609 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_0_111_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_EE4END_inbuf_1__0_ net44 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/EE4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1550_ Tile_X0Y1_DSP_bot/C12 Tile_X0Y1_DSP_bot_Inst_MULADD__1754_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1551_/B
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1481_ Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1733_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/X sky130_fd_sc_hd__and2_1
XFILLER_0_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__53_ net300 VGND VGND VPWR VPWR Tile_X0Y1_N2BEGb\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit3 net254 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[67\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/JS2BEG\[5\] Tile_X0Y1_DSP_bot/JS2BEG\[7\] Tile_X0Y1_DSP_bot/JW2BEG\[5\]
+ Tile_X0Y1_DSP_bot/JW2BEG\[7\] Tile_X0Y1_DSP_bot/ConfigBits\[153\] Tile_X0Y1_DSP_bot/ConfigBits\[154\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_N4BEG_outbuf_0__0_ Tile_X0Y1_DSP_bot/N4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N4BEG\[0\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1748_ net333 Tile_X0Y1_DSP_bot/C6 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1748_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1679_ Tile_X0Y1_DSP_bot_Inst_MULADD__1674_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1679_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1680_/A sky130_fd_sc_hd__and2b_1
XANTENNA_207 ANTENNA_207/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_218 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit11 net51 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[257\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_121_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit22 net63 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[268\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2
+ net764 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[352\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[353\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[338\] Tile_X0Y0_DSP_top/ConfigBits\[339\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0981_ Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/A Tile_X0Y1_DSP_bot/B4
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1299_/D VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/D
+ sky130_fd_sc_hd__o21ai_4
Xoutput406 net406 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[2] sky130_fd_sc_hd__buf_2
Xoutput417 net417 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[12] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot0 Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[0\]
+ Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[0\] Tile_X0Y0_DSP_top/J2END_AB_BEG\[0\] ANTENNA_65/DIODE
+ Tile_X0Y0_DSP_top/ConfigBits\[112\] Tile_X0Y0_DSP_top/ConfigBits\[113\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_124_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[0\] Tile_X0Y1_N2BEGb\[2\] Tile_X0Y1_N4BEG\[2\] net7 Tile_X0Y0_DSP_top/ConfigBits\[282\]
+ Tile_X0Y0_DSP_top/ConfigBits\[283\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
Xoutput439 net439 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput428 net428 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG3 net42
+ net101 net172 Tile_X0Y0_DSP_top/JW2BEG\[3\] Tile_X0Y0_DSP_top/ConfigBits\[396\]
+ Tile_X0Y0_DSP_top/ConfigBits\[397\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_EF_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1602_ Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/X
+ sky130_fd_sc_hd__and3_1
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1533_ Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/D sky130_fd_sc_hd__nand4_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit6 net257 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[102\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit5 net76 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[283\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1464_ Tile_X0Y1_DSP_bot_Inst_MULADD__1471_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1471_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1471_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1604_/A
+ sky130_fd_sc_hd__nand3_2
XTile_X0Y0_DSP_top_E6BEG_outbuf_5__0_ Tile_X0Y0_DSP_top/E6BEG_i\[5\] VGND VGND VPWR
+ VPWR net409 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1395_ Tile_X0Y1_DSP_bot_Inst_MULADD__1421_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1421_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1395_/Y
+ sky130_fd_sc_hd__a21boi_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit2 net71 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[24\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_EE4BEG_outbuf_7__0_ Tile_X0Y1_DSP_bot/EE4BEG_i\[7\] VGND VGND VPWR
+ VPWR net628 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__36_ net199 VGND VGND VPWR VPWR net601
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_W6BEG_outbuf_0__0_ Tile_X0Y1_DSP_bot/W6BEG_i\[0\] VGND VGND VPWR
+ VPWR net735 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_inbuf_31__0_ net73 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_31__0_/X
+ sky130_fd_sc_hd__buf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0
+ net3 net135 Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y0_DSP_top/ConfigBits\[108\]
+ Tile_X0Y0_DSP_top/ConfigBits\[109\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit15 net55 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[165\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit26 net67 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[176\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1
+ net204 Tile_X0Y0_S2BEGb\[3\] net341 net373 Tile_X0Y1_DSP_bot/ConfigBits\[264\] Tile_X0Y1_DSP_bot/ConfigBits\[265\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_data_inbuf_22__0_ net63 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_22__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1180_ Tile_X0Y1_DSP_bot_Inst_MULADD__1034_/X Tile_X0Y1_DSP_bot/B7
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1175_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1180_/Y
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_86_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__0964_ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1201_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0963_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0875_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/B sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0895_ Tile_X0Y1_DSP_bot_Inst_MULADD__0895_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/A sky130_fd_sc_hd__buf_4
XFILLER_0_57_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_data_inbuf_13__0_ net53 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_13__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1516_ Tile_X0Y1_DSP_bot_Inst_MULADD__1523_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1523_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1523_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1605_/B
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit11 net231 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[11\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit22 net243 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[22\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_156_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1447_ Tile_X0Y1_DSP_bot_Inst_MULADD__1386_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1386_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1366_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1370_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1390_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1447_/Y sky130_fd_sc_hd__o221ai_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[2\] Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2END_AB_BEG\[0\] Tile_X0Y1_DSP_bot/ConfigBits\[51\] Tile_X0Y1_DSP_bot/ConfigBits\[52\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit21 net62 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[299\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit10 net50 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[288\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1378_ Tile_X0Y1_DSP_bot_Inst_MULADD__1378_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1379_/B sky130_fd_sc_hd__nand4_1
XFILLER_0_77_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__19_ Tile_X0Y0_top2bot\[15\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[304\] Tile_X0Y0_DSP_top/ConfigBits\[305\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JE2BEG\[6\] sky130_fd_sc_hd__mux4_2
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0
+ net282 net290 net182 net190 Tile_X0Y1_DSP_bot/ConfigBits\[304\] Tile_X0Y1_DSP_bot/ConfigBits\[305\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_data_inbuf_31__0_ net253 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_31__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG3 Tile_X0Y1_N2BEGb\[0\]
+ net40 net85 net137 Tile_X0Y0_DSP_top/ConfigBits\[228\] Tile_X0Y0_DSP_top/ConfigBits\[229\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_CD_BEG\[3\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG3 net293
+ Tile_X0Y0_S2BEG\[0\] net346 Tile_X0Y1_DSP_bot/JW2BEG\[4\] Tile_X0Y1_DSP_bot/ConfigBits\[174\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[175\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_data_outbuf_20__0_ Tile_X0Y1_DSP_bot_data_inbuf_20__0_/X VGND VGND
+ VPWR VPWR net643 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit9 net260 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[201\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1301_ Tile_X0Y1_DSP_bot_Inst_MULADD__1034_/X Tile_X0Y1_DSP_bot/B6
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1378_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1121_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1301_/X sky130_fd_sc_hd__o211a_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit8 net79 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[382\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_data_inbuf_22__0_ net243 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_22__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1232_ Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1163_ Tile_X0Y1_DSP_bot_Inst_MULADD__1165_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1165_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1164_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1164_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1166_/A sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y1_DSP_bot_data_outbuf_11__0_ Tile_X0Y1_DSP_bot_data_inbuf_11__0_/X VGND VGND
+ VPWR VPWR net633 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1094_ Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1732_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1095_/A sky130_fd_sc_hd__and2_1
XFILLER_0_144_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_data_inbuf_4__0_ net75 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_4__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit25 net66 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[207\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_125_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit14 net54 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[196\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_S4BEG_outbuf_0__0_ Tile_X0Y1_DSP_bot/S4BEG_i\[0\] VGND VGND VPWR
+ VPWR net683 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit0 net49 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[86\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0947_ Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0946_/C Tile_X0Y1_DSP_bot_Inst_MULADD__0946_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/B sky130_fd_sc_hd__a22o_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0878_ Tile_X0Y1_DSP_bot_Inst_MULADD__0878_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0906_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0878_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0880_/A
+ sky130_fd_sc_hd__and3_1
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_data_inbuf_13__0_ net233 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_13__0_/X
+ sky130_fd_sc_hd__buf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[2\] Tile_X0Y1_N2BEGb\[4\] net9 net21 Tile_X0Y0_DSP_top/ConfigBits\[354\]
+ Tile_X0Y0_DSP_top/ConfigBits\[355\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG2 net308
+ net204 net357 Tile_X0Y1_DSP_bot/JS2BEG\[1\] Tile_X0Y1_DSP_bot/ConfigBits\[388\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[389\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_AB_BEG\[2\]
+ sky130_fd_sc_hd__mux4_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit10 net230 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[42\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit21 net242 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[53\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_NN4END_inbuf_10__0_ net322 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/NN4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_122_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit20 net61 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[330\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit31 net73 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[341\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG0 net292
+ net221 Tile_X0Y0_S2BEGb\[7\] net345 Tile_X0Y1_DSP_bot/ConfigBits\[240\] Tile_X0Y1_DSP_bot/ConfigBits\[241\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_EF_BEG\[0\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit18 net58 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[104\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit29 net70 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[115\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1215_ Tile_X0Y1_DSP_bot_Inst_MULADD__1054_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1103_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1215_/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1146_ Tile_X0Y1_DSP_bot_Inst_MULADD__1131_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1146_/Y sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_157_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1077_ Tile_X0Y1_DSP_bot_Inst_MULADD__1074_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1073_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1073_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1167_/A
+ sky130_fd_sc_hd__o21bai_4
XFILLER_0_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput317 Tile_X0Y1_NN4END[0] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__buf_1
Xinput306 Tile_X0Y1_N4END[14] VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_1
Xinput339 Tile_X0Y1_W2END[1] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_NN4END_inbuf_6__0_ net318 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/NN4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
Xinput328 Tile_X0Y1_NN4END[5] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_N4BEG_outbuf_9__0_ Tile_X0Y0_DSP_top/N4BEG_i\[9\] VGND VGND VPWR
+ VPWR net517 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[7\] Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[2\] Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2END_EF_BEG\[1\] Tile_X0Y0_DSP_top/ConfigBits\[19\] Tile_X0Y0_DSP_top/ConfigBits\[20\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit13 net53 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[227\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit24 net65 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[238\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1000_ Tile_X0Y1_DSP_bot_Inst_MULADD__1002_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1002_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1002_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1001_/A
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[1\] net82 net134 Tile_X0Y1_bot2top\[5\] Tile_X0Y0_DSP_top/ConfigBits\[101\]
+ Tile_X0Y0_DSP_top/ConfigBits\[102\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0
+ net284 net292 net184 net192 Tile_X0Y1_DSP_bot/ConfigBits\[376\] Tile_X0Y1_DSP_bot/ConfigBits\[377\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit3 net74 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[185\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1695_ Tile_X0Y1_DSP_bot_Inst_MULADD__1695_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1129_ Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1043_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_118_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0
+ Tile_X0Y1_NN4BEG\[3\] net2 net8 net24 Tile_X0Y0_DSP_top/ConfigBits\[318\] Tile_X0Y0_DSP_top/ConfigBits\[319\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput125 Tile_X0Y0_SS4END[2] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_2
Xinput103 Tile_X0Y0_S4END[11] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
Xinput114 Tile_X0Y0_S4END[7] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
Xinput136 Tile_X0Y0_W1END[3] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_4
Xinput158 Tile_X0Y0_W6END[3] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
Xinput169 Tile_X0Y0_WW4END[13] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
Xinput147 Tile_X0Y0_W2MID[2] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit31 net253 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[95\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit20 net241 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[84\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_W6BEG_outbuf_9__0_ Tile_X0Y0_DSP_top/W6BEG_i\[9\] VGND VGND VPWR
+ VPWR net566 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit1 net240 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[321\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit30 net72 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[372\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit19 net239 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[403\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit28 net69 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[146\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit17 net57 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[135\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1480_ Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/A Tile_X0Y1_DSP_bot/A7
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1480_/X sky130_fd_sc_hd__and2b_1
XTile_X0Y0_DSP_top_strobe_outbuf_0__0_ Tile_X0Y0_DSP_top_strobe_inbuf_0__0_/X VGND
+ VGND VPWR VPWR net462 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__52_ net299 VGND VGND VPWR VPWR Tile_X0Y1_N2BEGb\[6\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit4 net255 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[68\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1747_ net333 Tile_X0Y1_DSP_bot/C5 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1747_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1678_ Tile_X0Y1_DSP_bot_Inst_MULADD__1678_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1709_/D sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_NN4END_inbuf_2__0_ Tile_X0Y1_NN4BEG\[6\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/NN4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA_219 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_208 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit23 net64 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[269\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit12 net52 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[258\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_E6END_inbuf_7__0_ net32 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/E6BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[352\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[353\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_strobe_inbuf_15__0_ Tile_X0Y1_FrameStrobe_O\[15\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_15__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[340\] Tile_X0Y0_DSP_top/ConfigBits\[341\] VGND VGND
+ VPWR VPWR ANTENNA_179/DIODE sky130_fd_sc_hd__mux4_2
XFILLER_0_124_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0980_ Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0925_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0926_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/C
+ sky130_fd_sc_hd__o21a_2
XFILLER_0_81_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput407 net407 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot1 Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[1\] Tile_X0Y0_DSP_top/J2END_AB_BEG\[1\] Tile_X0Y0_DSP_top/J_l_AB_BEG\[1\]
+ Tile_X0Y0_DSP_top/ConfigBits\[114\] Tile_X0Y0_DSP_top/ConfigBits\[115\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[1\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1
+ net21 net87 net139 net174 Tile_X0Y0_DSP_top/ConfigBits\[282\] Tile_X0Y0_DSP_top/ConfigBits\[283\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput418 net418 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput429 net429 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[9] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0
+ net283 net291 net183 net191 Tile_X0Y1_DSP_bot/ConfigBits\[340\] Tile_X0Y1_DSP_bot/ConfigBits\[341\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_data_outbuf_29__0_ Tile_X0Y0_DSP_top_data_inbuf_29__0_/X VGND VGND
+ VPWR VPWR net451 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1601_ Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1620_/A sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1532_ Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/C sky130_fd_sc_hd__a22o_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit7 net258 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[103\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit6 net77 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[284\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1463_ Tile_X0Y1_DSP_bot_Inst_MULADD__1463_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1463_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1471_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_89_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1394_ Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/A
+ sky130_fd_sc_hd__a21boi_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit3 net74 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[25\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_159_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[3\] net4 net136 Tile_X0Y1_bot2top\[3\] Tile_X0Y0_DSP_top/ConfigBits\[75\]
+ Tile_X0Y0_DSP_top/ConfigBits\[76\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__35_ net198 VGND VGND VPWR VPWR net600
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[5\]
+ Tile_X0Y0_DSP_top/ConfigBits\[108\] Tile_X0Y0_DSP_top/ConfigBits\[109\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit16 net56 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[166\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit27 net68 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[177\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_S4BEG_outbuf_9__0_ ANTENNA_93/DIODE VGND VGND VPWR VPWR Tile_X0Y0_S4BEG\[9\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 net764 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[264\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[265\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_51_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_E6END_inbuf_7__0_ net212 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/E6BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0963_ Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/A Tile_X0Y1_DSP_bot/A4
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0962_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0963_/Y
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0894_ Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0892_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0893_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0895_/A
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1515_ Tile_X0Y1_DSP_bot_Inst_MULADD__1513_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1717_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1664_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1523_/C
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit12 net232 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[12\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit23 net244 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[23\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_156_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1446_ Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1452_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1446_/Y
+ sky130_fd_sc_hd__a21boi_4
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit22 net63 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[300\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit11 net51 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[289\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1377_ Tile_X0Y1_DSP_bot_Inst_MULADD__1378_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1379_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__18_ Tile_X0Y0_top2bot\[14\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput760 net760 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[7] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[1\] Tile_X0Y0_S1BEG\[3\] Tile_X0Y0_S2BEGb\[5\] net335 Tile_X0Y1_DSP_bot/ConfigBits\[304\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[305\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_inbuf_1__0_ net272 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_1__0_/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_outbuf_6__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_6__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[6\] sky130_fd_sc_hd__buf_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1300_ Tile_X0Y1_DSP_bot_Inst_MULADD__1203_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1299_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1300_/Y
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit9 net80 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[383\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1231_ Tile_X0Y1_DSP_bot_Inst_MULADD__1211_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1210_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1212_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1231_/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1162_ Tile_X0Y1_DSP_bot_Inst_MULADD__1712_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1252_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1164_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_157_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1093_ Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/A Tile_X0Y1_DSP_bot/A6
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1093_/Y sky130_fd_sc_hd__nor2b_4
XFILLER_0_157_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit26 net67 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[208\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit15 net55 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[197\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit1 net60 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[87\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0946_ Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0946_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0946_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/A sky130_fd_sc_hd__nand4_4
XFILLER_0_2_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0877_ Tile_X0Y1_DSP_bot_Inst_MULADD__0876_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1707_/Q
+ Tile_X0Y1_DSP_bot/ConfigBits\[3\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0878_/C
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1429_ Tile_X0Y1_DSP_bot_Inst_MULADD__1501_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0933_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1180_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/A sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_92_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1
+ net89 net101 net141 net153 Tile_X0Y0_DSP_top/ConfigBits\[354\] Tile_X0Y0_DSP_top/ConfigBits\[355\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG3 net301
+ net201 Tile_X0Y0_S4BEG\[0\] Tile_X0Y1_DSP_bot/JW2BEG\[1\] Tile_X0Y1_DSP_bot/ConfigBits\[390\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[391\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_AB_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
Xoutput590 net590 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_WW4BEG_outbuf_4__0_ ANTENNA_113/DIODE VGND VGND VPWR VPWR net757
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit11 net231 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[43\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit22 net243 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[54\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit10 net50 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[320\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit21 net62 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[331\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_122_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG1 net288
+ net188 Tile_X0Y0_S2BEGb\[3\] net373 Tile_X0Y1_DSP_bot/ConfigBits\[242\] Tile_X0Y1_DSP_bot/ConfigBits\[243\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_EF_BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_137_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit19 net59 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[105\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1214_ Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/X sky130_fd_sc_hd__and4_1
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1145_ Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_157_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1076_ Tile_X0Y1_DSP_bot_Inst_MULADD__1076_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q5 sky130_fd_sc_hd__buf_12
XFILLER_0_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[2\] Tile_X0Y1_N2BEGb\[6\] net3 net11 Tile_X0Y0_DSP_top/ConfigBits\[266\]
+ Tile_X0Y0_DSP_top/ConfigBits\[267\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0929_ Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1378_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0929_/Y sky130_fd_sc_hd__nand2_1
Xinput307 Tile_X0Y1_N4END[15] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_1
Xinput318 Tile_X0Y1_NN4END[10] VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_1
Xinput329 Tile_X0Y1_NN4END[6] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit14 net54 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[228\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit25 net66 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[239\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_146_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_WW4END_inbuf_7__0_ net368 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/WW4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[9\] Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[2\] Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2END_AB_BEG\[2\] Tile_X0Y0_DSP_top/ConfigBits\[101\] Tile_X0Y0_DSP_top/ConfigBits\[102\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[1\] Tile_X0Y0_S1BEG\[3\] Tile_X0Y0_S2BEGb\[7\] net337 Tile_X0Y1_DSP_bot/ConfigBits\[376\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[377\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_107_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_NN4BEG_outbuf_1__0_ Tile_X0Y0_DSP_top/NN4BEG_i\[1\] VGND VGND VPWR
+ VPWR net525 sky130_fd_sc_hd__clkbuf_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit4 net75 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[186\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1694_ Tile_X0Y1_DSP_bot_Inst_MULADD__1674_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1694_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1695_/A sky130_fd_sc_hd__and2b_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1128_ Tile_X0Y1_DSP_bot_Inst_MULADD__1128_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1
+ net88 net110 net140 net156 Tile_X0Y0_DSP_top/ConfigBits\[318\] Tile_X0Y0_DSP_top/ConfigBits\[319\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1059_ Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1016_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1059_/X sky130_fd_sc_hd__a41o_1
XTile_X0Y0_DSP_top_SS4BEG_outbuf_4__0_ Tile_X0Y0_DSP_top/SS4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_SS4BEG\[4\] sky130_fd_sc_hd__buf_4
XFILLER_0_43_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput126 Tile_X0Y0_SS4END[3] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_1
Xinput115 Tile_X0Y0_S4END[8] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_1
Xinput104 Tile_X0Y0_S4END[12] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
Xinput159 Tile_X0Y0_W6END[4] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_1
Xinput137 Tile_X0Y0_W2END[0] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_2
Xinput148 Tile_X0Y0_W2MID[3] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit10 net230 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[74\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit21 net242 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[85\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit2 net251 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[322\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit20 net61 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[362\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_85_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit31 net73 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[373\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[47\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__o21ai_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit18 net58 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[136\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit29 net70 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[147\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__49_ Tile_X0Y0_DSP_top/JW2BEG\[1\] VGND
+ VGND VPWR VPWR net540 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__51_ net298 VGND VGND VPWR VPWR Tile_X0Y1_N2BEGb\[5\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_150_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit5 net256 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[69\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1746_ net333 Tile_X0Y1_DSP_bot/C4 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1677_ Tile_X0Y1_DSP_bot_Inst_MULADD__1674_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1677_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1678_/A sky130_fd_sc_hd__and2b_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit24 net65 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[270\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_133_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit13 net53 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[259\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[354\] Tile_X0Y1_DSP_bot/ConfigBits\[355\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JW2BEG\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_156_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_WW4END_inbuf_3__0_ net178 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/WW4BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_2
Xoutput408 net408 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[4] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot2 Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[2\] Tile_X0Y0_DSP_top/J2END_AB_BEG\[2\] Tile_X0Y0_DSP_top/J_l_AB_BEG\[2\]
+ Tile_X0Y0_DSP_top/ConfigBits\[116\] Tile_X0Y0_DSP_top/ConfigBits\[117\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[2\] sky130_fd_sc_hd__mux4_1
Xoutput419 net419 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[14] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[282\] Tile_X0Y0_DSP_top/ConfigBits\[283\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[2\] Tile_X0Y0_S2BEGb\[6\] net334 net336 Tile_X0Y1_DSP_bot/ConfigBits\[340\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[341\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1600_ Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/B
+ sky130_fd_sc_hd__nand3_2
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1531_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/C
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit8 net259 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[104\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit7 net78 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[285\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_145_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1462_ Tile_X0Y1_DSP_bot_Inst_MULADD__1471_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1471_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1463_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1463_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1465_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_145_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1393_ Tile_X0Y1_DSP_bot_Inst_MULADD__1314_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1389_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1391_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1392_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1421_/C sky130_fd_sc_hd__o211ai_4
XFILLER_0_145_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit4 net75 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[26\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_159_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_161_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[7\] Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[2\] Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2END_EF_BEG\[3\] Tile_X0Y0_DSP_top/ConfigBits\[75\] Tile_X0Y0_DSP_top/ConfigBits\[76\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__34_ net197 VGND VGND VPWR VPWR net599
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit30 net72 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[404\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1729_ net333 Tile_X0Y1_DSP_bot/A3 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1729_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[108\] Tile_X0Y0_DSP_top/ConfigBits\[109\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit17 net57 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[167\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit28 net69 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[178\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[264\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[265\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[53\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_NN4BEG_outbuf_7__0_ Tile_X0Y1_DSP_bot/NN4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y1_NN4BEG\[7\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0962_ Tile_X0Y1_DSP_bot_Inst_MULADD__1730_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0962_/X sky130_fd_sc_hd__or2b_2
XTile_X0Y1_DSP_bot_SS4END_inbuf_9__0_ Tile_X0Y0_SS4BEG\[13\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/SS4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0893_ Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1736_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0893_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_120_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit13 net233 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[13\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit24 net245 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[24\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1514_ Tile_X0Y1_DSP_bot_Inst_MULADD__1614_/S VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1664_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1445_ Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1452_/A
+ sky130_fd_sc_hd__a21boi_2
XFILLER_0_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit12 net52 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[290\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1376_ Tile_X0Y1_DSP_bot_Inst_MULADD__0933_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1128_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1275_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1375_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/B sky130_fd_sc_hd__o221ai_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit23 net64 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[301\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__17_ Tile_X0Y0_top2bot\[13\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_S4END_inbuf_1__0_ net112 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/S4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput761 net761 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput750 net750 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[12] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[304\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[305\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1230_ Tile_X0Y1_DSP_bot_Inst_MULADD__1243_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1243_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1243_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1230_/Y
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1161_ Tile_X0Y1_DSP_bot_Inst_MULADD__1252_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1161_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1164_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_59_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1092_ Tile_X0Y1_DSP_bot_Inst_MULADD__1089_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1091_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1092_/Y
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_W6END_inbuf_5__0_ net162 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/W6BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_WW4BEG_outbuf_10__0_ Tile_X0Y1_DSP_bot/WW4BEG_i\[10\] VGND VGND
+ VPWR VPWR net748 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_EE4END_inbuf_8__0_ net216 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/EE4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_70_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit16 net56 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[198\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit27 net68 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[209\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0945_ Tile_X0Y1_DSP_bot_Inst_MULADD__0943_/X Tile_X0Y1_DSP_bot_Inst_MULADD__0944_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0942_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0946_/C
+ sky130_fd_sc_hd__o21bai_2
XFILLER_0_140_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit2 net71 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[88\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0876_ Tile_X0Y1_DSP_bot/C1 Tile_X0Y1_DSP_bot_Inst_MULADD__1743_/Q
+ Tile_X0Y1_DSP_bot/ConfigBits\[2\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0876_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1428_ Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/A Tile_X0Y1_DSP_bot/A4
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0962_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1427_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/B sky130_fd_sc_hd__o2111ai_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1359_ Tile_X0Y1_DSP_bot_Inst_MULADD__1019_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1358_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1356_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1354_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1359_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_148_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_EE4BEG_outbuf_4__0_ Tile_X0Y0_DSP_top/EE4BEG_i\[4\] VGND VGND VPWR
+ VPWR net424 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[354\] Tile_X0Y0_DSP_top/ConfigBits\[355\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_S4END_inbuf_1__0_ Tile_X0Y0_S4BEG\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/S4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
Xoutput580 net580 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput591 net591 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[4] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit0 net229 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[224\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit12 net232 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[44\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit23 net244 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[55\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_107_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_SS4END_inbuf_5__0_ net132 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/SS4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit22 net63 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[332\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit11 net51 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[321\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[94\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG2 net290
+ net190 Tile_X0Y0_SS4BEG\[1\] net343 Tile_X0Y1_DSP_bot/ConfigBits\[244\] Tile_X0Y1_DSP_bot/ConfigBits\[245\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_EF_BEG\[2\] sky130_fd_sc_hd__mux4_1
XFILLER_0_137_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_strobe_outbuf_16__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_16__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[16\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1213_ Tile_X0Y1_DSP_bot_Inst_MULADD__1210_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1211_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1212_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1213_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1144_ Tile_X0Y1_DSP_bot_Inst_MULADD__1144_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1144_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1144_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1075_ Tile_X0Y1_DSP_bot_Inst_MULADD__1681_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1711_/Q
+ Tile_X0Y1_DSP_bot/ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1076_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_W6END_inbuf_5__0_ net363 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/W6BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0928_ Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/A sky130_fd_sc_hd__buf_4
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1
+ net83 net91 net133 net135 Tile_X0Y0_DSP_top/ConfigBits\[266\] Tile_X0Y0_DSP_top/ConfigBits\[267\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0859_ Tile_X0Y1_DSP_bot_Inst_MULADD__1706_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0858_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q0
+ sky130_fd_sc_hd__a21bo_4
Xinput308 Tile_X0Y1_N4END[1] VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput319 Tile_X0Y1_NN4END[11] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_WW4END_inbuf_10__0_ net371 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/WW4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit26 net67 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[240\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit15 net55 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[229\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[376\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[377\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_EE4END_inbuf_4__0_ net47 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/EE4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_150_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_N4BEG_outbuf_11__0_ ANTENNA_185/DIODE VGND VGND VPWR VPWR Tile_X0Y1_N4BEG\[11\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1693_ Tile_X0Y1_DSP_bot_Inst_MULADD__1693_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1717_/D sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit5 net76 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[187\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[0\] Tile_X0Y1_N2BEGb\[0\] net1 net5 Tile_X0Y0_DSP_top/ConfigBits\[306\]
+ Tile_X0Y0_DSP_top/ConfigBits\[307\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1127_ Tile_X0Y1_DSP_bot_Inst_MULADD__1034_/X Tile_X0Y1_DSP_bot/B6
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1121_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1128_/A
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1058_ Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/A sky130_fd_sc_hd__buf_4
XFILLER_0_145_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[318\] Tile_X0Y0_DSP_top/ConfigBits\[319\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_NN4BEG_outbuf_11__0_ ANTENNA_78/DIODE VGND VGND VPWR VPWR net520
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_N4BEG_outbuf_3__0_ Tile_X0Y1_DSP_bot/N4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N4BEG\[3\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput127 Tile_X0Y0_SS4END[4] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
Xinput116 Tile_X0Y0_S4END[9] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
Xinput105 Tile_X0Y0_S4END[13] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
Xinput138 Tile_X0Y0_W2END[1] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_2
Xinput149 Tile_X0Y0_W2MID[4] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit11 net231 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[75\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit22 net243 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[86\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit3 net254 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[323\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit21 net62 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[363\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit10 net50 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[352\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[47\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit19 net59 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[137\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__48_ net137 VGND VGND VPWR VPWR net539
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__50_ net297 VGND VGND VPWR VPWR Tile_X0Y1_N2BEGb\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit6 net257 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[70\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[100\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1745_ net333 Tile_X0Y1_DSP_bot/C3 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1676_ Tile_X0Y1_DSP_bot_Inst_MULADD__1676_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1708_/D sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_E6BEG_outbuf_8__0_ Tile_X0Y0_DSP_top/E6BEG_i\[8\] VGND VGND VPWR
+ VPWR net412 sky130_fd_sc_hd__clkbuf_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_strobe_outbuf_11__0_ Tile_X0Y0_DSP_top_strobe_inbuf_11__0_/X VGND
+ VGND VPWR VPWR net464 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_W6BEG_outbuf_3__0_ Tile_X0Y1_DSP_bot/W6BEG_i\[3\] VGND VGND VPWR
+ VPWR net740 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_SS4END_inbuf_10__0_ net122 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/SS4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_data_outbuf_1__0_ Tile_X0Y0_DSP_top_data_inbuf_1__0_/X VGND VGND
+ VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit25 net66 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[271\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit14 net54 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[260\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot3 Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[3\]
+ Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[3\] Tile_X0Y0_DSP_top/J2END_AB_BEG\[3\] Tile_X0Y0_DSP_top/J_l_AB_BEG\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[118\] Tile_X0Y0_DSP_top/ConfigBits\[119\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[3\] sky130_fd_sc_hd__mux4_1
Xoutput409 net409 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[5] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[282\] Tile_X0Y0_DSP_top/ConfigBits\[283\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_data_inbuf_25__0_ net66 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_25__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[340\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[341\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_129_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1530_ Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/B sky130_fd_sc_hd__or2_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit9 net260 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[105\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1461_ Tile_X0Y1_DSP_bot_Inst_MULADD__1716_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1614_/S
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1463_/B sky130_fd_sc_hd__and2b_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit8 net79 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[286\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1392_ Tile_X0Y1_DSP_bot_Inst_MULADD__1386_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1386_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1382_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1365_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1392_/Y sky130_fd_sc_hd__o22ai_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit5 net76 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[27\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__33_ net196 VGND VGND VPWR VPWR net598
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_data_inbuf_16__0_ net56 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_16__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit31 net73 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[405\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit20 net61 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[394\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot10 Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2MID_EFb_BEG\[2\] Tile_X0Y0_DSP_top/J2END_EF_BEG\[2\] Tile_X0Y0_DSP_top/J_l_EF_BEG\[2\]
+ Tile_X0Y0_DSP_top/ConfigBits\[132\] Tile_X0Y0_DSP_top/ConfigBits\[133\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[10\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1728_ net333 Tile_X0Y1_DSP_bot/A2 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1728_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[2\] Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[2\] Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[2\] Tile_X0Y0_DSP_top/ConfigBits\[108\] Tile_X0Y0_DSP_top/ConfigBits\[109\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1659_ Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1659_/X sky130_fd_sc_hd__a31o_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit18 net58 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[168\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit29 net70 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[179\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[266\] Tile_X0Y1_DSP_bot/ConfigBits\[267\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JN2BEG\[2\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_data_outbuf_1__0_ Tile_X0Y1_DSP_bot_data_inbuf_1__0_/X VGND VGND
+ VPWR VPWR net642 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[53\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_data_outbuf_23__0_ Tile_X0Y1_DSP_bot_data_inbuf_23__0_/X VGND VGND
+ VPWR VPWR net646 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__0961_ Tile_X0Y1_DSP_bot_Inst_MULADD__0959_/X Tile_X0Y1_DSP_bot_Inst_MULADD__0960_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0946_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/A
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_152_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0892_ ANTENNA_97/DIODE VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0892_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1513_ Tile_X0Y1_DSP_bot/C11 Tile_X0Y1_DSP_bot_Inst_MULADD__1753_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1513_/X
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit14 net234 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[14\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_data_inbuf_25__0_ net246 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_25__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1444_ Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/C
+ sky130_fd_sc_hd__nand3_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit25 net246 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[25\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1375_ Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/D Tile_X0Y1_DSP_bot_Inst_MULADD__0963_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1371_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1375_/X
+ sky130_fd_sc_hd__o21a_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit13 net53 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[291\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_data_outbuf_14__0_ Tile_X0Y1_DSP_bot_data_inbuf_14__0_/X VGND VGND
+ VPWR VPWR net636 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit24 net65 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[302\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_147_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__16_ Tile_X0Y0_top2bot\[12\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_S4BEG_outbuf_3__0_ ANTENNA_108/DIODE VGND VGND VPWR VPWR net692
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_data_inbuf_7__0_ net78 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_7__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput751 net751 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput762 net762 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput740 net740 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[304\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[305\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_data_inbuf_16__0_ net236 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_16__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1160_ Tile_X0Y1_DSP_bot/C6 Tile_X0Y1_DSP_bot_Inst_MULADD__1748_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1459_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1161_/B
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1091_ Tile_X0Y1_DSP_bot_Inst_MULADD__1091_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1091_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit17 net57 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[199\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit28 net69 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[210\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0944_ Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0934_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0944_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_140_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit3 net74 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[89\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0875_ Tile_X0Y1_DSP_bot_Inst_MULADD__0875_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0906_/C sky130_fd_sc_hd__or4_4
XFILLER_0_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1427_ Tile_X0Y1_DSP_bot_Inst_MULADD__1356_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1354_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1019_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1358_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1427_/Y sky130_fd_sc_hd__o2bb2ai_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1358_ Tile_X0Y1_DSP_bot_Inst_MULADD__1093_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1095_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1358_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1289_ Tile_X0Y1_DSP_bot_Inst_MULADD__1289_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1289_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1289_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[354\] Tile_X0Y0_DSP_top/ConfigBits\[355\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_135_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput570 net570 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput581 net581 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[8] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_NN4END_inbuf_9__0_ net321 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/NN4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
Xoutput592 net592 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[5] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit1 net240 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[225\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit24 net245 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[56\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit13 net233 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[45\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_134_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit23 net64 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[333\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit12 net52 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[322\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[94\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG3 net325
+ net186 Tile_X0Y0_S2BEGb\[1\] net339 Tile_X0Y1_DSP_bot/ConfigBits\[246\] Tile_X0Y1_DSP_bot/ConfigBits\[247\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_EF_BEG\[3\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1212_ Tile_X0Y1_DSP_bot_Inst_MULADD__1378_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1204_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1201_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1212_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1143_ Tile_X0Y1_DSP_bot_Inst_MULADD__1133_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1141_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1142_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1144_/B
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y0_DSP_top_data_outbuf_10__0_ Tile_X0Y0_DSP_top_data_inbuf_10__0_/X VGND VGND
+ VPWR VPWR net431 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_190 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1074_ Tile_X0Y1_DSP_bot_Inst_MULADD__1074_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1074_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1681_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0927_ Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0925_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0926_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/A
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[266\] Tile_X0Y0_DSP_top/ConfigBits\[267\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0858_ Tile_X0Y1_DSP_bot/ConfigBits\[5\] Tile_X0Y1_DSP_bot_Inst_MULADD__1672_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1672_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0858_/X
+ sky130_fd_sc_hd__or3_1
Xinput309 Tile_X0Y1_N4END[2] VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_EE4END_inbuf_10__0_ net38 VGND VGND VPWR VPWR ANTENNA_175/DIODE
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit27 net68 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[241\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit16 net56 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[230\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/Q5 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9
+ Tile_X0Y1_DSP_bot/ConfigBits\[376\] Tile_X0Y1_DSP_bot/ConfigBits\[377\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1761_ net333 Tile_X0Y1_DSP_bot/C19 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1761_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit6 net77 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[188\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1692_ Tile_X0Y1_DSP_bot_Inst_MULADD__1674_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1692_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1693_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_strobe_outbuf_3__0_ Tile_X0Y0_DSP_top_strobe_inbuf_3__0_/X VGND
+ VGND VPWR VPWR net475 sky130_fd_sc_hd__clkbuf_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1
+ net81 net83 net117 net165 Tile_X0Y0_DSP_top/ConfigBits\[306\] Tile_X0Y0_DSP_top/ConfigBits\[307\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1126_ Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/A
+ sky130_fd_sc_hd__and3_2
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1057_ Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/D sky130_fd_sc_hd__buf_4
XFILLER_0_16_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[318\] Tile_X0Y0_DSP_top/ConfigBits\[319\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_data_inbuf_0__0_ net229 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_0__0_/X
+ sky130_fd_sc_hd__clkbuf_1
Xinput117 Tile_X0Y0_SS4END[0] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
Xinput106 Tile_X0Y0_S4END[14] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
Xinput128 Tile_X0Y0_SS4END[5] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
Xinput139 Tile_X0Y0_W2END[2] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_NN4END_inbuf_5__0_ Tile_X0Y1_NN4BEG\[9\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/NN4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit12 net232 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[76\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit23 net244 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[87\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_S1BEG0 Tile_X0Y1_DSP_bot/Q4
+ Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[3\] Tile_X0Y1_DSP_bot/JE2BEG\[3\] Tile_X0Y1_DSP_bot/J_l_CD_BEG\[1\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[62\] Tile_X0Y1_DSP_bot/ConfigBits\[63\] VGND VGND
+ VPWR VPWR net663 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit4 net255 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[324\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit11 net51 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[353\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit22 net63 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[364\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_90 ANTENNA_91/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__47_ net100 VGND VGND VPWR VPWR Tile_X0Y0_S2BEGb\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_SS4BEG_outbuf_10__0_ Tile_X0Y1_DSP_bot/SS4BEG_i\[10\] VGND VGND
+ VPWR VPWR net700 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_WW4BEG_outbuf_1__0_ Tile_X0Y0_DSP_top/WW4BEG_i\[1\] VGND VGND VPWR
+ VPWR net574 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_strobe_inbuf_18__0_ Tile_X0Y1_FrameStrobe_O\[18\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_18__0_/X sky130_fd_sc_hd__clkbuf_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit7 net258 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[71\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[100\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1744_ net333 Tile_X0Y1_DSP_bot/C2 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1675_ Tile_X0Y1_DSP_bot_Inst_MULADD__1674_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1675_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1676_/A sky130_fd_sc_hd__and2b_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1109_ Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/Y
+ sky130_fd_sc_hd__nand3_2
XFILLER_0_63_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_inbuf_11__0_ net263 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_11__0_/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_133_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit26 net67 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[272\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit15 net55 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[261\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_N4END_inbuf_1__0_ Tile_X0Y1_N4BEG\[5\] VGND VGND VPWR VPWR ANTENNA_74/DIODE
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot4 Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[0\]
+ Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[0\] Tile_X0Y0_DSP_top/J2END_CD_BEG\[0\] Tile_X0Y0_DSP_top/J_l_CD_BEG\[0\]
+ Tile_X0Y0_DSP_top/ConfigBits\[120\] Tile_X0Y0_DSP_top/ConfigBits\[121\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[4\] sky130_fd_sc_hd__mux4_2
XFILLER_0_105_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst0
+ net283 net183 net336 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/ConfigBits\[22\] Tile_X0Y1_DSP_bot/ConfigBits\[23\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[284\] Tile_X0Y0_DSP_top/ConfigBits\[285\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JE2BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q4 wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[340\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[341\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1460_ Tile_X0Y1_DSP_bot_Inst_MULADD__1614_/S Tile_X0Y1_DSP_bot_Inst_MULADD__1460_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1463_/A sky130_fd_sc_hd__nor2_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit9 net80 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[287\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1391_ Tile_X0Y1_DSP_bot_Inst_MULADD__1366_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1370_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1386_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1390_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1391_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_89_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit6 net77 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[28\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_89_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__32_ net195 VGND VGND VPWR VPWR net597
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit10 net50 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[384\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot11 Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[3\]
+ Tile_X0Y0_DSP_top/J2MID_EFb_BEG\[3\] Tile_X0Y0_DSP_top/J2END_EF_BEG\[3\] Tile_X0Y0_DSP_top/J_l_EF_BEG\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[134\] Tile_X0Y0_DSP_top/ConfigBits\[135\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[11\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit21 net62 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[395\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1727_ net333 Tile_X0Y1_DSP_bot/A1 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1727_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[110\] Tile_X0Y0_DSP_top/ConfigBits\[111\] VGND VGND
+ VPWR VPWR net557 sky130_fd_sc_hd__mux4_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1658_ Tile_X0Y1_DSP_bot_Inst_MULADD__1658_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1658_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/C sky130_fd_sc_hd__nor2_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit19 net59 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[169\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1589_ Tile_X0Y1_DSP_bot_Inst_MULADD__1589_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1589_/Y sky130_fd_sc_hd__inv_2
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_strobe_inbuf_4__0_ net275 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_4__0_/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[83\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR Tile_X0Y0_SS4BEG\[15\] sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0960_ Tile_X0Y1_DSP_bot_Inst_MULADD__0942_/B Tile_X0Y1_DSP_bot_Inst_MULADD__0942_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0942_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0960_/Y
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot_strobe_outbuf_9__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_9__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[9\] sky130_fd_sc_hd__buf_8
XTile_X0Y1_DSP_bot_Inst_MULADD__0891_ Tile_X0Y1_DSP_bot/ConfigBits\[1\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/A sky130_fd_sc_hd__buf_4
XTile_X0Y1_DSP_bot_N4END_inbuf_1__0_ net312 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/N4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1512_ Tile_X0Y1_DSP_bot_Inst_MULADD__1446_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1450_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1458_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1458_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1511_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1523_/B sky130_fd_sc_hd__o221ai_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit15 net235 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[15\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1443_ Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/B
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit26 net247 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[26\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1374_ Tile_X0Y1_DSP_bot_Inst_MULADD__1371_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1372_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1373_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/A
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit25 net66 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[303\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit14 net54 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[292\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_105_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__15_ Tile_X0Y0_top2bot\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput730 net730 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput752 net752 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput741 net741 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[4] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[306\] Tile_X0Y1_DSP_bot/ConfigBits\[307\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JE2BEG\[4\] sky130_fd_sc_hd__mux4_2
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_WW4BEG_outbuf_7__0_ Tile_X0Y1_DSP_bot/WW4BEG_i\[7\] VGND VGND VPWR
+ VPWR net760 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1090_ Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/A Tile_X0Y1_DSP_bot/A5
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1091_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_142_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit18 net58 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[200\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_82_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit29 net70 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[211\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0943_ Tile_X0Y1_DSP_bot_Inst_MULADD__0888_/X Tile_X0Y1_DSP_bot_Inst_MULADD__0889_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0934_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0943_/X sky130_fd_sc_hd__o2111a_1
XFILLER_0_140_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit4 net75 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[90\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0874_ Tile_X0Y1_DSP_bot/A0 Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0849_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/A
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1426_ Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1354_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1356_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1425_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1501_/A sky130_fd_sc_hd__a221o_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1357_ Tile_X0Y1_DSP_bot_Inst_MULADD__1354_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1356_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1357_/Y
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1288_ Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1283_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1288_/X sky130_fd_sc_hd__a22o_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[356\] Tile_X0Y0_DSP_top/ConfigBits\[357\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JW2BEG\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_108_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0
+ net281 net287 net187 net201 Tile_X0Y1_DSP_bot/ConfigBits\[356\] Tile_X0Y1_DSP_bot/ConfigBits\[357\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0
+ net184 net337 Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/ConfigBits\[110\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[111\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput560 net560 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput571 net571 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput582 net582 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput593 net593 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[6] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit2 net251 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[226\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_158_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_strobe_inbuf_0__0_ Tile_X0Y1_FrameStrobe_O\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_0__0_/X sky130_fd_sc_hd__buf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit25 net246 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[57\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit14 net234 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[46\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_108_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit24 net65 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[334\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit13 net53 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[323\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1211_ Tile_X0Y1_DSP_bot_Inst_MULADD__0933_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0963_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1211_/X sky130_fd_sc_hd__o22a_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1142_ Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1064_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1079_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1142_/Y
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_153_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_180 ANTENNA_180/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1073_ Tile_X0Y1_DSP_bot_Inst_MULADD__1073_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1073_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1074_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_145_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[89\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__o21ai_2
XFILLER_0_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_NN4BEG_outbuf_4__0_ Tile_X0Y0_DSP_top/NN4BEG_i\[4\] VGND VGND VPWR
+ VPWR net528 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__0926_ Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1737_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0926_/Y sky130_fd_sc_hd__nand2_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[266\] Tile_X0Y0_DSP_top/ConfigBits\[267\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0857_ Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/D Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0856_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1672_/C
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1409_ Tile_X0Y1_DSP_bot_Inst_MULADD__1408_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1715_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1614_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1412_/B
+ sky130_fd_sc_hd__mux2_1
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_SS4BEG_outbuf_7__0_ Tile_X0Y0_DSP_top/SS4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_SS4BEG\[7\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__63_ net152 VGND VGND VPWR VPWR net554
+ sky130_fd_sc_hd__clkbuf_1
Xoutput390 net390 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[4] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_S4BEG_outbuf_11__0_ Tile_X0Y0_DSP_top/S4BEG_i\[11\] VGND VGND VPWR
+ VPWR Tile_X0Y0_S4BEG\[11\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit17 net57 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[231\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit28 net69 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[242\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[378\] Tile_X0Y1_DSP_bot/ConfigBits\[379\] VGND VGND
+ VPWR VPWR ANTENNA_184/DIODE sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_E1BEG0 Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[3\] Tile_X0Y0_DSP_top/JN2BEG\[3\] Tile_X0Y0_DSP_top/J_l_CD_BEG\[1\]
+ Tile_X0Y0_DSP_top/ConfigBits\[28\] Tile_X0Y0_DSP_top/ConfigBits\[29\] VGND VGND
+ VPWR VPWR net382 sky130_fd_sc_hd__mux4_1
XFILLER_0_12_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1760_ net333 Tile_X0Y1_DSP_bot/C18 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_SS4BEG_outbuf_0__0_ Tile_X0Y1_DSP_bot/SS4BEG_i\[0\] VGND VGND VPWR
+ VPWR net699 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1691_ Tile_X0Y1_DSP_bot_Inst_MULADD__1691_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit7 net78 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[189\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[306\] Tile_X0Y0_DSP_top/ConfigBits\[307\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1125_ Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1124_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/C sky130_fd_sc_hd__a31oi_4
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1056_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0963_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1019_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0875_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1056_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_22_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[320\] Tile_X0Y0_DSP_top/ConfigBits\[321\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JS2BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_160_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0
+ net324 net184 net186 net204 Tile_X0Y1_DSP_bot/ConfigBits\[320\] Tile_X0Y1_DSP_bot/ConfigBits\[321\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__0909_ Tile_X0Y1_DSP_bot/ConfigBits\[3\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1252_/A sky130_fd_sc_hd__clkbuf_4
Xinput118 Tile_X0Y0_SS4END[10] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
Xinput107 Tile_X0Y0_S4END[15] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
Xinput129 Tile_X0Y0_SS4END[6] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit13 net233 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[77\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit24 net245 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[88\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_S1BEG1 Tile_X0Y1_DSP_bot/Q5
+ Tile_X0Y1_DSP_bot/J2MID_EFb_BEG\[0\] Tile_X0Y1_DSP_bot/JE2BEG\[0\] Tile_X0Y1_DSP_bot/J_l_EF_BEG\[2\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[64\] Tile_X0Y1_DSP_bot/ConfigBits\[65\] VGND VGND
+ VPWR VPWR net664 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit5 net256 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[325\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit12 net52 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[354\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit23 net64 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[365\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_93_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_80 ANTENNA_86/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 ANTENNA_91/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__46_ net99 VGND VGND VPWR VPWR Tile_X0Y0_S2BEGb\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_WW4END_inbuf_6__0_ net166 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/WW4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1743_ net333 Tile_X0Y1_DSP_bot/C1 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1743_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit8 net259 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[72\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_0_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1674_ Tile_X0Y1_DSP_bot/clr VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1674_/X
+ sky130_fd_sc_hd__buf_2
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1108_ Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1106_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1107_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/C sky130_fd_sc_hd__o2bb2ai_2
XFILLER_0_158_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1039_ Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1739_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_133_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit16 net56 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[262\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit27 net68 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[273\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_98_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot5 Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[1\] Tile_X0Y0_DSP_top/J2END_CD_BEG\[1\] Tile_X0Y0_DSP_top/J_l_CD_BEG\[1\]
+ Tile_X0Y0_DSP_top/ConfigBits\[122\] Tile_X0Y0_DSP_top/ConfigBits\[123\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[5\] sky130_fd_sc_hd__mux4_1
XFILLER_0_22_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst1
+ net763 ANTENNA_101/DIODE Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[1\] Tile_X0Y1_DSP_bot/J2END_GH_BEG\[1\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[22\] Tile_X0Y1_DSP_bot/ConfigBits\[23\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[342\] Tile_X0Y1_DSP_bot/ConfigBits\[343\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JS2BEG\[5\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__29_ Tile_X0Y1_N2BEG\[5\] VGND VGND
+ VPWR VPWR net499 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1390_ Tile_X0Y1_DSP_bot_Inst_MULADD__1293_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1273_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1390_/X sky130_fd_sc_hd__a221o_2
XFILLER_0_89_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit7 net78 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[29\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_89_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst0
+ net281 Tile_X0Y0_S1BEG\[0\] net334 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[104\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[105\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_E6BEG_outbuf_2__0_ Tile_X0Y1_DSP_bot/E6BEG_i\[2\] VGND VGND VPWR
+ VPWR net607 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__31_ net194 VGND VGND VPWR VPWR net596
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[2\] net3 net83 Tile_X0Y1_bot2top\[2\] Tile_X0Y0_DSP_top/ConfigBits\[36\]
+ Tile_X0Y0_DSP_top/ConfigBits\[37\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot12 Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[0\]
+ Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[0\] Tile_X0Y0_DSP_top/J2END_GH_BEG\[0\] Tile_X0Y0_DSP_top/J_l_GH_BEG\[0\]
+ Tile_X0Y0_DSP_top/ConfigBits\[136\] Tile_X0Y0_DSP_top/ConfigBits\[137\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[12\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit11 net51 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[385\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit22 net63 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[396\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1726_ net333 Tile_X0Y1_DSP_bot/A0 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1657_ Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1657_/B
+ Tile_X0Y1_DSP_bot/ConfigBits\[4\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1658_/B
+ sky130_fd_sc_hd__and3_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1588_ Tile_X0Y1_DSP_bot_Inst_MULADD__1588_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1593_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1589_/A sky130_fd_sc_hd__nor2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_S4END_inbuf_4__0_ net115 VGND VGND VPWR VPWR ANTENNA_87/DIODE sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit0 net229 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[128\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[83\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0890_ Tile_X0Y1_DSP_bot_Inst_MULADD__0888_/X Tile_X0Y1_DSP_bot_Inst_MULADD__0889_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0890_/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1511_ Tile_X0Y1_DSP_bot_Inst_MULADD__1511_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1511_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1442_ Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1440_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1441_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/C sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit16 net236 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[16\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit27 net248 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[27\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput290 Tile_X0Y1_N2END[5] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1373_ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1373_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1373_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1373_/X
+ sky130_fd_sc_hd__and3_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit26 net67 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[304\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit15 net55 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[293\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_W6END_inbuf_8__0_ net154 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/W6BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__14_ Tile_X0Y0_top2bot\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput720 net720 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput753 net753 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput731 net731 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[4] sky130_fd_sc_hd__clkbuf_4
Xoutput742 net742 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[5] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1709_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1709_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1709_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_EE4BEG_outbuf_7__0_ Tile_X0Y0_DSP_top/EE4BEG_i\[7\] VGND VGND VPWR
+ VPWR net427 sky130_fd_sc_hd__clkbuf_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG0 Tile_X0Y1_N2BEG\[7\]
+ net20 net100 net152 Tile_X0Y0_DSP_top/ConfigBits\[198\] Tile_X0Y0_DSP_top/ConfigBits\[199\]
+ VGND VGND VPWR VPWR ANTENNA_177/DIODE sky130_fd_sc_hd__mux4_2
XFILLER_0_83_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_S4END_inbuf_4__0_ Tile_X0Y0_S4BEG\[8\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/S4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0
+ Tile_X0Y1_N2BEGb\[1\] Tile_X0Y1_N4BEG\[1\] net4 net6 Tile_X0Y0_DSP_top/ConfigBits\[246\]
+ Tile_X0Y0_DSP_top/ConfigBits\[247\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_EE4BEG_outbuf_0__0_ Tile_X0Y1_DSP_bot/EE4BEG_i\[0\] VGND VGND VPWR
+ VPWR net615 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_SS4END_inbuf_8__0_ net120 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/SS4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit19 net59 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[201\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0942_ Tile_X0Y1_DSP_bot_Inst_MULADD__0942_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0942_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0942_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0946_/B
+ sky130_fd_sc_hd__nand3_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0873_ Tile_X0Y1_DSP_bot_Inst_MULADD__1175_/B Tile_X0Y1_DSP_bot/B1
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0866_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/A
+ sky130_fd_sc_hd__a21boi_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit5 net76 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[91\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_strobe_outbuf_19__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_19__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[19\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1425_ Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1425_/X sky130_fd_sc_hd__and4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1356_ Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/A Tile_X0Y1_DSP_bot/A4
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0962_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1275_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1356_/X sky130_fd_sc_hd__o211a_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst0
+ net283 net183 net336 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/ConfigBits\[78\] Tile_X0Y1_DSP_bot/ConfigBits\[79\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1287_ Tile_X0Y1_DSP_bot_Inst_MULADD__1197_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1195_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1286_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/B sky130_fd_sc_hd__o211ai_4
XFILLER_0_148_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_W6END_inbuf_8__0_ net355 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/W6BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1
+ Tile_X0Y0_S2BEGb\[2\] Tile_X0Y0_S4BEG\[2\] net340 net354 Tile_X0Y1_DSP_bot/ConfigBits\[356\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[357\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/Q5
+ Tile_X0Y1_DSP_bot/ConfigBits\[110\] Tile_X0Y1_DSP_bot/ConfigBits\[111\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
Xoutput572 net572 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput561 net561 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput550 net550 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput583 net583 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput594 net594 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[7] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit3 net254 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[227\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_96_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit15 net235 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[47\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit26 net247 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[58\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit25 net66 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[335\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit14 net54 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[324\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1210_ Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1210_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1141_ Tile_X0Y1_DSP_bot_Inst_MULADD__1135_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1137_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1140_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1141_/Y
+ sky130_fd_sc_hd__o21bai_4
XANTENNA_170 Tile_X0Y1_FrameStrobe_O\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1072_ Tile_X0Y1_DSP_bot_Inst_MULADD__1070_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1072_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1072_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1073_/B
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_62_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_181 ANTENNA_181/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_192 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[89\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top_EE4END_inbuf_7__0_ net35 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/EE4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_153_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__0925_ Tile_X0Y1_DSP_bot/B3 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0925_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[268\] Tile_X0Y0_DSP_top/ConfigBits\[269\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JN2BEG\[5\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0856_ Tile_X0Y1_DSP_bot_Inst_MULADD__0856_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1672_/B
+ sky130_fd_sc_hd__and3_2
XFILLER_0_121_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0
+ net289 net301 net183 net189 Tile_X0Y1_DSP_bot/ConfigBits\[268\] Tile_X0Y1_DSP_bot/ConfigBits\[269\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1408_ Tile_X0Y1_DSP_bot/C9 Tile_X0Y1_DSP_bot_Inst_MULADD__1751_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1459_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1408_/X
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1339_ Tile_X0Y1_DSP_bot_Inst_MULADD__1339_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1339_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1339_/Y sky130_fd_sc_hd__nand2_1
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__62_ net151 VGND VGND VPWR VPWR net553
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_N4BEG_outbuf_6__0_ Tile_X0Y1_DSP_bot/N4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N4BEG\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput391 net391 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[5] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit18 net58 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[232\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit29 net70 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[243\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_E1BEG1 Tile_X0Y1_bot2top\[4\]
+ ANTENNA_177/DIODE Tile_X0Y0_DSP_top/JN2BEG\[0\] Tile_X0Y0_DSP_top/J_l_EF_BEG\[2\]
+ Tile_X0Y0_DSP_top/ConfigBits\[30\] Tile_X0Y0_DSP_top/ConfigBits\[31\] VGND VGND
+ VPWR VPWR net383 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1690_ Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1690_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1690_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1691_/A
+ sky130_fd_sc_hd__and3b_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit8 net79 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[190\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[306\] Tile_X0Y0_DSP_top/ConfigBits\[307\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1124_ Tile_X0Y1_DSP_bot_Inst_MULADD__1124_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1124_/X sky130_fd_sc_hd__and4_1
XFILLER_0_118_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1055_ Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1025_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1055_/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1
+ Tile_X0Y0_S2BEGb\[1\] Tile_X0Y0_S4BEG\[1\] net339 net357 Tile_X0Y1_DSP_bot/ConfigBits\[320\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[321\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_NN4END_inbuf_10__0_ Tile_X0Y1_NN4BEG\[14\] VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top/NN4BEG_i\[10\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0908_ Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/D Tile_X0Y1_DSP_bot_Inst_MULADD__0907_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0915_/A sky130_fd_sc_hd__or2b_1
Xinput108 Tile_X0Y0_S4END[1] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_4
Xinput119 Tile_X0Y0_SS4END[11] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_strobe_outbuf_14__0_ Tile_X0Y0_DSP_top_strobe_inbuf_14__0_/X VGND
+ VGND VPWR VPWR net467 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit14 net234 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[78\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit25 net246 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[89\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit6 net257 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[326\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_S1BEG2 net763 Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[1\]
+ Tile_X0Y1_DSP_bot/JE2BEG\[1\] Tile_X0Y1_DSP_bot/J_l_GH_BEG\[3\] Tile_X0Y1_DSP_bot/ConfigBits\[66\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[67\] VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit24 net65 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[366\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_109_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit13 net53 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[355\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_W6BEG_outbuf_6__0_ Tile_X0Y1_DSP_bot/W6BEG_i\[6\] VGND VGND VPWR
+ VPWR net743 sky130_fd_sc_hd__clkbuf_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_data_outbuf_4__0_ Tile_X0Y0_DSP_top_data_inbuf_4__0_/X VGND VGND
+ VPWR VPWR net456 sky130_fd_sc_hd__clkbuf_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_70 ANTENNA_73/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_81 ANTENNA_86/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 ANTENNA_92/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__45_ net98 VGND VGND VPWR VPWR Tile_X0Y0_S2BEGb\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_159_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_data_inbuf_28__0_ net69 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_28__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1742_ net333 Tile_X0Y1_DSP_bot/C0 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1742_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit9 net260 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[73\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1673_ Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1673_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1707_/D sky130_fd_sc_hd__nor2_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1107_ Tile_X0Y1_DSP_bot_Inst_MULADD__1034_/X ANTENNA_97/DIODE
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/D VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1107_/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1038_ Tile_X0Y1_DSP_bot/B5 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1038_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit17 net57 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[263\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_data_inbuf_19__0_ net59 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_19__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput90 Tile_X0Y0_S2END[5] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_N4BEG_outbuf_2__0_ Tile_X0Y0_DSP_top/N4BEG_i\[2\] VGND VGND VPWR
+ VPWR net510 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit28 net69 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[274\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_data_outbuf_4__0_ Tile_X0Y1_DSP_bot_data_inbuf_4__0_/X VGND VGND
+ VPWR VPWR net657 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot6 Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[2\] Tile_X0Y0_DSP_top/J2END_CD_BEG\[2\] Tile_X0Y0_DSP_top/J_l_CD_BEG\[2\]
+ Tile_X0Y0_DSP_top/ConfigBits\[124\] Tile_X0Y0_DSP_top/ConfigBits\[125\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[6\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__28_ Tile_X0Y1_N2BEG\[4\] VGND VGND
+ VPWR VPWR net498 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_data_outbuf_26__0_ Tile_X0Y1_DSP_bot_data_inbuf_26__0_/X VGND VGND
+ VPWR VPWR net649 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit8 net79 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[30\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_147_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q8 ANTENNA_105/DIODE Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[1\] Tile_X0Y1_DSP_bot/J2END_CD_BEG\[2\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[104\] Tile_X0Y1_DSP_bot/ConfigBits\[105\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__30_ net193 VGND VGND VPWR VPWR net595
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[6\] Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[1\] Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2END_GH_BEG\[0\] Tile_X0Y0_DSP_top/ConfigBits\[36\] Tile_X0Y0_DSP_top/ConfigBits\[37\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit23 net64 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[397\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_data_inbuf_28__0_ net249 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_28__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1725_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1725_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1725_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit12 net52 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[386\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot13 Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[1\] Tile_X0Y0_DSP_top/J2END_GH_BEG\[1\] Tile_X0Y0_DSP_top/J_l_GH_BEG\[1\]
+ Tile_X0Y0_DSP_top/ConfigBits\[138\] Tile_X0Y0_DSP_top/ConfigBits\[139\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[13\] sky130_fd_sc_hd__mux4_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1656_ Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/A Tile_X0Y1_DSP_bot/ConfigBits\[4\]
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1657_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1658_/A
+ sky130_fd_sc_hd__a21oi_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1587_ Tile_X0Y1_DSP_bot_Inst_MULADD__1587_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1587_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1595_/B sky130_fd_sc_hd__nor2_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_data_outbuf_17__0_ Tile_X0Y1_DSP_bot_data_inbuf_17__0_/X VGND VGND
+ VPWR VPWR net639 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[0\] net1 net133 Tile_X0Y1_bot2top\[4\] Tile_X0Y0_DSP_top/ConfigBits\[22\]
+ Tile_X0Y0_DSP_top/ConfigBits\[23\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_S4BEG_outbuf_6__0_ Tile_X0Y1_DSP_bot/S4BEG_i\[6\] VGND VGND VPWR
+ VPWR net695 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_W6BEG_outbuf_2__0_ ANTENNA_95/DIODE VGND VGND VPWR VPWR net559
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG0 net19
+ net99 net151 Tile_X0Y0_DSP_top/JN2BEG\[4\] Tile_X0Y0_DSP_top/ConfigBits\[158\] Tile_X0Y0_DSP_top/ConfigBits\[159\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[0\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0
+ net4 net136 Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y0_DSP_top/ConfigBits\[48\]
+ Tile_X0Y0_DSP_top/ConfigBits\[49\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_data_inbuf_19__0_ net239 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_19__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit1 net240 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[129\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit0 net49 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[310\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_86_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_152_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1510_ Tile_X0Y1_DSP_bot_Inst_MULADD__1510_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1511_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1523_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1441_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1435_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1441_/Y
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit28 net249 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[28\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit17 net237 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[17\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput280 Tile_X0Y1_FrameStrobe[9] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__buf_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1372_ Tile_X0Y1_DSP_bot_Inst_MULADD__1371_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1371_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1275_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1372_/Y
+ sky130_fd_sc_hd__a21oi_1
Xinput291 Tile_X0Y1_N2END[6] VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit27 net68 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[305\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit16 net56 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[294\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__13_ Tile_X0Y0_top2bot\[9\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C11 sky130_fd_sc_hd__buf_1
XFILLER_0_92_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput721 net721 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput710 net710 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput754 net754 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput732 net732 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput743 net743 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[6] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1708_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1708_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1708_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1639_ Tile_X0Y1_DSP_bot/C17 Tile_X0Y1_DSP_bot_Inst_MULADD__1759_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1640_/B
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y0_DSP_top_E6END_inbuf_0__0_ net25 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/E6BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_data_outbuf_31__0_ Tile_X0Y0_DSP_top_data_inbuf_31__0_/X VGND VGND
+ VPWR VPWR net454 sky130_fd_sc_hd__clkbuf_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top/JN2BEG\[4\] Tile_X0Y0_DSP_top/JN2BEG\[6\] Tile_X0Y0_DSP_top/JE2BEG\[4\]
+ Tile_X0Y0_DSP_top/JE2BEG\[6\] Tile_X0Y0_DSP_top/ConfigBits\[144\] Tile_X0Y0_DSP_top/ConfigBits\[145\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG1 Tile_X0Y1_N2BEG\[3\]
+ net16 net96 net148 Tile_X0Y0_DSP_top/ConfigBits\[200\] Tile_X0Y0_DSP_top/ConfigBits\[201\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_EFb_BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_64_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1
+ net24 net124 net138 net156 Tile_X0Y0_DSP_top/ConfigBits\[246\] Tile_X0Y0_DSP_top/ConfigBits\[247\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_outbuf_22__0_ Tile_X0Y0_DSP_top_data_inbuf_22__0_/X VGND VGND
+ VPWR VPWR net444 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__0941_ Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0934_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0942_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_50_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0872_ Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0889_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0862_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/B
+ sky130_fd_sc_hd__o21a_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit6 net77 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[92\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_92_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1424_ Tile_X0Y1_DSP_bot_Inst_MULADD__1424_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1424_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1424_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top_data_outbuf_13__0_ Tile_X0Y0_DSP_top_data_inbuf_13__0_/X VGND VGND
+ VPWR VPWR net434 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1355_ Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/Y sky130_fd_sc_hd__nand4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst1
+ net763 ANTENNA_101/DIODE Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[1\] Tile_X0Y1_DSP_bot/J2END_GH_BEG\[3\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[78\] Tile_X0Y1_DSP_bot/ConfigBits\[79\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1286_ Tile_X0Y1_DSP_bot_Inst_MULADD__1268_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1269_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1270_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1286_/Y
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_25_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_S4BEG_outbuf_2__0_ Tile_X0Y0_DSP_top/S4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_S4BEG\[2\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4
+ Tile_X0Y1_DSP_bot/ConfigBits\[356\] Tile_X0Y1_DSP_bot/ConfigBits\[357\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2
+ wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[110\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[111\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
Xoutput562 net562 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput551 net551 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[4] sky130_fd_sc_hd__clkbuf_4
Xoutput540 net540 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput573 net573 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput584 net584 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput595 net595 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit4 net255 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[228\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[1\] Tile_X0Y1_N2BEGb\[3\] Tile_X0Y1_N4BEG\[3\] net8 Tile_X0Y0_DSP_top/ConfigBits\[286\]
+ Tile_X0Y0_DSP_top/ConfigBits\[287\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_E6END_inbuf_0__0_ net205 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/E6BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit16 net236 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[48\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit27 net248 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[59\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_107_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit15 net55 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[325\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit26 net67 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[336\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_130_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1140_ Tile_X0Y1_DSP_bot_Inst_MULADD__1140_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1140_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1140_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_160 Tile_X0Y0_SS4BEG\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1071_ Tile_X0Y1_DSP_bot_Inst_MULADD__1072_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1072_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1070_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1073_/A
+ sky130_fd_sc_hd__a21boi_1
XANTENNA_193 Tile_X0Y0_SS4BEG\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 ANTENNA_183/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_171 Tile_X0Y1_N1BEG\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_28_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0924_ Tile_X0Y1_DSP_bot_Inst_MULADD__1252_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0922_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0923_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0950_/A
+ sky130_fd_sc_hd__o21a_1
XTile_X0Y0_DSP_top_strobe_outbuf_6__0_ Tile_X0Y0_DSP_top_strobe_inbuf_6__0_/X VGND
+ VGND VPWR VPWR net478 sky130_fd_sc_hd__buf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0855_ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1
+ net201 Tile_X0Y0_S2BEGb\[4\] net342 net354 Tile_X0Y1_DSP_bot/ConfigBits\[268\] Tile_X0Y1_DSP_bot/ConfigBits\[269\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1407_ Tile_X0Y1_DSP_bot_Inst_MULADD__1407_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1407_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1407_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1411_/B
+ sky130_fd_sc_hd__and3_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1338_ Tile_X0Y1_DSP_bot_Inst_MULADD__1249_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1337_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1339_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1338_/Y
+ sky130_fd_sc_hd__a21oi_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1269_ Tile_X0Y1_DSP_bot_Inst_MULADD__1093_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1095_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/B Tile_X0Y1_DSP_bot_Inst_MULADD__0895_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1269_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_108_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__61_ net150 VGND VGND VPWR VPWR net552
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_data_inbuf_3__0_ net254 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_3__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_NN4END_inbuf_8__0_ Tile_X0Y1_NN4BEG\[12\] VGND VGND VPWR VPWR ANTENNA_79/DIODE
+ sky130_fd_sc_hd__buf_2
Xoutput392 net392 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[6] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_S4BEG0 net204 Tile_X0Y0_S2BEGb\[2\]
+ Tile_X0Y0_S4BEG\[1\] Tile_X0Y1_DSP_bot/Q0 Tile_X0Y1_DSP_bot/ConfigBits\[70\] Tile_X0Y1_DSP_bot/ConfigBits\[71\]
+ VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit19 net59 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[233\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_E1BEG2 Tile_X0Y1_bot2top\[5\]
+ Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[1\] ANTENNA_61/DIODE Tile_X0Y0_DSP_top/J_l_GH_BEG\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[32\] Tile_X0Y0_DSP_top/ConfigBits\[33\] VGND VGND
+ VPWR VPWR net384 sky130_fd_sc_hd__mux4_1
XFILLER_0_103_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit9 net80 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[191\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_WW4BEG_outbuf_4__0_ Tile_X0Y0_DSP_top/WW4BEG_i\[4\] VGND VGND VPWR
+ VPWR net577 sky130_fd_sc_hd__clkbuf_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[308\] Tile_X0Y0_DSP_top/ConfigBits\[309\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JE2BEG\[7\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1123_ Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/A sky130_fd_sc_hd__buf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0
+ net283 net291 net183 net191 Tile_X0Y1_DSP_bot/ConfigBits\[308\] Tile_X0Y1_DSP_bot/ConfigBits\[309\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1054_ Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1054_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1054_/X
+ sky130_fd_sc_hd__and3_1
XFILLER_0_75_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2
+ net764 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[320\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[321\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap764 max_cap764/A VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__clkbuf_8
XTile_X0Y1_DSP_bot_Inst_MULADD__0907_ Tile_X0Y1_DSP_bot_Inst_MULADD__0906_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0906_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0906_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0907_/Y
+ sky130_fd_sc_hd__o21ai_1
Xinput109 Tile_X0Y0_S4END[2] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG0 net300
+ net200 Tile_X0Y0_S2BEG\[7\] net353 Tile_X0Y1_DSP_bot/ConfigBits\[216\] Tile_X0Y1_DSP_bot/ConfigBits\[217\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[0\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit15 net235 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[79\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit26 net247 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[90\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit7 net258 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[327\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_S1BEG3 Tile_X0Y1_DSP_bot/Q7
+ Tile_X0Y1_DSP_bot/J2MID_ABb_BEG\[2\] Tile_X0Y1_DSP_bot/JE2BEG\[2\] Tile_X0Y1_DSP_bot/J_l_AB_BEG\[0\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[68\] Tile_X0Y1_DSP_bot/ConfigBits\[69\] VGND VGND
+ VPWR VPWR net666 sky130_fd_sc_hd__mux4_1
XFILLER_0_2_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit25 net66 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[367\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit14 net54 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[356\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_inbuf_14__0_ net266 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_14__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_60 ANTENNA_60/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_71 ANTENNA_73/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 ANTENNA_86/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 ANTENNA_93/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__44_ net97 VGND VGND VPWR VPWR Tile_X0Y0_S2BEGb\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_N4END_inbuf_4__0_ Tile_X0Y1_N4BEG\[8\] VGND VGND VPWR VPWR ANTENNA_207/DIODE
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_159_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1741_ net333 Tile_X0Y1_DSP_bot/B7 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1741_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[1\] Tile_X0Y1_N2BEGb\[5\] net2 net10 Tile_X0Y0_DSP_top/ConfigBits\[358\]
+ Tile_X0Y0_DSP_top/ConfigBits\[359\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1672_ Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1672_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1672_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1706_/D
+ sky130_fd_sc_hd__nor3_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1106_ Tile_X0Y1_DSP_bot_Inst_MULADD__1736_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1175_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1106_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_118_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1037_ Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1036_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1043_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput91 Tile_X0Y0_S2END[6] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit18 net58 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[264\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit29 net70 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[275\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput80 Tile_X0Y0_FrameData[9] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_4
XFILLER_0_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot7 Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[3\]
+ Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[3\] Tile_X0Y0_DSP_top/J2END_CD_BEG\[3\] Tile_X0Y0_DSP_top/J_l_CD_BEG\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[126\] Tile_X0Y0_DSP_top/ConfigBits\[127\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[7\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_WW4END_inbuf_0__0_ net376 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/WW4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__27_ Tile_X0Y1_N2BEG\[3\] VGND VGND
+ VPWR VPWR net497 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit9 net80 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[31\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_strobe_inbuf_7__0_ net278 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_7__0_/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_N4END_inbuf_4__0_ net315 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/N4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_130_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit24 net65 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[398\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_95_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1724_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1724_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1724_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit13 net53 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[387\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot14 Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[2\] ANTENNA_206/DIODE Tile_X0Y0_DSP_top/J_l_GH_BEG\[2\]
+ Tile_X0Y0_DSP_top/ConfigBits\[140\] Tile_X0Y0_DSP_top/ConfigBits\[141\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[14\] sky130_fd_sc_hd__mux4_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1655_ Tile_X0Y1_DSP_bot_Inst_MULADD__1651_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1652_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/C sky130_fd_sc_hd__a22oi_2
XFILLER_0_95_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1586_ Tile_X0Y1_DSP_bot_Inst_MULADD__1587_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1587_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1595_/A sky130_fd_sc_hd__and2_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[8\] Tile_X0Y0_DSP_top/J2MID_EFb_BEG\[1\] Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2END_CD_BEG\[1\] Tile_X0Y0_DSP_top/ConfigBits\[22\] Tile_X0Y0_DSP_top/ConfigBits\[23\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__89_ Tile_X0Y1_DSP_bot/Q13 VGND VGND
+ VPWR VPWR Tile_X0Y1_bot2top\[3\] sky130_fd_sc_hd__buf_12
XFILLER_0_44_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG1 Tile_X0Y1_N2BEG\[2\]
+ net15 net147 Tile_X0Y0_DSP_top/JE2BEG\[4\] Tile_X0Y0_DSP_top/ConfigBits\[160\] Tile_X0Y0_DSP_top/ConfigBits\[161\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[1\] sky130_fd_sc_hd__mux4_1
XFILLER_0_161_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[5\]
+ Tile_X0Y0_DSP_top/ConfigBits\[48\] Tile_X0Y0_DSP_top/ConfigBits\[49\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit2 net251 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[130\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit1 net60 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[311\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0
+ net281 net285 net181 net185 Tile_X0Y1_DSP_bot/ConfigBits\[380\] Tile_X0Y1_DSP_bot/ConfigBits\[381\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1440_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1269_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1435_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1440_/X sky130_fd_sc_hd__o211a_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0
+ Tile_X0Y1_N2BEGb\[4\] net3 net9 net21 Tile_X0Y0_DSP_top/ConfigBits\[322\] Tile_X0Y0_DSP_top/ConfigBits\[323\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit18 net238 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[18\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit29 net250 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[29\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput281 Tile_X0Y1_N1END[0] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__buf_4
Xinput270 Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1371_ Tile_X0Y1_DSP_bot_Inst_MULADD__1371_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1371_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1371_/Y sky130_fd_sc_hd__nor2_1
Xinput292 Tile_X0Y1_N2END[7] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__buf_2
XFILLER_0_157_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit17 net57 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[295\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit28 net69 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[306\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__12_ Tile_X0Y0_top2bot\[8\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput700 net700 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput711 net711 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput733 net733 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[6] sky130_fd_sc_hd__clkbuf_4
Xoutput722 net722 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput744 net744 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput755 net755 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1707_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1707_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1707_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1638_ Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1700_/B sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1569_ Tile_X0Y1_DSP_bot_Inst_MULADD__1541_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1545_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1565_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1567_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1593_/B sky130_fd_sc_hd__o211a_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top/JS2BEG\[4\] Tile_X0Y0_DSP_top/JS2BEG\[6\] Tile_X0Y0_DSP_top/JW2BEG\[4\]
+ Tile_X0Y0_DSP_top/JW2BEG\[6\] Tile_X0Y0_DSP_top/ConfigBits\[144\] Tile_X0Y0_DSP_top/ConfigBits\[145\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG2 Tile_X0Y1_N2BEG\[5\]
+ net18 net98 net150 Tile_X0Y0_DSP_top/ConfigBits\[202\] Tile_X0Y0_DSP_top/ConfigBits\[203\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_EFb_BEG\[2\] sky130_fd_sc_hd__mux4_1
XFILLER_0_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[246\] Tile_X0Y0_DSP_top/ConfigBits\[247\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_strobe_inbuf_3__0_ Tile_X0Y1_FrameStrobe_O\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_3__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0940_ Tile_X0Y1_DSP_bot_Inst_MULADD__0888_/X Tile_X0Y1_DSP_bot_Inst_MULADD__0889_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0934_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0942_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_0_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__0871_ Tile_X0Y1_DSP_bot_Inst_MULADD__1175_/B Tile_X0Y1_DSP_bot/B0
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0854_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0875_/A
+ sky130_fd_sc_hd__a21boi_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit7 net78 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[93\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1423_ Tile_X0Y1_DSP_bot_Inst_MULADD__1403_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1422_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1407_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1424_/B
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1354_ Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/C Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1354_/Y sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1285_ Tile_X0Y1_DSP_bot_Inst_MULADD__1285_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1285_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_58_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_NN4BEG_outbuf_7__0_ ANTENNA_181/DIODE VGND VGND VPWR VPWR net531
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[356\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[357\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput530 net530 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput563 net563 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput552 net552 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput541 net541 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3
+ ANTENNA_101/DIODE Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[1\] ANTENNA_105/DIODE Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[1\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[110\] Tile_X0Y1_DSP_bot/ConfigBits\[111\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
Xoutput574 net574 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput585 net585 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput596 net596 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_157_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit5 net256 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[229\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1
+ net24 net88 net140 net156 Tile_X0Y0_DSP_top/ConfigBits\[286\] Tile_X0Y0_DSP_top/ConfigBits\[287\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0
+ net284 net292 net184 net192 Tile_X0Y1_DSP_bot/ConfigBits\[344\] Tile_X0Y1_DSP_bot/ConfigBits\[345\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit17 net237 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[49\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_64_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit28 net249 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[60\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_134_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit16 net56 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[326\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit27 net68 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[337\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[0\] net1 net133 Tile_X0Y1_bot2top\[4\] Tile_X0Y0_DSP_top/ConfigBits\[78\]
+ Tile_X0Y0_DSP_top/ConfigBits\[79\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_NN4BEG_outbuf_0__0_ Tile_X0Y1_DSP_bot/NN4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y1_NN4BEG\[0\] sky130_fd_sc_hd__buf_1
XTile_X0Y1_DSP_bot_SS4END_inbuf_2__0_ Tile_X0Y0_SS4BEG\[6\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/SS4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_161 Tile_X0Y0_SS4BEG\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_150 net482 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1070_ Tile_X0Y1_DSP_bot_Inst_MULADD__1069_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1711_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1252_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1070_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_194 Tile_X0Y0_SS4BEG\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_172 Tile_X0Y1_N1BEG\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_183 ANTENNA_183/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_SS4BEG_outbuf_3__0_ Tile_X0Y1_DSP_bot/SS4BEG_i\[3\] VGND VGND VPWR
+ VPWR net708 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0923_ Tile_X0Y1_DSP_bot_Inst_MULADD__1252_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1709_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0923_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_51_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0854_ Tile_X0Y1_DSP_bot_Inst_MULADD__0854_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0854_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_11_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[268\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[269\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 Tile_X0Y0_E1END[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1406_ Tile_X0Y1_DSP_bot_Inst_MULADD__1407_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1407_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1407_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1411_/A
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG0 net299
+ net199 net352 Tile_X0Y1_DSP_bot/JN2BEG\[5\] Tile_X0Y1_DSP_bot/ConfigBits\[176\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[177\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1337_ Tile_X0Y1_DSP_bot_Inst_MULADD__1147_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1336_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1171_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1337_/X
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1268_ Tile_X0Y1_DSP_bot_Inst_MULADD__1268_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/D sky130_fd_sc_hd__buf_4
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1199_ Tile_X0Y1_DSP_bot_Inst_MULADD__0895_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1189_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1289_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_116_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__60_ net149 VGND VGND VPWR VPWR net551
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput393 net393 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput382 net382 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[0] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_S4BEG1 net201 Tile_X0Y0_S2BEGb\[3\]
+ Tile_X0Y0_S4BEG\[2\] net764 Tile_X0Y1_DSP_bot/ConfigBits\[72\] Tile_X0Y1_DSP_bot/ConfigBits\[73\]
+ VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__mux4_1
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_E1BEG3 Tile_X0Y1_bot2top\[6\]
+ Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[2\] Tile_X0Y0_DSP_top/JN2BEG\[2\] ANTENNA_65/DIODE
+ Tile_X0Y0_DSP_top/ConfigBits\[34\] Tile_X0Y0_DSP_top/ConfigBits\[35\] VGND VGND
+ VPWR VPWR net385 sky130_fd_sc_hd__mux4_1
XFILLER_0_33_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_EE4END_inbuf_1__0_ net224 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/EE4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_WW4END_inbuf_9__0_ net169 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/WW4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1122_ Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/A Tile_X0Y1_DSP_bot/B6
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1121_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/C
+ sky130_fd_sc_hd__o21a_4
XFILLER_0_28_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[0\] Tile_X0Y0_S1BEG\[2\] Tile_X0Y0_S2BEGb\[6\] net336 Tile_X0Y1_DSP_bot/ConfigBits\[308\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[309\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1053_ Tile_X0Y1_DSP_bot_Inst_MULADD__1051_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1052_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1053_/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[320\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[321\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0906_ Tile_X0Y1_DSP_bot_Inst_MULADD__0906_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0906_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0906_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/D
+ sky130_fd_sc_hd__nor3_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG1 net296
+ net196 Tile_X0Y0_S2BEG\[3\] net349 Tile_X0Y1_DSP_bot/ConfigBits\[218\] Tile_X0Y1_DSP_bot/ConfigBits\[219\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit27 net248 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[91\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit16 net236 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[80\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit8 net259 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[328\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit26 net67 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[368\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit15 net55 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[357\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_50 Tile_X0Y1_FrameStrobe_O\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 ANTENNA_86/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 ANTENNA_61/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_72 ANTENNA_73/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_94 ANTENNA_94/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__43_ net96 VGND VGND VPWR VPWR Tile_X0Y0_S2BEGb\[3\]
+ sky130_fd_sc_hd__clkbuf_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1740_ net333 Tile_X0Y1_DSP_bot/B6 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1740_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1
+ net82 net84 net90 net134 Tile_X0Y0_DSP_top/ConfigBits\[358\] Tile_X0Y0_DSP_top/ConfigBits\[359\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1671_ Tile_X0Y1_DSP_bot/clr VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/A
+ sky130_fd_sc_hd__clkbuf_4
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_WW4END_inbuf_10__0_ net170 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/WW4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_E6BEG_outbuf_5__0_ Tile_X0Y1_DSP_bot/E6BEG_i\[5\] VGND VGND VPWR
+ VPWR net610 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1105_ Tile_X0Y1_DSP_bot_Inst_MULADD__1092_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1096_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1100_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/B
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_158_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1036_ Tile_X0Y1_DSP_bot_Inst_MULADD__1034_/X Tile_X0Y1_DSP_bot/B5
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1035_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1036_/Y
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_114_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput81 Tile_X0Y0_S1END[0] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_4
Xinput70 Tile_X0Y0_FrameData[29] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit19 net59 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[265\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput92 Tile_X0Y0_S2END[7] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_N4BEG_outbuf_11__0_ ANTENNA_73/DIODE VGND VGND VPWR VPWR net504
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_S4END_inbuf_7__0_ net103 VGND VGND VPWR VPWR ANTENNA_92/DIODE sky130_fd_sc_hd__buf_2
XFILLER_0_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot8 Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[0\]
+ ANTENNA_177/DIODE Tile_X0Y0_DSP_top/J2END_EF_BEG\[0\] Tile_X0Y0_DSP_top/J_l_EF_BEG\[0\]
+ Tile_X0Y0_DSP_top/ConfigBits\[128\] Tile_X0Y0_DSP_top/ConfigBits\[129\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[8\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__26_ Tile_X0Y1_N2BEG\[2\] VGND VGND
+ VPWR VPWR net496 sky130_fd_sc_hd__buf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[3\] Tile_X0Y1_N2BEGb\[7\] net4 net12 Tile_X0Y0_DSP_top/ConfigBits\[270\]
+ Tile_X0Y0_DSP_top/ConfigBits\[271\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit14 net54 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[388\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1723_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1723_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1723_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit25 net66 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[399\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot15 Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[3\]
+ Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[3\] Tile_X0Y0_DSP_top/J2END_GH_BEG\[3\] Tile_X0Y0_DSP_top/J_l_GH_BEG\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[142\] Tile_X0Y0_DSP_top/ConfigBits\[143\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[15\] sky130_fd_sc_hd__mux4_1
XFILLER_0_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1654_ Tile_X0Y1_DSP_bot_Inst_MULADD__1665_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1643_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1645_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/B
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_EE4BEG_outbuf_10__0_ ANTENNA_175/DIODE VGND VGND VPWR VPWR net415
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1585_ Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1565_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1587_/B
+ sky130_fd_sc_hd__o21ai_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__88_ Tile_X0Y1_DSP_bot/Q12 VGND VGND
+ VPWR VPWR Tile_X0Y1_bot2top\[2\] sky130_fd_sc_hd__buf_12
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1019_ Tile_X0Y1_DSP_bot_Inst_MULADD__1018_/Y Tile_X0Y1_DSP_bot/A5
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1014_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1019_/Y
+ sky130_fd_sc_hd__a21boi_4
XFILLER_0_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG2 Tile_X0Y1_N2BEG\[4\]
+ net17 net97 Tile_X0Y0_DSP_top/JS2BEG\[4\] Tile_X0Y0_DSP_top/ConfigBits\[162\] Tile_X0Y0_DSP_top/ConfigBits\[163\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[48\] Tile_X0Y0_DSP_top/ConfigBits\[49\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit3 net254 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[131\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit2 net71 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[312\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[0\] Tile_X0Y0_S1BEG\[2\] Tile_X0Y0_S2BEGb\[0\] net334 Tile_X0Y1_DSP_bot/ConfigBits\[380\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[381\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_S4END_inbuf_7__0_ Tile_X0Y0_S4BEG\[11\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/S4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_105_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst0
+ net299 net193 net199 Tile_X0Y0_S2BEG\[0\] Tile_X0Y1_DSP_bot/ConfigBits\[156\] Tile_X0Y1_DSP_bot/ConfigBits\[157\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit30 net72 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[20\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__09_ net14 VGND VGND VPWR VPWR net395
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1
+ net89 net101 net141 net173 Tile_X0Y0_DSP_top/ConfigBits\[322\] Tile_X0Y0_DSP_top/ConfigBits\[323\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit19 net239 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[19\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput271 Tile_X0Y1_FrameStrobe[19] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_1
Xinput260 Tile_X0Y1_FrameData[9] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1370_ Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1284_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1368_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1369_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1370_/Y sky130_fd_sc_hd__o2bb2ai_4
Xinput293 Tile_X0Y1_N2MID[0] VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_4
Xinput282 Tile_X0Y1_N1END[1] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__buf_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit18 net58 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[296\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit29 net70 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[307\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_E6BEG_outbuf_1__0_ Tile_X0Y0_DSP_top/E6BEG_i\[1\] VGND VGND VPWR
+ VPWR net405 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__11_ Tile_X0Y0_top2bot\[7\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/B7 sky130_fd_sc_hd__buf_2
XFILLER_0_73_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_EE4BEG_outbuf_3__0_ ANTENNA_100/DIODE VGND VGND VPWR VPWR net624
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG0 Tile_X0Y1_N4BEG\[3\]
+ net33 net110 Tile_X0Y0_DSP_top/JN2BEG\[4\] Tile_X0Y0_DSP_top/ConfigBits\[398\] Tile_X0Y0_DSP_top/ConfigBits\[399\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_GH_BEG\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_121_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput701 net701 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput712 net712 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput734 net734 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput723 net723 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput745 net745 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput756 net756 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1706_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1706_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1706_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1637_ Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1637_/B
+ Tile_X0Y1_DSP_bot/ConfigBits\[4\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1645_/A
+ sky130_fd_sc_hd__nand3_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1568_ Tile_X0Y1_DSP_bot_Inst_MULADD__1565_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1567_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1541_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1545_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1593_/A sky130_fd_sc_hd__a211oi_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1499_ Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1441_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1499_/Y sky130_fd_sc_hd__a31oi_2
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG3 Tile_X0Y1_N2BEG\[1\]
+ net14 net94 net146 Tile_X0Y0_DSP_top/ConfigBits\[204\] Tile_X0Y0_DSP_top/ConfigBits\[205\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_EFb_BEG\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[246\] Tile_X0Y0_DSP_top/ConfigBits\[247\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0870_ Tile_X0Y1_DSP_bot/ConfigBits\[1\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1175_/B sky130_fd_sc_hd__inv_2
XFILLER_0_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit8 net79 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[94\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1422_ Tile_X0Y1_DSP_bot_Inst_MULADD__1422_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1422_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1422_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1353_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1353_/Y
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1284_ Tile_X0Y1_DSP_bot_Inst_MULADD__1285_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1285_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1283_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1284_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_116_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[358\] Tile_X0Y1_DSP_bot/ConfigBits\[359\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JW2BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_61_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput520 net520 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput531 net531 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput553 net553 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[6] sky130_fd_sc_hd__clkbuf_4
Xoutput542 net542 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[112\] Tile_X0Y1_DSP_bot/ConfigBits\[113\] VGND VGND
+ VPWR VPWR net736 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0999_ Tile_X0Y1_DSP_bot_Inst_MULADD__0998_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1710_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1252_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1002_/C
+ sky130_fd_sc_hd__mux2_1
Xoutput564 net564 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput575 net575 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput586 net586 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[3] sky130_fd_sc_hd__buf_2
Xoutput597 net597 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_157_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit6 net257 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[230\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[286\] Tile_X0Y0_DSP_top/ConfigBits\[287\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[3\] Tile_X0Y0_S2BEGb\[7\] net335 net337 Tile_X0Y1_DSP_bot/ConfigBits\[344\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[345\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_WW4BEG_outbuf_11__0_ Tile_X0Y0_DSP_top/WW4BEG_i\[11\] VGND VGND
+ VPWR VPWR net569 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit18 net238 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[50\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_64_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_N4BEG_outbuf_9__0_ Tile_X0Y1_DSP_bot/N4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N4BEG\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit29 net250 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[61\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit17 net57 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[327\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit28 net69 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[338\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[8\] Tile_X0Y0_DSP_top/J2MID_EFb_BEG\[1\] Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2END_CD_BEG\[3\] Tile_X0Y0_DSP_top/ConfigBits\[78\] Tile_X0Y0_DSP_top/ConfigBits\[79\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG0 Tile_X0Y1_N2BEGb\[7\]
+ net41 net92 net144 Tile_X0Y0_DSP_top/ConfigBits\[230\] Tile_X0Y0_DSP_top/ConfigBits\[231\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_EF_BEG\[0\] sky130_fd_sc_hd__mux4_1
XANTENNA_151 net495 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_140 net314 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 Tile_X0Y1_N2BEG\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_184 ANTENNA_184/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_162 Tile_X0Y0_SS4BEG\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_195 Tile_X0Y0_SS4BEG\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0922_ Tile_X0Y1_DSP_bot_Inst_MULADD__1459_/S Tile_X0Y1_DSP_bot/C3
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0921_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0922_/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_140_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0853_ Tile_X0Y1_DSP_bot/ConfigBits\[1\] Tile_X0Y1_DSP_bot/B0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0854_/B sky130_fd_sc_hd__or2b_4
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_inbuf_0__0_ net49 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_0__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[268\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[269\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
Xinput2 Tile_X0Y0_E1END[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1405_ Tile_X0Y1_DSP_bot_Inst_MULADD__1395_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1397_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1424_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1407_/C
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[149\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR Tile_X0Y0_top2bot\[17\] sky130_fd_sc_hd__o21ai_4
XFILLER_0_127_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG1 net295
+ net195 Tile_X0Y0_S2BEG\[2\] Tile_X0Y1_DSP_bot/JE2BEG\[5\] Tile_X0Y1_DSP_bot/ConfigBits\[178\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[179\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1336_ Tile_X0Y1_DSP_bot_Inst_MULADD__1239_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1335_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1248_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1336_/Y
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1267_ Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1228_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1220_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1313_/A
+ sky130_fd_sc_hd__a21oi_1
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1198_ Tile_X0Y1_DSP_bot_Inst_MULADD__1099_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1192_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/D VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1289_/A
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_116_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_strobe_outbuf_17__0_ Tile_X0Y0_DSP_top_strobe_inbuf_17__0_/X VGND
+ VGND VPWR VPWR net470 sky130_fd_sc_hd__clkbuf_1
Xoutput394 net394 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput383 net383 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[1] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_S4BEG2 Tile_X0Y0_S2BEGb\[0\]
+ Tile_X0Y0_S4BEG\[3\] net357 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/ConfigBits\[74\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[75\] VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_W6BEG_outbuf_9__0_ Tile_X0Y1_DSP_bot/W6BEG_i\[9\] VGND VGND VPWR
+ VPWR net746 sky130_fd_sc_hd__clkbuf_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_data_outbuf_7__0_ Tile_X0Y0_DSP_top_data_inbuf_7__0_/X VGND VGND
+ VPWR VPWR net459 sky130_fd_sc_hd__clkbuf_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1121_ Tile_X0Y1_DSP_bot_Inst_MULADD__1740_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1121_/X sky130_fd_sc_hd__or2b_2
XFILLER_0_75_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 net764 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[308\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[309\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1052_ Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0989_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0984_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1052_/X
+ sky130_fd_sc_hd__o21a_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[322\] Tile_X0Y1_DSP_bot/ConfigBits\[323\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JS2BEG\[0\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0905_ Tile_X0Y1_DSP_bot_Inst_MULADD__0900_/X Tile_X0Y1_DSP_bot_Inst_MULADD__0902_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0906_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG2 net298
+ net198 Tile_X0Y0_S2BEG\[5\] net351 Tile_X0Y1_DSP_bot/ConfigBits\[220\] Tile_X0Y1_DSP_bot/ConfigBits\[221\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[2\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit28 net249 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[92\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit17 net237 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[81\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit9 net260 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[329\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_NN4END_inbuf_2__0_ net329 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/NN4BEG_i\[2\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_78_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1319_ Tile_X0Y1_DSP_bot_Inst_MULADD__1306_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1306_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1291_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1297_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1319_/X sky130_fd_sc_hd__a22o_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit27 net68 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[369\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit16 net56 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[358\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_93_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_40 Tile_X0Y1_FrameStrobe_O\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 ANTENNA_86/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 Tile_X0Y1_FrameStrobe_O\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_N4BEG_outbuf_5__0_ ANTENNA_76/DIODE VGND VGND VPWR VPWR net513
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_73 ANTENNA_73/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 ANTENNA_63/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[41\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__o21ai_1
XANTENNA_95 ANTENNA_95/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__42_ net95 VGND VGND VPWR VPWR Tile_X0Y0_S2BEGb\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit0 net49 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[214\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_data_outbuf_7__0_ Tile_X0Y1_DSP_bot_data_inbuf_7__0_/X VGND VGND
+ VPWR VPWR net660 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[358\] Tile_X0Y0_DSP_top/ConfigBits\[359\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1670_ Tile_X0Y1_DSP_bot_Inst_MULADD__1258_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1661_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1669_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q19
+ sky130_fd_sc_hd__o21ai_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_data_outbuf_29__0_ Tile_X0Y1_DSP_bot_data_inbuf_29__0_/X VGND VGND
+ VPWR VPWR net652 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1104_ Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1100_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1103_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1104_/Y
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_75_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1035_ Tile_X0Y1_DSP_bot_Inst_MULADD__1739_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1175_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1035_/X sky130_fd_sc_hd__or2_2
XFILLER_0_133_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput82 Tile_X0Y0_S1END[1] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
Xinput60 Tile_X0Y0_FrameData[1] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_8
Xinput71 Tile_X0Y0_FrameData[2] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_8
Xinput93 Tile_X0Y0_S2MID[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_S4BEG_outbuf_9__0_ ANTENNA_110/DIODE VGND VGND VPWR VPWR net698
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_W6BEG_outbuf_5__0_ Tile_X0Y0_DSP_top/W6BEG_i\[5\] VGND VGND VPWR
+ VPWR net562 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_top2bot9 Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2MID_EFb_BEG\[1\] Tile_X0Y0_DSP_top/J2END_EF_BEG\[1\] Tile_X0Y0_DSP_top/J_l_EF_BEG\[1\]
+ Tile_X0Y0_DSP_top/ConfigBits\[130\] Tile_X0Y0_DSP_top/ConfigBits\[131\] VGND VGND
+ VPWR VPWR Tile_X0Y0_top2bot\[9\] sky130_fd_sc_hd__mux4_1
XFILLER_0_132_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__25_ Tile_X0Y1_N2BEG\[1\] VGND VGND
+ VPWR VPWR net495 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1
+ net84 net92 net134 net136 Tile_X0Y0_DSP_top/ConfigBits\[270\] Tile_X0Y0_DSP_top/ConfigBits\[271\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1722_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1722_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1722_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit15 net55 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[389\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit26 net67 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[400\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1653_ Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/A
+ sky130_fd_sc_hd__nand3_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1584_ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1180_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1587_/A sky130_fd_sc_hd__a211o_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__87_ Tile_X0Y1_DSP_bot/Q11 VGND VGND
+ VPWR VPWR Tile_X0Y1_bot2top\[1\] sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1018_ Tile_X0Y1_DSP_bot/ConfigBits\[0\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1018_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_161_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG3 Tile_X0Y1_N2BEG\[0\]
+ net93 net145 Tile_X0Y0_DSP_top/JW2BEG\[4\] Tile_X0Y0_DSP_top/ConfigBits\[164\] Tile_X0Y0_DSP_top/ConfigBits\[165\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[3\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[1\] Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[1\] Tile_X0Y0_DSP_top/J2MID_EFb_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[1\] Tile_X0Y0_DSP_top/ConfigBits\[48\] Tile_X0Y0_DSP_top/ConfigBits\[49\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_E6END_inbuf_3__0_ net28 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/E6BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit4 net255 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[132\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 net764 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[380\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[381\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit3 net74 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[313\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit0 net49 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[54\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_strobe_inbuf_11__0_ Tile_X0Y1_FrameStrobe_O\[11\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_11__0_/X sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[47\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst1
+ net346 Tile_X0Y1_DSP_bot/JN2BEG\[2\] Tile_X0Y1_DSP_bot/JN2BEG\[3\] Tile_X0Y1_DSP_bot/JE2BEG\[2\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[156\] Tile_X0Y1_DSP_bot/ConfigBits\[157\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__08_ net13 VGND VGND VPWR VPWR net394
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit31 net73 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[21\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit20 net61 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[10\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_156_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[322\] Tile_X0Y0_DSP_top/ConfigBits\[323\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_data_outbuf_25__0_ Tile_X0Y0_DSP_top_data_inbuf_25__0_/X VGND VGND
+ VPWR VPWR net447 sky130_fd_sc_hd__clkbuf_1
Xinput261 Tile_X0Y1_FrameStrobe[0] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__buf_8
Xinput272 Tile_X0Y1_FrameStrobe[1] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_16
Xinput250 Tile_X0Y1_FrameData[29] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_8
Xinput294 Tile_X0Y1_N2MID[1] VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__buf_2
Xinput283 Tile_X0Y1_N1END[2] VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__buf_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit19 net59 Tile_X0Y1_FrameStrobe_O\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[297\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame3_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__10_ Tile_X0Y0_top2bot\[6\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/B6 sky130_fd_sc_hd__buf_2
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput702 net702 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG1 Tile_X0Y1_N4BEG\[2\]
+ net125 net139 Tile_X0Y0_DSP_top/JE2BEG\[4\] Tile_X0Y0_DSP_top/ConfigBits\[400\]
+ Tile_X0Y0_DSP_top/ConfigBits\[401\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_GH_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput724 net724 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput713 net713 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput735 net735 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput757 net757 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput746 net746 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1705_ Tile_X0Y1_DSP_bot_Inst_MULADD__1666_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1668_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1725_/D
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1636_ Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1722_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1700_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1635_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q16 sky130_fd_sc_hd__a22o_1
XTile_X0Y0_DSP_top_data_outbuf_16__0_ Tile_X0Y0_DSP_top_data_inbuf_16__0_/X VGND VGND
+ VPWR VPWR net437 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1567_ Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1567_/X sky130_fd_sc_hd__a311o_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1498_ Tile_X0Y1_DSP_bot_Inst_MULADD__1490_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1491_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1494_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1498_/Y sky130_fd_sc_hd__a22oi_2
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_S4BEG_outbuf_5__0_ ANTENNA_89/DIODE VGND VGND VPWR VPWR Tile_X0Y0_S4BEG\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[248\] Tile_X0Y0_DSP_top/ConfigBits\[249\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JN2BEG\[0\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_E6END_inbuf_3__0_ net208 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/E6BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_157_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit9 net80 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[95\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1421_ Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1421_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1421_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1422_/B
+ sky130_fd_sc_hd__nand3b_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1352_ Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/B sky130_fd_sc_hd__buf_4
XFILLER_0_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1283_ Tile_X0Y1_DSP_bot_Inst_MULADD__1373_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1373_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1283_/X sky130_fd_sc_hd__a32o_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[24\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput510 net510 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_strobe_outbuf_9__0_ Tile_X0Y0_DSP_top_strobe_inbuf_9__0_/X VGND
+ VGND VPWR VPWR net481 sky130_fd_sc_hd__buf_1
Xoutput532 net532 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput521 net521 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput554 net554 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput543 net543 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[4] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0998_ Tile_X0Y1_DSP_bot/C4 Tile_X0Y1_DSP_bot_Inst_MULADD__1746_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1459_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0998_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput565 net565 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput576 net576 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput587 net587 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput598 net598 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1619_ Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1619_/Y sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit7 net258 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[231\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[286\] Tile_X0Y0_DSP_top/ConfigBits\[287\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[344\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[345\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit30 net72 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[52\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit19 net239 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[51\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_data_inbuf_6__0_ net257 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_6__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit18 net58 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[328\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit29 net70 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[339\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_outbuf_2__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_2__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[2\] sky130_fd_sc_hd__buf_8
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG1 Tile_X0Y1_N2BEGb\[3\]
+ net8 net88 net172 Tile_X0Y0_DSP_top/ConfigBits\[232\] Tile_X0Y0_DSP_top/ConfigBits\[233\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_EF_BEG\[1\] sky130_fd_sc_hd__mux4_1
XANTENNA_152 net703 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_141 net314 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_130 net184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_174 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_163 Tile_X0Y0_SS4BEG\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_185 ANTENNA_185/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_196 Tile_X0Y0_SS4BEG\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0921_ Tile_X0Y1_DSP_bot_Inst_MULADD__1745_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1459_/S
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0921_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0852_ Tile_X0Y1_DSP_bot_Inst_MULADD__1734_/Q Tile_X0Y1_DSP_bot/ConfigBits\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0854_/A sky130_fd_sc_hd__nand2_4
XTile_X0Y0_DSP_top_WW4BEG_outbuf_7__0_ Tile_X0Y0_DSP_top/WW4BEG_i\[7\] VGND VGND VPWR
+ VPWR net580 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[270\] Tile_X0Y1_DSP_bot/ConfigBits\[271\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JN2BEG\[3\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1404_ Tile_X0Y1_DSP_bot_Inst_MULADD__1395_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1403_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1424_/A
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[149\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
Xinput3 Tile_X0Y0_E1END[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG2 net297
+ Tile_X0Y0_S2BEG\[4\] net350 Tile_X0Y1_DSP_bot/JS2BEG\[5\] Tile_X0Y1_DSP_bot/ConfigBits\[180\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[181\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[2\]
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1335_ Tile_X0Y1_DSP_bot_Inst_MULADD__1135_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1242_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1244_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1335_/Y
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_143_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1266_ Tile_X0Y1_DSP_bot_Inst_MULADD__1261_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1238_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1260_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1230_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/A sky130_fd_sc_hd__o32ai_4
XFILLER_0_52_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1197_ Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1197_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_0_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput395 net395 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput384 net384 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[2] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_S4BEG3 Tile_X0Y0_S2BEGb\[1\]
+ Tile_X0Y0_S4BEG\[0\] net354 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[76\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[77\] VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_WW4BEG_outbuf_0__0_ Tile_X0Y1_DSP_bot/WW4BEG_i\[0\] VGND VGND VPWR
+ VPWR net747 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_strobe_inbuf_17__0_ net269 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_17__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG0 net188
+ Tile_X0Y0_SS4BEG\[3\] net374 Tile_X0Y1_DSP_bot/JN2BEG\[2\] Tile_X0Y1_DSP_bot/ConfigBits\[392\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[393\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_CD_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1120_ Tile_X0Y1_DSP_bot_Inst_MULADD__1026_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1062_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1120_/Y
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1051_ Tile_X0Y1_DSP_bot_Inst_MULADD__1026_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1044_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1048_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1051_/Y
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q4 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[308\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[309\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_N4END_inbuf_7__0_ Tile_X0Y1_N4BEG\[11\] VGND VGND VPWR VPWR ANTENNA_77/DIODE
+ sky130_fd_sc_hd__buf_2
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0904_ Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0892_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0893_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/B
+ sky130_fd_sc_hd__o21a_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG3 net294
+ net194 Tile_X0Y0_S2BEG\[1\] net347 Tile_X0Y1_DSP_bot/ConfigBits\[222\] Tile_X0Y1_DSP_bot/ConfigBits\[223\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_47_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit29 net250 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[93\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit18 net238 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[82\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[30\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_NN4BEG\[14\] sky130_fd_sc_hd__o21ai_2
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1318_ Tile_X0Y1_DSP_bot_Inst_MULADD__1317_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1296_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1306_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1318_/X
+ sky130_fd_sc_hd__a21o_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit17 net57 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[359\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit28 net69 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[370\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1249_ Tile_X0Y1_DSP_bot_Inst_MULADD__1246_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1248_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1171_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1249_/Y
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_41 Tile_X0Y1_FrameStrobe_O\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_30 Tile_X0Y1_FrameStrobe_O\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 ANTENNA_74/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 Tile_X0Y1_FrameStrobe_O\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_63 ANTENNA_63/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_85 ANTENNA_86/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[41\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XANTENNA_96 ANTENNA_96/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__41_ net94 VGND VGND VPWR VPWR Tile_X0Y0_S2BEGb\[1\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit1 net60 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[215\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_WW4END_inbuf_3__0_ net379 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/WW4BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_150_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[358\] Tile_X0Y0_DSP_top/ConfigBits\[359\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1103_ Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1103_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_0_158_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1034_ Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1034_/X sky130_fd_sc_hd__buf_4
XFILLER_0_16_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_N4END_inbuf_7__0_ net303 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/N4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_SS4BEG_outbuf_11__0_ Tile_X0Y0_DSP_top/SS4BEG_i\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y0_SS4BEG\[11\] sky130_fd_sc_hd__clkbuf_4
Xinput72 Tile_X0Y0_FrameData[30] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_8
Xinput50 Tile_X0Y0_FrameData[10] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_8
Xinput61 Tile_X0Y0_FrameData[20] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_6
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput94 Tile_X0Y0_S2MID[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_4
Xinput83 Tile_X0Y0_S1END[2] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_SS4BEG_outbuf_0__0_ Tile_X0Y0_DSP_top/SS4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y0_SS4BEG\[0\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_N4END_inbuf_11__0_ Tile_X0Y1_N4BEG\[15\] VGND VGND VPWR VPWR ANTENNA_73/DIODE
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__24_ Tile_X0Y1_N2BEG\[0\] VGND VGND
+ VPWR VPWR net494 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[103\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[270\] Tile_X0Y0_DSP_top/ConfigBits\[271\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1721_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1721_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit16 net56 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[390\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit27 net68 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[401\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1652_ Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1665_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1652_/X sky130_fd_sc_hd__or2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1583_ Tile_X0Y1_DSP_bot_Inst_MULADD__1583_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q13 sky130_fd_sc_hd__buf_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1017_ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1016_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1045_/A sky130_fd_sc_hd__a41oi_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__86_ Tile_X0Y1_DSP_bot/Q10 VGND VGND
+ VPWR VPWR Tile_X0Y1_bot2top\[0\] sky130_fd_sc_hd__clkbuf_16
XFILLER_0_146_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[50\] Tile_X0Y0_DSP_top/ConfigBits\[51\] VGND VGND
+ VPWR VPWR net403 sky130_fd_sc_hd__mux4_1
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit5 net256 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[133\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit4 net75 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[314\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[380\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[381\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit1 net60 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[55\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_156_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[47\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/JE2BEG\[3\] Tile_X0Y1_DSP_bot/JS2BEG\[2\] Tile_X0Y1_DSP_bot/JS2BEG\[3\]
+ Tile_X0Y1_DSP_bot/JW2BEG\[2\] Tile_X0Y1_DSP_bot/ConfigBits\[156\] Tile_X0Y1_DSP_bot/ConfigBits\[157\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__07_ Tile_X0Y0_DSP_top/JE2BEG\[7\] VGND
+ VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit21 net62 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[11\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit10 net50 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[0\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[322\] Tile_X0Y0_DSP_top/ConfigBits\[323\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
Xinput262 Tile_X0Y1_FrameStrobe[10] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__buf_8
Xinput251 Tile_X0Y1_FrameData[2] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_6
Xinput240 Tile_X0Y1_FrameData[1] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_8
Xinput295 Tile_X0Y1_N2MID[2] VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkbuf_4
Xinput284 Tile_X0Y1_N1END[3] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__buf_4
Xinput273 Tile_X0Y1_FrameStrobe[2] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__buf_8
XTile_X0Y0_DSP_top_strobe_inbuf_6__0_ Tile_X0Y1_FrameStrobe_O\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_6__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput703 net703 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG2 net24
+ net108 net174 Tile_X0Y0_DSP_top/JS2BEG\[4\] Tile_X0Y0_DSP_top/ConfigBits\[402\]
+ Tile_X0Y0_DSP_top/ConfigBits\[403\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_GH_BEG\[2\]
+ sky130_fd_sc_hd__mux4_1
Xoutput725 net725 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput714 net714 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput736 net736 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput758 net758 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput747 net747 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[0] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1704_ Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1724_/D
+ sky130_fd_sc_hd__nor3_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1635_ Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1635_/Y
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1566_ Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/Y sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1497_ Tile_X0Y1_DSP_bot_Inst_MULADD__1477_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1478_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1490_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1491_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1536_/C sky130_fd_sc_hd__o211a_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__69_ Tile_X0Y0_S2BEG\[7\] VGND VGND
+ VPWR VPWR net682 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_NN4BEG_outbuf_3__0_ Tile_X0Y1_DSP_bot/NN4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y1_NN4BEG\[3\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[109\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_SS4END_inbuf_5__0_ Tile_X0Y0_SS4BEG\[9\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/SS4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1420_ Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1422_/A
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1351_ Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1407_/B sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1282_ Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/Y sky130_fd_sc_hd__nand4_4
XFILLER_0_148_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[24\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_SS4BEG_outbuf_6__0_ Tile_X0Y1_DSP_bot/SS4BEG_i\[6\] VGND VGND VPWR
+ VPWR net711 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput500 net500 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput511 net511 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput522 net522 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput533 net533 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput544 net544 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[5] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0997_ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/C Tile_X0Y1_DSP_bot_Inst_MULADD__0995_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0996_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1002_/B sky130_fd_sc_hd__a311o_1
Xoutput566 net566 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput555 net555 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput577 net577 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput588 net588 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput599 net599 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[4] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1618_ Tile_X0Y1_DSP_bot_Inst_MULADD__1620_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1620_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1622_/A sky130_fd_sc_hd__o2111a_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1549_ Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1554_/B
+ sky130_fd_sc_hd__nand3_1
XTile_X0Y1_DSP_bot_S4BEG_outbuf_10__0_ ANTENNA_187/DIODE VGND VGND VPWR VPWR net684
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit8 net259 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[232\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst0
+ net284 net184 net337 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[25\] Tile_X0Y1_DSP_bot/ConfigBits\[26\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[288\] Tile_X0Y0_DSP_top/ConfigBits\[289\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JE2BEG\[2\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/Q5 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8
+ Tile_X0Y1_DSP_bot/ConfigBits\[344\] Tile_X0Y1_DSP_bot/ConfigBits\[345\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0
+ net284 net286 net308 net220 Tile_X0Y1_DSP_bot/ConfigBits\[288\] Tile_X0Y1_DSP_bot/ConfigBits\[289\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_S4END_inbuf_11__0_ net107 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/S4BEG_i\[11\]
+ sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit20 net61 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[42\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit31 net73 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[53\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit19 net59 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[329\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_120 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG2 Tile_X0Y1_N2BEGb\[5\]
+ net10 net124 net142 Tile_X0Y0_DSP_top/ConfigBits\[234\] Tile_X0Y0_DSP_top/ConfigBits\[235\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_EF_BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_87_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_142 net314 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_131 net184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_153 Tile_X0Y0_SS4BEG\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_175 ANTENNA_175/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 Tile_X0Y0_SS4BEG\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_197 Tile_X0Y0_SS4BEG\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_186 ANTENNA_187/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_W6END_inbuf_1__0_ net158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/W6BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__0920_ Tile_X0Y1_DSP_bot_Inst_MULADD__0920_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q2 sky130_fd_sc_hd__buf_12
XFILLER_0_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_EE4END_inbuf_4__0_ net227 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/EE4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0851_ Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/D sky130_fd_sc_hd__buf_4
XFILLER_0_87_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1403_ Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1403_/Y
+ sky130_fd_sc_hd__a21boi_4
Xinput4 Tile_X0Y0_E1END[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG3 net193
+ Tile_X0Y0_S2BEG\[0\] net346 Tile_X0Y1_DSP_bot/JW2BEG\[5\] Tile_X0Y1_DSP_bot/ConfigBits\[182\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[183\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG0 Tile_X0Y1_NN4BEG\[3\]
+ net110 net165 ANTENNA_61/DIODE Tile_X0Y0_DSP_top/ConfigBits\[374\] Tile_X0Y0_DSP_top/ConfigBits\[375\]
+ VGND VGND VPWR VPWR ANTENNA_65/DIODE sky130_fd_sc_hd__mux4_2
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1334_ Tile_X0Y1_DSP_bot_Inst_MULADD__1334_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1334_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1342_/B sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1265_ Tile_X0Y1_DSP_bot_Inst_MULADD__1264_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1248_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1171_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1246_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/A sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_19_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1196_ Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1195_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1196_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_EE4BEG_outbuf_0__0_ Tile_X0Y0_DSP_top/EE4BEG_i\[0\] VGND VGND VPWR
+ VPWR net414 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput396 net396 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[2] sky130_fd_sc_hd__clkbuf_4
Xoutput385 net385 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG1 net309
+ net187 net345 Tile_X0Y1_DSP_bot/JE2BEG\[2\] Tile_X0Y1_DSP_bot/ConfigBits\[394\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[395\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_CD_BEG\[1\]
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit0 net229 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[0\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_SS4END_inbuf_1__0_ net128 VGND VGND VPWR VPWR ANTENNA_94/DIODE
+ sky130_fd_sc_hd__buf_2
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_outbuf_12__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_12__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[12\] sky130_fd_sc_hd__clkbuf_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1050_ Tile_X0Y1_DSP_bot_Inst_MULADD__1026_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1044_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1048_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1049_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1050_/X sky130_fd_sc_hd__o211a_4
XFILLER_0_75_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[310\] Tile_X0Y1_DSP_bot/ConfigBits\[311\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JE2BEG\[5\] sky130_fd_sc_hd__mux4_2
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0903_ Tile_X0Y1_DSP_bot/ConfigBits\[1\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/A sky130_fd_sc_hd__buf_4
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_W6END_inbuf_1__0_ net359 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/W6BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit30 net72 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[84\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_44_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit19 net239 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[83\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame10_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_E6BEG_outbuf_8__0_ Tile_X0Y1_DSP_bot/E6BEG_i\[8\] VGND VGND VPWR
+ VPWR net613 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[30\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1317_ Tile_X0Y1_DSP_bot_Inst_MULADD__1315_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1284_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1273_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1317_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_154_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit18 net58 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[360\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_63_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit29 net70 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[371\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_93_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1248_ Tile_X0Y1_DSP_bot_Inst_MULADD__1248_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1248_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1248_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1248_/X
+ sky130_fd_sc_hd__and3_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1179_ Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/X sky130_fd_sc_hd__and4b_1
XANTENNA_31 Tile_X0Y1_FrameStrobe_O\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 Tile_X0Y0_SS4BEG\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_75 ANTENNA_75/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 ANTENNA_64/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 Tile_X0Y1_FrameStrobe_O\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 Tile_X0Y1_FrameStrobe_O\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_86 ANTENNA_86/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__40_ net93 VGND VGND VPWR VPWR Tile_X0Y0_S2BEGb\[0\]
+ sky130_fd_sc_hd__buf_2
XANTENNA_97 ANTENNA_97/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit2 net71 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[216\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[360\] Tile_X0Y0_DSP_top/ConfigBits\[361\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JW2BEG\[4\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_EE4END_inbuf_0__0_ net43 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/EE4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0
+ net282 net288 net188 net204 Tile_X0Y1_DSP_bot/ConfigBits\[360\] Tile_X0Y1_DSP_bot/ConfigBits\[361\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0
+ net183 net336 Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/ConfigBits\[114\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[115\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit0 net229 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[352\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1102_ Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/C Tile_X0Y1_DSP_bot_Inst_MULADD__0875_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/C sky130_fd_sc_hd__o2bb2ai_2
XFILLER_0_124_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1033_ Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/D Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/A sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_8_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput40 Tile_X0Y0_EE4END[1] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
Xinput73 Tile_X0Y0_FrameData[31] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_8
Xinput62 Tile_X0Y0_FrameData[21] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_6
Xinput51 Tile_X0Y0_FrameData[11] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput95 Tile_X0Y0_S2MID[2] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_4
Xinput84 Tile_X0Y0_S1END[3] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_2
XFILLER_0_12_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__23_ Tile_X0Y0_DSP_top/JN2BEG\[7\] VGND
+ VGND VPWR VPWR net493 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[103\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[270\] Tile_X0Y0_DSP_top/ConfigBits\[271\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1720_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1720_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit17 net57 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[391\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit28 net69 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[402\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1651_ Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/A Tile_X0Y1_DSP_bot/ConfigBits\[4\]
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1657_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1651_/X
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1582_ Tile_X0Y1_DSP_bot_Inst_MULADD__1696_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1719_/Q
+ Tile_X0Y1_DSP_bot/ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1583_/A
+ sky130_fd_sc_hd__mux2_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_E6BEG_outbuf_4__0_ Tile_X0Y0_DSP_top/E6BEG_i\[4\] VGND VGND VPWR
+ VPWR net408 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_EE4BEG_outbuf_6__0_ Tile_X0Y1_DSP_bot/EE4BEG_i\[6\] VGND VGND VPWR
+ VPWR net627 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__85_ net353 VGND VGND VPWR VPWR net734
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1016_ Tile_X0Y1_DSP_bot_Inst_MULADD__0968_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0969_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1201_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1016_/Y
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_151_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_data_inbuf_30__0_ net72 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_30__0_/X
+ sky130_fd_sc_hd__buf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit6 net257 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[134\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit5 net76 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[315\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[382\] Tile_X0Y1_DSP_bot/ConfigBits\[383\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JW2BEG\[7\] sky130_fd_sc_hd__mux4_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit2 net71 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[56\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_94_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/JW2BEG\[3\] Tile_X0Y1_DSP_bot/JW2BEG\[5\] net765 net766 Tile_X0Y1_DSP_bot/ConfigBits\[156\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[157\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_160_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__06_ Tile_X0Y0_DSP_top/JE2BEG\[6\] VGND
+ VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit22 net63 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[12\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit11 net51 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[1\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[77\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR Tile_X0Y0_SS4BEG\[13\] sky130_fd_sc_hd__o21ai_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[324\] Tile_X0Y0_DSP_top/ConfigBits\[325\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JS2BEG\[3\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_data_inbuf_21__0_ net62 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_21__0_/X
+ sky130_fd_sc_hd__clkbuf_1
Xinput263 Tile_X0Y1_FrameStrobe[11] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_8
Xinput230 Tile_X0Y1_FrameData[10] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_8
Xinput241 Tile_X0Y1_FrameData[20] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_8
Xinput252 Tile_X0Y1_FrameData[30] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0
+ net325 net181 net221 net201 Tile_X0Y1_DSP_bot/ConfigBits\[324\] Tile_X0Y1_DSP_bot/ConfigBits\[325\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
Xinput285 Tile_X0Y1_N2END[0] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_4
Xinput296 Tile_X0Y1_N2MID[3] VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkbuf_4
Xinput274 Tile_X0Y1_FrameStrobe[3] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG3 Tile_X0Y1_NN4BEG\[0\]
+ net21 net137 Tile_X0Y0_DSP_top/JW2BEG\[4\] Tile_X0Y0_DSP_top/ConfigBits\[404\] Tile_X0Y0_DSP_top/ConfigBits\[405\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_GH_BEG\[3\] sky130_fd_sc_hd__mux4_2
Xoutput726 net726 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput715 net715 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput704 net704 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput748 net748 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput759 net759 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput737 net737 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[11] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1703_ Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/B
+ sky130_fd_sc_hd__and3_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1634_ Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1700_/C sky130_fd_sc_hd__or2_1
XFILLER_0_39_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_inbuf_12__0_ net52 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_12__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1565_ Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1565_/X
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_146_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1496_ Tile_X0Y1_DSP_bot_Inst_MULADD__1496_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1496_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1496_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1505_/B
+ sky130_fd_sc_hd__nand3_2
XFILLER_0_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__68_ Tile_X0Y0_S2BEG\[6\] VGND VGND
+ VPWR VPWR net681 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_data_inbuf_30__0_ net252 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_30__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[109\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1350_ Tile_X0Y1_DSP_bot_Inst_MULADD__1348_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1349_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/B
+ sky130_fd_sc_hd__a21oi_4
XTile_X0Y1_DSP_bot_data_inbuf_21__0_ net242 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_21__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1281_ Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot_data_outbuf_10__0_ Tile_X0Y1_DSP_bot_data_inbuf_10__0_/X VGND VGND
+ VPWR VPWR net632 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput501 net501 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[7] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_data_inbuf_3__0_ net74 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_3__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0996_ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0996_/Y
+ sky130_fd_sc_hd__a21oi_1
Xoutput534 net534 VGND VGND VPWR VPWR Tile_X0Y0_UserCLKo sky130_fd_sc_hd__clkbuf_4
Xoutput523 net523 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput512 net512 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput545 net545 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput556 net556 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput578 net578 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput567 net567 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput589 net589 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1617_ Tile_X0Y1_DSP_bot_Inst_MULADD__1180_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1611_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1616_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/D sky130_fd_sc_hd__o311ai_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1548_ Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1554_/A
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit9 net260 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[233\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[2\] Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2END_EF_BEG\[1\] Tile_X0Y1_DSP_bot/ConfigBits\[25\] Tile_X0Y1_DSP_bot/ConfigBits\[26\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_data_inbuf_12__0_ net232 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_12__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[346\] Tile_X0Y1_DSP_bot/ConfigBits\[347\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JS2BEG\[6\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1479_ Tile_X0Y1_DSP_bot_Inst_MULADD__1093_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1095_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1479_/Y
+ sky130_fd_sc_hd__o21ai_2
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1
+ net204 Tile_X0Y0_S2BEGb\[1\] net339 net357 Tile_X0Y1_DSP_bot/ConfigBits\[288\] Tile_X0Y1_DSP_bot/ConfigBits\[289\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit10 net50 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[32\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit21 net62 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[43\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst0
+ net282 Tile_X0Y0_S1BEG\[1\] net335 Tile_X0Y1_DSP_bot/Q5 Tile_X0Y1_DSP_bot/ConfigBits\[107\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[108\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit0 net49 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[118\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[3\] net4 net84 Tile_X0Y1_bot2top\[3\] Tile_X0Y0_DSP_top/ConfigBits\[39\]
+ Tile_X0Y0_DSP_top/ConfigBits\[40\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_157_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_110 ANTENNA_110/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG3 Tile_X0Y1_NN4BEG\[2\]
+ net6 net86 net138 Tile_X0Y0_DSP_top/ConfigBits\[236\] Tile_X0Y0_DSP_top/ConfigBits\[237\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_EF_BEG\[3\] sky130_fd_sc_hd__mux4_1
XANTENNA_143 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 net184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_165 Tile_X0Y1_FrameStrobe_O\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_154 Tile_X0Y0_SS4BEG\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_176 ANTENNA_206/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 ANTENNA_187/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_198 Tile_X0Y0_SS4BEG\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__0850_ Tile_X0Y1_DSP_bot/A0 Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0849_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/B
+ sky130_fd_sc_hd__o21a_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[83\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1402_ Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/Y
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 Tile_X0Y0_E2END[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1333_ Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1334_/B
+ sky130_fd_sc_hd__or3_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG1 net41
+ net109 net144 Tile_X0Y0_DSP_top/JE2BEG\[1\] Tile_X0Y0_DSP_top/ConfigBits\[376\]
+ Tile_X0Y0_DSP_top/ConfigBits\[377\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_AB_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1264_ Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1263_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1147_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1264_/Y
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1195_ Tile_X0Y1_DSP_bot_Inst_MULADD__1089_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1091_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0895_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1195_/Y
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0979_ Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1299_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1299_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1124_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/B sky130_fd_sc_hd__a32o_1
Xoutput386 net386 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput397 net397 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_77_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_NN4END_inbuf_5__0_ net332 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/NN4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_N4BEG_outbuf_8__0_ ANTENNA_180/DIODE VGND VGND VPWR VPWR net516
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit1 net240 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[1\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG2 net324
+ net220 Tile_X0Y0_S4BEG\[1\] Tile_X0Y1_DSP_bot/JS2BEG\[2\] Tile_X0Y1_DSP_bot/ConfigBits\[396\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[397\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_CD_BEG\[2\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__0902_ Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1378_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0902_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG0 net292
+ net192 Tile_X0Y0_S2BEGb\[7\] net366 Tile_X0Y1_DSP_bot/ConfigBits\[248\] Tile_X0Y1_DSP_bot/ConfigBits\[249\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_GH_BEG\[0\] sky130_fd_sc_hd__mux4_2
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit20 net61 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[74\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit31 net73 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[85\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0
+ Tile_X0Y1_N2BEGb\[2\] Tile_X0Y1_N4BEG\[2\] net1 net7 Tile_X0Y0_DSP_top/ConfigBits\[250\]
+ Tile_X0Y0_DSP_top/ConfigBits\[251\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_154_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1316_ Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_154_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit19 net59 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[361\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1247_ Tile_X0Y1_DSP_bot_Inst_MULADD__1050_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1078_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1135_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1146_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1141_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1248_/C sky130_fd_sc_hd__o221a_1
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1178_ Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1113_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1172_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/C sky130_fd_sc_hd__o211ai_4
XANTENNA_32 Tile_X0Y1_FrameStrobe_O\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 Tile_X0Y0_SS4BEG\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 Tile_X0Y0_SS4BEG\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 Tile_X0Y1_FrameStrobe_O\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_65 ANTENNA_65/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_54 Tile_X0Y1_FrameStrobe_O\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 ANTENNA_76/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 ANTENNA_87/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 ANTENNA_98/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit3 net74 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[217\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_100_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_W6BEG_outbuf_8__0_ Tile_X0Y0_DSP_top/W6BEG_i\[8\] VGND VGND VPWR
+ VPWR net565 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst0
+ net284 net184 net337 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[81\] Tile_X0Y1_DSP_bot/ConfigBits\[82\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1
+ Tile_X0Y0_S2BEGb\[3\] Tile_X0Y0_S4BEG\[3\] net341 net357 Tile_X0Y1_DSP_bot/ConfigBits\[360\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[361\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit1 net240 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[353\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/Q5
+ Tile_X0Y1_DSP_bot/ConfigBits\[114\] Tile_X0Y1_DSP_bot/ConfigBits\[115\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1101_ Tile_X0Y1_DSP_bot_Inst_MULADD__1018_/Y Tile_X0Y1_DSP_bot/A6
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/C
+ sky130_fd_sc_hd__a21boi_4
XFILLER_0_158_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1032_ Tile_X0Y1_DSP_bot_Inst_MULADD__1124_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1032_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/C sky130_fd_sc_hd__nand4_4
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG0 net300
+ net200 Tile_X0Y0_S2BEG\[7\] net353 Tile_X0Y1_DSP_bot/ConfigBits\[192\] Tile_X0Y1_DSP_bot/ConfigBits\[193\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_ABb_BEG\[0\] sky130_fd_sc_hd__mux4_1
Xinput30 Tile_X0Y0_E6END[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput63 Tile_X0Y0_FrameData[22] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_6
Xinput52 Tile_X0Y0_FrameData[12] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput41 Tile_X0Y0_EE4END[2] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput96 Tile_X0Y0_S2MID[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_4
Xinput85 Tile_X0Y0_S2END[0] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
Xinput74 Tile_X0Y0_FrameData[3] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_6
XFILLER_0_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_NN4END_inbuf_1__0_ Tile_X0Y1_NN4BEG\[5\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/NN4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_149_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__22_ Tile_X0Y0_DSP_top/JN2BEG\[6\] VGND
+ VGND VPWR VPWR net492 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_E6END_inbuf_6__0_ net31 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/E6BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_100_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[272\] Tile_X0Y0_DSP_top/ConfigBits\[273\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JN2BEG\[6\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_strobe_inbuf_14__0_ Tile_X0Y1_FrameStrobe_O\[14\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_14__0_/X sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0
+ net282 net290 net182 net190 Tile_X0Y1_DSP_bot/ConfigBits\[272\] Tile_X0Y1_DSP_bot/ConfigBits\[273\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_123_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1650_ Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1657_/B sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit18 net58 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[392\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit29 net70 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[403\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_data_outbuf_28__0_ Tile_X0Y0_DSP_top_data_inbuf_28__0_/X VGND VGND
+ VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1581_ Tile_X0Y1_DSP_bot_Inst_MULADD__1581_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1581_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1696_/B sky130_fd_sc_hd__xor2_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__84_ net352 VGND VGND VPWR VPWR net733
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1015_ Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1013_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1014_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/C
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_151_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_outbuf_19__0_ Tile_X0Y0_DSP_top_data_inbuf_19__0_/X VGND VGND
+ VPWR VPWR net440 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit7 net258 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[135\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit6 net77 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[316\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_S4BEG_outbuf_8__0_ Tile_X0Y0_DSP_top/S4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_S4BEG\[8\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit3 net74 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[57\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_79_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[158\] Tile_X0Y1_DSP_bot/ConfigBits\[159\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/clr sky130_fd_sc_hd__mux4_2
XFILLER_0_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__05_ Tile_X0Y0_DSP_top/JE2BEG\[5\] VGND
+ VGND VPWR VPWR net391 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit23 net64 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[13\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit12 net52 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[2\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[77\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
Xinput220 Tile_X0Y1_EE4END[1] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_E6END_inbuf_6__0_ net211 VGND VGND VPWR VPWR ANTENNA_98/DIODE sky130_fd_sc_hd__clkbuf_2
Xinput231 Tile_X0Y1_FrameData[11] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_8
Xinput242 Tile_X0Y1_FrameData[21] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__buf_6
Xinput253 Tile_X0Y1_FrameData[31] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__buf_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1
+ Tile_X0Y0_S4BEG\[2\] Tile_X0Y0_SS4BEG\[2\] net340 net354 Tile_X0Y1_DSP_bot/ConfigBits\[324\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[325\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
Xinput286 Tile_X0Y1_N2END[1] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_2
Xinput297 Tile_X0Y1_N2MID[4] VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__buf_2
Xinput264 Tile_X0Y1_FrameStrobe[12] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_16
Xinput275 Tile_X0Y1_FrameStrobe[4] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput727 net727 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput716 net716 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput705 net705 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput749 net749 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput738 net738 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[1] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1702_ Tile_X0Y1_DSP_bot_Inst_MULADD__1644_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1645_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1723_/D
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1633_ Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1631_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1606_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/A sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1564_ Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_146_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1495_ Tile_X0Y1_DSP_bot_Inst_MULADD__1490_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1491_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1494_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1496_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_159_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__67_ Tile_X0Y0_S2BEG\[5\] VGND VGND
+ VPWR VPWR net680 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_data_inbuf_9__0_ net260 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_9__0_/X
+ sky130_fd_sc_hd__buf_1
XFILLER_0_118_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_inbuf_0__0_ net261 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_0__0_/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_outbuf_5__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_5__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[5\] sky130_fd_sc_hd__buf_8
XFILLER_0_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1280_ Tile_X0Y1_DSP_bot_Inst_MULADD__1371_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1371_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_25_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput502 net502 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[0] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0995_ Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0995_/Y
+ sky130_fd_sc_hd__nand3_1
Xoutput524 net524 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput513 net513 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput535 net535 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput557 net557 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput568 net568 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput546 net546 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput579 net579 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1616_ Tile_X0Y1_DSP_bot_Inst_MULADD__1616_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1616_/Y sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1547_ Tile_X0Y1_DSP_bot_Inst_MULADD__1547_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1547_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/A sky130_fd_sc_hd__nand2_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1478_ Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1478_/X sky130_fd_sc_hd__o211a_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit11 net51 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[33\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2
+ net764 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[288\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[289\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit22 net63 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[44\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[2\] Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2END_AB_BEG\[2\] Tile_X0Y1_DSP_bot/ConfigBits\[107\] Tile_X0Y1_DSP_bot/ConfigBits\[108\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit1 net60 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[119\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_WW4BEG_outbuf_3__0_ Tile_X0Y1_DSP_bot/WW4BEG_i\[3\] VGND VGND VPWR
+ VPWR net756 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[7\] Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[2\] Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2END_EF_BEG\[0\] Tile_X0Y0_DSP_top/ConfigBits\[39\] Tile_X0Y0_DSP_top/ConfigBits\[40\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_100 ANTENNA_100/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_122 net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 ANTENNA_111/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_166 Tile_X0Y1_FrameStrobe_O\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_155 Tile_X0Y0_SS4BEG\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_144 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_199 Tile_X0Y0_SS4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_188 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_177 ANTENNA_177/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[1\] net2 net134 Tile_X0Y1_bot2top\[5\] Tile_X0Y0_DSP_top/ConfigBits\[25\]
+ Tile_X0Y0_DSP_top/ConfigBits\[26\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[83\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1401_ Tile_X0Y1_DSP_bot_Inst_MULADD__1314_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1389_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1391_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1392_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/C sky130_fd_sc_hd__o211a_2
Xinput6 Tile_X0Y0_E2END[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1332_ Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1334_/A
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0
+ net3 net135 Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y0_DSP_top/ConfigBits\[52\]
+ Tile_X0Y0_DSP_top/ConfigBits\[53\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG2 Tile_X0Y1_N4BEG\[1\]
+ net24 net156 ANTENNA_63/DIODE Tile_X0Y0_DSP_top/ConfigBits\[378\] Tile_X0Y0_DSP_top/ConfigBits\[379\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_AB_BEG\[2\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1263_ Tile_X0Y1_DSP_bot_Inst_MULADD__1263_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1263_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1263_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1194_ Tile_X0Y1_DSP_bot_Inst_MULADD__1190_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1191_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1193_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/A
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_19_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0978_ Tile_X0Y1_DSP_bot_Inst_MULADD__1738_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1299_/D sky130_fd_sc_hd__or2b_2
Xoutput387 net387 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput398 net398 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_96_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit2 net251 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[2\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG3 net301
+ Tile_X0Y0_SS4BEG\[0\] net354 Tile_X0Y1_DSP_bot/JW2BEG\[2\] Tile_X0Y1_DSP_bot/ConfigBits\[398\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[399\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_CD_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_N1BEG0 Tile_X0Y1_bot2top\[2\]
+ Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[3\] Tile_X0Y0_DSP_top/JW2BEG\[3\] Tile_X0Y0_DSP_top/J_l_CD_BEG\[1\]
+ Tile_X0Y0_DSP_top/ConfigBits\[0\] Tile_X0Y0_DSP_top/ConfigBits\[1\] VGND VGND VPWR
+ VPWR net482 sky130_fd_sc_hd__mux4_2
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_WW4END_inbuf_6__0_ net367 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/WW4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_153_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0901_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0887_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0890_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0896_/X Tile_X0Y1_DSP_bot_Inst_MULADD__0900_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0906_/A sky130_fd_sc_hd__o311a_1
XFILLER_0_106_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top/JN2BEG\[5\] Tile_X0Y0_DSP_top/JN2BEG\[7\] Tile_X0Y0_DSP_top/JE2BEG\[5\]
+ Tile_X0Y0_DSP_top/JE2BEG\[7\] Tile_X0Y0_DSP_top/ConfigBits\[147\] Tile_X0Y0_DSP_top/ConfigBits\[148\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG1 net288
+ net188 Tile_X0Y0_SS4BEG\[0\] net341 Tile_X0Y1_DSP_bot/ConfigBits\[250\] Tile_X0Y1_DSP_bot/ConfigBits\[251\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_GH_BEG\[1\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_NN4BEG_outbuf_0__0_ Tile_X0Y0_DSP_top/NN4BEG_i\[0\] VGND VGND VPWR
+ VPWR net518 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit10 net50 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[64\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit21 net62 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[75\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1
+ net21 net87 net139 net153 Tile_X0Y0_DSP_top/ConfigBits\[250\] Tile_X0Y0_DSP_top/ConfigBits\[251\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_154_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1315_ Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1292_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1315_/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1246_ Tile_X0Y1_DSP_bot_Inst_MULADD__1133_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1157_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1248_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1248_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1246_/Y sky130_fd_sc_hd__a22oi_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1177_ Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/A sky130_fd_sc_hd__buf_4
XFILLER_0_144_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_22 Tile_X0Y0_SS4BEG\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 Tile_X0Y0_SS4BEG\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 Tile_X0Y1_FrameStrobe_O\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 ANTENNA_68/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 Tile_X0Y1_FrameStrobe_O\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_55 Tile_X0Y1_FrameStrobe_O\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 ANTENNA_77/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_99 ANTENNA_99/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 ANTENNA_89/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_SS4BEG_outbuf_3__0_ Tile_X0Y0_DSP_top/SS4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_SS4BEG\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit4 net75 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[218\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_100_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[2\] Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2END_EF_BEG\[3\] Tile_X0Y1_DSP_bot/ConfigBits\[81\] Tile_X0Y1_DSP_bot/ConfigBits\[82\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 net764 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[360\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[361\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit2 net251 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[354\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2
+ wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[114\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[115\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1100_ Tile_X0Y1_DSP_bot_Inst_MULADD__1092_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1096_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1099_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1100_/Y
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_158_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1031_ Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1029_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1030_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/B
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_33_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG1 net296
+ net196 Tile_X0Y0_S2BEG\[3\] net349 Tile_X0Y1_DSP_bot/ConfigBits\[194\] Tile_X0Y1_DSP_bot/ConfigBits\[195\]
+ VGND VGND VPWR VPWR ANTENNA_101/DIODE sky130_fd_sc_hd__mux4_2
Xinput31 Tile_X0Y0_E6END[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput20 Tile_X0Y0_E2MID[7] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[2\] Tile_X0Y1_N2BEGb\[4\] Tile_X0Y1_N4BEG\[0\] net9 Tile_X0Y0_DSP_top/ConfigBits\[290\]
+ Tile_X0Y0_DSP_top/ConfigBits\[291\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_83_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput64 Tile_X0Y0_FrameData[23] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_6
Xinput53 Tile_X0Y0_FrameData[13] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_8
Xinput42 Tile_X0Y0_EE4END[3] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput97 Tile_X0Y0_S2MID[4] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_4
Xinput86 Tile_X0Y0_S2END[1] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_4
Xinput75 Tile_X0Y0_FrameData[4] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1229_ Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1137_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1149_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1243_/A
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_117_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__21_ Tile_X0Y0_DSP_top/JN2BEG\[5\] VGND
+ VGND VPWR VPWR net491 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[1\] Tile_X0Y0_S2BEGb\[5\] net335 net337 Tile_X0Y1_DSP_bot/ConfigBits\[272\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[273\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_WW4END_inbuf_2__0_ net177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/WW4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit19 net59 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[393\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1580_ Tile_X0Y1_DSP_bot_Inst_MULADD__1557_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1556_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1556_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1581_/B
+ sky130_fd_sc_hd__a21bo_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_strobe_inbuf_9__0_ Tile_X0Y1_FrameStrobe_O\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_9__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__83_ net351 VGND VGND VPWR VPWR net732
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1014_ Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1731_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1014_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit8 net259 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[136\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit7 net78 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[317\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit4 net75 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[58\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_94_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__04_ Tile_X0Y0_DSP_top/JE2BEG\[4\] VGND
+ VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit13 net53 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[3\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit24 net65 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[14\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0
+ net284 net292 net184 net192 Tile_X0Y1_DSP_bot/ConfigBits\[312\] Tile_X0Y1_DSP_bot/ConfigBits\[313\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
Xinput210 Tile_X0Y1_E6END[7] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
Xinput221 Tile_X0Y1_EE4END[2] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_2
Xinput254 Tile_X0Y1_FrameData[3] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__buf_6
Xinput232 Tile_X0Y1_FrameData[12] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_8
Xinput243 Tile_X0Y1_FrameData[22] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_8
Xinput265 Tile_X0Y1_FrameStrobe[13] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_1
Xinput287 Tile_X0Y1_N2END[2] VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__buf_2
Xinput276 Tile_X0Y1_FrameStrobe[5] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__buf_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4
+ Tile_X0Y1_DSP_bot/ConfigBits\[324\] Tile_X0Y1_DSP_bot/ConfigBits\[325\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
Xinput298 Tile_X0Y1_N2MID[5] VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__buf_2
XFILLER_0_105_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_NN4BEG_outbuf_6__0_ Tile_X0Y1_DSP_bot/NN4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y1_NN4BEG\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_SS4END_inbuf_8__0_ Tile_X0Y0_SS4BEG\[12\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/SS4BEG_i\[8\]
+ sky130_fd_sc_hd__buf_2
Xoutput717 net717 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput706 net706 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[1] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1701_ Tile_X0Y1_DSP_bot_Inst_MULADD__1701_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1722_/D sky130_fd_sc_hd__clkbuf_1
Xoutput728 net728 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput739 net739 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1632_ Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/Y sky130_fd_sc_hd__nand4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1563_ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1562_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/B
+ sky130_fd_sc_hd__a21bo_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1494_ Tile_X0Y1_DSP_bot_Inst_MULADD__1299_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1299_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1494_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_SS4BEG_outbuf_9__0_ Tile_X0Y1_DSP_bot/SS4BEG_i\[9\] VGND VGND VPWR
+ VPWR net714 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__66_ Tile_X0Y0_S2BEG\[4\] VGND VGND
+ VPWR VPWR net679 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_S4END_inbuf_0__0_ net111 VGND VGND VPWR VPWR ANTENNA_86/DIODE sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[152\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/C8 sky130_fd_sc_hd__o21ai_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[2\] Tile_X0Y1_N2BEGb\[6\] net3 net11 Tile_X0Y0_DSP_top/ConfigBits\[362\]
+ Tile_X0Y0_DSP_top/ConfigBits\[363\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_W6END_inbuf_4__0_ net161 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/W6BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_73_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_EE4END_inbuf_7__0_ net215 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/EE4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0994_ Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/C
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1002_/A sky130_fd_sc_hd__a32o_1
Xoutput514 net514 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput503 net503 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput525 net525 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput536 net536 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput558 net558 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput569 net569 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput547 net547 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1615_ Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1616_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/C sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1546_ Tile_X0Y1_DSP_bot_Inst_MULADD__1588_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1547_/B sky130_fd_sc_hd__inv_2
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1477_ Tile_X0Y1_DSP_bot_Inst_MULADD__1036_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1477_/X sky130_fd_sc_hd__o211a_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[288\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[289\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit12 net52 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[34\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit23 net64 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[45\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_49_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_EE4BEG_outbuf_3__0_ ANTENNA_60/DIODE VGND VGND VPWR VPWR net423
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__49_ net296 VGND VGND VPWR VPWR Tile_X0Y1_N2BEGb\[3\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit2 net71 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[120\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_S4END_inbuf_0__0_ Tile_X0Y0_S4BEG\[4\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/S4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_123 net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 ANTENNA_112/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_101 ANTENNA_101/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_134 net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 Tile_X0Y0_SS4BEG\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_167 Tile_X0Y1_FrameStrobe_O\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_145 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_189 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_178 ANTENNA_64/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[9\] Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[2\] Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2END_AB_BEG\[1\] Tile_X0Y0_DSP_top/ConfigBits\[25\] Tile_X0Y0_DSP_top/ConfigBits\[26\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top_SS4END_inbuf_4__0_ net131 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/SS4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1400_ Tile_X0Y1_DSP_bot_Inst_MULADD__1391_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1392_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1399_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/B
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput7 Tile_X0Y0_E2END[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1331_ Tile_X0Y1_DSP_bot_Inst_MULADD__1614_/S Tile_X0Y1_DSP_bot_Inst_MULADD__1329_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1330_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/A
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[5\]
+ Tile_X0Y0_DSP_top/ConfigBits\[52\] Tile_X0Y0_DSP_top/ConfigBits\[53\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG3 Tile_X0Y1_N4BEG\[0\]
+ net21 net101 Tile_X0Y0_DSP_top/JW2BEG\[1\] Tile_X0Y0_DSP_top/ConfigBits\[380\] Tile_X0Y0_DSP_top/ConfigBits\[381\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_AB_BEG\[3\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit0 net229 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[256\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_strobe_outbuf_15__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_15__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[15\] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1262_ Tile_X0Y1_DSP_bot_Inst_MULADD__1238_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1260_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1261_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1263_/A
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1193_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1019_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1096_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1099_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1192_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1193_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_W6END_inbuf_4__0_ net362 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/W6BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0977_ Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/A Tile_X0Y1_DSP_bot/B4
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1299_/C sky130_fd_sc_hd__or2_1
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput399 net399 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput388 net388 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[2] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1529_ Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1424_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1424_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1528_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/C sky130_fd_sc_hd__a31oi_4
XFILLER_0_139_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[1\] Tile_X0Y1_N2BEGb\[5\] net2 net10 Tile_X0Y0_DSP_top/ConfigBits\[326\]
+ Tile_X0Y0_DSP_top/ConfigBits\[327\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit3 net254 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[3\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_N1BEG1 Tile_X0Y1_bot2top\[3\]
+ ANTENNA_177/DIODE Tile_X0Y0_DSP_top/JW2BEG\[0\] Tile_X0Y0_DSP_top/J_l_EF_BEG\[2\]
+ Tile_X0Y0_DSP_top/ConfigBits\[2\] Tile_X0Y0_DSP_top/ConfigBits\[3\] VGND VGND VPWR
+ VPWR net483 sky130_fd_sc_hd__mux4_2
XFILLER_0_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0900_ Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1378_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0900_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_EE4END_inbuf_3__0_ net46 VGND VGND VPWR VPWR ANTENNA_60/DIODE sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_cus_mux41_buf_inst1
+ ANTENNA_64/DIODE ANTENNA_179/DIODE Tile_X0Y0_DSP_top/JW2BEG\[5\] Tile_X0Y0_DSP_top/JW2BEG\[7\]
+ Tile_X0Y0_DSP_top/ConfigBits\[147\] Tile_X0Y0_DSP_top/ConfigBits\[148\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot17_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG2 net324
+ net190 Tile_X0Y0_S2BEGb\[5\] net343 Tile_X0Y1_DSP_bot/ConfigBits\[252\] Tile_X0Y1_DSP_bot/ConfigBits\[253\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_GH_BEG\[2\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit11 net51 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[65\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit22 net63 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[76\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_N4BEG_outbuf_10__0_ Tile_X0Y1_DSP_bot/N4BEG_i\[10\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N4BEG\[10\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[250\] Tile_X0Y0_DSP_top/ConfigBits\[251\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1314_ Tile_X0Y1_DSP_bot_Inst_MULADD__1273_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1284_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1288_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1290_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1314_/X sky130_fd_sc_hd__o211a_2
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1245_ Tile_X0Y1_DSP_bot_Inst_MULADD__1135_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1242_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1263_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1244_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1248_/B sky130_fd_sc_hd__o211ai_4
XFILLER_0_59_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1176_ Tile_X0Y1_DSP_bot_Inst_MULADD__1034_/X Tile_X0Y1_DSP_bot/B7
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1175_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/C
+ sky130_fd_sc_hd__o21a_4
XANTENNA_23 Tile_X0Y0_SS4BEG\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 Tile_X0Y0_SS4BEG\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 Tile_X0Y1_FrameStrobe_O\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 Tile_X0Y1_N1BEG\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 Tile_X0Y1_FrameStrobe_O\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 ANTENNA_78/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_67 ANTENNA_68/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 ANTENNA_89/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_NN4BEG_outbuf_10__0_ Tile_X0Y0_DSP_top/NN4BEG_i\[10\] VGND VGND
+ VPWR VPWR net519 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_N4BEG_outbuf_2__0_ Tile_X0Y1_DSP_bot/N4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N4BEG\[2\] sky130_fd_sc_hd__buf_2
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit5 net76 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[219\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_97_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[360\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[361\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit3 net254 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[355\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[2\] Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[2\] Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[2\] Tile_X0Y1_DSP_bot/ConfigBits\[114\] Tile_X0Y1_DSP_bot/ConfigBits\[115\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1030_ Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1738_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1030_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_75_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG2 net298
+ net198 Tile_X0Y0_S2BEG\[5\] net351 Tile_X0Y1_DSP_bot/ConfigBits\[196\] Tile_X0Y1_DSP_bot/ConfigBits\[197\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_ABb_BEG\[2\] sky130_fd_sc_hd__mux4_2
Xinput21 Tile_X0Y0_E6END[0] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
Xinput10 Tile_X0Y0_E2END[5] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1
+ net21 net89 net141 net153 Tile_X0Y0_DSP_top/ConfigBits\[290\] Tile_X0Y0_DSP_top/ConfigBits\[291\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
Xinput54 Tile_X0Y0_FrameData[14] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_6
Xinput32 Tile_X0Y0_E6END[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 Tile_X0Y0_EE4END[4] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0
+ net281 net285 net181 net185 Tile_X0Y1_DSP_bot/ConfigBits\[348\] Tile_X0Y1_DSP_bot/ConfigBits\[349\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
Xinput87 Tile_X0Y0_S2END[2] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
Xinput98 Tile_X0Y0_S2MID[5] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_4
Xinput65 Tile_X0Y0_FrameData[24] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_8
Xinput76 Tile_X0Y0_FrameData[5] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_6
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_E6BEG_outbuf_7__0_ Tile_X0Y0_DSP_top/E6BEG_i\[7\] VGND VGND VPWR
+ VPWR net411 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_strobe_outbuf_10__0_ Tile_X0Y0_DSP_top_strobe_inbuf_10__0_/X VGND
+ VGND VPWR VPWR net463 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[1\] net2 net134 Tile_X0Y1_bot2top\[5\] Tile_X0Y0_DSP_top/ConfigBits\[81\]
+ Tile_X0Y0_DSP_top/ConfigBits\[82\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_EE4BEG_outbuf_9__0_ Tile_X0Y1_DSP_bot/EE4BEG_i\[9\] VGND VGND VPWR
+ VPWR net630 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1228_ Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1228_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1243_/C
+ sky130_fd_sc_hd__nand3_2
XFILLER_0_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1159_ Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1165_/B sky130_fd_sc_hd__nand4_4
XFILLER_0_114_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_W6BEG_outbuf_2__0_ Tile_X0Y1_DSP_bot/W6BEG_i\[2\] VGND VGND VPWR
+ VPWR net739 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__20_ Tile_X0Y0_DSP_top/JN2BEG\[4\] VGND
+ VGND VPWR VPWR net490 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_data_outbuf_0__0_ Tile_X0Y0_DSP_top_data_inbuf_0__0_/X VGND VGND
+ VPWR VPWR net430 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[272\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[273\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_data_inbuf_24__0_ net65 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_24__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG0 net291
+ net191 Tile_X0Y0_SS4BEG\[3\] net344 Tile_X0Y1_DSP_bot/ConfigBits\[224\] Tile_X0Y1_DSP_bot/ConfigBits\[225\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_AB_BEG\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_48_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__82_ net350 VGND VGND VPWR VPWR net731
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1013_ Tile_X0Y1_DSP_bot/A5 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1013_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_data_inbuf_15__0_ net55 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_15__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit9 net260 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[137\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit8 net79 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[318\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit5 net76 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[59\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_data_outbuf_31__0_ Tile_X0Y1_DSP_bot_data_inbuf_31__0_/X VGND VGND
+ VPWR VPWR net655 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__03_ Tile_X0Y0_DSP_top/JE2BEG\[3\] VGND
+ VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit14 net54 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[4\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_data_outbuf_0__0_ Tile_X0Y1_DSP_bot_data_inbuf_0__0_/X VGND VGND
+ VPWR VPWR net631 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[1\] Tile_X0Y0_S1BEG\[3\] Tile_X0Y0_S2BEGb\[7\] net337 Tile_X0Y1_DSP_bot/ConfigBits\[312\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[313\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit25 net66 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[15\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput200 Tile_X0Y1_E2MID[7] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_2
Xinput211 Tile_X0Y1_E6END[8] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
Xinput222 Tile_X0Y1_EE4END[3] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__buf_1
Xinput233 Tile_X0Y1_FrameData[13] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_8
Xinput244 Tile_X0Y1_FrameData[23] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_8
Xinput277 Tile_X0Y1_FrameStrobe[6] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__buf_8
Xinput288 Tile_X0Y1_N2END[3] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_4
Xinput266 Tile_X0Y1_FrameStrobe[14] VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_1
Xinput255 Tile_X0Y1_FrameData[4] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__buf_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[324\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[325\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
Xinput299 Tile_X0Y1_N2MID[6] VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__buf_4
XTile_X0Y1_DSP_bot_data_outbuf_22__0_ Tile_X0Y1_DSP_bot_data_inbuf_22__0_/X VGND VGND
+ VPWR VPWR net645 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput718 net718 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput707 net707 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1700_ Tile_X0Y1_DSP_bot_Inst_MULADD__1674_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1700_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1700_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1701_/A
+ sky130_fd_sc_hd__and3b_1
Xoutput729 net729 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1631_ Tile_X0Y1_DSP_bot_Inst_MULADD__1631_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1631_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1631_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1562_ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1562_/X sky130_fd_sc_hd__a22o_1
XTile_X0Y1_DSP_bot_data_inbuf_24__0_ net245 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_24__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1493_ Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/B sky130_fd_sc_hd__nand4_4
XTile_X0Y1_DSP_bot_data_outbuf_13__0_ Tile_X0Y1_DSP_bot_data_inbuf_13__0_/X VGND VGND
+ VPWR VPWR net635 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__65_ Tile_X0Y0_S2BEG\[3\] VGND VGND
+ VPWR VPWR net678 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_inbuf_6__0_ net77 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_6__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_S4BEG_outbuf_2__0_ ANTENNA_107/DIODE VGND VGND VPWR VPWR net691
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit30 net252 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[126\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_96_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_data_inbuf_15__0_ net235 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_15__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[152\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1
+ net81 net83 net91 net135 Tile_X0Y0_DSP_top/ConfigBits\[362\] Tile_X0Y0_DSP_top/ConfigBits\[363\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__0993_ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/C
+ sky130_fd_sc_hd__a21o_1
Xoutput526 net526 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput515 net515 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput504 net504 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput559 net559 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput548 net548 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput537 net537 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1614_ Tile_X0Y1_DSP_bot_Inst_MULADD__1613_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1721_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1614_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1616_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1545_ Tile_X0Y1_DSP_bot_Inst_MULADD__1545_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1545_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1545_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1588_/A
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1476_ Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1441_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1496_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[290\] Tile_X0Y1_DSP_bot/ConfigBits\[291\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JE2BEG\[0\] sky130_fd_sc_hd__mux4_2
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit24 net65 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[46\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit13 net53 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[35\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__48_ net295 VGND VGND VPWR VPWR Tile_X0Y1_N2BEGb\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_134_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[0\] Tile_X0Y1_N2BEGb\[0\] net1 net33 Tile_X0Y0_DSP_top/ConfigBits\[274\]
+ Tile_X0Y0_DSP_top/ConfigBits\[275\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit3 net74 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[121\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_NN4END_inbuf_8__0_ net320 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/NN4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_124 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_113 ANTENNA_113/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_102 ANTENNA_105/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 Tile_X0Y0_SS4BEG\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_146 net343 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_168 Tile_X0Y1_FrameStrobe_O\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_179 ANTENNA_179/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 Tile_X0Y0_E2END[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_0_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1330_ Tile_X0Y1_DSP_bot_Inst_MULADD__1714_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1614_/S
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1330_/X sky130_fd_sc_hd__or2b_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[52\] Tile_X0Y0_DSP_top/ConfigBits\[53\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit1 net240 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[257\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1261_ Tile_X0Y1_DSP_bot_Inst_MULADD__1114_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1120_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1137_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1261_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1192_ Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1192_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_0_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0976_ Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/Y sky130_fd_sc_hd__nand2_2
Xoutput389 net389 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_0_10_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1528_ Tile_X0Y1_DSP_bot_Inst_MULADD__1503_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1506_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1527_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1474_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1528_/Y sky130_fd_sc_hd__o22ai_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1459_ Tile_X0Y1_DSP_bot/C10 Tile_X0Y1_DSP_bot_Inst_MULADD__1752_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1459_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1460_/B
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1
+ net82 net90 net134 net136 Tile_X0Y0_DSP_top/ConfigBits\[326\] Tile_X0Y0_DSP_top/ConfigBits\[327\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit4 net255 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[4\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_N1BEG2 Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[1\] Tile_X0Y0_DSP_top/JW2BEG\[1\] Tile_X0Y0_DSP_top/J_l_GH_BEG\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[4\] Tile_X0Y0_DSP_top/ConfigBits\[5\] VGND VGND VPWR
+ VPWR net484 sky130_fd_sc_hd__mux4_2
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG3 net286
+ net222 Tile_X0Y0_S2BEGb\[1\] net339 Tile_X0Y1_DSP_bot/ConfigBits\[254\] Tile_X0Y1_DSP_bot/ConfigBits\[255\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_GH_BEG\[3\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit12 net52 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[66\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit23 net64 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[77\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_138_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_strobe_outbuf_2__0_ Tile_X0Y0_DSP_top_strobe_inbuf_2__0_/X VGND
+ VGND VPWR VPWR net474 sky130_fd_sc_hd__buf_1
XFILLER_0_47_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1313_ Tile_X0Y1_DSP_bot_Inst_MULADD__1313_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1313_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1313_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/A
+ sky130_fd_sc_hd__nand3_4
XFILLER_0_154_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[250\] Tile_X0Y0_DSP_top/ConfigBits\[251\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1244_ Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1043_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1244_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1175_ Tile_X0Y1_DSP_bot_Inst_MULADD__1741_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1175_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1175_/X sky130_fd_sc_hd__or2_2
XFILLER_0_74_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_13 Tile_X0Y0_SS4BEG\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_46 Tile_X0Y1_FrameStrobe_O\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_57 Tile_X0Y1_N1BEG\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 Tile_X0Y0_SS4BEG\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 Tile_X0Y1_FrameStrobe_O\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 ANTENNA_79/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 ANTENNA_68/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__0959_ Tile_X0Y1_DSP_bot_Inst_MULADD__0926_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0958_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0959_/X
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit6 net77 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[220\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_NN4END_inbuf_4__0_ Tile_X0Y1_NN4BEG\[8\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/NN4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_E6END_inbuf_9__0_ net23 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/E6BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[362\] Tile_X0Y1_DSP_bot/ConfigBits\[363\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JW2BEG\[2\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_WW4BEG_outbuf_0__0_ Tile_X0Y0_DSP_top/WW4BEG_i\[0\] VGND VGND VPWR
+ VPWR net567 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_strobe_inbuf_17__0_ Tile_X0Y1_FrameStrobe_O\[17\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_17__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit4 net255 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[356\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[116\] Tile_X0Y1_DSP_bot/ConfigBits\[117\] VGND VGND
+ VPWR VPWR net737 sky130_fd_sc_hd__mux4_1
XFILLER_0_158_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG3 net294
+ net194 Tile_X0Y0_S2BEG\[1\] net347 Tile_X0Y1_DSP_bot/ConfigBits\[198\] Tile_X0Y1_DSP_bot/ConfigBits\[199\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_ABb_BEG\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput22 Tile_X0Y0_E6END[10] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 Tile_X0Y0_E2END[6] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[290\] Tile_X0Y0_DSP_top/ConfigBits\[291\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
Xinput55 Tile_X0Y0_FrameData[15] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput33 Tile_X0Y0_EE4END[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
Xinput44 Tile_X0Y0_EE4END[5] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[0\] Tile_X0Y0_S2BEGb\[0\] net334 net336 Tile_X0Y1_DSP_bot/ConfigBits\[348\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[349\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
Xinput88 Tile_X0Y0_S2END[3] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
Xinput66 Tile_X0Y0_FrameData[25] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_8
Xinput77 Tile_X0Y0_FrameData[6] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput99 Tile_X0Y0_S2MID[6] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_2
XFILLER_0_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[9\] Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[2\] Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2END_AB_BEG\[3\] Tile_X0Y0_DSP_top/ConfigBits\[81\] Tile_X0Y0_DSP_top/ConfigBits\[82\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1227_ Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1183_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1228_/C
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1158_ Tile_X0Y1_DSP_bot_Inst_MULADD__1133_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1157_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1144_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/C
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_74_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1089_ Tile_X0Y1_DSP_bot_Inst_MULADD__1089_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1089_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_inbuf_10__0_ net262 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_10__0_/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_132_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[272\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[273\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_N4END_inbuf_0__0_ Tile_X0Y1_N4BEG\[4\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/N4BEG_i\[0\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_E6END_inbuf_9__0_ net203 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/E6BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG1 net317
+ net187 Tile_X0Y0_S2BEGb\[2\] net340 Tile_X0Y1_DSP_bot/ConfigBits\[226\] Tile_X0Y1_DSP_bot/ConfigBits\[227\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_AB_BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_158_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__81_ net349 VGND VGND VPWR VPWR net730
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1012_ Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1012_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/A sky130_fd_sc_hd__and4_2
XFILLER_0_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit9 net80 Tile_X0Y1_FrameStrobe_O\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[319\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame2_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit6 net77 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[60\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_149_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__02_ Tile_X0Y0_DSP_top/JE2BEG\[2\] VGND
+ VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit15 net55 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[5\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[312\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[313\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit26 net67 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[16\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput201 Tile_X0Y1_E6END[0] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__buf_4
Xinput223 Tile_X0Y1_EE4END[4] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_1
Xinput212 Tile_X0Y1_E6END[9] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
Xinput234 Tile_X0Y1_FrameData[14] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_8
Xinput245 Tile_X0Y1_FrameData[24] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_8
Xinput278 Tile_X0Y1_FrameStrobe[7] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__buf_8
Xinput267 Tile_X0Y1_FrameStrobe[15] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_1
Xinput256 Tile_X0Y1_FrameData[5] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__buf_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[326\] Tile_X0Y1_DSP_bot/ConfigBits\[327\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JS2BEG\[1\] sky130_fd_sc_hd__mux4_2
Xinput289 Tile_X0Y1_N2END[4] VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_inbuf_3__0_ net274 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_3__0_/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput708 net708 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput719 net719 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[0] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_strobe_outbuf_8__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_8__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[8\] sky130_fd_sc_hd__clkbuf_16
XTile_X0Y1_DSP_bot_N4END_inbuf_0__0_ net311 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/N4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1630_ Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1616_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1631_/B sky130_fd_sc_hd__a32oi_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1561_ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/X
+ sky130_fd_sc_hd__and3_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1492_ Tile_X0Y1_DSP_bot_Inst_MULADD__1477_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1478_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1490_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1491_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1496_/B sky130_fd_sc_hd__o211ai_1
XFILLER_0_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__64_ Tile_X0Y0_S2BEG\[2\] VGND VGND
+ VPWR VPWR net677 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit20 net241 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[116\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_142_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit31 net253 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[127\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_142_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_E1BEG0 Tile_X0Y1_DSP_bot/Q3
+ Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[3\] Tile_X0Y1_DSP_bot/JN2BEG\[3\] Tile_X0Y1_DSP_bot/J_l_CD_BEG\[1\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[34\] Tile_X0Y1_DSP_bot/ConfigBits\[35\] VGND VGND
+ VPWR VPWR net583 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1759_ net333 Tile_X0Y1_DSP_bot/C17 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1759_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[362\] Tile_X0Y0_DSP_top/ConfigBits\[363\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_WW4BEG_outbuf_6__0_ Tile_X0Y1_DSP_bot/WW4BEG_i\[6\] VGND VGND VPWR
+ VPWR net759 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0992_ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/D
+ sky130_fd_sc_hd__nand3_2
Xoutput505 net505 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput516 net516 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput527 net527 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput549 net549 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[2] sky130_fd_sc_hd__clkbuf_4
Xoutput538 net538 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1613_ Tile_X0Y1_DSP_bot/C15 Tile_X0Y1_DSP_bot_Inst_MULADD__1757_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1613_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1544_ Tile_X0Y1_DSP_bot_Inst_MULADD__1545_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1545_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1545_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1547_/A
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1475_ Tile_X0Y1_DSP_bot_Inst_MULADD__1458_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1458_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1474_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1510_/A
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit14 net54 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[36\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit25 net66 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[47\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_119_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__47_ net294 VGND VGND VPWR VPWR Tile_X0Y1_N2BEGb\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1
+ net81 net85 net133 net135 Tile_X0Y0_DSP_top/ConfigBits\[274\] Tile_X0Y0_DSP_top/ConfigBits\[275\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit4 net75 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[122\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_125 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 ANTENNA_105/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_136 net295 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_158 Tile_X0Y0_SS4BEG\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_147 net343 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_169 Tile_X0Y1_FrameStrobe_O\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[2\] Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[2\] Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[2\] Tile_X0Y0_DSP_top/ConfigBits\[52\] Tile_X0Y0_DSP_top/ConfigBits\[53\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
Xinput9 Tile_X0Y0_E2END[4] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit2 net251 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[258\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit30 net252 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[158\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1260_ Tile_X0Y1_DSP_bot_Inst_MULADD__1234_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1222_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1223_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1228_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1260_/X sky130_fd_sc_hd__o311a_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG0 Tile_X0Y1_N2BEG\[7\]
+ net20 net100 net152 Tile_X0Y0_DSP_top/ConfigBits\[206\] Tile_X0Y0_DSP_top/ConfigBits\[207\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[0\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_N4BEG0 Tile_X0Y1_N2BEGb\[2\]
+ Tile_X0Y1_N4BEG\[1\] net24 Tile_X0Y1_bot2top\[4\] Tile_X0Y0_DSP_top/ConfigBits\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[9\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__mux4_2
XFILLER_0_52_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1191_ Tile_X0Y1_DSP_bot_Inst_MULADD__0968_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0969_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1189_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1191_/X sky130_fd_sc_hd__o2111a_2
XTile_X0Y1_DSP_bot_WW4END_inbuf_9__0_ net370 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/WW4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_NN4BEG_outbuf_3__0_ Tile_X0Y0_DSP_top/NN4BEG_i\[3\] VGND VGND VPWR
+ VPWR net527 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0975_ Tile_X0Y1_DSP_bot_Inst_MULADD__0888_/X Tile_X0Y1_DSP_bot_Inst_MULADD__0889_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0895_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0934_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/B sky130_fd_sc_hd__o211ai_4
XFILLER_0_10_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1527_ Tile_X0Y1_DSP_bot_Inst_MULADD__1507_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1506_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1506_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1527_/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1458_ Tile_X0Y1_DSP_bot_Inst_MULADD__1458_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1458_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1471_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1389_ Tile_X0Y1_DSP_bot_Inst_MULADD__1317_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1296_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1306_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1389_/Y
+ sky130_fd_sc_hd__a21oi_2
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[326\] Tile_X0Y0_DSP_top/ConfigBits\[327\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_SS4BEG_outbuf_6__0_ Tile_X0Y0_DSP_top/SS4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_SS4BEG\[6\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit5 net256 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[5\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_130_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_S4BEG_outbuf_10__0_ Tile_X0Y0_DSP_top/S4BEG_i\[10\] VGND VGND VPWR
+ VPWR Tile_X0Y0_S4BEG\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_N1BEG3 Tile_X0Y1_bot2top\[5\]
+ Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[2\] Tile_X0Y0_DSP_top/JW2BEG\[2\] ANTENNA_65/DIODE
+ Tile_X0Y0_DSP_top/ConfigBits\[6\] Tile_X0Y0_DSP_top/ConfigBits\[7\] VGND VGND VPWR
+ VPWR net485 sky130_fd_sc_hd__mux4_2
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit13 net53 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[67\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit24 net65 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[78\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1312_ Tile_X0Y1_DSP_bot_Inst_MULADD__1398_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1398_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1294_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1311_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1297_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1313_/C sky130_fd_sc_hd__o221ai_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[252\] Tile_X0Y0_DSP_top/ConfigBits\[253\] VGND VGND
+ VPWR VPWR ANTENNA_61/DIODE sky130_fd_sc_hd__mux4_2
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1243_ Tile_X0Y1_DSP_bot_Inst_MULADD__1243_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1243_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1243_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1263_/B
+ sky130_fd_sc_hd__nand3_4
XFILLER_0_59_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1174_ Tile_X0Y1_DSP_bot_Inst_MULADD__1113_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1172_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1173_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/A
+ sky130_fd_sc_hd__a21oi_4
XANTENNA_14 Tile_X0Y0_SS4BEG\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 Tile_X0Y1_FrameStrobe_O\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 Tile_X0Y1_FrameStrobe_O\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 Tile_X0Y1_FrameStrobe_O\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 ANTENNA_73/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0958_ Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/A Tile_X0Y1_DSP_bot/B3
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0958_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0889_ Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0889_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0889_/Y sky130_fd_sc_hd__nor2_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit7 net78 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[221\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst0
+ net283 net183 Tile_X0Y0_S1BEG\[2\] Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/ConfigBits\[42\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[43\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_EE4BEG_outbuf_11__0_ ANTENNA_99/DIODE VGND VGND VPWR VPWR net617
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit5 net256 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[357\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_WW4END_inbuf_5__0_ net180 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/WW4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 Tile_X0Y0_E2END[7] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[290\] Tile_X0Y0_DSP_top/ConfigBits\[291\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_141_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput23 Tile_X0Y0_E6END[11] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 Tile_X0Y0_EE4END[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput45 Tile_X0Y0_EE4END[6] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 net764 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[348\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[349\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
Xinput89 Tile_X0Y0_S2END[4] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xinput67 Tile_X0Y0_FrameData[26] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_4
Xinput56 Tile_X0Y0_FrameData[16] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_8
Xinput78 Tile_X0Y0_FrameData[7] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1226_ Tile_X0Y1_DSP_bot/A0 Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0849_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/C
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_0_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1157_ Tile_X0Y1_DSP_bot_Inst_MULADD__1050_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1078_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1156_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1157_/Y sky130_fd_sc_hd__a2bb2oi_4
XFILLER_0_74_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1088_ Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1731_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1089_/A sky130_fd_sc_hd__and2_1
XFILLER_0_117_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[274\] Tile_X0Y1_DSP_bot/ConfigBits\[275\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JN2BEG\[4\] sky130_fd_sc_hd__mux4_2
XFILLER_0_53_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG2 net289
+ net213 Tile_X0Y0_S2BEGb\[4\] net342 Tile_X0Y1_DSP_bot/ConfigBits\[228\] Tile_X0Y1_DSP_bot/ConfigBits\[229\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_AB_BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__80_ net348 VGND VGND VPWR VPWR net729
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_E6BEG_outbuf_1__0_ Tile_X0Y1_DSP_bot/E6BEG_i\[1\] VGND VGND VPWR
+ VPWR net606 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1011_ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/X
+ sky130_fd_sc_hd__and3_2
XFILLER_0_151_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_NN4BEG_outbuf_9__0_ Tile_X0Y1_DSP_bot/NN4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y1_NN4BEG\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit7 net78 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[61\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1209_ Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_149_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_S4END_inbuf_3__0_ net114 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/S4BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__01_ Tile_X0Y0_DSP_top/JE2BEG\[1\] VGND
+ VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/Q5 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9
+ Tile_X0Y1_DSP_bot/ConfigBits\[312\] Tile_X0Y1_DSP_bot/ConfigBits\[313\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit27 net68 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[17\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit16 net56 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[6\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput202 Tile_X0Y1_E6END[10] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
Xinput213 Tile_X0Y1_EE4END[0] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_2
Xinput224 Tile_X0Y1_EE4END[5] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_1
Xinput235 Tile_X0Y1_FrameData[15] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__buf_6
Xinput279 Tile_X0Y1_FrameStrobe[8] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_8
Xinput268 Tile_X0Y1_FrameStrobe[16] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_1
Xinput257 Tile_X0Y1_FrameData[6] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_8
Xinput246 Tile_X0Y1_FrameData[25] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput709 net709 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1560_ Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1560_/Y
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1491_ Tile_X0Y1_DSP_bot_Inst_MULADD__1489_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1485_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0963_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1180_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1491_/Y sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit0 net229 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[160\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_159_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_W6END_inbuf_7__0_ net164 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/W6BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__63_ Tile_X0Y0_S2BEG\[1\] VGND VGND
+ VPWR VPWR net676 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit10 net230 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[106\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit21 net242 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[117\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_E1BEG1 Tile_X0Y1_DSP_bot/Q4
+ Tile_X0Y1_DSP_bot/J2MID_EFb_BEG\[0\] Tile_X0Y1_DSP_bot/JN2BEG\[0\] Tile_X0Y1_DSP_bot/J_l_EF_BEG\[2\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[36\] Tile_X0Y1_DSP_bot/ConfigBits\[37\] VGND VGND
+ VPWR VPWR net584 sky130_fd_sc_hd__mux4_2
XFILLER_0_142_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1758_ net333 Tile_X0Y1_DSP_bot/C16 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1758_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1689_ Tile_X0Y1_DSP_bot_Inst_MULADD__1689_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1715_/D sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[362\] Tile_X0Y0_DSP_top/ConfigBits\[363\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_EE4BEG_outbuf_6__0_ Tile_X0Y0_DSP_top/EE4BEG_i\[6\] VGND VGND VPWR
+ VPWR net426 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_S4END_inbuf_3__0_ Tile_X0Y0_S4BEG\[7\] VGND VGND VPWR VPWR ANTENNA_108/DIODE
+ sky130_fd_sc_hd__buf_2
XFILLER_0_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG0 Tile_X0Y1_N2BEG\[6\]
+ net19 net151 Tile_X0Y0_DSP_top/JN2BEG\[5\] Tile_X0Y0_DSP_top/ConfigBits\[166\] Tile_X0Y0_DSP_top/ConfigBits\[167\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_54_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[18\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__o21ai_2
XFILLER_0_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0991_ Tile_X0Y1_DSP_bot_Inst_MULADD__0986_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0989_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/C
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y0_DSP_top_SS4END_inbuf_7__0_ net119 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/SS4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_1
Xoutput506 net506 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput517 net517 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput528 net528 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput539 net539 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1612_ Tile_X0Y1_DSP_bot_Inst_MULADD__1180_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1611_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/A sky130_fd_sc_hd__o31ai_4
XFILLER_0_157_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1543_ Tile_X0Y1_DSP_bot_Inst_MULADD__1502_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1542_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1505_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1545_/A
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_outbuf_18__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_18__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[18\] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1474_ Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1448_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1473_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1474_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_0_82_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit26 net67 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[48\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit15 net55 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[37\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__46_ net293 VGND VGND VPWR VPWR Tile_X0Y1_N2BEGb\[0\]
+ sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_W6END_inbuf_7__0_ net365 VGND VGND VPWR VPWR ANTENNA_112/DIODE
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[274\] Tile_X0Y0_DSP_top/ConfigBits\[275\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit5 net76 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[123\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 ANTENNA_105/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_137 net299 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_148 net345 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_159 Tile_X0Y0_SS4BEG\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[54\] Tile_X0Y0_DSP_top/ConfigBits\[55\] VGND VGND
+ VPWR VPWR net404 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit3 net254 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[259\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit31 net253 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[159\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit20 net241 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[148\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_N4BEG1 Tile_X0Y1_N2BEGb\[3\]
+ Tile_X0Y1_N4BEG\[2\] net21 Tile_X0Y1_bot2top\[5\] Tile_X0Y0_DSP_top/ConfigBits\[10\]
+ Tile_X0Y0_DSP_top/ConfigBits\[11\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG1 Tile_X0Y1_N2BEG\[3\]
+ net16 net96 net148 Tile_X0Y0_DSP_top/ConfigBits\[208\] Tile_X0Y0_DSP_top/ConfigBits\[209\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[1\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1190_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1019_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1189_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1190_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_EE4END_inbuf_6__0_ net34 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/EE4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_109_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0974_ Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/B Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0973_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0974_/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1526_ Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/B sky130_fd_sc_hd__nand4_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1457_ Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1424_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1424_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1458_/A sky130_fd_sc_hd__a32oi_4
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1388_ Tile_X0Y1_DSP_bot_Inst_MULADD__1365_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1387_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1291_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1318_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1421_/B sky130_fd_sc_hd__o2111ai_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[326\] Tile_X0Y0_DSP_top/ConfigBits\[327\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__29_ Tile_X0Y1_DSP_bot/JE2BEG\[7\] VGND
+ VGND VPWR VPWR net594 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_N4BEG_outbuf_5__0_ Tile_X0Y1_DSP_bot/N4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N4BEG\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit6 net257 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[6\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit14 net54 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[68\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit25 net66 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[79\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1311_ Tile_X0Y1_DSP_bot_Inst_MULADD__1273_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1284_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1290_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1311_/Y
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1242_ Tile_X0Y1_DSP_bot_Inst_MULADD__1236_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1235_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1242_/Y sky130_fd_sc_hd__a22oi_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1173_ Tile_X0Y1_DSP_bot_Inst_MULADD__0888_/X Tile_X0Y1_DSP_bot_Inst_MULADD__0889_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1173_/Y
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_117_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_37 Tile_X0Y1_FrameStrobe_O\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 Tile_X0Y1_FrameStrobe_O\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 Tile_X0Y0_SS4BEG\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_48 Tile_X0Y1_FrameStrobe_O\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[24\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_NN4BEG\[12\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_59 ANTENNA_59/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0957_ Tile_X0Y1_DSP_bot_Inst_MULADD__0957_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q3 sky130_fd_sc_hd__buf_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0888_ Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1727_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0888_/X sky130_fd_sc_hd__and2_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit8 net79 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[222\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1509_ Tile_X0Y1_DSP_bot_Inst_MULADD__1503_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1506_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1508_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1511_/A
+ sky130_fd_sc_hd__o21a_1
XTile_X0Y0_DSP_top_strobe_outbuf_13__0_ Tile_X0Y0_DSP_top_strobe_inbuf_13__0_/X VGND
+ VGND VPWR VPWR net466 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_W6BEG_outbuf_5__0_ Tile_X0Y1_DSP_bot/W6BEG_i\[5\] VGND VGND VPWR
+ VPWR net742 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_data_outbuf_3__0_ Tile_X0Y0_DSP_top_data_inbuf_3__0_/X VGND VGND
+ VPWR VPWR net455 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit30 net252 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[190\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst1
+ net763 ANTENNA_101/DIODE Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[1\] Tile_X0Y1_DSP_bot/J2END_GH_BEG\[0\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[42\] Tile_X0Y1_DSP_bot/ConfigBits\[43\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit6 net257 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[358\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_158_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst0
+ net281 net181 net334 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[28\] Tile_X0Y1_DSP_bot/ConfigBits\[29\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput13 Tile_X0Y0_E2MID[0] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[292\] Tile_X0Y0_DSP_top/ConfigBits\[293\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JE2BEG\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_83_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput24 Tile_X0Y0_E6END[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_4
Xinput46 Tile_X0Y0_EE4END[7] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput35 Tile_X0Y0_EE4END[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[348\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[349\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
Xinput68 Tile_X0Y0_FrameData[27] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_4
Xinput57 Tile_X0Y0_FrameData[17] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_8
Xinput79 Tile_X0Y0_FrameData[8] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_4
XTile_X0Y0_DSP_top_data_inbuf_27__0_ net68 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_27__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0
+ net281 net287 net309 net187 Tile_X0Y1_DSP_bot/ConfigBits\[292\] Tile_X0Y1_DSP_bot/ConfigBits\[293\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0
+ net184 net337 Tile_X0Y1_DSP_bot/Q0 net764 Tile_X0Y1_DSP_bot/ConfigBits\[54\] Tile_X0Y1_DSP_bot/ConfigBits\[55\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1225_ Tile_X0Y1_DSP_bot_Inst_MULADD__1219_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1218_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1207_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1216_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/B sky130_fd_sc_hd__o211ai_4
XFILLER_0_157_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1156_ Tile_X0Y1_DSP_bot_Inst_MULADD__1114_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1120_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1132_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1156_/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1087_ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/D sky130_fd_sc_hd__nand4_4
XFILLER_0_74_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_data_inbuf_18__0_ net58 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_18__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_N4BEG_outbuf_1__0_ ANTENNA_74/DIODE VGND VGND VPWR VPWR net509
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[97\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_data_outbuf_3__0_ Tile_X0Y1_DSP_bot_data_inbuf_3__0_/X VGND VGND
+ VPWR VPWR net656 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[3\] Tile_X0Y1_N2BEGb\[1\] net6 net24 Tile_X0Y0_DSP_top/ConfigBits\[342\]
+ Tile_X0Y0_DSP_top/ConfigBits\[343\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_data_outbuf_25__0_ Tile_X0Y1_DSP_bot_data_inbuf_25__0_/X VGND VGND
+ VPWR VPWR net648 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG3 net285
+ net185 Tile_X0Y0_S2BEGb\[0\] net375 Tile_X0Y1_DSP_bot/ConfigBits\[230\] Tile_X0Y1_DSP_bot/ConfigBits\[231\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_AB_BEG\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_158_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1010_ Tile_X0Y1_DSP_bot_Inst_MULADD__1006_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1001_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1006_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1074_/A
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_data_inbuf_27__0_ net248 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_27__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_data_outbuf_16__0_ Tile_X0Y1_DSP_bot_data_inbuf_16__0_/X VGND VGND
+ VPWR VPWR net638 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit8 net79 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[62\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1208_ Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/A sky130_fd_sc_hd__buf_4
XTile_X0Y0_DSP_top_data_inbuf_9__0_ net80 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_9__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_S4BEG_outbuf_5__0_ Tile_X0Y1_DSP_bot/S4BEG_i\[5\] VGND VGND VPWR
+ VPWR net694 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1139_ Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1043_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1140_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_W6BEG_outbuf_1__0_ Tile_X0Y0_DSP_top/W6BEG_i\[1\] VGND VGND VPWR
+ VPWR net558 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__00_ Tile_X0Y0_DSP_top/JE2BEG\[0\] VGND
+ VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit28 net69 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[18\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit17 net57 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[7\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[314\] Tile_X0Y1_DSP_bot/ConfigBits\[315\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JE2BEG\[6\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_data_inbuf_18__0_ net238 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_18__0_/X
+ sky130_fd_sc_hd__clkbuf_1
Xinput214 Tile_X0Y1_EE4END[10] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
Xinput225 Tile_X0Y1_EE4END[6] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_1
Xinput203 Tile_X0Y1_E6END[11] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
Xinput236 Tile_X0Y1_FrameData[16] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__buf_4
Xinput269 Tile_X0Y1_FrameStrobe[17] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
Xinput258 Tile_X0Y1_FrameData[7] VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_8
Xinput247 Tile_X0Y1_FrameData[26] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1490_ Tile_X0Y1_DSP_bot_Inst_MULADD__1097_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1485_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1489_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1490_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_0_146_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit1 net240 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[161\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit0 net49 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[342\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__62_ Tile_X0Y0_S2BEG\[0\] VGND VGND
+ VPWR VPWR net675 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit11 net231 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[107\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit22 net243 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[118\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_E1BEG2 Tile_X0Y1_DSP_bot/Q5
+ Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[1\] ANTENNA_106/DIODE Tile_X0Y1_DSP_bot/J_l_GH_BEG\[3\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[38\] Tile_X0Y1_DSP_bot/ConfigBits\[39\] VGND VGND
+ VPWR VPWR net585 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1757_ net333 Tile_X0Y1_DSP_bot/C15 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1688_ Tile_X0Y1_DSP_bot_Inst_MULADD__1674_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1688_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1689_/A sky130_fd_sc_hd__and2b_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_outbuf_30__0_ Tile_X0Y0_DSP_top_data_inbuf_30__0_/X VGND VGND
+ VPWR VPWR net453 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[364\] Tile_X0Y0_DSP_top/ConfigBits\[365\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JW2BEG\[5\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[2\] net83 net135 Tile_X0Y1_bot2top\[2\] Tile_X0Y0_DSP_top/ConfigBits\[92\]
+ Tile_X0Y0_DSP_top/ConfigBits\[93\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0
+ net283 net289 net189 net201 Tile_X0Y1_DSP_bot/ConfigBits\[364\] Tile_X0Y1_DSP_bot/ConfigBits\[365\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_160_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[103\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__o21ai_1
XTile_X0Y0_DSP_top_data_outbuf_21__0_ Tile_X0Y0_DSP_top_data_inbuf_21__0_/X VGND VGND
+ VPWR VPWR net443 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG1 Tile_X0Y1_N2BEG\[2\]
+ net15 net95 Tile_X0Y0_DSP_top/JE2BEG\[5\] Tile_X0Y0_DSP_top/ConfigBits\[168\] Tile_X0Y0_DSP_top/ConfigBits\[169\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[1\] sky130_fd_sc_hd__mux4_1
XFILLER_0_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0990_ Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_81_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[18\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
Xoutput518 net518 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput507 net507 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput529 net529 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[5] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1611_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1564_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1565_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1611_/X sky130_fd_sc_hd__o221a_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1542_ Tile_X0Y1_DSP_bot_Inst_MULADD__1536_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1498_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1499_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1542_/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1473_ Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1452_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1473_/X
+ sky130_fd_sc_hd__a21bo_1
XTile_X0Y0_DSP_top_data_outbuf_12__0_ Tile_X0Y0_DSP_top_data_inbuf_12__0_/X VGND VGND
+ VPWR VPWR net433 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit16 net56 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[38\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit27 net68 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[49\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__45_ ANTENNA_183/DIODE VGND VGND VPWR
+ VPWR Tile_X0Y1_N2BEG\[7\] sky130_fd_sc_hd__buf_2
XFILLER_0_72_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_S4BEG_outbuf_1__0_ Tile_X0Y0_DSP_top/S4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y0_S4BEG\[1\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[274\] Tile_X0Y0_DSP_top/ConfigBits\[275\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit6 net77 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[124\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_105 ANTENNA_105/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_149 net366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_138 net299 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit4 net255 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[260\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit21 net242 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[149\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit10 net230 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[138\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_N4BEG2 Tile_X0Y1_N2BEGb\[0\]
+ Tile_X0Y1_N4BEG\[3\] net156 Tile_X0Y1_bot2top\[6\] Tile_X0Y0_DSP_top/ConfigBits\[12\]
+ Tile_X0Y0_DSP_top/ConfigBits\[13\] VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG2 Tile_X0Y1_N2BEG\[5\]
+ net18 net98 net150 Tile_X0Y0_DSP_top/ConfigBits\[210\] Tile_X0Y0_DSP_top/ConfigBits\[211\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[2\] sky130_fd_sc_hd__mux4_1
XFILLER_0_156_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0973_ Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0973_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_0_112_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_strobe_outbuf_5__0_ Tile_X0Y0_DSP_top_strobe_inbuf_5__0_/X VGND
+ VGND VPWR VPWR net477 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1525_ Tile_X0Y1_DSP_bot_Inst_MULADD__1503_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1506_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1508_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1474_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1454_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/D sky130_fd_sc_hd__o2111a_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1456_ Tile_X0Y1_DSP_bot_Inst_MULADD__1419_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1424_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1458_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1471_/A
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1387_ Tile_X0Y1_DSP_bot_Inst_MULADD__1382_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1365_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1386_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1387_/Y
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_77_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[328\] Tile_X0Y0_DSP_top/ConfigBits\[329\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JS2BEG\[4\] sky130_fd_sc_hd__mux4_2
XFILLER_0_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__28_ Tile_X0Y1_DSP_bot/JE2BEG\[6\] VGND
+ VGND VPWR VPWR net593 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0
+ net326 net182 net188 net204 Tile_X0Y1_DSP_bot/ConfigBits\[328\] Tile_X0Y1_DSP_bot/ConfigBits\[329\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit7 net258 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[7\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_data_inbuf_2__0_ net251 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_2__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_NN4END_inbuf_7__0_ Tile_X0Y1_NN4BEG\[11\] VGND VGND VPWR VPWR ANTENNA_181/DIODE
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit15 net55 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[69\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit26 net67 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[80\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_WW4BEG_outbuf_3__0_ Tile_X0Y0_DSP_top/WW4BEG_i\[3\] VGND VGND VPWR
+ VPWR net576 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1310_ Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1398_/B
+ sky130_fd_sc_hd__and3_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1241_ Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1172_ Tile_X0Y1_DSP_bot_Inst_MULADD__1034_/X Tile_X0Y1_DSP_bot/B5
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1035_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1113_/C
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1172_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_0_86_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_27 Tile_X0Y1_FrameStrobe_O\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 Tile_X0Y1_FrameStrobe_O\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_16 Tile_X0Y0_SS4BEG\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[24\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XANTENNA_49 Tile_X0Y1_FrameStrobe_O\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0956_ Tile_X0Y1_DSP_bot_Inst_MULADD__1677_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1709_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0957_/A
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0887_ Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0885_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0886_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0887_/X
+ sky130_fd_sc_hd__o21a_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit9 net80 Tile_X0Y1_FrameStrobe_O\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[223\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame5_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1508_ Tile_X0Y1_DSP_bot_Inst_MULADD__1507_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1506_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1506_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1508_/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1439_ Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/B sky130_fd_sc_hd__nand4_4
XFILLER_0_144_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_strobe_inbuf_13__0_ net265 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_13__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_N4END_inbuf_11__0_ net307 VGND VGND VPWR VPWR ANTENNA_185/DIODE
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit31 net253 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[191\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit20 net241 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[180\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput690 net690 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[1] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG0 net299
+ net199 Tile_X0Y0_S2BEG\[6\] Tile_X0Y1_DSP_bot/JN2BEG\[6\] Tile_X0Y1_DSP_bot/ConfigBits\[184\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[185\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit7 net258 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[359\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_68_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q8 ANTENNA_105/DIODE Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[1\] Tile_X0Y1_DSP_bot/J2END_CD_BEG\[1\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[28\] Tile_X0Y1_DSP_bot/ConfigBits\[29\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_N4END_inbuf_3__0_ Tile_X0Y1_N4BEG\[7\] VGND VGND VPWR VPWR ANTENNA_75/DIODE
+ sky130_fd_sc_hd__buf_2
Xinput25 Tile_X0Y0_E6END[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 Tile_X0Y0_EE4END[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput14 Tile_X0Y0_E2MID[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
XFILLER_0_107_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput69 Tile_X0Y0_FrameData[28] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_8
Xinput58 Tile_X0Y0_FrameData[18] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_6
XFILLER_0_134_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput47 Tile_X0Y0_EE4END[8] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[350\] Tile_X0Y1_DSP_bot/ConfigBits\[351\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JS2BEG\[7\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1
+ net201 Tile_X0Y0_S2BEGb\[2\] net340 net375 Tile_X0Y1_DSP_bot/ConfigBits\[292\] Tile_X0Y1_DSP_bot/ConfigBits\[293\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/Q5
+ Tile_X0Y1_DSP_bot/ConfigBits\[54\] Tile_X0Y1_DSP_bot/ConfigBits\[55\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1224_ Tile_X0Y1_DSP_bot_Inst_MULADD__1222_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1223_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1216_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/A
+ sky130_fd_sc_hd__o21bai_4
XFILLER_0_90_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1155_ Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[0\] net1 net81 Tile_X0Y1_bot2top\[4\] Tile_X0Y0_DSP_top/ConfigBits\[42\]
+ Tile_X0Y0_DSP_top/ConfigBits\[43\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1086_ Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1084_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/C
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_15_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0939_ Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/A sky130_fd_sc_hd__nand4_4
XFILLER_0_139_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[97\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1
+ net86 net108 net138 net156 Tile_X0Y0_DSP_top/ConfigBits\[342\] Tile_X0Y0_DSP_top/ConfigBits\[343\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_strobe_inbuf_6__0_ net277 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_6__0_/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_N4END_inbuf_3__0_ net314 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/N4BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit30 net252 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[222\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_149_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit9 net80 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[63\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_149_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1207_ Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1218_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1207_/X
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1138_ Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1140_/A sky130_fd_sc_hd__inv_2
XFILLER_0_145_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1069_ Tile_X0Y1_DSP_bot/C5 Tile_X0Y1_DSP_bot_Inst_MULADD__1747_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1459_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1069_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit29 net70 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[19\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit18 net58 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[8\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput226 Tile_X0Y1_EE4END[7] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
Xinput215 Tile_X0Y1_EE4END[11] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_1
Xinput204 Tile_X0Y1_E6END[1] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__buf_4
Xinput259 Tile_X0Y1_FrameData[8] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_8
Xinput237 Tile_X0Y1_FrameData[17] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__buf_4
Xinput248 Tile_X0Y1_FrameData[27] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0
+ Tile_X0Y1_N2BEGb\[3\] Tile_X0Y1_N4BEG\[3\] net2 net8 Tile_X0Y0_DSP_top/ConfigBits\[254\]
+ Tile_X0Y0_DSP_top/ConfigBits\[255\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_WW4BEG_outbuf_9__0_ Tile_X0Y1_DSP_bot/WW4BEG_i\[9\] VGND VGND VPWR
+ VPWR net762 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__59_ net148 VGND VGND VPWR VPWR net550
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit2 net251 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[162\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit1 net60 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[343\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__61_ Tile_X0Y1_DSP_bot/JS2BEG\[7\] VGND
+ VGND VPWR VPWR net674 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit23 net244 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[119\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit12 net232 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[108\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_E1BEG3 net763 Tile_X0Y1_DSP_bot/J2MID_ABb_BEG\[2\]
+ Tile_X0Y1_DSP_bot/JN2BEG\[2\] Tile_X0Y1_DSP_bot/J_l_AB_BEG\[0\] Tile_X0Y1_DSP_bot/ConfigBits\[40\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[41\] VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__mux4_2
XFILLER_0_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1756_ net333 Tile_X0Y1_DSP_bot/C14 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1756_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1687_ Tile_X0Y1_DSP_bot_Inst_MULADD__1687_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1714_/D sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst0
+ net281 net181 net334 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[84\] Tile_X0Y1_DSP_bot/ConfigBits\[85\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[6\] Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[1\] Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[1\]
+ ANTENNA_206/DIODE Tile_X0Y0_DSP_top/ConfigBits\[92\] Tile_X0Y0_DSP_top/ConfigBits\[93\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1
+ Tile_X0Y0_S2BEGb\[4\] Tile_X0Y0_S4BEG\[0\] net342 net354 Tile_X0Y1_DSP_bot/ConfigBits\[364\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[365\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_S4END_inbuf_11__0_ Tile_X0Y0_S4BEG\[15\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/S4BEG_i\[11\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_63_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[103\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top_strobe_inbuf_2__0_ Tile_X0Y1_FrameStrobe_O\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_2__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG2 Tile_X0Y1_N2BEG\[4\]
+ net97 net149 ANTENNA_64/DIODE Tile_X0Y0_DSP_top/ConfigBits\[170\] Tile_X0Y0_DSP_top/ConfigBits\[171\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_26_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
Xoutput508 net508 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput519 net519 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1610_ Tile_X0Y1_DSP_bot_Inst_MULADD__1608_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1698_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1720_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q14 sky130_fd_sc_hd__a2bb2o_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1541_ Tile_X0Y1_DSP_bot_Inst_MULADD__1541_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1541_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1541_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1545_/C
+ sky130_fd_sc_hd__nor3_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1472_ Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1465_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1518_/B
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit17 net57 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[39\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit28 net69 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[50\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_119_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__44_ Tile_X0Y1_DSP_bot/JN2BEG\[6\] VGND
+ VGND VPWR VPWR Tile_X0Y1_N2BEG\[6\] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_NN4BEG_outbuf_6__0_ Tile_X0Y0_DSP_top/NN4BEG_i\[6\] VGND VGND VPWR
+ VPWR net530 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[276\] Tile_X0Y0_DSP_top/ConfigBits\[277\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JN2BEG\[7\] sky130_fd_sc_hd__mux4_2
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0
+ net283 net291 net183 net191 Tile_X0Y1_DSP_bot/ConfigBits\[276\] Tile_X0Y1_DSP_bot/ConfigBits\[277\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit7 net78 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[125\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1739_ net333 Tile_X0Y1_DSP_bot/B5 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1739_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 ANTENNA_106/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 net314 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_SS4BEG_outbuf_9__0_ Tile_X0Y0_DSP_top/SS4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_SS4BEG\[9\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit5 net256 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[261\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_SS4END_inbuf_1__0_ Tile_X0Y0_SS4BEG\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/SS4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit11 net231 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[139\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit22 net243 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[150\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG3 Tile_X0Y1_N2BEG\[1\]
+ net14 net94 net146 Tile_X0Y0_DSP_top/ConfigBits\[212\] Tile_X0Y0_DSP_top/ConfigBits\[213\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[3\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_N4BEG3 Tile_X0Y1_N2BEGb\[1\]
+ Tile_X0Y1_N4BEG\[0\] net153 Tile_X0Y1_bot2top\[7\] Tile_X0Y0_DSP_top/ConfigBits\[14\]
+ Tile_X0Y0_DSP_top/ConfigBits\[15\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__mux4_2
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_SS4BEG_outbuf_2__0_ Tile_X0Y1_DSP_bot/SS4BEG_i\[2\] VGND VGND VPWR
+ VPWR net707 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0972_ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/A sky130_fd_sc_hd__nand4_4
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1524_ Tile_X0Y1_DSP_bot_Inst_MULADD__1604_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1690_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1604_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1605_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1557_/A sky130_fd_sc_hd__a31oi_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1455_ Tile_X0Y1_DSP_bot_Inst_MULADD__1446_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1450_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1454_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1458_/B
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1386_ Tile_X0Y1_DSP_bot_Inst_MULADD__1386_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1386_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1386_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__27_ Tile_X0Y1_DSP_bot/JE2BEG\[5\] VGND
+ VGND VPWR VPWR net592 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1
+ Tile_X0Y0_S2BEGb\[3\] Tile_X0Y0_S4BEG\[3\] net341 net357 Tile_X0Y1_DSP_bot/ConfigBits\[328\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[329\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit8 net259 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[8\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_5_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit27 net68 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[81\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit16 net56 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[70\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_EE4END_inbuf_0__0_ net223 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/EE4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_47_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1240_ Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1230_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1239_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1248_/A sky130_fd_sc_hd__o32ai_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1171_ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1171_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_WW4END_inbuf_8__0_ net168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/WW4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_39 Tile_X0Y1_FrameStrobe_O\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_17 Tile_X0Y0_SS4BEG\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 Tile_X0Y1_FrameStrobe_O\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_15_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0955_ Tile_X0Y1_DSP_bot_Inst_MULADD__0955_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0954_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1677_/B sky130_fd_sc_hd__or2b_1
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__0886_ Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1728_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0886_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1507_ Tile_X0Y1_DSP_bot_Inst_MULADD__1505_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1505_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1502_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1507_/X
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1438_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1435_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/D
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1369_ Tile_X0Y1_DSP_bot_Inst_MULADD__1369_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1369_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1369_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_53_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit10 net230 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[170\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit21 net242 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[181\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput680 net680 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput691 net691 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG1 net295
+ Tile_X0Y0_S2BEG\[2\] net348 Tile_X0Y1_DSP_bot/JE2BEG\[6\] Tile_X0Y1_DSP_bot/ConfigBits\[186\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[187\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit8 net259 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[360\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput26 Tile_X0Y0_E6END[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput37 Tile_X0Y0_EE4END[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput15 Tile_X0Y0_E2MID[2] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
XFILLER_0_24_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput59 Tile_X0Y0_FrameData[19] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_6
XFILLER_0_134_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput48 Tile_X0Y0_EE4END[9] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire763 wire763/A VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__buf_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4
+ Tile_X0Y1_DSP_bot/ConfigBits\[292\] Tile_X0Y1_DSP_bot/ConfigBits\[293\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2
+ net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[54\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[55\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_E6BEG_outbuf_4__0_ Tile_X0Y1_DSP_bot/E6BEG_i\[4\] VGND VGND VPWR
+ VPWR net609 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1223_ Tile_X0Y1_DSP_bot_Inst_MULADD__1210_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1211_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1212_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1223_/X sky130_fd_sc_hd__o2111a_1
XFILLER_0_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1154_ Tile_X0Y1_DSP_bot_Inst_MULADD__1154_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/B sky130_fd_sc_hd__inv_2
XFILLER_0_157_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[8\] Tile_X0Y0_DSP_top/J2MID_EFb_BEG\[1\] Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2END_CD_BEG\[0\] Tile_X0Y0_DSP_top/ConfigBits\[42\] Tile_X0Y0_DSP_top/ConfigBits\[43\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1085_ Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1732_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_62_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0938_ Tile_X0Y1_DSP_bot_Inst_MULADD__1201_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/A sky130_fd_sc_hd__buf_6
XTile_X0Y0_DSP_top_N4BEG_outbuf_10__0_ ANTENNA_68/DIODE VGND VGND VPWR VPWR net503
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0869_ Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/D Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0878_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_155_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_93_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_S4END_inbuf_6__0_ net102 VGND VGND VPWR VPWR ANTENNA_91/DIODE sky130_fd_sc_hd__clkbuf_2
XFILLER_0_148_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[342\] Tile_X0Y0_DSP_top/ConfigBits\[343\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit31 net253 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[223\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit20 net241 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[212\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1206_ Tile_X0Y1_DSP_bot_Inst_MULADD__1202_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1204_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1205_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1218_/B
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_125_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1137_ Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1136_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1137_/Y
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_157_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1068_ Tile_X0Y1_DSP_bot_Inst_MULADD__1050_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1053_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1081_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1002_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1072_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_0_145_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit19 net59 Tile_X0Y1_FrameStrobe_O\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[9\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame12_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput227 Tile_X0Y1_EE4END[8] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_1
Xinput205 Tile_X0Y1_E6END[2] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_1
Xinput216 Tile_X0Y1_EE4END[12] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_1
Xinput238 Tile_X0Y1_FrameData[18] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_8
Xinput249 Tile_X0Y1_FrameData[28] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_8
XTile_X0Y0_DSP_top_EE4BEG_outbuf_9__0_ Tile_X0Y0_DSP_top/EE4BEG_i\[9\] VGND VGND VPWR
+ VPWR net429 sky130_fd_sc_hd__clkbuf_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_C0 Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[0\]
+ Tile_X0Y1_DSP_bot/J2MID_EFb_BEG\[0\] Tile_X0Y1_DSP_bot/J2END_EF_BEG\[0\] Tile_X0Y1_DSP_bot/J_l_EF_BEG\[0\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[134\] Tile_X0Y1_DSP_bot/ConfigBits\[135\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C0 sky130_fd_sc_hd__mux4_1
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1
+ net24 net88 net140 net172 Tile_X0Y0_DSP_top/ConfigBits\[254\] Tile_X0Y0_DSP_top/ConfigBits\[255\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_S4END_inbuf_6__0_ Tile_X0Y0_S4BEG\[10\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/S4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_104_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__58_ net147 VGND VGND VPWR VPWR net549
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit3 net254 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[163\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit2 net71 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[344\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_159_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_E6BEG_outbuf_0__0_ Tile_X0Y0_DSP_top/E6BEG_i\[0\] VGND VGND VPWR
+ VPWR net402 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__60_ Tile_X0Y1_DSP_bot/JS2BEG\[6\] VGND
+ VGND VPWR VPWR net673 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_EE4BEG_outbuf_2__0_ Tile_X0Y1_DSP_bot/EE4BEG_i\[2\] VGND VGND VPWR
+ VPWR net623 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit24 net245 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[120\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit13 net233 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[109\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1755_ net333 Tile_X0Y1_DSP_bot/C13 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1686_ Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1686_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1686_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1687_/A
+ sky130_fd_sc_hd__and3b_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q8 ANTENNA_105/DIODE Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[1\] Tile_X0Y1_DSP_bot/J2END_CD_BEG\[3\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[84\] Tile_X0Y1_DSP_bot/ConfigBits\[85\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[364\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[365\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[1\] Tile_X0Y1_N2BEGb\[5\] net2 net10 Tile_X0Y0_DSP_top/ConfigBits\[294\]
+ Tile_X0Y0_DSP_top/ConfigBits\[295\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG3 net13
+ net93 net145 Tile_X0Y0_DSP_top/JW2BEG\[5\] Tile_X0Y0_DSP_top/ConfigBits\[172\] Tile_X0Y0_DSP_top/ConfigBits\[173\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_151_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput509 net509 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit30 net252 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[254\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_157_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1540_ Tile_X0Y1_DSP_bot_Inst_MULADD__1541_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1541_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1541_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1545_/B
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1471_ Tile_X0Y1_DSP_bot_Inst_MULADD__1471_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1471_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1471_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1518_/A
+ sky130_fd_sc_hd__and3_1
XFILLER_0_147_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit29 net70 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[51\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit18 net58 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[40\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__43_ Tile_X0Y1_DSP_bot/JN2BEG\[5\] VGND
+ VGND VPWR VPWR Tile_X0Y1_N2BEG\[5\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_EE4END_inbuf_9__0_ net37 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/EE4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit8 net79 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[126\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[2\] Tile_X0Y0_S2BEGb\[6\] net334 net336 Tile_X0Y1_DSP_bot/ConfigBits\[276\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[277\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1738_ net333 Tile_X0Y1_DSP_bot/B4 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1738_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1669_ Tile_X0Y1_DSP_bot_Inst_MULADD__1666_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1668_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1669_/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_107 ANTENNA_107/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_118 net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_129 net184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top_WW4BEG_outbuf_10__0_ Tile_X0Y0_DSP_top/WW4BEG_i\[10\] VGND VGND
+ VPWR VPWR net568 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_N4BEG_outbuf_8__0_ Tile_X0Y1_DSP_bot/N4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N4BEG\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit12 net232 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[140\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit23 net244 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[151\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit6 net257 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[262\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_129_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__0971_ Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/C Tile_X0Y1_DSP_bot_Inst_MULADD__0970_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/A sky130_fd_sc_hd__a41oi_4
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1523_ Tile_X0Y1_DSP_bot_Inst_MULADD__1523_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1523_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1523_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1604_/B
+ sky130_fd_sc_hd__nand3_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1454_ Tile_X0Y1_DSP_bot_Inst_MULADD__1446_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1452_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1453_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1454_/Y
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1385_ Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1386_/B
+ sky130_fd_sc_hd__and3_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0
+ net281 net285 net181 net185 Tile_X0Y1_DSP_bot/ConfigBits\[316\] Tile_X0Y1_DSP_bot/ConfigBits\[317\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__26_ Tile_X0Y1_DSP_bot/JE2BEG\[4\] VGND
+ VGND VPWR VPWR net591 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 net764 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[328\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[329\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit9 net260 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[9\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame12_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_strobe_outbuf_16__0_ Tile_X0Y0_DSP_top_strobe_inbuf_16__0_/X VGND
+ VGND VPWR VPWR net469 sky130_fd_sc_hd__clkbuf_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_W6BEG_outbuf_8__0_ Tile_X0Y1_DSP_bot/W6BEG_i\[8\] VGND VGND VPWR
+ VPWR net745 sky130_fd_sc_hd__clkbuf_1
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_data_outbuf_6__0_ Tile_X0Y0_DSP_top_data_inbuf_6__0_/X VGND VGND
+ VPWR VPWR net458 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit28 net69 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[82\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit17 net57 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[71\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG0 Tile_X0Y1_N2BEGb\[7\]
+ net12 net92 net165 Tile_X0Y0_DSP_top/ConfigBits\[238\] Tile_X0Y0_DSP_top/ConfigBits\[239\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_GH_BEG\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1170_ Tile_X0Y1_DSP_bot_Inst_MULADD__1165_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1165_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1165_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1167_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1166_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1255_/A sky130_fd_sc_hd__a32oi_4
XANTENNA_29 Tile_X0Y1_FrameStrobe_O\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_18 Tile_X0Y0_SS4BEG\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[3\] Tile_X0Y1_N2BEGb\[7\] net4 net12 Tile_X0Y0_DSP_top/ConfigBits\[366\]
+ Tile_X0Y0_DSP_top/ConfigBits\[367\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__0954_ Tile_X0Y1_DSP_bot_Inst_MULADD__0953_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0953_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0953_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0954_/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0885_ Tile_X0Y1_DSP_bot/A2 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0885_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1506_ Tile_X0Y1_DSP_bot_Inst_MULADD__1506_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1506_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1506_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1437_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/X sky130_fd_sc_hd__or4_1
XFILLER_0_144_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1368_ Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1368_/X sky130_fd_sc_hd__a211o_1
XTile_X0Y1_DSP_bot_NN4END_inbuf_1__0_ net328 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/NN4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1299_ Tile_X0Y1_DSP_bot_Inst_MULADD__1373_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1373_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1299_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1299_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1299_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_58_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__09_ Tile_X0Y0_top2bot\[5\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/B5 sky130_fd_sc_hd__buf_2
XFILLER_0_73_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_N4BEG_outbuf_4__0_ ANTENNA_207/DIODE VGND VGND VPWR VPWR net512
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit22 net243 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[182\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit11 net231 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[171\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput681 net681 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput670 net670 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput692 net692 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG2 net197
+ Tile_X0Y0_S2BEG\[4\] net350 Tile_X0Y1_DSP_bot/JS2BEG\[6\] Tile_X0Y1_DSP_bot/ConfigBits\[188\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[189\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[2\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_158_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit9 net260 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[361\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_data_outbuf_6__0_ Tile_X0Y1_DSP_bot_data_inbuf_6__0_/X VGND VGND
+ VPWR VPWR net659 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput27 Tile_X0Y0_E6END[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput16 Tile_X0Y0_E2MID[3] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
XFILLER_0_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput49 Tile_X0Y0_FrameData[0] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_8
Xinput38 Tile_X0Y0_EE4END[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[292\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[293\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit0 net49 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[246\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3
+ ANTENNA_101/DIODE Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[1\] ANTENNA_105/DIODE Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[1\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[54\] Tile_X0Y1_DSP_bot/ConfigBits\[55\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_data_outbuf_28__0_ Tile_X0Y1_DSP_bot_data_inbuf_28__0_/X VGND VGND
+ VPWR VPWR net651 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1222_ Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1218_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1222_/Y
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1153_ Tile_X0Y1_DSP_bot_Inst_MULADD__1080_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1081_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1144_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1152_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1165_/A sky130_fd_sc_hd__o22ai_4
XFILLER_0_157_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1084_ Tile_X0Y1_DSP_bot/A6 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1084_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0937_ Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0935_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0936_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1201_/B
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_140_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0868_ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0939_/B sky130_fd_sc_hd__buf_4
XFILLER_0_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_data_outbuf_19__0_ Tile_X0Y1_DSP_bot_data_inbuf_19__0_/X VGND VGND
+ VPWR VPWR net641 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_S4BEG_outbuf_8__0_ Tile_X0Y1_DSP_bot/S4BEG_i\[8\] VGND VGND VPWR
+ VPWR net697 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_W6BEG_outbuf_4__0_ Tile_X0Y0_DSP_top/W6BEG_i\[4\] VGND VGND VPWR
+ VPWR net561 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[342\] Tile_X0Y0_DSP_top/ConfigBits\[343\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[2\] Tile_X0Y1_N2BEGb\[6\] net3 net11 Tile_X0Y0_DSP_top/ConfigBits\[330\]
+ Tile_X0Y0_DSP_top/ConfigBits\[331\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit10 net230 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[202\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit21 net242 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[213\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_125_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1205_ Tile_X0Y1_DSP_bot_Inst_MULADD__1378_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1204_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1201_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1205_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_0_87_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1136_ Tile_X0Y1_DSP_bot_Inst_MULADD__1054_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1055_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1044_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1136_/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_157_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1067_ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1154_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1072_/C
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput217 Tile_X0Y1_EE4END[13] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_1
Xinput206 Tile_X0Y1_E6END[3] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_E6END_inbuf_2__0_ net27 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/E6BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
Xinput228 Tile_X0Y1_EE4END[9] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
Xinput239 Tile_X0Y1_FrameData[19] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_8
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_C1 Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[1\]
+ ANTENNA_105/DIODE Tile_X0Y1_DSP_bot/J2END_EF_BEG\[1\] Tile_X0Y1_DSP_bot/J_l_EF_BEG\[1\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[136\] Tile_X0Y1_DSP_bot/ConfigBits\[137\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C1 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_B0 Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[0\]
+ Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[0\] Tile_X0Y1_DSP_bot/J2END_CD_BEG\[0\] Tile_X0Y1_DSP_bot/J_l_CD_BEG\[0\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[126\] Tile_X0Y1_DSP_bot/ConfigBits\[127\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/B0 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_strobe_inbuf_10__0_ Tile_X0Y1_FrameStrobe_O\[10\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_10__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[254\] Tile_X0Y0_DSP_top/ConfigBits\[255\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__57_ net146 VGND VGND VPWR VPWR net548
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit4 net255 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[164\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_data_outbuf_24__0_ Tile_X0Y0_DSP_top_data_inbuf_24__0_/X VGND VGND
+ VPWR VPWR net446 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit3 net74 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[345\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_159_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit25 net246 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[121\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit14 net234 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[110\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1754_ net333 Tile_X0Y1_DSP_bot/C12 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1754_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1685_ Tile_X0Y1_DSP_bot_Inst_MULADD__1685_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1713_/D sky130_fd_sc_hd__clkbuf_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_data_outbuf_15__0_ Tile_X0Y0_DSP_top_data_inbuf_15__0_/X VGND VGND
+ VPWR VPWR net436 sky130_fd_sc_hd__clkbuf_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[364\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[365\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_S4BEG_outbuf_4__0_ ANTENNA_87/DIODE VGND VGND VPWR VPWR Tile_X0Y0_S4BEG\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1119_ Tile_X0Y1_DSP_bot_Inst_MULADD__1116_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1117_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/B
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_75_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1
+ net82 net84 net90 net134 Tile_X0Y0_DSP_top/ConfigBits\[294\] Tile_X0Y0_DSP_top/ConfigBits\[295\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_E6END_inbuf_2__0_ net207 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/E6BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit31 net253 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[255\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit20 net241 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[244\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_157_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1470_ Tile_X0Y1_DSP_bot_Inst_MULADD__1258_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1690_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1690_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1469_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q10 sky130_fd_sc_hd__a31o_1
XFILLER_0_89_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit19 net59 Tile_X0Y1_FrameStrobe_O\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[41\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame11_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__42_ Tile_X0Y1_DSP_bot/JN2BEG\[4\] VGND
+ VGND VPWR VPWR Tile_X0Y1_N2BEG\[4\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_strobe_outbuf_8__0_ Tile_X0Y0_DSP_top_strobe_inbuf_8__0_/X VGND
+ VGND VPWR VPWR net480 sky130_fd_sc_hd__buf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit9 net80 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[127\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[276\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[277\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1737_ net333 Tile_X0Y1_DSP_bot/B3 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1737_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1668_ Tile_X0Y1_DSP_bot_Inst_MULADD__1665_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1657_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1665_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1667_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1668_/Y sky130_fd_sc_hd__o211ai_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1599_ Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/A
+ sky130_fd_sc_hd__a21o_1
XANTENNA_119 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_108 ANTENNA_108/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_data_inbuf_5__0_ net256 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_5__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_strobe_outbuf_1__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_1__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[1\] sky130_fd_sc_hd__buf_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit13 net233 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[141\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit7 net258 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[263\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit24 net245 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[152\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_98_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0970_ Tile_X0Y1_DSP_bot_Inst_MULADD__0968_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0969_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0970_/Y
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_WW4BEG_outbuf_6__0_ Tile_X0Y0_DSP_top/WW4BEG_i\[6\] VGND VGND VPWR
+ VPWR net579 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1522_ Tile_X0Y1_DSP_bot_Inst_MULADD__1522_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q11 sky130_fd_sc_hd__buf_1
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1453_ Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1421_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1453_/X
+ sky130_fd_sc_hd__o21a_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1384_ Tile_X0Y1_DSP_bot_Inst_MULADD__1034_/X Tile_X0Y1_DSP_bot/B7
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1378_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1175_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/C sky130_fd_sc_hd__o211a_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[0\] Tile_X0Y0_S1BEG\[2\] Tile_X0Y0_SS4BEG\[0\] net366 Tile_X0Y1_DSP_bot/ConfigBits\[316\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[317\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_147_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__25_ Tile_X0Y1_DSP_bot/JE2BEG\[3\] VGND
+ VGND VPWR VPWR net590 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[328\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[329\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_strobe_inbuf_16__0_ net268 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_16__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit30 net252 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[286\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG0 Tile_X0Y1_N2BEG\[7\]
+ net20 net100 net152 Tile_X0Y0_DSP_top/ConfigBits\[182\] Tile_X0Y0_DSP_top/ConfigBits\[183\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit18 net58 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[72\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_102_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit29 net70 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[83\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_W1BEG0 Tile_X0Y1_bot2top\[5\]
+ Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[3\] Tile_X0Y0_DSP_top/JS2BEG\[3\] Tile_X0Y0_DSP_top/J_l_CD_BEG\[1\]
+ Tile_X0Y0_DSP_top/ConfigBits\[84\] Tile_X0Y0_DSP_top/ConfigBits\[85\] VGND VGND
+ VPWR VPWR net535 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG1 Tile_X0Y1_N2BEGb\[3\]
+ net8 net117 net140 Tile_X0Y0_DSP_top/ConfigBits\[240\] Tile_X0Y0_DSP_top/ConfigBits\[241\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_GH_BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_N4END_inbuf_6__0_ Tile_X0Y1_N4BEG\[10\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/N4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 Tile_X0Y0_SS4BEG\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1
+ net82 net84 net92 net136 Tile_X0Y0_DSP_top/ConfigBits\[366\] Tile_X0Y0_DSP_top/ConfigBits\[367\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0953_ Tile_X0Y1_DSP_bot_Inst_MULADD__0953_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0953_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0953_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0955_/A
+ sky130_fd_sc_hd__and3_1
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0884_ Tile_X0Y1_DSP_bot_Inst_MULADD__0878_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0906_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0878_/C Tile_X0Y1_DSP_bot_Inst_MULADD__0881_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1672_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0917_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1505_ Tile_X0Y1_DSP_bot_Inst_MULADD__1502_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1505_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1505_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1506_/B
+ sky130_fd_sc_hd__nand3b_1
XFILLER_0_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1436_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1269_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1435_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/C sky130_fd_sc_hd__o211ai_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1367_ Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1298_ Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/X sky130_fd_sc_hd__and4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__08_ Tile_X0Y0_top2bot\[4\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/B4 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit23 net244 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[183\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit12 net232 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[172\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput671 net671 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput660 net660 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[7] sky130_fd_sc_hd__buf_2
Xoutput682 net682 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput693 net693 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[4] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG3 net293
+ net193 net346 ANTENNA_184/DIODE Tile_X0Y1_DSP_bot/ConfigBits\[190\] Tile_X0Y1_DSP_bot/ConfigBits\[191\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput28 Tile_X0Y0_E6END[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput17 Tile_X0Y0_E2MID[4] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput39 Tile_X0Y0_EE4END[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_WW4END_inbuf_2__0_ net378 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/WW4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG0 net310
+ net188 net341 Tile_X0Y1_DSP_bot/JN2BEG\[3\] Tile_X0Y1_DSP_bot/ConfigBits\[400\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[401\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_EF_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[294\] Tile_X0Y1_DSP_bot/ConfigBits\[295\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JE2BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit1 net60 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[247\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[56\] Tile_X0Y1_DSP_bot/ConfigBits\[57\] VGND VGND
+ VPWR VPWR net604 sky130_fd_sc_hd__mux4_1
XFILLER_0_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_strobe_inbuf_9__0_ net280 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_9__0_/X
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1221_ Tile_X0Y1_DSP_bot_Inst_MULADD__1179_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1183_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1217_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1220_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1243_/B sky130_fd_sc_hd__o22ai_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1152_ Tile_X0Y1_DSP_bot_Inst_MULADD__1159_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1154_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1147_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1151_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1152_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1083_ Tile_X0Y1_DSP_bot_Inst_MULADD__1016_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1056_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1054_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/A
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_157_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_N4END_inbuf_6__0_ net302 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/N4BEG_i\[6\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_55_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_SS4BEG_outbuf_10__0_ Tile_X0Y0_DSP_top/SS4BEG_i\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y0_SS4BEG\[10\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0936_ Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1729_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0936_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0867_ Tile_X0Y1_DSP_bot/ConfigBits\[1\] Tile_X0Y1_DSP_bot_Inst_MULADD__0865_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0866_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/B
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_139_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1419_ Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1419_/Y
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_N4END_inbuf_10__0_ Tile_X0Y1_N4BEG\[14\] VGND VGND VPWR VPWR ANTENNA_68/DIODE
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput490 net490 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[4] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[344\] Tile_X0Y0_DSP_top/ConfigBits\[345\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JW2BEG\[0\] sky130_fd_sc_hd__mux4_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1
+ net83 net91 net133 net135 Tile_X0Y0_DSP_top/ConfigBits\[330\] Tile_X0Y0_DSP_top/ConfigBits\[331\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit11 net231 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[203\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit22 net243 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[214\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_79_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1204_ Tile_X0Y1_DSP_bot_Inst_MULADD__0933_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1203_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1204_/Y
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1135_ Tile_X0Y1_DSP_bot_Inst_MULADD__1026_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1062_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1135_/X sky130_fd_sc_hd__o211a_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1066_ Tile_X0Y1_DSP_bot_Inst_MULADD__1050_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1053_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1081_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1154_/A
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_28_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0919_ Tile_X0Y1_DSP_bot_Inst_MULADD__1675_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1708_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0920_/A
+ sky130_fd_sc_hd__mux2_1
Xinput218 Tile_X0Y1_EE4END[14] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_1
Xinput207 Tile_X0Y1_E6END[4] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_1
Xinput229 Tile_X0Y1_FrameData[0] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_A0 Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[0\]
+ Tile_X0Y1_DSP_bot/J2MID_ABb_BEG\[0\] Tile_X0Y1_DSP_bot/J2END_AB_BEG\[0\] Tile_X0Y1_DSP_bot/J_l_AB_BEG\[0\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[118\] Tile_X0Y1_DSP_bot/ConfigBits\[119\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/A0 sky130_fd_sc_hd__mux4_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_B1 Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[1\]
+ Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[1\] Tile_X0Y1_DSP_bot/J2END_CD_BEG\[1\] Tile_X0Y1_DSP_bot/J_l_CD_BEG\[1\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[128\] Tile_X0Y1_DSP_bot/ConfigBits\[129\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/B1 sky130_fd_sc_hd__mux4_2
XFILLER_0_46_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_C2 Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2MID_EFb_BEG\[2\] Tile_X0Y1_DSP_bot/J2END_EF_BEG\[2\] Tile_X0Y1_DSP_bot/J_l_EF_BEG\[2\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[138\] Tile_X0Y1_DSP_bot/ConfigBits\[139\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C2 sky130_fd_sc_hd__mux4_2
XFILLER_0_53_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[254\] Tile_X0Y0_DSP_top/ConfigBits\[255\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__56_ net145 VGND VGND VPWR VPWR net547
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit5 net256 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[165\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit4 net75 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[346\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_strobe_inbuf_5__0_ Tile_X0Y1_FrameStrobe_O\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_5__0_/X sky130_fd_sc_hd__buf_1
XFILLER_0_29_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit26 net247 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[122\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit15 net235 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[111\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1753_ net333 Tile_X0Y1_DSP_bot/C11 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1684_ Tile_X0Y1_DSP_bot_Inst_MULADD__1674_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1684_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1685_/A sky130_fd_sc_hd__and2b_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[366\] Tile_X0Y1_DSP_bot/ConfigBits\[367\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JW2BEG\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1118_ Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/Y sky130_fd_sc_hd__nand2_2
XTile_X0Y0_DSP_top_NN4BEG_outbuf_9__0_ Tile_X0Y0_DSP_top/NN4BEG_i\[9\] VGND VGND VPWR
+ VPWR net533 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1049_ Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0989_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0984_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1049_/Y
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[294\] Tile_X0Y0_DSP_top/ConfigBits\[295\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit10 net230 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[234\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit21 net242 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[245\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_NN4BEG_outbuf_2__0_ Tile_X0Y1_DSP_bot/NN4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y1_NN4BEG\[2\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__39_ ANTENNA_179/DIODE VGND VGND VPWR
+ VPWR Tile_X0Y0_S2BEG\[7\] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_SS4END_inbuf_4__0_ Tile_X0Y0_SS4BEG\[8\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/SS4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__41_ Tile_X0Y1_DSP_bot/JN2BEG\[3\] VGND
+ VGND VPWR VPWR Tile_X0Y1_N2BEG\[3\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_SS4BEG_outbuf_5__0_ Tile_X0Y1_DSP_bot/SS4BEG_i\[5\] VGND VGND VPWR
+ VPWR net710 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q4 wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[276\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[277\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1736_ net333 ANTENNA_97/DIODE VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1736_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1667_ Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1703_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1658_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1658_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1667_/Y sky130_fd_sc_hd__o2bb2ai_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1598_ Tile_X0Y1_DSP_bot_Inst_MULADD__1597_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1720_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1664_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/C
+ sky130_fd_sc_hd__mux2_1
XANTENNA_109 ANTENNA_110/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_S4END_inbuf_10__0_ net106 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/S4BEG_i\[10\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit14 net234 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[142\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_98_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit8 net259 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[264\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit25 net246 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[153\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_98_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_W6END_inbuf_0__0_ net157 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/W6BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_EE4END_inbuf_3__0_ net226 VGND VGND VPWR VPWR ANTENNA_100/DIODE
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_NN4BEG_outbuf_11__0_ Tile_X0Y1_DSP_bot/NN4BEG_i\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y1_NN4BEG\[11\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1521_ Tile_X0Y1_DSP_bot_Inst_MULADD__1692_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1717_/Q
+ Tile_X0Y1_DSP_bot/ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1522_/A
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1452_ Tile_X0Y1_DSP_bot_Inst_MULADD__1452_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1452_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1452_/Y
+ sky130_fd_sc_hd__nor3b_1
XFILLER_0_93_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1383_ Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1385_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0887_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1180_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1386_/A sky130_fd_sc_hd__o2bb2a_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 net764 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[316\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[317\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_147_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__24_ Tile_X0Y1_DSP_bot/JE2BEG\[2\] VGND
+ VGND VPWR VPWR net589 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[330\] Tile_X0Y1_DSP_bot/ConfigBits\[331\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JS2BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1719_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1719_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1719_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit20 net241 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[276\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit31 net253 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[287\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG1 Tile_X0Y1_N2BEG\[3\]
+ net16 net96 net148 Tile_X0Y0_DSP_top/ConfigBits\[184\] Tile_X0Y0_DSP_top/ConfigBits\[185\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[1\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit19 net59 Tile_X0Y1_FrameStrobe_O\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[73\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame10_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_102_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_SS4END_inbuf_0__0_ net127 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/SS4BEG_i\[0\]
+ sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_W1BEG1 Tile_X0Y1_bot2top\[6\]
+ ANTENNA_177/DIODE Tile_X0Y0_DSP_top/JS2BEG\[0\] Tile_X0Y0_DSP_top/J_l_EF_BEG\[2\]
+ Tile_X0Y0_DSP_top/ConfigBits\[86\] Tile_X0Y0_DSP_top/ConfigBits\[87\] VGND VGND
+ VPWR VPWR net536 sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG2 Tile_X0Y1_NN4BEG\[1\]
+ net10 net90 net142 Tile_X0Y0_DSP_top/ConfigBits\[242\] Tile_X0Y0_DSP_top/ConfigBits\[243\]
+ VGND VGND VPWR VPWR ANTENNA_206/DIODE sky130_fd_sc_hd__mux4_2
XFILLER_0_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_strobe_outbuf_11__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_11__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[11\] sky130_fd_sc_hd__buf_8
XFILLER_0_86_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[366\] Tile_X0Y0_DSP_top/ConfigBits\[367\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__0952_ Tile_X0Y1_DSP_bot_Inst_MULADD__0917_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0915_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0916_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0953_/C
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0883_ Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1673_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0882_/Y VGND VGND VPWR VPWR max_cap764/A sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit0 net229 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[32\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_W6END_inbuf_0__0_ net358 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/W6BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG0 net8
+ net126 net173 Tile_X0Y0_DSP_top/JN2BEG\[2\] Tile_X0Y0_DSP_top/ConfigBits\[382\]
+ Tile_X0Y0_DSP_top/ConfigBits\[383\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_CD_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_128_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1504_ Tile_X0Y1_DSP_bot_Inst_MULADD__1452_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1452_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1506_/A
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_E6BEG_outbuf_7__0_ Tile_X0Y1_DSP_bot/E6BEG_i\[7\] VGND VGND VPWR
+ VPWR net612 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1435_ Tile_X0Y1_DSP_bot_Inst_MULADD__1435_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1435_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1435_/Y sky130_fd_sc_hd__nand2_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1366_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1353_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1357_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1359_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1366_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1297_ Tile_X0Y1_DSP_bot_Inst_MULADD__1294_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1295_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1296_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1297_/Y
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_77_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__07_ Tile_X0Y0_top2bot\[3\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/A7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit13 net233 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[173\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit24 net245 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[184\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_103_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput672 net672 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput661 net661 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[8] sky130_fd_sc_hd__buf_2
Xoutput650 net650 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput683 net683 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput694 net694 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[5] sky130_fd_sc_hd__buf_2
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_S4END_inbuf_9__0_ net105 VGND VGND VPWR VPWR ANTENNA_93/DIODE sky130_fd_sc_hd__clkbuf_4
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput18 Tile_X0Y0_E2MID[5] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_4
Xinput29 Tile_X0Y0_E6END[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG1 net325
+ net187 Tile_X0Y0_S4BEG\[2\] Tile_X0Y1_DSP_bot/JE2BEG\[3\] Tile_X0Y1_DSP_bot/ConfigBits\[402\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[403\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_EF_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit2 net71 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[248\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1220_ Tile_X0Y1_DSP_bot_Inst_MULADD__1218_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1219_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1216_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1207_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1220_/X sky130_fd_sc_hd__o211a_2
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1151_ Tile_X0Y1_DSP_bot_Inst_MULADD__1148_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1150_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1142_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1151_/Y
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_157_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1082_ Tile_X0Y1_DSP_bot_Inst_MULADD__1050_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1053_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1081_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1144_/A sky130_fd_sc_hd__o211ai_1
XFILLER_0_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__0935_ Tile_X0Y1_DSP_bot/A3 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0935_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit30 net252 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[318\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0866_ Tile_X0Y1_DSP_bot/ConfigBits\[1\] Tile_X0Y1_DSP_bot_Inst_MULADD__1735_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0866_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_139_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1418_ Tile_X0Y1_DSP_bot_Inst_MULADD__1395_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1397_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1424_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/C
+ sky130_fd_sc_hd__o21a_2
XFILLER_0_64_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit0 net229 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[384\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1349_ Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1349_/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput480 net480 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[8] sky130_fd_sc_hd__clkbuf_4
Xoutput491 net491 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_S4END_inbuf_9__0_ Tile_X0Y0_S4BEG\[13\] VGND VGND VPWR VPWR ANTENNA_110/DIODE
+ sky130_fd_sc_hd__clkbuf_4
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG0 Tile_X0Y1_N2BEGb\[6\]
+ net11 net126 net143 Tile_X0Y0_DSP_top/ConfigBits\[214\] Tile_X0Y0_DSP_top/ConfigBits\[215\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_AB_BEG\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_107_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[330\] Tile_X0Y0_DSP_top/ConfigBits\[331\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_122_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit12 net232 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[204\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_E6BEG_outbuf_3__0_ Tile_X0Y0_DSP_top/E6BEG_i\[3\] VGND VGND VPWR
+ VPWR net407 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit23 net244 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[215\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1203_ Tile_X0Y1_DSP_bot_Inst_MULADD__1097_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1203_/Y
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1134_ Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1104_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1145_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_EE4BEG_outbuf_5__0_ Tile_X0Y1_DSP_bot/EE4BEG_i\[5\] VGND VGND VPWR
+ VPWR net626 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1065_ Tile_X0Y1_DSP_bot_Inst_MULADD__1050_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1064_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0990_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1081_/A
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_90_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0918_ Tile_X0Y1_DSP_bot/ConfigBits\[5\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput208 Tile_X0Y1_E6END[5] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0849_ Tile_X0Y1_DSP_bot_Inst_MULADD__1726_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0849_/X sky130_fd_sc_hd__or2b_2
Xinput219 Tile_X0Y1_EE4END[15] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG0 net300
+ net200 Tile_X0Y0_S2BEG\[7\] net353 Tile_X0Y1_DSP_bot/ConfigBits\[200\] Tile_X0Y1_DSP_bot/ConfigBits\[201\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[0\] sky130_fd_sc_hd__mux4_1
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_B2 Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[2\] Tile_X0Y1_DSP_bot/J2END_CD_BEG\[2\] Tile_X0Y1_DSP_bot/J_l_CD_BEG\[2\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[130\] Tile_X0Y1_DSP_bot/ConfigBits\[131\] VGND VGND
+ VPWR VPWR ANTENNA_97/DIODE sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_A1 Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[1\]
+ ANTENNA_101/DIODE Tile_X0Y1_DSP_bot/J2END_AB_BEG\[1\] Tile_X0Y1_DSP_bot/J_l_AB_BEG\[1\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[120\] Tile_X0Y1_DSP_bot/ConfigBits\[121\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/A1 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_C3 Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[3\]
+ Tile_X0Y1_DSP_bot/J2MID_EFb_BEG\[3\] Tile_X0Y1_DSP_bot/J2END_EF_BEG\[3\] Tile_X0Y1_DSP_bot/J_l_EF_BEG\[3\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[140\] Tile_X0Y1_DSP_bot/ConfigBits\[141\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C3 sky130_fd_sc_hd__mux4_2
XFILLER_0_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[256\] Tile_X0Y0_DSP_top/ConfigBits\[257\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JN2BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0
+ net286 net308 net184 net186 Tile_X0Y1_DSP_bot/ConfigBits\[256\] Tile_X0Y1_DSP_bot/ConfigBits\[257\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__55_ net144 VGND VGND VPWR VPWR net546
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_data_inbuf_20__0_ net61 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_20__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit6 net257 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[166\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit5 net76 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[347\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_159_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit27 net248 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[123\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit16 net236 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[112\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1752_ net333 Tile_X0Y1_DSP_bot/C10 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1683_ Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1683_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1712_/D sky130_fd_sc_hd__nor2_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_data_inbuf_11__0_ net51 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_11__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst0
+ net284 net184 Tile_X0Y0_S1BEG\[3\] Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[45\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[46\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_152_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1117_ Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1117_/Y
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1048_ Tile_X0Y1_DSP_bot_Inst_MULADD__1026_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1047_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1043_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1048_/Y
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[294\] Tile_X0Y0_DSP_top/ConfigBits\[295\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit11 net231 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[235\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit22 net243 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[246\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__38_ Tile_X0Y0_DSP_top/JS2BEG\[6\] VGND
+ VGND VPWR VPWR Tile_X0Y0_S2BEG\[6\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_data_inbuf_20__0_ net241 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_20__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__40_ Tile_X0Y1_DSP_bot/JN2BEG\[2\] VGND
+ VGND VPWR VPWR Tile_X0Y1_N2BEG\[2\] sky130_fd_sc_hd__buf_2
XFILLER_0_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_inbuf_2__0_ net71 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_2__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[278\] Tile_X0Y1_DSP_bot/ConfigBits\[279\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JN2BEG\[5\] sky130_fd_sc_hd__mux4_2
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1735_ net333 Tile_X0Y1_DSP_bot/B1 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1735_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1666_ Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1665_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1666_/Y
+ sky130_fd_sc_hd__o21bai_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1597_ Tile_X0Y1_DSP_bot/C14 Tile_X0Y1_DSP_bot_Inst_MULADD__1756_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1597_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_data_inbuf_11__0_ net231 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_11__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_strobe_outbuf_19__0_ Tile_X0Y0_DSP_top_strobe_inbuf_19__0_/X VGND
+ VGND VPWR VPWR net472 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit9 net260 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[265\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit26 net247 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[154\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit15 net235 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[143\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_data_outbuf_9__0_ Tile_X0Y0_DSP_top_data_inbuf_9__0_/X VGND VGND
+ VPWR VPWR net461 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit0 net49 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[150\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1520_ Tile_X0Y1_DSP_bot_Inst_MULADD__1520_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1520_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1692_/B sky130_fd_sc_hd__or2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1451_ Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1452_/B
+ sky130_fd_sc_hd__a21oi_1
Xinput380 Tile_X0Y1_WW4END[8] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1382_ Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1284_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1382_/Y
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_89_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[316\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[317\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__23_ Tile_X0Y1_DSP_bot/JE2BEG\[1\] VGND
+ VGND VPWR VPWR net588 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_SS4END_inbuf_11__0_ Tile_X0Y0_SS4BEG\[15\] VGND VGND VPWR VPWR
+ ANTENNA_111/DIODE sky130_fd_sc_hd__clkbuf_2
XFILLER_0_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1718_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1718_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1649_ Tile_X0Y1_DSP_bot_Inst_MULADD__1648_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1724_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1664_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/B
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot_NN4END_inbuf_4__0_ net331 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/NN4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit10 net230 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[266\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit21 net242 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[277\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_83_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_N4BEG_outbuf_7__0_ ANTENNA_77/DIODE VGND VGND VPWR VPWR net515
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG2 Tile_X0Y1_N2BEG\[5\]
+ net18 net98 net150 Tile_X0Y0_DSP_top/ConfigBits\[186\] Tile_X0Y0_DSP_top/ConfigBits\[187\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[2\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_W1BEG2 Tile_X0Y1_bot2top\[7\]
+ Tile_X0Y0_DSP_top/J2MID_GHb_BEG\[1\] ANTENNA_63/DIODE Tile_X0Y0_DSP_top/J_l_GH_BEG\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[88\] Tile_X0Y0_DSP_top/ConfigBits\[89\] VGND VGND
+ VPWR VPWR net537 sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG3 Tile_X0Y1_N2BEGb\[1\]
+ net42 net86 net138 Tile_X0Y0_DSP_top/ConfigBits\[244\] Tile_X0Y0_DSP_top/ConfigBits\[245\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_GH_BEG\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_86_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_data_outbuf_9__0_ Tile_X0Y1_DSP_bot_data_inbuf_9__0_/X VGND VGND
+ VPWR VPWR net662 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[366\] Tile_X0Y0_DSP_top/ConfigBits\[367\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0951_ Tile_X0Y1_DSP_bot_Inst_MULADD__0950_/C Tile_X0Y1_DSP_bot_Inst_MULADD__0950_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0950_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0953_/B
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0882_ Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1707_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0882_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit1 net240 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[33\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_120_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1503_ Tile_X0Y1_DSP_bot_Inst_MULADD__1505_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1505_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1502_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1503_/Y
+ sky130_fd_sc_hd__a21boi_2
XFILLER_0_128_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG1 Tile_X0Y1_N4BEG\[2\]
+ net7 net144 Tile_X0Y0_DSP_top/JE2BEG\[2\] Tile_X0Y0_DSP_top/ConfigBits\[384\] Tile_X0Y0_DSP_top/ConfigBits\[385\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_CD_BEG\[1\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1434_ Tile_X0Y1_DSP_bot_Inst_MULADD__1089_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1091_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1432_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1435_/B sky130_fd_sc_hd__o2111ai_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1365_ Tile_X0Y1_DSP_bot_Inst_MULADD__1293_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1273_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1365_/Y sky130_fd_sc_hd__a221oi_4
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1296_ Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1218_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1219_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1296_/Y
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_77_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__06_ Tile_X0Y0_top2bot\[2\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/A6 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_85_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit14 net234 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[174\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit25 net246 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[185\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_103_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput662 net662 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[9] sky130_fd_sc_hd__clkbuf_4
Xoutput640 net640 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput651 net651 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput673 net673 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput684 net684 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput695 net695 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[6] sky130_fd_sc_hd__clkbuf_4
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_W6BEG_outbuf_7__0_ Tile_X0Y0_DSP_top/W6BEG_i\[7\] VGND VGND VPWR
+ VPWR net564 sky130_fd_sc_hd__clkbuf_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 Tile_X0Y0_E2MID[6] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_0_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG2 net308
+ Tile_X0Y0_SS4BEG\[1\] net342 Tile_X0Y1_DSP_bot/JS2BEG\[3\] Tile_X0Y1_DSP_bot/ConfigBits\[404\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[405\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_EF_BEG\[2\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit3 net74 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[249\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1150_ Tile_X0Y1_DSP_bot_Inst_MULADD__1149_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1132_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1140_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1150_/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1081_ Tile_X0Y1_DSP_bot_Inst_MULADD__1081_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1081_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0934_ Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1032_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0933_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0875_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0934_/Y sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_100_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit31 net253 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[319\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit20 net241 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[308\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0865_ Tile_X0Y1_DSP_bot/B1 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0865_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_64_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1417_ Tile_X0Y1_DSP_bot_Inst_MULADD__1417_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q9 sky130_fd_sc_hd__buf_8
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1348_ Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1323_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1335_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1263_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1348_/Y sky130_fd_sc_hd__a32oi_4
XTile_X0Y0_DSP_top_NN4END_inbuf_0__0_ Tile_X0Y1_NN4BEG\[4\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/NN4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit1 net240 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[385\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1279_ Tile_X0Y1_DSP_bot_Inst_MULADD__0926_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0958_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1089_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1091_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1371_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_0_148_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG0 net299
+ Tile_X0Y0_S2BEG\[6\] net352 Tile_X0Y1_DSP_bot/JN2BEG\[3\] Tile_X0Y1_DSP_bot/ConfigBits\[160\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[161\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput470 net470 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[17] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_E6END_inbuf_5__0_ net30 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/E6BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
Xoutput492 net492 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput481 net481 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_strobe_inbuf_13__0_ Tile_X0Y1_FrameStrobe_O\[13\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_13__0_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG1 Tile_X0Y1_NN4BEG\[0\]
+ net7 net87 net139 Tile_X0Y0_DSP_top/ConfigBits\[216\] Tile_X0Y0_DSP_top/ConfigBits\[217\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_AB_BEG\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_52_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[330\] Tile_X0Y0_DSP_top/ConfigBits\[331\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_outbuf_27__0_ Tile_X0Y0_DSP_top_data_inbuf_27__0_/X VGND VGND
+ VPWR VPWR net449 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit13 net233 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[205\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit24 net245 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[216\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1202_ Tile_X0Y1_DSP_bot_Inst_MULADD__1034_/X Tile_X0Y1_DSP_bot/B5
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1035_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1201_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1202_/X sky130_fd_sc_hd__o2111a_1
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1133_ Tile_X0Y1_DSP_bot_Inst_MULADD__1114_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1120_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1155_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1132_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1133_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_0_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1064_ Tile_X0Y1_DSP_bot_Inst_MULADD__1063_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1048_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1049_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1064_/Y
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0917_ Tile_X0Y1_DSP_bot_Inst_MULADD__0917_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0917_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1675_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__0848_ Tile_X0Y1_DSP_bot/ConfigBits\[0\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/A sky130_fd_sc_hd__buf_2
Xinput209 Tile_X0Y1_E6END[6] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_data_outbuf_18__0_ Tile_X0Y0_DSP_top_data_inbuf_18__0_/X VGND VGND
+ VPWR VPWR net439 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_S4BEG_outbuf_7__0_ ANTENNA_92/DIODE VGND VGND VPWR VPWR Tile_X0Y0_S4BEG\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG1 net296
+ net196 Tile_X0Y0_S2BEG\[3\] net349 Tile_X0Y1_DSP_bot/ConfigBits\[202\] Tile_X0Y1_DSP_bot/ConfigBits\[203\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[1\] sky130_fd_sc_hd__mux4_2
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_B3 Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[3\]
+ Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[3\] Tile_X0Y1_DSP_bot/J2END_CD_BEG\[3\] Tile_X0Y1_DSP_bot/J_l_CD_BEG\[3\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[132\] Tile_X0Y1_DSP_bot/ConfigBits\[133\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/B3 sky130_fd_sc_hd__mux4_2
XFILLER_0_19_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_A2 Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2MID_ABb_BEG\[2\] Tile_X0Y1_DSP_bot/J2END_AB_BEG\[2\] Tile_X0Y1_DSP_bot/J_l_AB_BEG\[2\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[122\] Tile_X0Y1_DSP_bot/ConfigBits\[123\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/A2 sky130_fd_sc_hd__mux4_2
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_C4 Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[0\]
+ Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[0\] Tile_X0Y1_DSP_bot/J2END_GH_BEG\[0\] Tile_X0Y1_DSP_bot/J_l_GH_BEG\[0\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[142\] Tile_X0Y1_DSP_bot/ConfigBits\[143\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C4 sky130_fd_sc_hd__mux4_1
XFILLER_0_151_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1
+ net204 Tile_X0Y0_SS4BEG\[1\] net339 net357 Tile_X0Y1_DSP_bot/ConfigBits\[256\] Tile_X0Y1_DSP_bot/ConfigBits\[257\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__54_ Tile_X0Y0_DSP_top/JW2BEG\[6\] VGND
+ VGND VPWR VPWR net545 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit7 net258 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[167\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_E6END_inbuf_5__0_ net210 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/E6BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit6 net77 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[348\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_159_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit30 net252 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[350\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit17 net237 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[113\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_154_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit28 net249 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[124\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1751_ net333 Tile_X0Y1_DSP_bot/C9 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1751_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1682_ Tile_X0Y1_DSP_bot_Inst_MULADD__1682_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1711_/D sky130_fd_sc_hd__clkbuf_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[44\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__o21ai_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[2\] Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2END_EF_BEG\[0\] Tile_X0Y1_DSP_bot/ConfigBits\[45\] Tile_X0Y1_DSP_bot/ConfigBits\[46\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_N1BEG0 Tile_X0Y1_DSP_bot/Q2
+ Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[3\] Tile_X0Y1_DSP_bot/JW2BEG\[3\] Tile_X0Y1_DSP_bot/J_l_CD_BEG\[1\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[6\] Tile_X0Y1_DSP_bot/ConfigBits\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N1BEG\[0\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_EE4END_inbuf_11__0_ net219 VGND VGND VPWR VPWR ANTENNA_99/DIODE
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1116_ Tile_X0Y1_DSP_bot_Inst_MULADD__1100_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1214_/D
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1054_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1103_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1116_/Y sky130_fd_sc_hd__a221oi_4
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1047_ Tile_X0Y1_DSP_bot_Inst_MULADD__1045_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1046_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1047_/Y
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_160_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst0
+ net282 net182 net335 Tile_X0Y1_DSP_bot/Q5 Tile_X0Y1_DSP_bot/ConfigBits\[31\] Tile_X0Y1_DSP_bot/ConfigBits\[32\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[296\] Tile_X0Y0_DSP_top/ConfigBits\[297\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JE2BEG\[4\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0
+ net282 net288 net310 net188 Tile_X0Y1_DSP_bot/ConfigBits\[296\] Tile_X0Y1_DSP_bot/ConfigBits\[297\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0
+ net183 net336 Tile_X0Y1_DSP_bot/Q0 net764 Tile_X0Y1_DSP_bot/ConfigBits\[58\] Tile_X0Y1_DSP_bot/ConfigBits\[59\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst3_765
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst3_765/HI
+ net765 sky130_fd_sc_hd__conb_1
XTile_X0Y1_DSP_bot_data_inbuf_8__0_ net259 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_8__0_/X
+ sky130_fd_sc_hd__buf_1
XFILLER_0_124_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit12 net232 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[236\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit23 net244 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[247\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__37_ ANTENNA_64/DIODE VGND VGND VPWR
+ VPWR Tile_X0Y0_S2BEG\[5\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_strobe_outbuf_4__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_4__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[4\] sky130_fd_sc_hd__buf_8
XFILLER_0_159_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_WW4BEG_outbuf_9__0_ Tile_X0Y0_DSP_top/WW4BEG_i\[9\] VGND VGND VPWR
+ VPWR net582 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1734_ net333 Tile_X0Y1_DSP_bot/B0 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1734_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1665_ Tile_X0Y1_DSP_bot_Inst_MULADD__1665_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1665_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1665_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1596_ Tile_X0Y1_DSP_bot_Inst_MULADD__1593_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1589_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1594_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1595_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/B sky130_fd_sc_hd__o211ai_4
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[0\] Tile_X0Y1_N2BEGb\[2\] net7 net21 Tile_X0Y0_DSP_top/ConfigBits\[346\]
+ Tile_X0Y0_DSP_top/ConfigBits\[347\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_WW4BEG_outbuf_2__0_ Tile_X0Y1_DSP_bot/WW4BEG_i\[2\] VGND VGND VPWR
+ VPWR net755 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit27 net248 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[155\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit16 net236 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[144\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_strobe_inbuf_19__0_ net271 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_19__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit1 net60 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[151\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1450_ Tile_X0Y1_DSP_bot_Inst_MULADD__1402_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1448_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1449_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1450_/Y
+ sky130_fd_sc_hd__o21ai_4
Xinput381 Tile_X0Y1_WW4END[9] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkbuf_1
Xinput370 Tile_X0Y1_WW4END[13] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1381_ Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[318\] Tile_X0Y1_DSP_bot/ConfigBits\[319\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JE2BEG\[7\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_N4END_inbuf_9__0_ Tile_X0Y1_N4BEG\[13\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/N4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__22_ Tile_X0Y1_DSP_bot/JE2BEG\[0\] VGND
+ VGND VPWR VPWR net587 sky130_fd_sc_hd__buf_1
XFILLER_0_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1717_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1717_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[50\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__o21ai_1
XFILLER_0_158_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1648_ Tile_X0Y1_DSP_bot/C18 Tile_X0Y1_DSP_bot_Inst_MULADD__1760_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1648_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1579_ Tile_X0Y1_DSP_bot_Inst_MULADD__1629_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1579_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1581_/A sky130_fd_sc_hd__and2_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit11 net231 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[267\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit22 net243 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[278\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG3 Tile_X0Y1_N2BEG\[1\]
+ net14 net94 net146 Tile_X0Y0_DSP_top/ConfigBits\[188\] Tile_X0Y0_DSP_top/ConfigBits\[189\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_W1BEG3 Tile_X0Y1_bot2top\[0\]
+ Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[2\] Tile_X0Y0_DSP_top/JS2BEG\[2\] ANTENNA_65/DIODE
+ Tile_X0Y0_DSP_top/ConfigBits\[90\] Tile_X0Y0_DSP_top/ConfigBits\[91\] VGND VGND
+ VPWR VPWR net538 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_WW4END_inbuf_5__0_ net381 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/WW4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[368\] Tile_X0Y0_DSP_top/ConfigBits\[369\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JW2BEG\[6\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[3\] net84 net136 Tile_X0Y1_bot2top\[3\] Tile_X0Y0_DSP_top/ConfigBits\[95\]
+ Tile_X0Y0_DSP_top/ConfigBits\[96\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0950_ Tile_X0Y1_DSP_bot_Inst_MULADD__0950_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0950_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0950_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0953_/A
+ sky130_fd_sc_hd__or3_1
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0881_ Tile_X0Y1_DSP_bot_Inst_MULADD__1672_/B Tile_X0Y1_DSP_bot_Inst_MULADD__0881_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1673_/B sky130_fd_sc_hd__xnor2_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit2 net251 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[34\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0
+ net282 net290 net182 net190 Tile_X0Y1_DSP_bot/ConfigBits\[368\] Tile_X0Y1_DSP_bot/ConfigBits\[369\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1502_ Tile_X0Y1_DSP_bot_Inst_MULADD__0933_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1501_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1502_/X
+ sky130_fd_sc_hd__o21a_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG2 Tile_X0Y1_NN4BEG\[1\]
+ net40 net108 Tile_X0Y0_DSP_top/JS2BEG\[2\] Tile_X0Y0_DSP_top/ConfigBits\[386\] Tile_X0Y0_DSP_top/ConfigBits\[387\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_CD_BEG\[2\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1433_ Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1432_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1435_/A sky130_fd_sc_hd__a22o_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1364_ Tile_X0Y1_DSP_bot_Inst_MULADD__1369_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1369_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1364_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/B
+ sky130_fd_sc_hd__nand3_4
XFILLER_0_77_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1295_ Tile_X0Y1_DSP_bot_Inst_MULADD__1285_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1285_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1283_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1295_/X sky130_fd_sc_hd__o2111a_1
XFILLER_0_77_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_N4END_inbuf_9__0_ net305 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/N4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__05_ Tile_X0Y0_top2bot\[1\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/A5 sky130_fd_sc_hd__buf_2
XFILLER_0_73_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit15 net235 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[175\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit26 net247 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[186\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_SS4BEG_outbuf_2__0_ Tile_X0Y0_DSP_top/SS4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_SS4BEG\[2\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0
+ Tile_X0Y1_NN4BEG\[1\] net4 net6 net24 Tile_X0Y0_DSP_top/ConfigBits\[310\] Tile_X0Y0_DSP_top/ConfigBits\[311\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
Xoutput663 net663 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput630 net630 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput641 net641 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput652 net652 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[29] sky130_fd_sc_hd__clkbuf_4
Xoutput674 net674 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput685 net685 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput696 net696 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[7] sky130_fd_sc_hd__clkbuf_4
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG3 net222
+ Tile_X0Y0_S4BEG\[0\] net373 Tile_X0Y1_DSP_bot/JW2BEG\[3\] Tile_X0Y1_DSP_bot/ConfigBits\[406\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[407\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J_l_EF_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[27\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__o21ai_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit4 net75 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[250\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1080_ Tile_X0Y1_DSP_bot_Inst_MULADD__1078_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1079_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1011_/X Tile_X0Y1_DSP_bot_Inst_MULADD__0995_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0996_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1080_/X sky130_fd_sc_hd__a2111o_1
XFILLER_0_157_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0933_ Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/A Tile_X0Y1_DSP_bot/A3
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1373_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0933_/Y
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit10 net230 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[298\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit21 net242 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[309\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0864_ Tile_X0Y1_DSP_bot_Inst_MULADD__1124_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/A sky130_fd_sc_hd__buf_4
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1416_ Tile_X0Y1_DSP_bot_Inst_MULADD__1688_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1715_/Q
+ Tile_X0Y1_DSP_bot/ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1417_/A
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1347_ Tile_X0Y1_DSP_bot_Inst_MULADD__1345_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1334_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/A
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1278_ Tile_X0Y1_DSP_bot_Inst_MULADD__1030_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1097_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1371_/A sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit2 net251 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[386\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG1 net195
+ Tile_X0Y0_S2BEG\[2\] net348 Tile_X0Y1_DSP_bot/JE2BEG\[3\] Tile_X0Y1_DSP_bot/ConfigBits\[162\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[163\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[1\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput471 net471 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput460 net460 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[8] sky130_fd_sc_hd__buf_2
Xoutput482 net482 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput493 net493 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG2 Tile_X0Y1_N2BEGb\[4\]
+ net33 net89 net141 Tile_X0Y0_DSP_top/ConfigBits\[218\] Tile_X0Y0_DSP_top/ConfigBits\[219\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_AB_BEG\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_WW4END_inbuf_1__0_ net176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/WW4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[332\] Tile_X0Y0_DSP_top/ConfigBits\[333\] VGND VGND
+ VPWR VPWR ANTENNA_64/DIODE sky130_fd_sc_hd__mux4_2
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0
+ net289 net183 net189 net201 Tile_X0Y1_DSP_bot/ConfigBits\[332\] Tile_X0Y1_DSP_bot/ConfigBits\[333\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_strobe_inbuf_8__0_ Tile_X0Y1_FrameStrobe_O\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_8__0_/X sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit14 net234 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[206\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit25 net246 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[217\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1201_ Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1201_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1201_/Y sky130_fd_sc_hd__nand4_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1132_ Tile_X0Y1_DSP_bot_Inst_MULADD__1114_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1130_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1131_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1132_/Y
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1063_ Tile_X0Y1_DSP_bot_Inst_MULADD__1054_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1055_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1062_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1063_/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_145_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0916_ Tile_X0Y1_DSP_bot_Inst_MULADD__0916_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0915_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0917_/B sky130_fd_sc_hd__or2b_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0847_ Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1481_/A sky130_fd_sc_hd__buf_4
XFILLER_0_78_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG2 net298
+ net198 Tile_X0Y0_S2BEG\[5\] net351 Tile_X0Y1_DSP_bot/ConfigBits\[204\] Tile_X0Y1_DSP_bot/ConfigBits\[205\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[2\] sky130_fd_sc_hd__mux4_1
XFILLER_0_148_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_A3 Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[3\]
+ Tile_X0Y1_DSP_bot/J2MID_ABb_BEG\[3\] Tile_X0Y1_DSP_bot/J2END_AB_BEG\[3\] Tile_X0Y1_DSP_bot/J_l_AB_BEG\[3\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[124\] Tile_X0Y1_DSP_bot/ConfigBits\[125\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/A3 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_C5 Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[1\]
+ Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[1\] Tile_X0Y1_DSP_bot/J2END_GH_BEG\[1\] Tile_X0Y1_DSP_bot/J_l_GH_BEG\[1\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[144\] Tile_X0Y1_DSP_bot/ConfigBits\[145\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C5 sky130_fd_sc_hd__mux4_1
XFILLER_0_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__53_ Tile_X0Y0_DSP_top/JW2BEG\[5\] VGND
+ VGND VPWR VPWR net544 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2
+ net764 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[256\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[257\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit8 net259 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[168\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit7 net78 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[349\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_159_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit20 net241 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[340\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_84_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit31 net253 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[351\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit18 net238 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[114\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[33\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_NN4BEG\[15\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit29 net250 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[125\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_NN4BEG_outbuf_5__0_ Tile_X0Y1_DSP_bot/NN4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y1_NN4BEG\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1750_ net333 Tile_X0Y1_DSP_bot/C8 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_SS4END_inbuf_7__0_ Tile_X0Y0_SS4BEG\[11\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/SS4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1681_ Tile_X0Y1_DSP_bot_Inst_MULADD__1674_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1681_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1682_/A sky130_fd_sc_hd__and2b_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[44\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_N1BEG1 Tile_X0Y1_DSP_bot/Q3
+ Tile_X0Y1_DSP_bot/J2MID_EFb_BEG\[0\] Tile_X0Y1_DSP_bot/JW2BEG\[0\] Tile_X0Y1_DSP_bot/J_l_EF_BEG\[2\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[8\] Tile_X0Y1_DSP_bot/ConfigBits\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N1BEG\[1\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1115_ Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_SS4BEG_outbuf_8__0_ Tile_X0Y1_DSP_bot/SS4BEG_i\[8\] VGND VGND VPWR
+ VPWR net713 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1046_ Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1054_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1046_/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[2\] Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2END_AB_BEG\[1\] Tile_X0Y1_DSP_bot/ConfigBits\[31\] Tile_X0Y1_DSP_bot/ConfigBits\[32\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1
+ net204 Tile_X0Y0_S2BEGb\[3\] net341 net357 Tile_X0Y1_DSP_bot/ConfigBits\[296\] Tile_X0Y1_DSP_bot/ConfigBits\[297\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/Q5
+ Tile_X0Y1_DSP_bot/ConfigBits\[58\] Tile_X0Y1_DSP_bot/ConfigBits\[59\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_109_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst3_766
+ VGND VGND VPWR VPWR net766 Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_clr_cus_mux41_buf_inst3_766/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit13 net233 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[237\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit24 net245 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[248\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__36_ Tile_X0Y0_DSP_top/JS2BEG\[4\] VGND
+ VGND VPWR VPWR Tile_X0Y0_S2BEG\[4\] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[1\] net2 net82 Tile_X0Y1_bot2top\[5\] Tile_X0Y0_DSP_top/ConfigBits\[45\]
+ Tile_X0Y0_DSP_top/ConfigBits\[46\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_W6END_inbuf_3__0_ net160 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/W6BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_EE4END_inbuf_6__0_ net214 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/EE4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1733_ net333 Tile_X0Y1_DSP_bot/A7 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1733_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1664_ Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1725_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1664_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1665_/B
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1595_ Tile_X0Y1_DSP_bot_Inst_MULADD__1595_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1595_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1595_/Y sky130_fd_sc_hd__nor2_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_EE4BEG_outbuf_2__0_ ANTENNA_59/DIODE VGND VGND VPWR VPWR net422
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1
+ net87 net109 net139 net153 Tile_X0Y0_DSP_top/ConfigBits\[346\] Tile_X0Y0_DSP_top/ConfigBits\[347\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1029_ Tile_X0Y1_DSP_bot/B4 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1029_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_44_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit30 net252 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[382\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit28 net249 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[156\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit17 net237 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[145\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__19_ Tile_X0Y0_DSP_top/JN2BEG\[3\] VGND
+ VGND VPWR VPWR net489 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit2 net71 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[152\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_SS4END_inbuf_3__0_ net130 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/SS4BEG_i\[3\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_117_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1380_ Tile_X0Y1_DSP_bot_Inst_MULADD__1366_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1370_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1379_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1365_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1444_/A sky130_fd_sc_hd__o22ai_4
Xinput371 Tile_X0Y1_WW4END[14] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_1
Xinput360 Tile_X0Y1_W6END[4] VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_strobe_outbuf_14__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_14__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[14\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__21_ Tile_X0Y0_top2bot\[17\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_W6END_inbuf_3__0_ net361 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/W6BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_158_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[50\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1716_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1716_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1716_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0
+ Tile_X0Y1_N2BEGb\[4\] Tile_X0Y1_N4BEG\[0\] net3 net9 Tile_X0Y0_DSP_top/ConfigBits\[258\]
+ Tile_X0Y0_DSP_top/ConfigBits\[259\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1647_ Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1723_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1646_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q17
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1578_ Tile_X0Y1_DSP_bot_Inst_MULADD__1578_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1578_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1578_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1579_/B
+ sky130_fd_sc_hd__nand3_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit0 net229 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[288\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit12 net232 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[268\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit23 net244 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[279\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst0
+ net282 net182 net335 Tile_X0Y1_DSP_bot/Q5 Tile_X0Y1_DSP_bot/ConfigBits\[87\] Tile_X0Y1_DSP_bot/ConfigBits\[88\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[7\] Tile_X0Y0_DSP_top/J2MID_ABa_BEG\[2\] Tile_X0Y0_DSP_top/J2MID_CDa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2END_EF_BEG\[2\] Tile_X0Y0_DSP_top/ConfigBits\[95\] Tile_X0Y0_DSP_top/ConfigBits\[96\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0880_ Tile_X0Y1_DSP_bot_Inst_MULADD__0880_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0880_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0881_/B sky130_fd_sc_hd__nor2_1
XTile_X0Y0_DSP_top_EE4END_inbuf_2__0_ net45 VGND VGND VPWR VPWR ANTENNA_59/DIODE sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit3 net254 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[35\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[1\] Tile_X0Y0_S1BEG\[3\] Tile_X0Y0_S2BEGb\[5\] net335 Tile_X0Y1_DSP_bot/ConfigBits\[368\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[369\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1501_ Tile_X0Y1_DSP_bot_Inst_MULADD__1501_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1501_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG3 Tile_X0Y1_N4BEG\[0\]
+ net117 net153 Tile_X0Y0_DSP_top/JW2BEG\[2\] Tile_X0Y0_DSP_top/ConfigBits\[388\]
+ Tile_X0Y0_DSP_top/ConfigBits\[389\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J_l_CD_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1432_ Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1268_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/C VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1432_/Y sky130_fd_sc_hd__o2bb2ai_1
Xinput190 Tile_X0Y1_E2END[5] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1363_ Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1364_/C
+ sky130_fd_sc_hd__and3_1
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1294_ Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1316_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1293_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1294_/Y
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_58_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__04_ Tile_X0Y0_top2bot\[0\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/A4 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit16 net236 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[176\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit27 net248 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[187\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1
+ net86 net108 net138 net156 Tile_X0Y0_DSP_top/ConfigBits\[310\] Tile_X0Y0_DSP_top/ConfigBits\[311\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput620 net620 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput631 net631 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[0] sky130_fd_sc_hd__buf_2
Xoutput642 net642 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput653 net653 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput664 net664 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput675 net675 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput697 net697 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput686 net686 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_N4BEG_outbuf_1__0_ Tile_X0Y1_DSP_bot/N4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N4BEG\[1\] sky130_fd_sc_hd__clkbuf_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[27\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit5 net76 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[251\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_99_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0
+ net284 net292 net184 net192 Tile_X0Y1_DSP_bot/ConfigBits\[280\] Tile_X0Y1_DSP_bot/ConfigBits\[281\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0932_ Tile_X0Y1_DSP_bot_Inst_MULADD__1729_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1373_/B sky130_fd_sc_hd__or2b_2
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit11 net231 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[299\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit22 net243 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[310\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0863_ Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0889_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0862_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1124_/A
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_139_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_E6BEG_outbuf_6__0_ Tile_X0Y0_DSP_top/E6BEG_i\[6\] VGND VGND VPWR
+ VPWR net410 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1415_ Tile_X0Y1_DSP_bot_Inst_MULADD__1415_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1415_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1688_/B sky130_fd_sc_hd__or2_1
XTile_X0Y1_DSP_bot_EE4BEG_outbuf_8__0_ Tile_X0Y1_DSP_bot/EE4BEG_i\[8\] VGND VGND VPWR
+ VPWR net629 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1346_ Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/Y
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_148_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1277_ Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/A Tile_X0Y1_DSP_bot/B4
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/X sky130_fd_sc_hd__or2b_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit3 net254 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[387\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_93_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_W6BEG_outbuf_1__0_ Tile_X0Y1_DSP_bot/W6BEG_i\[1\] VGND VGND VPWR
+ VPWR net738 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG2 net297
+ net197 net350 Tile_X0Y1_DSP_bot/JS2BEG\[3\] Tile_X0Y1_DSP_bot/ConfigBits\[164\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[165\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[2\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_46_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput450 net450 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[28] sky130_fd_sc_hd__clkbuf_4
Xoutput461 net461 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[9] sky130_fd_sc_hd__buf_2
Xoutput494 net494 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput472 net472 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput483 net483 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG3 Tile_X0Y1_N2BEGb\[0\]
+ net5 net85 net174 Tile_X0Y0_DSP_top/ConfigBits\[220\] Tile_X0Y0_DSP_top/ConfigBits\[221\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2END_AB_BEG\[3\] sky130_fd_sc_hd__mux4_2
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_data_inbuf_23__0_ net64 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_23__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1
+ Tile_X0Y0_S2BEGb\[4\] Tile_X0Y0_S4BEG\[0\] net342 net374 Tile_X0Y1_DSP_bot/ConfigBits\[332\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[333\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit15 net235 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[207\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit26 net247 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[218\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1200_ Tile_X0Y1_DSP_bot_Inst_MULADD__1196_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1197_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1289_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1289_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/B sky130_fd_sc_hd__o211ai_4
XFILLER_0_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1131_ Tile_X0Y1_DSP_bot_Inst_MULADD__1054_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1055_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1043_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1047_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1131_/X sky130_fd_sc_hd__o22a_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1062_ Tile_X0Y1_DSP_bot_Inst_MULADD__1060_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1061_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1043_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1062_/Y
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_28_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0915_ Tile_X0Y1_DSP_bot_Inst_MULADD__0915_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0915_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0915_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0846_ Tile_X0Y1_DSP_bot/ConfigBits\[0\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/A sky130_fd_sc_hd__clkbuf_8
XTile_X0Y0_DSP_top_data_inbuf_14__0_ net54 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_14__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1329_ Tile_X0Y1_DSP_bot/C8 Tile_X0Y1_DSP_bot_Inst_MULADD__1750_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1329_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG3 net294
+ net194 Tile_X0Y0_S2BEG\[1\] net347 Tile_X0Y1_DSP_bot/ConfigBits\[206\] Tile_X0Y1_DSP_bot/ConfigBits\[207\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_38_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_data_outbuf_30__0_ Tile_X0Y1_DSP_bot_data_inbuf_30__0_/X VGND VGND
+ VPWR VPWR net654 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_C6 Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[2\] Tile_X0Y1_DSP_bot/J2END_GH_BEG\[2\] Tile_X0Y1_DSP_bot/J_l_GH_BEG\[2\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[146\] Tile_X0Y1_DSP_bot/ConfigBits\[147\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C6 sky130_fd_sc_hd__mux4_1
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__52_ net141 VGND VGND VPWR VPWR net543
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/ConfigBits\[256\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[257\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit9 net260 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[169\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit8 net79 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[350\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_159_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit10 net230 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[330\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_data_outbuf_21__0_ Tile_X0Y1_DSP_bot_data_inbuf_21__0_/X VGND VGND
+ VPWR VPWR net644 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit21 net242 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[341\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_127_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[33\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit19 net239 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[115\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1680_ Tile_X0Y1_DSP_bot_Inst_MULADD__1680_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1710_/D sky130_fd_sc_hd__clkbuf_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG0 net326
+ net191 Tile_X0Y0_S2BEGb\[6\] net344 Tile_X0Y1_DSP_bot/ConfigBits\[232\] Tile_X0Y1_DSP_bot/ConfigBits\[233\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_CD_BEG\[0\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_data_inbuf_23__0_ net244 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_23__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_data_outbuf_12__0_ Tile_X0Y1_DSP_bot_data_inbuf_12__0_/X VGND VGND
+ VPWR VPWR net634 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_N1BEG2 Tile_X0Y1_DSP_bot/Q4
+ Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[1\] Tile_X0Y1_DSP_bot/JW2BEG\[1\] Tile_X0Y1_DSP_bot/J_l_GH_BEG\[3\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[10\] Tile_X0Y1_DSP_bot/ConfigBits\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y1_N1BEG\[2\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1114_ Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1104_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1109_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1114_/X sky130_fd_sc_hd__o2111a_2
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1045_ Tile_X0Y1_DSP_bot_Inst_MULADD__1045_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1045_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_145_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_S4BEG_outbuf_1__0_ Tile_X0Y1_DSP_bot/S4BEG_i\[1\] VGND VGND VPWR
+ VPWR net690 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_data_inbuf_5__0_ net76 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_5__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_data_inbuf_14__0_ net234 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_14__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 net764 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[296\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[297\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2
+ net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[58\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[59\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit14 net234 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[238\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit25 net246 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[249\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__35_ Tile_X0Y0_DSP_top/JS2BEG\[3\] VGND
+ VGND VPWR VPWR Tile_X0Y0_S2BEG\[3\] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[9\] Tile_X0Y0_DSP_top/J2MID_EFa_BEG\[2\] Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[2\]
+ Tile_X0Y0_DSP_top/J2END_AB_BEG\[0\] Tile_X0Y0_DSP_top/ConfigBits\[45\] Tile_X0Y0_DSP_top/ConfigBits\[46\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_NN4END_inbuf_11__0_ net323 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/NN4BEG_i\[11\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1732_ net333 Tile_X0Y1_DSP_bot/A6 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1663_ Tile_X0Y1_DSP_bot/C19 Tile_X0Y1_DSP_bot_Inst_MULADD__1761_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/X
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1594_ Tile_X0Y1_DSP_bot_Inst_MULADD__1594_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1594_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1594_/Y sky130_fd_sc_hd__nand2_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1028_ Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1045_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1025_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1028_/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[346\] Tile_X0Y0_DSP_top/ConfigBits\[347\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit31 net253 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[383\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit20 net241 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[372\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_NN4END_inbuf_7__0_ net319 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/NN4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit29 net250 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[157\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit18 net238 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[146\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__18_ Tile_X0Y0_DSP_top/JN2BEG\[2\] VGND
+ VGND VPWR VPWR net488 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit3 net74 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[153\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_93_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput350 Tile_X0Y1_W2MID[4] VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkbuf_4
Xinput372 Tile_X0Y1_WW4END[15] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkbuf_1
Xinput361 Tile_X0Y1_W6END[5] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__20_ Tile_X0Y0_top2bot\[16\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1715_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1715_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1646_ Tile_X0Y1_DSP_bot_Inst_MULADD__1644_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1645_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1646_/Y
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1
+ net21 net89 net141 net153 Tile_X0Y0_DSP_top/ConfigBits\[258\] Tile_X0Y0_DSP_top/ConfigBits\[259\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1577_ Tile_X0Y1_DSP_bot_Inst_MULADD__1577_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1577_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1578_/C sky130_fd_sc_hd__nor2_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit1 net240 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[289\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[80\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR Tile_X0Y0_SS4BEG\[14\] sky130_fd_sc_hd__o21ai_4
XFILLER_0_95_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit13 net233 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[269\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit24 net245 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[280\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[2\] Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2END_AB_BEG\[3\] Tile_X0Y1_DSP_bot/ConfigBits\[87\] Tile_X0Y1_DSP_bot/ConfigBits\[88\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit4 net255 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[36\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[368\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[369\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1500_ Tile_X0Y1_DSP_bot_Inst_MULADD__1536_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1498_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1499_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1505_/C
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1431_ Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/Y sky130_fd_sc_hd__nand4_4
XTile_X0Y0_DSP_top_strobe_outbuf_1__0_ Tile_X0Y0_DSP_top_strobe_inbuf_1__0_/X VGND
+ VGND VPWR VPWR net473 sky130_fd_sc_hd__clkbuf_1
Xinput180 Tile_X0Y0_WW4END[9] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1362_ Tile_X0Y1_DSP_bot_Inst_MULADD__1019_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1358_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1535_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1354_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1369_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_0_144_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput191 Tile_X0Y1_E2END[6] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1293_ Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1292_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1293_/Y
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_144_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[2\] Tile_X0Y1_N2BEGb\[6\] net3 net11 Tile_X0Y0_DSP_top/ConfigBits\[298\]
+ Tile_X0Y0_DSP_top/ConfigBits\[299\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit30 net252 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[414\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit17 net237 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[177\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_131_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit28 net249 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[188\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[310\] Tile_X0Y0_DSP_top/ConfigBits\[311\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
Xoutput610 net610 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput621 net621 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput632 net632 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[10] sky130_fd_sc_hd__buf_2
Xoutput643 net643 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[20] sky130_fd_sc_hd__clkbuf_4
Xoutput654 net654 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput665 net665 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput676 net676 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput687 net687 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput698 net698 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[9] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1629_ Tile_X0Y1_DSP_bot_Inst_MULADD__1629_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1632_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1629_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1631_/A sky130_fd_sc_hd__nand4_1
XTile_X0Y0_DSP_top_NN4END_inbuf_3__0_ Tile_X0Y1_NN4BEG\[7\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/NN4BEG_i\[3\]
+ sky130_fd_sc_hd__buf_2
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top_E6END_inbuf_8__0_ net22 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/E6BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit6 net77 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[252\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_99_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1
+ Tile_X0Y0_S1BEG\[3\] Tile_X0Y0_S2BEGb\[7\] net335 net337 Tile_X0Y1_DSP_bot/ConfigBits\[280\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[281\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_strobe_inbuf_16__0_ Tile_X0Y1_FrameStrobe_O\[16\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_16__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__0931_ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/B sky130_fd_sc_hd__buf_6
XFILLER_0_70_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0862_ Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1727_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0862_/Y sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit12 net232 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[300\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit23 net244 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[311\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1414_ Tile_X0Y1_DSP_bot_Inst_MULADD__1465_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1415_/B
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1345_ Tile_X0Y1_DSP_bot_Inst_MULADD__1255_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1338_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1339_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1345_/Y
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit4 net255 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[388\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1276_ Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1533_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1275_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/A sky130_fd_sc_hd__a41oi_4
XFILLER_0_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG3 net293
+ net193 Tile_X0Y0_S2BEG\[0\] Tile_X0Y1_DSP_bot/JW2BEG\[3\] Tile_X0Y1_DSP_bot/ConfigBits\[166\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[167\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput462 net462 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput451 net451 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput440 net440 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[19] sky130_fd_sc_hd__buf_2
Xoutput473 net473 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[1] sky130_fd_sc_hd__clkbuf_4
Xoutput484 net484 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput495 net495 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[1] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[86\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__o21ai_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_E6END_inbuf_8__0_ net202 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/E6BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[332\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[333\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit27 net248 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[219\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit16 net236 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[208\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1130_ Tile_X0Y1_DSP_bot_Inst_MULADD__1116_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1117_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1130_/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1061_ Tile_X0Y1_DSP_bot_Inst_MULADD__0875_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0933_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0963_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1061_/X sky130_fd_sc_hd__o41a_1
XFILLER_0_157_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__0914_ Tile_X0Y1_DSP_bot_Inst_MULADD__0915_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0915_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0916_/A sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0845_ Tile_X0Y1_DSP_bot_Inst_MULADD__0844_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1706_/Q
+ Tile_X0Y1_DSP_bot/ConfigBits\[3\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0856_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_N4BEG0 net287 net308
+ net204 Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[14\] Tile_X0Y1_DSP_bot/ConfigBits\[15\]
+ VGND VGND VPWR VPWR Tile_X0Y1_N4BEG\[12\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1328_ Tile_X0Y1_DSP_bot_Inst_MULADD__1459_/S VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/S sky130_fd_sc_hd__buf_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_MULADD__1259_ Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1566_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1259_/X
+ sky130_fd_sc_hd__or3_2
XFILLER_0_148_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_C7 Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[3\]
+ Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[3\] Tile_X0Y1_DSP_bot/J2END_GH_BEG\[3\] Tile_X0Y1_DSP_bot/J_l_GH_BEG\[3\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[148\] Tile_X0Y1_DSP_bot/ConfigBits\[149\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/C7 sky130_fd_sc_hd__mux4_2
XFILLER_0_151_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__51_ net140 VGND VGND VPWR VPWR net542
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[258\] Tile_X0Y1_DSP_bot/ConfigBits\[259\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JN2BEG\[0\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[0\] Tile_X0Y1_N2BEGb\[0\] net1 net5 Tile_X0Y0_DSP_top/ConfigBits\[370\]
+ Tile_X0Y0_DSP_top/ConfigBits\[371\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit9 net80 Tile_X0Y1_FrameStrobe_O\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[351\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame1_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_69_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit11 net231 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[331\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit22 net243 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[342\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot_strobe_inbuf_2__0_ net273 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_2__0_/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_strobe_outbuf_7__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_7__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[7\] sky130_fd_sc_hd__buf_8
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG1 net287
+ net187 Tile_X0Y0_S2BEGb\[2\] net374 Tile_X0Y1_DSP_bot/ConfigBits\[234\] Tile_X0Y1_DSP_bot/ConfigBits\[235\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_CD_BEG\[1\] sky130_fd_sc_hd__mux4_1
XFILLER_0_45_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1113_ Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1113_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1113_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/B sky130_fd_sc_hd__nand4_4
XFILLER_0_158_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_N1BEG3 Tile_X0Y1_DSP_bot/Q5
+ Tile_X0Y1_DSP_bot/J2MID_ABb_BEG\[2\] Tile_X0Y1_DSP_bot/JW2BEG\[2\] Tile_X0Y1_DSP_bot/J_l_AB_BEG\[0\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[12\] Tile_X0Y1_DSP_bot/ConfigBits\[13\] VGND VGND
+ VPWR VPWR Tile_X0Y1_N1BEG\[3\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1044_ Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1028_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1043_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1044_/Y
+ sky130_fd_sc_hd__o21bai_4
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 net763 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[296\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[297\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/J2MID_ABa_BEG\[2\] Tile_X0Y1_DSP_bot/J2MID_CDa_BEG\[2\] Tile_X0Y1_DSP_bot/J2MID_EFa_BEG\[2\]
+ Tile_X0Y1_DSP_bot/J2MID_GHa_BEG\[2\] Tile_X0Y1_DSP_bot/ConfigBits\[58\] Tile_X0Y1_DSP_bot/ConfigBits\[59\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit15 net235 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[239\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit26 net247 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[250\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__34_ Tile_X0Y0_DSP_top/JS2BEG\[2\] VGND
+ VGND VPWR VPWR Tile_X0Y0_S2BEG\[2\] sky130_fd_sc_hd__buf_2
XFILLER_0_100_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_WW4BEG_outbuf_5__0_ Tile_X0Y1_DSP_bot/WW4BEG_i\[5\] VGND VGND VPWR
+ VPWR net758 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1731_ net333 Tile_X0Y1_DSP_bot/A5 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1731_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1662_ Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/B
+ Tile_X0Y1_DSP_bot/ConfigBits\[4\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/X
+ sky130_fd_sc_hd__and3_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1593_ Tile_X0Y1_DSP_bot_Inst_MULADD__1593_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1593_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1594_/B
+ sky130_fd_sc_hd__nor3_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1027_ Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[346\] Tile_X0Y0_DSP_top/ConfigBits\[347\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit10 net230 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[362\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit21 net242 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[373\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit30 net72 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[116\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit19 net239 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[147\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame8_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[3\] Tile_X0Y1_N2BEGb\[7\] net4 net12 Tile_X0Y0_DSP_top/ConfigBits\[334\]
+ Tile_X0Y0_DSP_top/ConfigBits\[335\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__17_ ANTENNA_61/DIODE VGND VGND VPWR
+ VPWR net487 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit4 net75 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[154\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput340 Tile_X0Y1_W2END[2] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_2
Xinput351 Tile_X0Y1_W2MID[5] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_4
Xinput362 Tile_X0Y1_W6END[6] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_1
Xinput373 Tile_X0Y1_WW4END[1] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_WW4END_inbuf_8__0_ net369 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/WW4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_NN4BEG_outbuf_2__0_ Tile_X0Y0_DSP_top/NN4BEG_i\[2\] VGND VGND VPWR
+ VPWR net526 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1714_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1714_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1645_ Tile_X0Y1_DSP_bot_Inst_MULADD__1645_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1700_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1645_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1645_/Y sky130_fd_sc_hd__nand4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/ConfigBits\[258\] Tile_X0Y0_DSP_top/ConfigBits\[259\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1576_ Tile_X0Y1_DSP_bot_Inst_MULADD__1578_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1578_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1577_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1577_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1629_/A sky130_fd_sc_hd__o2bb2ai_2
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG0 Tile_X0Y1_N2BEG\[6\]
+ net19 net99 Tile_X0Y0_DSP_top/JN2BEG\[6\] Tile_X0Y0_DSP_top/ConfigBits\[174\] Tile_X0Y0_DSP_top/ConfigBits\[175\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[0\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit2 net251 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[290\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__3_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__3_/A
+ Tile_X0Y0_DSP_top/ConfigBits\[80\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit14 net234 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[270\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit25 net246 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[281\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_138_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_SS4BEG_outbuf_5__0_ Tile_X0Y0_DSP_top/SS4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_SS4BEG\[5\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__79_ net347 VGND VGND VPWR VPWR net728
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit5 net256 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[37\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[368\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[369\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1430_ Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1501_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1439_/B sky130_fd_sc_hd__nand4_4
Xinput170 Tile_X0Y0_WW4END[14] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_1
Xinput181 Tile_X0Y1_E1END[0] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1361_ Tile_X0Y1_DSP_bot_Inst_MULADD__1298_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1354_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1369_/A sky130_fd_sc_hd__a22o_1
Xinput192 Tile_X0Y1_E2END[7] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1292_ Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1281_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1292_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1
+ net81 net83 net91 net135 Tile_X0Y0_DSP_top/ConfigBits\[298\] Tile_X0Y0_DSP_top/ConfigBits\[299\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit20 net241 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[404\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit31 net253 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[415\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_131_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit29 net250 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[189\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit18 net238 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[178\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[310\] Tile_X0Y0_DSP_top/ConfigBits\[311\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
Xoutput600 net600 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput611 net611 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput622 net622 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput633 net633 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[11] sky130_fd_sc_hd__buf_2
Xoutput644 net644 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput677 net677 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput666 net666 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[3] sky130_fd_sc_hd__buf_2
Xoutput688 net688 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput655 net655 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[31] sky130_fd_sc_hd__buf_2
Xoutput699 net699 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[0] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1628_ Tile_X0Y1_DSP_bot_Inst_MULADD__1665_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1637_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/B sky130_fd_sc_hd__xnor2_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1559_ Tile_X0Y1_DSP_bot_Inst_MULADD__1559_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q12 sky130_fd_sc_hd__buf_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit7 net78 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[253\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_EE4BEG_outbuf_10__0_ Tile_X0Y1_DSP_bot/EE4BEG_i\[10\] VGND VGND
+ VPWR VPWR net616 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 max_cap764/A Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/ConfigBits\[280\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[281\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_220 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_WW4END_inbuf_4__0_ net179 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/WW4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0930_ Tile_X0Y1_DSP_bot_Inst_MULADD__0896_/X Tile_X0Y1_DSP_bot_Inst_MULADD__0900_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0929_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__0890_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0942_/A sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0861_ Tile_X0Y1_DSP_bot/A1 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0889_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_0_140_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit13 net233 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[301\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit24 net245 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[312\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_48_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1413_ Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1465_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1415_/A
+ sky130_fd_sc_hd__and3_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1344_ Tile_X0Y1_DSP_bot_Inst_MULADD__1258_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1686_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1686_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1343_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q8 sky130_fd_sc_hd__a31o_4
XFILLER_0_78_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit5 net256 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[389\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1275_ Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1275_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1275_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_86_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput452 net452 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[2] sky130_fd_sc_hd__clkbuf_4
Xoutput441 net441 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[1] sky130_fd_sc_hd__clkbuf_4
Xoutput430 net430 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput463 net463 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[10] sky130_fd_sc_hd__clkbuf_4
Xoutput474 net474 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[2] sky130_fd_sc_hd__clkbuf_4
Xoutput485 net485 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput496 net496 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[86\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q5 wire763/A Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q9 Tile_X0Y1_DSP_bot/ConfigBits\[332\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[333\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit28 net249 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[220\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit17 net237 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[209\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_140_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1060_ Tile_X0Y1_DSP_bot_Inst_MULADD__1056_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1059_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1046_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1060_/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_157_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_E6BEG_outbuf_0__0_ Tile_X0Y1_DSP_bot/E6BEG_i\[0\] VGND VGND VPWR
+ VPWR net603 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_NN4BEG_outbuf_8__0_ Tile_X0Y1_DSP_bot/NN4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y1_NN4BEG\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__0913_ Tile_X0Y1_DSP_bot_Inst_MULADD__1252_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0911_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0912_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0915_/B
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0844_ Tile_X0Y1_DSP_bot/C0 Tile_X0Y1_DSP_bot_Inst_MULADD__1742_/Q
+ Tile_X0Y1_DSP_bot/ConfigBits\[2\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0844_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_N4BEG1 net288 net309
+ net201 Tile_X0Y1_DSP_bot/Q5 Tile_X0Y1_DSP_bot/ConfigBits\[16\] Tile_X0Y1_DSP_bot/ConfigBits\[17\]
+ VGND VGND VPWR VPWR Tile_X0Y1_N4BEG\[13\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1327_ Tile_X0Y1_DSP_bot_Inst_MULADD__1407_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1326_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/B
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1258_ Tile_X0Y1_DSP_bot/ConfigBits\[5\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1258_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1189_ Tile_X0Y1_DSP_bot_Inst_MULADD__1087_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1268_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0875_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1189_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_144_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_S4END_inbuf_2__0_ net113 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/S4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__50_ Tile_X0Y0_DSP_top/JW2BEG\[2\] VGND
+ VGND VPWR VPWR net541 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1
+ net81 net83 net85 net133 Tile_X0Y0_DSP_top/ConfigBits\[370\] Tile_X0Y0_DSP_top/ConfigBits\[371\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit12 net232 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[332\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit23 net244 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[343\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG2 net289
+ net189 Tile_X0Y0_SS4BEG\[2\] net342 Tile_X0Y1_DSP_bot/ConfigBits\[236\] Tile_X0Y1_DSP_bot/ConfigBits\[237\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_CD_BEG\[2\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1112_ Tile_X0Y1_DSP_bot_Inst_MULADD__1124_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1113_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1113_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1118_/A sky130_fd_sc_hd__a22o_2
XFILLER_0_158_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_W6END_inbuf_6__0_ net163 VGND VGND VPWR VPWR ANTENNA_96/DIODE sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_WW4BEG_outbuf_11__0_ Tile_X0Y1_DSP_bot/WW4BEG_i\[11\] VGND VGND
+ VPWR VPWR net749 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1043_ Tile_X0Y1_DSP_bot_Inst_MULADD__1043_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1043_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1043_/Y sky130_fd_sc_hd__nand2_2
XTile_X0Y1_DSP_bot_EE4END_inbuf_9__0_ net217 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/EE4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_126_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit0 net229 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[192\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[298\] Tile_X0Y1_DSP_bot/ConfigBits\[299\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JE2BEG\[2\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_EE4BEG_outbuf_5__0_ Tile_X0Y0_DSP_top/EE4BEG_i\[5\] VGND VGND VPWR
+ VPWR net425 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[60\] Tile_X0Y1_DSP_bot/ConfigBits\[61\] VGND VGND
+ VPWR VPWR net605 sky130_fd_sc_hd__mux4_1
XFILLER_0_132_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit16 net236 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[240\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__33_ ANTENNA_63/DIODE VGND VGND VPWR
+ VPWR Tile_X0Y0_S2BEG\[1\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit27 net248 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[251\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_S4END_inbuf_2__0_ Tile_X0Y0_S4BEG\[6\] VGND VGND VPWR VPWR ANTENNA_107/DIODE
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1730_ net333 Tile_X0Y1_DSP_bot/A4 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1730_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top_SS4END_inbuf_6__0_ net118 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/SS4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1661_ Tile_X0Y1_DSP_bot_Inst_MULADD__1725_/Q VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1661_/Y sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1592_ Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1602_/C
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1594_/A sky130_fd_sc_hd__nand2_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_strobe_outbuf_17__0_ Tile_X0Y1_DSP_bot_strobe_inbuf_17__0_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_FrameStrobe_O\[17\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1026_ Tile_X0Y1_DSP_bot_Inst_MULADD__1045_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1025_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1026_/Y sky130_fd_sc_hd__a221oi_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__95_ Tile_X0Y1_DSP_bot/Q19 VGND VGND
+ VPWR VPWR Tile_X0Y1_bot2top\[9\] sky130_fd_sc_hd__buf_8
XFILLER_0_118_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[348\] Tile_X0Y0_DSP_top/ConfigBits\[349\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JW2BEG\[1\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_W6END_inbuf_6__0_ net364 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/W6BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_126_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit11 net231 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[363\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit22 net243 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[374\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit20 net61 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[106\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit31 net73 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[117\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1
+ net84 net92 net134 net136 Tile_X0Y0_DSP_top/ConfigBits\[334\] Tile_X0Y0_DSP_top/ConfigBits\[335\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__16_ Tile_X0Y0_DSP_top/JN2BEG\[0\] VGND
+ VGND VPWR VPWR net486 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit5 net76 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[155\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_WW4END_inbuf_11__0_ net372 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/WW4BEG_i\[11\]
+ sky130_fd_sc_hd__clkbuf_2
Xinput330 Tile_X0Y1_NN4END[7] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_1
Xinput341 Tile_X0Y1_W2END[3] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_4
Xinput352 Tile_X0Y1_W2MID[6] VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkbuf_4
Xinput363 Tile_X0Y1_W6END[7] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_1
Xinput374 Tile_X0Y1_WW4END[2] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__buf_2
XFILLER_0_26_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_EE4END_inbuf_5__0_ net48 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/EE4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1 Tile_X0Y0_S1BEG\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1713_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1713_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1713_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1644_ Tile_X0Y1_DSP_bot_Inst_MULADD__1645_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1700_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1645_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1644_/X sky130_fd_sc_hd__a22o_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[8\]
+ Tile_X0Y0_DSP_top/ConfigBits\[258\] Tile_X0Y0_DSP_top/ConfigBits\[259\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1575_ Tile_X0Y1_DSP_bot_Inst_MULADD__1719_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1664_/S
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1577_/B sky130_fd_sc_hd__and2b_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit3 net254 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[291\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG1 Tile_X0Y1_N2BEG\[2\]
+ net95 net147 Tile_X0Y0_DSP_top/JE2BEG\[6\] Tile_X0Y0_DSP_top/ConfigBits\[176\] Tile_X0Y0_DSP_top/ConfigBits\[177\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[1\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit15 net235 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[271\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit26 net247 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[282\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_83_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__78_ net346 VGND VGND VPWR VPWR net727
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1009_ Tile_X0Y1_DSP_bot_Inst_MULADD__1009_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q4 sky130_fd_sc_hd__buf_12
XFILLER_0_142_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_N4BEG_outbuf_4__0_ Tile_X0Y1_DSP_bot/N4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N4BEG\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit6 net257 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[38\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[370\] Tile_X0Y1_DSP_bot/ConfigBits\[371\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JW2BEG\[4\] sky130_fd_sc_hd__mux4_2
XFILLER_0_120_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput160 Tile_X0Y0_W6END[5] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
Xinput171 Tile_X0Y0_WW4END[15] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1360_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1353_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1357_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1359_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1381_/A sky130_fd_sc_hd__o22ai_4
Xinput182 Tile_X0Y1_E1END[1] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_4
Xinput193 Tile_X0Y1_E2MID[0] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1291_ Tile_X0Y1_DSP_bot_Inst_MULADD__1273_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1284_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1288_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1290_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1291_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_144_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit10 net230 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[394\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[155\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/C9 sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[298\] Tile_X0Y0_DSP_top/ConfigBits\[299\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit21 net242 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[405\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit30 net72 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[148\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit19 net239 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[179\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame7_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[312\] Tile_X0Y0_DSP_top/ConfigBits\[313\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JS2BEG\[0\] sky130_fd_sc_hd__mux4_2
Xoutput601 net601 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput623 net623 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_0_41_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput612 net612 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput634 net634 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[12] sky130_fd_sc_hd__buf_2
Xoutput645 net645 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput678 net678 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput667 net667 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput656 net656 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_E6BEG_outbuf_9__0_ Tile_X0Y0_DSP_top/E6BEG_i\[9\] VGND VGND VPWR
+ VPWR net413 sky130_fd_sc_hd__clkbuf_1
Xoutput689 net689 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1627_ Tile_X0Y1_DSP_bot_Inst_MULADD__1626_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1722_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1664_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1637_/B
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1558_ Tile_X0Y1_DSP_bot_Inst_MULADD__1694_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1718_/Q
+ Tile_X0Y1_DSP_bot/ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1559_/A
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y0_DSP_top_strobe_outbuf_12__0_ Tile_X0Y0_DSP_top_strobe_inbuf_12__0_/X VGND
+ VGND VPWR VPWR net465 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1489_ Tile_X0Y1_DSP_bot_Inst_MULADD__1486_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1487_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1488_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1489_/Y
+ sky130_fd_sc_hd__o21bai_4
XFILLER_0_68_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_W6BEG_outbuf_4__0_ Tile_X0Y1_DSP_bot/W6BEG_i\[4\] VGND VGND VPWR
+ VPWR net741 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_SS4END_inbuf_11__0_ net123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/SS4BEG_i\[11\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_data_outbuf_2__0_ Tile_X0Y0_DSP_top_data_inbuf_2__0_/X VGND VGND
+ VPWR VPWR net452 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit8 net79 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[254\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/Q5 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/Q8
+ Tile_X0Y1_DSP_bot/ConfigBits\[280\] Tile_X0Y1_DSP_bot/ConfigBits\[281\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_157_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_210 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_221 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__0860_ Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/A sky130_fd_sc_hd__buf_6
XTile_X0Y0_DSP_top_data_inbuf_26__0_ net67 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_26__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit14 net234 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[302\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit25 net246 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[313\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_139_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1412_ Tile_X0Y1_DSP_bot_Inst_MULADD__1412_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1412_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1467_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_155_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1343_ Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1714_/Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1343_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit6 net257 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[390\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1274_ Tile_X0Y1_DSP_bot_Inst_MULADD__1268_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1269_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1270_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1285_/B
+ sky130_fd_sc_hd__o21a_2
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_inbuf_17__0_ net57 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_17__0_/X
+ sky130_fd_sc_hd__buf_1
Xoutput420 net420 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[15] sky130_fd_sc_hd__buf_2
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_N4BEG_outbuf_0__0_ Tile_X0Y0_DSP_top/N4BEG_i\[0\] VGND VGND VPWR
+ VPWR net502 sky130_fd_sc_hd__clkbuf_1
Xoutput453 net453 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput442 net442 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput431 net431 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[10] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0989_ Tile_X0Y1_DSP_bot_Inst_MULADD__0987_/X Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0976_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0989_/Y
+ sky130_fd_sc_hd__a21oi_2
Xoutput464 net464 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[11] sky130_fd_sc_hd__clkbuf_4
Xoutput475 net475 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[3] sky130_fd_sc_hd__clkbuf_4
Xoutput486 net486 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput497 net497 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_data_outbuf_2__0_ Tile_X0Y1_DSP_bot_data_inbuf_2__0_/X VGND VGND
+ VPWR VPWR net653 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[334\] Tile_X0Y1_DSP_bot/ConfigBits\[335\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JS2BEG\[3\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit18 net238 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[210\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit29 net250 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[221\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_data_outbuf_24__0_ Tile_X0Y1_DSP_bot_data_inbuf_24__0_/X VGND VGND
+ VPWR VPWR net647 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst0
+ net283 Tile_X0Y0_S1BEG\[2\] net336 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/ConfigBits\[98\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[99\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__0912_ Tile_X0Y1_DSP_bot_Inst_MULADD__1708_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1252_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0912_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0843_ Tile_X0Y1_DSP_bot/ConfigBits\[5\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/A sky130_fd_sc_hd__buf_4
XTile_X0Y1_DSP_bot_data_inbuf_26__0_ net247 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_26__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_data_outbuf_15__0_ Tile_X0Y1_DSP_bot_data_inbuf_15__0_/X VGND VGND
+ VPWR VPWR net637 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_N4BEG2 net285 net310
+ net357 net763 Tile_X0Y1_DSP_bot/ConfigBits\[18\] Tile_X0Y1_DSP_bot/ConfigBits\[19\]
+ VGND VGND VPWR VPWR Tile_X0Y1_N4BEG\[14\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1326_ Tile_X0Y1_DSP_bot_Inst_MULADD__1526_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1407_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1326_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1346_/C
+ sky130_fd_sc_hd__and3_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1257_ Tile_X0Y1_DSP_bot_Inst_MULADD__1257_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q7 sky130_fd_sc_hd__buf_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1188_ Tile_X0Y1_DSP_bot_Inst_MULADD__1018_/Y Tile_X0Y1_DSP_bot/A7
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1268_/A
+ sky130_fd_sc_hd__a21boi_4
XTile_X0Y0_DSP_top_data_inbuf_8__0_ net79 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_8__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_S4BEG_outbuf_4__0_ Tile_X0Y1_DSP_bot/S4BEG_i\[4\] VGND VGND VPWR
+ VPWR net693 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_W6BEG_outbuf_0__0_ Tile_X0Y0_DSP_top/W6BEG_i\[0\] VGND VGND VPWR
+ VPWR net555 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_data_inbuf_17__0_ net237 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_17__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[370\] Tile_X0Y0_DSP_top/ConfigBits\[371\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit13 net233 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[333\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit24 net245 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[344\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_127_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG3 net285
+ net220 Tile_X0Y0_S2BEGb\[0\] net338 Tile_X0Y1_DSP_bot/ConfigBits\[238\] Tile_X0Y1_DSP_bot/ConfigBits\[239\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/J2END_CD_BEG\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1111_ Tile_X0Y1_DSP_bot_Inst_MULADD__1209_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1355_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1113_/D sky130_fd_sc_hd__nand4_4
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1042_ Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1042_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1043_/B sky130_fd_sc_hd__nand4_4
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit1 net240 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[193\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit0 net49 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[374\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1309_ Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1398_/A
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__32_ Tile_X0Y0_DSP_top/JS2BEG\[0\] VGND
+ VGND VPWR VPWR Tile_X0Y0_S2BEG\[0\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit28 net249 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[252\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit17 net237 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[241\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_data_outbuf_20__0_ Tile_X0Y0_DSP_top_data_inbuf_20__0_/X VGND VGND
+ VPWR VPWR net442 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_cus_mux41_buf_inst0
+ Tile_X0Y1_DSP_bot/JN2BEG\[4\] Tile_X0Y1_DSP_bot/JN2BEG\[6\] Tile_X0Y1_DSP_bot/JE2BEG\[4\]
+ Tile_X0Y1_DSP_bot/JE2BEG\[6\] Tile_X0Y1_DSP_bot/ConfigBits\[150\] Tile_X0Y1_DSP_bot/ConfigBits\[151\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1660_ Tile_X0Y1_DSP_bot_Inst_MULADD__1704_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1659_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1724_/Q VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q18 sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1591_ Tile_X0Y1_DSP_bot_Inst_MULADD__1595_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1595_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1589_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1560_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1590_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1600_/A sky130_fd_sc_hd__o221ai_4
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_data_outbuf_11__0_ Tile_X0Y0_DSP_top_data_inbuf_11__0_/X VGND VGND
+ VPWR VPWR net432 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1025_ Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1054_/C
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1025_/Y
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__94_ Tile_X0Y1_DSP_bot/Q18 VGND VGND
+ VPWR VPWR Tile_X0Y1_bot2top\[8\] sky130_fd_sc_hd__buf_8
XFILLER_0_16_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_161_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_S4BEG_outbuf_0__0_ ANTENNA_86/DIODE VGND VGND VPWR VPWR Tile_X0Y0_S4BEG\[0\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_126_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit12 net232 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[364\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit23 net244 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[375\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit10 net50 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[96\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit21 net62 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[107\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2
+ Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\]
+ Tile_X0Y0_DSP_top/ConfigBits\[334\] Tile_X0Y0_DSP_top/ConfigBits\[335\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_EE4END_inbuf_11__0_ net39 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/EE4BEG_i\[11\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__15_ net20 VGND VGND VPWR VPWR net401
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit6 net77 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[156\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput320 Tile_X0Y1_NN4END[12] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_1
Xinput342 Tile_X0Y1_W2END[4] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_4
Xinput353 Tile_X0Y1_W2MID[7] VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__clkbuf_4
Xinput331 Tile_X0Y1_NN4END[8] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_1
Xinput375 Tile_X0Y1_WW4END[3] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_2
Xinput364 Tile_X0Y1_W6END[8] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_2 Tile_X0Y0_S1BEG\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1712_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1712_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1712_/Q sky130_fd_sc_hd__dfxtp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1643_ Tile_X0Y1_DSP_bot_Inst_MULADD__1665_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1643_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1645_/D sky130_fd_sc_hd__or2_1
XTile_X0Y0_DSP_top_strobe_outbuf_4__0_ Tile_X0Y0_DSP_top_strobe_inbuf_4__0_/X VGND
+ VGND VPWR VPWR net476 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[260\] Tile_X0Y0_DSP_top/ConfigBits\[261\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JN2BEG\[3\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1574_ Tile_X0Y1_DSP_bot_Inst_MULADD__1664_/S Tile_X0Y1_DSP_bot_Inst_MULADD__1574_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1577_/A sky130_fd_sc_hd__nor2_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0
+ net287 net309 net181 net187 Tile_X0Y1_DSP_bot/ConfigBits\[260\] Tile_X0Y1_DSP_bot/ConfigBits\[261\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit4 net255 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[292\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG2 net17
+ net97 net149 Tile_X0Y0_DSP_top/JS2BEG\[6\] Tile_X0Y0_DSP_top/ConfigBits\[178\] Tile_X0Y0_DSP_top/ConfigBits\[179\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[2\] sky130_fd_sc_hd__mux4_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit16 net236 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[272\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit27 net248 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[283\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__77_ net345 VGND VGND VPWR VPWR net726
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1008_ Tile_X0Y1_DSP_bot_Inst_MULADD__1679_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1710_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/A VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1009_/A
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_data_inbuf_1__0_ net240 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_data_inbuf_1__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_NN4END_inbuf_6__0_ Tile_X0Y1_NN4BEG\[10\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/NN4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst0
+ net281 net181 Tile_X0Y0_S1BEG\[0\] Tile_X0Y1_DSP_bot/Q4 Tile_X0Y1_DSP_bot/ConfigBits\[48\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[49\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_SS4BEG_outbuf_11__0_ ANTENNA_111/DIODE VGND VGND VPWR VPWR net701
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit7 net258 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[39\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_120_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_WW4BEG_outbuf_2__0_ Tile_X0Y0_DSP_top/WW4BEG_i\[2\] VGND VGND VPWR
+ VPWR net575 sky130_fd_sc_hd__clkbuf_1
Xinput161 Tile_X0Y0_W6END[6] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
Xinput172 Tile_X0Y0_WW4END[1] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
Xinput150 Tile_X0Y0_W2MID[5] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_2
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_strobe_inbuf_19__0_ Tile_X0Y1_FrameStrobe_O\[19\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_19__0_/X sky130_fd_sc_hd__clkbuf_1
Xinput183 Tile_X0Y1_E1END[2] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_4
Xinput194 Tile_X0Y1_E2MID[1] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1290_ Tile_X0Y1_DSP_bot_Inst_MULADD__1218_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1232_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1289_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1191_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1290_/Y sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_my_mux2_inst__3_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_my_mux2_inst__3_/A
+ Tile_X0Y1_DSP_bot/ConfigBits\[155\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_my_mux2_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[298\] Tile_X0Y0_DSP_top/ConfigBits\[299\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit11 net231 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[395\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit22 net243 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[406\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_160_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit20 net61 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[138\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit31 net73 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[149\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput602 net602 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput624 net624 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput613 net613 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[8] sky130_fd_sc_hd__buf_2
Xoutput635 net635 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput679 net679 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[4] sky130_fd_sc_hd__clkbuf_4
Xoutput668 net668 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput657 net657 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[4] sky130_fd_sc_hd__clkbuf_4
Xoutput646 net646 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[23] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1626_ Tile_X0Y1_DSP_bot/C16 Tile_X0Y1_DSP_bot_Inst_MULADD__1758_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1626_/X
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1557_ Tile_X0Y1_DSP_bot_Inst_MULADD__1557_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1605_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1694_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1488_ Tile_X0Y1_DSP_bot_Inst_MULADD__1089_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1091_/X
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1561_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1488_/Y
+ sky130_fd_sc_hd__o21ai_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_strobe_inbuf_12__0_ net264 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_12__0_/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_N4END_inbuf_10__0_ net306 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/N4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit9 net80 Tile_X0Y1_FrameStrobe_O\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[255\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame4_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_200 Tile_X0Y0_SS4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2/X
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3/X
+ Tile_X0Y1_DSP_bot/ConfigBits\[282\] Tile_X0Y1_DSP_bot/ConfigBits\[283\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/JN2BEG\[6\] sky130_fd_sc_hd__mux4_2
XANTENNA_211 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_N4END_inbuf_2__0_ Tile_X0Y1_N4BEG\[6\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/N4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_106_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit15 net235 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[303\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit26 net247 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[314\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_155_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1411_ Tile_X0Y1_DSP_bot_Inst_MULADD__1411_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1411_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1412_/A sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1342_ Tile_X0Y1_DSP_bot_Inst_MULADD__1342_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1342_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1686_/C sky130_fd_sc_hd__or2_1
XFILLER_0_161_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1273_ Tile_X0Y1_DSP_bot_Inst_MULADD__1437_/D Tile_X0Y1_DSP_bot_Inst_MULADD__1269_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1270_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1285_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1273_/X sky130_fd_sc_hd__o211a_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit7 net258 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[391\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_6_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput410 net410 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_0_120_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput443 net443 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[21] sky130_fd_sc_hd__clkbuf_4
Xoutput432 net432 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[11] sky130_fd_sc_hd__clkbuf_4
Xoutput421 net421 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[1] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0988_ Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/A Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/Y sky130_fd_sc_hd__nand2_1
Xoutput465 net465 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput476 net476 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[4] sky130_fd_sc_hd__clkbuf_4
Xoutput487 net487 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput454 net454 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[31] sky130_fd_sc_hd__clkbuf_4
Xoutput498 net498 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[4] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_MULADD__1609_ Tile_X0Y1_DSP_bot_Inst_MULADD__1620_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1620_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1698_/C sky130_fd_sc_hd__and2_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit30 net72 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[180\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit19 net239 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[211\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_strobe_inbuf_5__0_ net276 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_strobe_inbuf_5__0_/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_68_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst1
+ wire763/A ANTENNA_101/DIODE Tile_X0Y1_DSP_bot/J2MID_CDb_BEG\[1\] Tile_X0Y1_DSP_bot/J2END_GH_BEG\[2\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[98\] Tile_X0Y1_DSP_bot/ConfigBits\[99\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_153_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot_Inst_MULADD__0911_ Tile_X0Y1_DSP_bot/C2 Tile_X0Y1_DSP_bot_Inst_MULADD__1744_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1459_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0911_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_N4END_inbuf_2__0_ net313 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/N4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_S1BEG0 Tile_X0Y1_bot2top\[4\]
+ Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[3\] Tile_X0Y0_DSP_top/JE2BEG\[3\] Tile_X0Y0_DSP_top/J_l_CD_BEG\[1\]
+ Tile_X0Y0_DSP_top/ConfigBits\[56\] Tile_X0Y0_DSP_top/ConfigBits\[57\] VGND VGND
+ VPWR VPWR Tile_X0Y0_S1BEG\[0\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1325_ Tile_X0Y1_DSP_bot_Inst_MULADD__1244_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1263_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1239_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1326_/C sky130_fd_sc_hd__a221o_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux41_buf_N4BEG3 net286 net301
+ net354 Tile_X0Y1_DSP_bot/Q7 Tile_X0Y1_DSP_bot/ConfigBits\[20\] Tile_X0Y1_DSP_bot/ConfigBits\[21\]
+ VGND VGND VPWR VPWR Tile_X0Y1_N4BEG\[15\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1256_ Tile_X0Y1_DSP_bot_Inst_MULADD__1684_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1713_/Q
+ Tile_X0Y1_DSP_bot/ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1257_/A
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[2\] net3 net135 Tile_X0Y1_bot2top\[2\] Tile_X0Y0_DSP_top/ConfigBits\[16\]
+ Tile_X0Y0_DSP_top/ConfigBits\[17\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1187_ Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/C Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/D VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1187_/Y sky130_fd_sc_hd__nand4_4
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[6\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[370\] Tile_X0Y0_DSP_top/ConfigBits\[371\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit14 net234 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[334\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit25 net246 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[345\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_WW4BEG_outbuf_8__0_ Tile_X0Y1_DSP_bot/WW4BEG_i\[8\] VGND VGND VPWR
+ VPWR net761 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1110_ Tile_X0Y1_DSP_bot_Inst_MULADD__1282_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1430_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0982_/D Tile_X0Y1_DSP_bot_Inst_MULADD__0887_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1113_/C sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_158_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1041_ Tile_X0Y1_DSP_bot_Inst_MULADD__1275_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1493_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit2 net251 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[194\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit1 net60 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[375\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1308_ Tile_X0Y1_DSP_bot_Inst_MULADD__1034_/X Tile_X0Y1_DSP_bot/B7
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1305_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1175_/X VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1310_/B sky130_fd_sc_hd__o211a_2
XFILLER_0_35_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_MULADD__1239_ Tile_X0Y1_DSP_bot_Inst_MULADD__1236_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1146_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1149_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1238_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1239_/Y sky130_fd_sc_hd__a221oi_4
XTile_X0Y1_DSP_bot_S4END_inbuf_10__0_ Tile_X0Y0_S4BEG\[14\] VGND VGND VPWR VPWR ANTENNA_187/DIODE
+ sky130_fd_sc_hd__buf_2
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__31_ Tile_X0Y1_N2BEG\[7\] VGND VGND
+ VPWR VPWR net501 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit18 net238 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[242\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit29 net250 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[253\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_97_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/JS2BEG\[4\] Tile_X0Y1_DSP_bot/JS2BEG\[6\] Tile_X0Y1_DSP_bot/JW2BEG\[4\]
+ ANTENNA_184/DIODE Tile_X0Y1_DSP_bot/ConfigBits\[150\] Tile_X0Y1_DSP_bot/ConfigBits\[151\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C8_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_strobe_inbuf_1__0_ Tile_X0Y1_FrameStrobe_O\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top_strobe_inbuf_1__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1590_ Tile_X0Y1_DSP_bot_Inst_MULADD__1593_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1590_/Y sky130_fd_sc_hd__inv_2
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1024_ Tile_X0Y1_DSP_bot_Inst_MULADD__1729_/Q Tile_X0Y1_DSP_bot_Inst_MULADD__1018_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1373_/C Tile_X0Y1_DSP_bot_Inst_MULADD__0895_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1115_/B sky130_fd_sc_hd__o211a_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__93_ Tile_X0Y1_DSP_bot/Q17 VGND VGND
+ VPWR VPWR Tile_X0Y1_bot2top\[7\] sky130_fd_sc_hd__buf_12
XFILLER_0_16_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_NN4BEG_outbuf_5__0_ Tile_X0Y0_DSP_top/NN4BEG_i\[5\] VGND VGND VPWR
+ VPWR net529 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit13 net233 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[365\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit24 net245 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[376\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit11 net51 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[97\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit22 net63 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[108\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3
+ Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[5\] Tile_X0Y1_bot2top\[7\] Tile_X0Y1_bot2top\[9\]
+ Tile_X0Y0_DSP_top/ConfigBits\[334\] Tile_X0Y0_DSP_top/ConfigBits\[335\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[3\] Tile_X0Y1_N2BEGb\[1\] Tile_X0Y1_N4BEG\[1\] net40 Tile_X0Y0_DSP_top/ConfigBits\[278\]
+ Tile_X0Y0_DSP_top/ConfigBits\[279\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_SS4BEG_outbuf_8__0_ Tile_X0Y0_DSP_top/SS4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_SS4BEG\[8\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__14_ net19 VGND VGND VPWR VPWR net400
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit7 net78 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[157\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput321 Tile_X0Y1_NN4END[13] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_1
Xinput310 Tile_X0Y1_N4END[3] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__buf_2
Xinput343 Tile_X0Y1_W2END[5] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_2
Xinput332 Tile_X0Y1_NN4END[9] VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_1
Xinput354 Tile_X0Y1_W6END[0] VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__clkbuf_4
Xinput376 Tile_X0Y1_WW4END[4] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_SS4END_inbuf_0__0_ Tile_X0Y0_SS4BEG\[4\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/SS4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xinput365 Tile_X0Y1_W6END[9] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0
+ net4 net136 Tile_X0Y1_bot2top\[0\] Tile_X0Y1_bot2top\[1\] Tile_X0Y0_DSP_top/ConfigBits\[104\]
+ Tile_X0Y0_DSP_top/ConfigBits\[105\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_3 Tile_X0Y0_S1BEG\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_SS4BEG_outbuf_1__0_ Tile_X0Y1_DSP_bot/SS4BEG_i\[1\] VGND VGND VPWR
+ VPWR net706 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1711_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1711_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1642_ Tile_X0Y1_DSP_bot_Inst_MULADD__1664_/S Tile_X0Y1_DSP_bot_Inst_MULADD__1723_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1640_/X VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1643_/B
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1573_ Tile_X0Y1_DSP_bot/C13 Tile_X0Y1_DSP_bot_Inst_MULADD__1755_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1663_/S VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1574_/B
+ sky130_fd_sc_hd__mux2_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1
+ net201 Tile_X0Y0_S2BEGb\[2\] net340 net354 Tile_X0Y1_DSP_bot/ConfigBits\[260\] Tile_X0Y1_DSP_bot/ConfigBits\[261\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit5 net256 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[293\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG3 Tile_X0Y1_N2BEG\[0\]
+ net13 net145 Tile_X0Y0_DSP_top/JW2BEG\[6\] Tile_X0Y0_DSP_top/ConfigBits\[180\] Tile_X0Y0_DSP_top/ConfigBits\[181\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/J2MID_GHa_BEG\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_107_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit28 net249 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[284\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit17 net237 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[273\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__76_ ANTENNA_184/DIODE VGND VGND VPWR
+ VPWR net725 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1007_ Tile_X0Y1_DSP_bot_Inst_MULADD__1007_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1007_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1679_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_161_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot/Q8 ANTENNA_105/DIODE Tile_X0Y1_DSP_bot/J2MID_GHb_BEG\[1\] Tile_X0Y1_DSP_bot/J2END_CD_BEG\[0\]
+ Tile_X0Y1_DSP_bot/ConfigBits\[48\] Tile_X0Y1_DSP_bot/ConfigBits\[49\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit8 net259 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[40\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput162 Tile_X0Y0_W6END[7] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
Xinput140 Tile_X0Y0_W2END[3] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__buf_4
Xinput151 Tile_X0Y0_W2MID[6] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_4
Xinput173 Tile_X0Y0_WW4END[2] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_2
Xinput184 Tile_X0Y1_E1END[3] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_4
Xinput195 Tile_X0Y1_E2MID[2] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_2
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_WW4END_inbuf_7__0_ net167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/WW4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_my_mux2_inst__2_
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_my_mux2_inst__2_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_C9_my_mux2_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_160_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[300\] Tile_X0Y0_DSP_top/ConfigBits\[301\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JE2BEG\[5\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit12 net232 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[396\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit23 net244 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[407\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit10 net50 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[128\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit21 net62 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[139\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0
+ net283 net289 net301 net189 Tile_X0Y1_DSP_bot/ConfigBits\[300\] Tile_X0Y1_DSP_bot/ConfigBits\[301\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput625 net625 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput603 net603 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput614 net614 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput636 net636 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[14] sky130_fd_sc_hd__clkbuf_4
Xoutput669 net669 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput658 net658 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[5] sky130_fd_sc_hd__buf_2
Xoutput647 net647 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1625_ Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/A Tile_X0Y1_DSP_bot/ConfigBits\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1665_/A sky130_fd_sc_hd__nand2_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1556_ Tile_X0Y1_DSP_bot_Inst_MULADD__1556_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1556_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1605_/A sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1487_ Tile_X0Y1_DSP_bot_Inst_MULADD__1479_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1482_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1483_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1487_/Y
+ sky130_fd_sc_hd__a21oi_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__59_ Tile_X0Y1_DSP_bot/JS2BEG\[5\] VGND
+ VGND VPWR VPWR net672 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_201 Tile_X0Y0_SS4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_212 Tile_X0Y1_bot2top\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit16 net236 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[304\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit27 net248 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[315\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[1\] Tile_X0Y1_N2BEGb\[3\] net8 net24 Tile_X0Y0_DSP_top/ConfigBits\[350\]
+ Tile_X0Y0_DSP_top/ConfigBits\[351\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1410_ Tile_X0Y1_DSP_bot_Inst_MULADD__1411_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1411_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1412_/B VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1465_/A
+ sky130_fd_sc_hd__o21bai_2
XFILLER_0_155_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_MULADD__1341_ Tile_X0Y1_DSP_bot_Inst_MULADD__1342_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1342_/A
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1686_/B sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1272_ Tile_X0Y1_DSP_bot_Inst_MULADD__0875_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1268_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1195_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1197_/Y
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1285_/A sky130_fd_sc_hd__o32ai_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit8 net259 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[392\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_E6BEG_outbuf_3__0_ Tile_X0Y1_DSP_bot/E6BEG_i\[3\] VGND VGND VPWR
+ VPWR net608 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput411 net411 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput400 net400 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput444 net444 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[22] sky130_fd_sc_hd__clkbuf_4
Xoutput433 net433 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput422 net422 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[2] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__0987_ Tile_X0Y1_DSP_bot_Inst_MULADD__1363_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1378_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__0988_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1027_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__0987_/X sky130_fd_sc_hd__a22o_1
Xoutput466 net466 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[13] sky130_fd_sc_hd__clkbuf_4
Xoutput477 net477 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[5] sky130_fd_sc_hd__clkbuf_4
Xoutput455 net455 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput488 net488 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput499 net499 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[5] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit0 net229 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[96\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame9_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1608_ Tile_X0Y1_DSP_bot_Inst_MULADD__1620_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1620_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1258_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1608_/Y
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1539_ Tile_X0Y1_DSP_bot_Inst_MULADD__0963_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1180_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1538_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1489_/Y VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1541_/A sky130_fd_sc_hd__o31a_1
XFILLER_0_96_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_S4END_inbuf_5__0_ net116 VGND VGND VPWR VPWR ANTENNA_89/DIODE sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[146\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_top2bot16_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR Tile_X0Y0_top2bot\[16\] sky130_fd_sc_hd__o21ai_2
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit31 net73 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[181\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit20 net61 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[170\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__0910_ Tile_X0Y1_DSP_bot/ConfigBits\[2\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1459_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux41_buf_S1BEG1 Tile_X0Y1_bot2top\[5\]
+ ANTENNA_177/DIODE Tile_X0Y0_DSP_top/JE2BEG\[0\] Tile_X0Y0_DSP_top/J_l_EF_BEG\[2\]
+ Tile_X0Y0_DSP_top/ConfigBits\[58\] Tile_X0Y0_DSP_top/ConfigBits\[59\] VGND VGND
+ VPWR VPWR Tile_X0Y0_S1BEG\[1\] sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1324_ Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1324_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1407_/A
+ sky130_fd_sc_hd__nand3_4
XFILLER_0_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_W6END_inbuf_9__0_ net155 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/W6BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1255_ Tile_X0Y1_DSP_bot_Inst_MULADD__1255_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1255_/B
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1684_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_59_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[6\] Tile_X0Y0_DSP_top/J2MID_ABb_BEG\[1\] Tile_X0Y0_DSP_top/J2MID_CDb_BEG\[1\]
+ Tile_X0Y0_DSP_top/J2END_GH_BEG\[1\] Tile_X0Y0_DSP_top/ConfigBits\[16\] Tile_X0Y0_DSP_top/ConfigBits\[17\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__3_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1186_ Tile_X0Y1_DSP_bot_Inst_MULADD__1098_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1184_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1185_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1431_/D
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_144_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top_inst_clk_buf Tile_X0Y1_UserCLKo VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[0\] net81 net133 Tile_X0Y1_bot2top\[4\] Tile_X0Y0_DSP_top/ConfigBits\[98\]
+ Tile_X0Y0_DSP_top/ConfigBits\[99\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[372\] Tile_X0Y0_DSP_top/ConfigBits\[373\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JW2BEG\[7\] sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_EE4BEG_outbuf_8__0_ Tile_X0Y0_DSP_top/EE4BEG_i\[8\] VGND VGND VPWR
+ VPWR net428 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0
+ net283 net291 net183 net191 Tile_X0Y1_DSP_bot/ConfigBits\[372\] Tile_X0Y1_DSP_bot/ConfigBits\[373\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit15 net235 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[335\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit26 net247 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[346\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame2_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_S4END_inbuf_5__0_ Tile_X0Y0_S4BEG\[9\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/S4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_150_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0
+ Tile_X0Y1_NN4BEG\[2\] net1 net41 net21 Tile_X0Y0_DSP_top/ConfigBits\[314\] Tile_X0Y0_DSP_top/ConfigBits\[315\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1040_ Tile_X0Y1_DSP_bot_Inst_MULADD__1277_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1038_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1039_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1275_/B
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__4_
+ Tile_X0Y0_DSP_top/ConfigBits\[38\] Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_/Y
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__o21ai_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_EE4BEG_outbuf_1__0_ Tile_X0Y1_DSP_bot/EE4BEG_i\[1\] VGND VGND VPWR
+ VPWR net622 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_SS4END_inbuf_9__0_ net121 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/SS4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit3 net254 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[195\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame6_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit2 net71 Tile_X0Y1_FrameStrobe_O\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[376\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame0_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1307_ Tile_X0Y1_DSP_bot_Inst_MULADD__1291_/Y Tile_X0Y1_DSP_bot_Inst_MULADD__1297_/Y
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1306_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1313_/B
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1238_ Tile_X0Y1_DSP_bot_Inst_MULADD__1237_/X Tile_X0Y1_DSP_bot_Inst_MULADD__1183_/A
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1241_/B VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1238_/Y sky130_fd_sc_hd__a22oi_4
XTile_X0Y1_DSP_bot_W6END_inbuf_9__0_ net356 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/W6BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1169_ Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1683_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/Y VGND VGND VPWR VPWR wire763/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_129_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__30_ Tile_X0Y1_N2BEG\[6\] VGND VGND
+ VPWR VPWR net500 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit30 net72 Tile_X0Y1_FrameStrobe_O\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[212\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame6_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit19 net239 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[243\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame5_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1023_ Tile_X0Y1_DSP_bot_Inst_MULADD__1085_/A Tile_X0Y1_DSP_bot/A3
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1373_/C sky130_fd_sc_hd__or2_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__92_ Tile_X0Y1_DSP_bot/Q16 VGND VGND
+ VPWR VPWR Tile_X0Y1_bot2top\[6\] sky130_fd_sc_hd__buf_12
XTile_X0Y0_DSP_top_EE4END_inbuf_8__0_ net36 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/EE4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit14 net234 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[366\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit25 net246 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[377\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame1_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit23 net64 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[109\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit12 net52 Tile_X0Y1_FrameStrobe_O\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[98\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame9_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2/X
+ Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3/X
+ Tile_X0Y0_DSP_top/ConfigBits\[336\] Tile_X0Y0_DSP_top/ConfigBits\[337\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top/JS2BEG\[6\] sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1
+ net24 net86 net138 net156 Tile_X0Y0_DSP_top/ConfigBits\[278\] Tile_X0Y0_DSP_top/ConfigBits\[279\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_153_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0
+ net282 net290 net182 net190 Tile_X0Y1_DSP_bot/ConfigBits\[336\] Tile_X0Y1_DSP_bot/ConfigBits\[337\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot_N4BEG_outbuf_7__0_ Tile_X0Y1_DSP_bot/N4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y1_N4BEG\[7\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix__13_ net18 VGND VGND VPWR VPWR net399
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit8 net79 Tile_X0Y1_FrameStrobe_O\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[158\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame7_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst0
+ Tile_X0Y1_N1BEG\[2\] net3 net135 Tile_X0Y1_bot2top\[2\] Tile_X0Y0_DSP_top/ConfigBits\[72\]
+ Tile_X0Y0_DSP_top/ConfigBits\[73\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__2_/A
+ sky130_fd_sc_hd__mux4_1
Xinput300 Tile_X0Y1_N2MID[7] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkbuf_4
Xinput311 Tile_X0Y1_N4END[4] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_1
Xinput344 Tile_X0Y1_W2END[6] VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput322 Tile_X0Y1_NN4END[14] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_1
Xinput333 Tile_X0Y1_UserCLK VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__buf_12
Xinput377 Tile_X0Y1_WW4END[5] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkbuf_1
Xinput366 Tile_X0Y1_WW4END[0] VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__buf_2
Xinput355 Tile_X0Y1_W6END[10] VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1
+ Tile_X0Y1_bot2top\[2\] Tile_X0Y1_bot2top\[3\] Tile_X0Y1_bot2top\[4\] Tile_X0Y1_bot2top\[5\]
+ Tile_X0Y0_DSP_top/ConfigBits\[104\] Tile_X0Y0_DSP_top/ConfigBits\[105\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top_Inst_DSP_top_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_4 Tile_X0Y0_S1BEG\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot_Inst_MULADD__1710_ net333 Tile_X0Y1_DSP_bot_Inst_MULADD__1710_/D
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot_Inst_MULADD__1641_ Tile_X0Y1_DSP_bot_Inst_MULADD__1664_/S Tile_X0Y1_DSP_bot_Inst_MULADD__1723_/Q
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1662_/A Tile_X0Y1_DSP_bot/ConfigBits\[4\] Tile_X0Y1_DSP_bot_Inst_MULADD__1640_/X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1653_/C sky130_fd_sc_hd__a221o_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1572_ Tile_X0Y1_DSP_bot_Inst_MULADD__1593_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1593_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1547_/B Tile_X0Y1_DSP_bot_Inst_MULADD__1554_/A VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1578_/B sky130_fd_sc_hd__o211ai_2
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot/Q0 Tile_X0Y1_DSP_bot/Q2 Tile_X0Y1_DSP_bot/Q3 Tile_X0Y1_DSP_bot/Q4
+ Tile_X0Y1_DSP_bot/ConfigBits\[260\] Tile_X0Y1_DSP_bot/ConfigBits\[261\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit6 net257 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[294\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame3_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__4_
+ Tile_X0Y1_DSP_bot/ConfigBits\[44\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__2_/Y
+ Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__3_/Y
+ VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit18 net238 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[274\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_88_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit29 net250 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[285\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame4_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_119_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix__75_ Tile_X0Y1_DSP_bot/JW2BEG\[5\] VGND
+ VGND VPWR VPWR net724 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1006_ Tile_X0Y1_DSP_bot_Inst_MULADD__1006_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1006_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1006_/C VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_MULADD__1007_/B
+ sky130_fd_sc_hd__or3_1
XFILLER_0_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top_NN4END_inbuf_11__0_ Tile_X0Y1_NN4BEG\[15\] VGND VGND VPWR VPWR
+ ANTENNA_78/DIODE sky130_fd_sc_hd__buf_2
XFILLER_0_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_strobe_outbuf_15__0_ Tile_X0Y0_DSP_top_strobe_inbuf_15__0_/X VGND
+ VGND VPWR VPWR net468 sky130_fd_sc_hd__clkbuf_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_W6BEG_outbuf_7__0_ ANTENNA_112/DIODE VGND VGND VPWR VPWR net744
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top_data_outbuf_5__0_ Tile_X0Y0_DSP_top_data_inbuf_5__0_/X VGND VGND
+ VPWR VPWR net457 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit9 net260 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[41\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame11_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput130 Tile_X0Y0_SS4END[7] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
Xinput163 Tile_X0Y0_W6END[8] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_1
Xinput141 Tile_X0Y0_W2END[4] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_4
Xinput152 Tile_X0Y0_W2MID[7] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_4
Xinput174 Tile_X0Y0_WW4END[3] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
Xinput196 Tile_X0Y1_E2MID[3] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_2
Xinput185 Tile_X0Y1_E2END[0] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_85_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit13 net233 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[397\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit24 net245 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot/ConfigBits\[408\] Tile_X0Y1_DSP_bot_Inst_DSP_bot_ConfigMem_Inst_frame0_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit11 net51 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[129\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1
+ net201 Tile_X0Y0_S2BEGb\[4\] net342 net354 Tile_X0Y1_DSP_bot/ConfigBits\[300\] Tile_X0Y1_DSP_bot/ConfigBits\[301\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot_Inst_DSP_bot_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit22 net63 Tile_X0Y1_FrameStrobe_O\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top/ConfigBits\[140\] Tile_X0Y0_DSP_top_Inst_DSP_top_ConfigMem_Inst_frame8_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top_data_inbuf_29__0_ net70 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top_data_inbuf_29__0_/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput615 net615 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput626 net626 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput604 net604 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput659 net659 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[6] sky130_fd_sc_hd__buf_2
Xoutput637 net637 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[15] sky130_fd_sc_hd__clkbuf_4
Xoutput648 net648 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[25] sky130_fd_sc_hd__buf_2
XFILLER_0_1_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot_Inst_MULADD__1624_ Tile_X0Y1_DSP_bot_Inst_MULADD__1168_/A Tile_X0Y1_DSP_bot_Inst_MULADD__1699_/B
+ Tile_X0Y1_DSP_bot_Inst_MULADD__1623_/Y VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot/Q15
+ sky130_fd_sc_hd__o21ai_1
.ends

