magic
tech sky130A
magscale 1 2
timestamp 1733394400
<< viali >>
rect 1685 8585 1719 8619
rect 2789 8585 2823 8619
rect 3157 8585 3191 8619
rect 3525 8585 3559 8619
rect 4261 8585 4295 8619
rect 4629 8585 4663 8619
rect 5181 8585 5215 8619
rect 6101 8585 6135 8619
rect 6837 8585 6871 8619
rect 7389 8585 7423 8619
rect 7757 8585 7791 8619
rect 8309 8585 8343 8619
rect 8677 8585 8711 8619
rect 9229 8585 9263 8619
rect 9781 8585 9815 8619
rect 10149 8585 10183 8619
rect 10701 8585 10735 8619
rect 11253 8585 11287 8619
rect 11805 8585 11839 8619
rect 12357 8585 12391 8619
rect 12909 8585 12943 8619
rect 13277 8585 13311 8619
rect 13829 8585 13863 8619
rect 14381 8585 14415 8619
rect 14749 8585 14783 8619
rect 15301 8585 15335 8619
rect 15853 8585 15887 8619
rect 16405 8585 16439 8619
rect 17141 8585 17175 8619
rect 17509 8585 17543 8619
rect 17877 8585 17911 8619
rect 18245 8585 18279 8619
rect 18981 8585 19015 8619
rect 19533 8585 19567 8619
rect 20085 8585 20119 8619
rect 22201 8585 22235 8619
rect 22477 8585 22511 8619
rect 23029 8585 23063 8619
rect 24041 8585 24075 8619
rect 27997 8585 28031 8619
rect 30205 8585 30239 8619
rect 30941 8585 30975 8619
rect 32321 8585 32355 8619
rect 32597 8585 32631 8619
rect 34437 8585 34471 8619
rect 34897 8585 34931 8619
rect 35173 8585 35207 8619
rect 36277 8585 36311 8619
rect 37013 8585 37047 8619
rect 37473 8585 37507 8619
rect 37749 8585 37783 8619
rect 38853 8585 38887 8619
rect 39221 8585 39255 8619
rect 39589 8585 39623 8619
rect 40049 8585 40083 8619
rect 40601 8585 40635 8619
rect 41521 8585 41555 8619
rect 42625 8585 42659 8619
rect 42993 8585 43027 8619
rect 44465 8585 44499 8619
rect 45201 8585 45235 8619
rect 3985 8517 4019 8551
rect 4905 8517 4939 8551
rect 10425 8517 10459 8551
rect 40509 8517 40543 8551
rect 41429 8517 41463 8551
rect 1501 8449 1535 8483
rect 2145 8449 2179 8483
rect 2513 8449 2547 8483
rect 2973 8449 3007 8483
rect 3341 8449 3375 8483
rect 4445 8449 4479 8483
rect 5917 8449 5951 8483
rect 6561 8449 6595 8483
rect 7205 8449 7239 8483
rect 7573 8449 7607 8483
rect 8033 8449 8067 8483
rect 8493 8449 8527 8483
rect 9045 8449 9079 8483
rect 9505 8449 9539 8483
rect 9965 8449 9999 8483
rect 10977 8449 11011 8483
rect 11621 8449 11655 8483
rect 12081 8449 12115 8483
rect 12725 8449 12759 8483
rect 13093 8449 13127 8483
rect 13553 8449 13587 8483
rect 14197 8449 14231 8483
rect 14565 8449 14599 8483
rect 15025 8449 15059 8483
rect 15669 8449 15703 8483
rect 16129 8449 16163 8483
rect 16957 8449 16991 8483
rect 17325 8449 17359 8483
rect 17693 8449 17727 8483
rect 18153 8449 18187 8483
rect 18797 8449 18831 8483
rect 19441 8449 19475 8483
rect 19993 8449 20027 8483
rect 20821 8449 20855 8483
rect 21097 8449 21131 8483
rect 21373 8449 21407 8483
rect 21649 8449 21683 8483
rect 22109 8449 22143 8483
rect 22385 8449 22419 8483
rect 22661 8449 22695 8483
rect 22937 8449 22971 8483
rect 23213 8449 23247 8483
rect 23489 8449 23523 8483
rect 23581 8449 23615 8483
rect 23857 8449 23891 8483
rect 24593 8449 24627 8483
rect 24869 8449 24903 8483
rect 25237 8449 25271 8483
rect 25605 8449 25639 8483
rect 25973 8449 26007 8483
rect 26341 8449 26375 8483
rect 26709 8449 26743 8483
rect 27169 8449 27203 8483
rect 27445 8449 27479 8483
rect 27813 8449 27847 8483
rect 28181 8449 28215 8483
rect 28549 8449 28583 8483
rect 28917 8449 28951 8483
rect 29285 8449 29319 8483
rect 29745 8449 29779 8483
rect 30021 8449 30055 8483
rect 30389 8449 30423 8483
rect 30757 8449 30791 8483
rect 31125 8449 31159 8483
rect 31493 8449 31527 8483
rect 31677 8449 31711 8483
rect 32137 8449 32171 8483
rect 32413 8449 32447 8483
rect 32781 8449 32815 8483
rect 33149 8449 33183 8483
rect 33517 8449 33551 8483
rect 33885 8449 33919 8483
rect 34253 8449 34287 8483
rect 34713 8449 34747 8483
rect 34989 8449 35023 8483
rect 35357 8449 35391 8483
rect 35725 8449 35759 8483
rect 36093 8449 36127 8483
rect 36461 8449 36495 8483
rect 36829 8449 36863 8483
rect 37289 8449 37323 8483
rect 37565 8449 37599 8483
rect 37933 8449 37967 8483
rect 38301 8449 38335 8483
rect 38669 8449 38703 8483
rect 39037 8449 39071 8483
rect 39405 8449 39439 8483
rect 39957 8449 39991 8483
rect 40969 8449 41003 8483
rect 41889 8449 41923 8483
rect 42441 8449 42475 8483
rect 42901 8449 42935 8483
rect 43453 8449 43487 8483
rect 43913 8449 43947 8483
rect 44373 8449 44407 8483
rect 45109 8449 45143 8483
rect 5641 8381 5675 8415
rect 21925 8313 21959 8347
rect 23765 8313 23799 8347
rect 24409 8313 24443 8347
rect 26525 8313 26559 8347
rect 27629 8313 27663 8347
rect 30573 8313 30607 8347
rect 31861 8313 31895 8347
rect 34069 8313 34103 8347
rect 35541 8313 35575 8347
rect 35909 8313 35943 8347
rect 36645 8313 36679 8347
rect 38117 8313 38151 8347
rect 38485 8313 38519 8347
rect 41153 8313 41187 8347
rect 42073 8313 42107 8347
rect 43637 8313 43671 8347
rect 44097 8313 44131 8347
rect 20637 8245 20671 8279
rect 20913 8245 20947 8279
rect 21189 8245 21223 8279
rect 21465 8245 21499 8279
rect 22753 8245 22787 8279
rect 23305 8245 23339 8279
rect 24685 8245 24719 8279
rect 25053 8245 25087 8279
rect 25421 8245 25455 8279
rect 25789 8245 25823 8279
rect 26157 8245 26191 8279
rect 26985 8245 27019 8279
rect 27261 8245 27295 8279
rect 28365 8245 28399 8279
rect 28733 8245 28767 8279
rect 29101 8245 29135 8279
rect 29561 8245 29595 8279
rect 29837 8245 29871 8279
rect 31309 8245 31343 8279
rect 32965 8245 32999 8279
rect 33333 8245 33367 8279
rect 33701 8245 33735 8279
rect 1869 8041 1903 8075
rect 2973 8041 3007 8075
rect 4629 8041 4663 8075
rect 5733 8041 5767 8075
rect 6653 8041 6687 8075
rect 7205 8041 7239 8075
rect 9229 8041 9263 8075
rect 10149 8041 10183 8075
rect 11805 8041 11839 8075
rect 12725 8041 12759 8075
rect 14381 8041 14415 8075
rect 15669 8041 15703 8075
rect 17877 8041 17911 8075
rect 18613 8041 18647 8075
rect 19625 8041 19659 8075
rect 21005 8041 21039 8075
rect 21281 8041 21315 8075
rect 21833 8041 21867 8075
rect 22569 8041 22603 8075
rect 22845 8041 22879 8075
rect 23121 8041 23155 8075
rect 23949 8041 23983 8075
rect 24225 8041 24259 8075
rect 24777 8041 24811 8075
rect 25881 8041 25915 8075
rect 26157 8041 26191 8075
rect 26709 8041 26743 8075
rect 27077 8041 27111 8075
rect 27813 8041 27847 8075
rect 28917 8041 28951 8075
rect 41153 8041 41187 8075
rect 45201 8041 45235 8075
rect 2513 7973 2547 8007
rect 4169 7973 4203 8007
rect 18153 7973 18187 8007
rect 22109 7973 22143 8007
rect 27445 7973 27479 8007
rect 44557 7973 44591 8007
rect 1777 7837 1811 7871
rect 2789 7837 2823 7871
rect 4445 7837 4479 7871
rect 6561 7837 6595 7871
rect 7021 7837 7055 7871
rect 9965 7837 9999 7871
rect 12541 7837 12575 7871
rect 15485 7837 15519 7871
rect 17785 7837 17819 7871
rect 18061 7837 18095 7871
rect 18337 7837 18371 7871
rect 18429 7837 18463 7871
rect 18889 7837 18923 7871
rect 19349 7837 19383 7871
rect 19809 7837 19843 7871
rect 19901 7837 19935 7871
rect 20177 7837 20211 7871
rect 20453 7837 20487 7871
rect 20729 7837 20763 7871
rect 21189 7837 21223 7871
rect 21465 7837 21499 7871
rect 21557 7837 21591 7871
rect 22017 7837 22051 7871
rect 22293 7837 22327 7871
rect 22385 7837 22419 7871
rect 22661 7837 22695 7871
rect 22937 7837 22971 7871
rect 23213 7837 23247 7871
rect 23489 7837 23523 7871
rect 23765 7837 23799 7871
rect 24041 7837 24075 7871
rect 24593 7837 24627 7871
rect 24869 7837 24903 7871
rect 25145 7837 25179 7871
rect 25421 7837 25455 7871
rect 25697 7837 25731 7871
rect 25973 7837 26007 7871
rect 26249 7837 26283 7871
rect 26525 7837 26559 7871
rect 26893 7837 26927 7871
rect 27261 7837 27295 7871
rect 27629 7837 27663 7871
rect 27997 7837 28031 7871
rect 28365 7837 28399 7871
rect 28733 7837 28767 7871
rect 40969 7837 41003 7871
rect 44097 7837 44131 7871
rect 2329 7769 2363 7803
rect 3985 7769 4019 7803
rect 5457 7769 5491 7803
rect 9137 7769 9171 7803
rect 11713 7769 11747 7803
rect 14289 7769 14323 7803
rect 43729 7769 43763 7803
rect 44281 7769 44315 7803
rect 45109 7769 45143 7803
rect 17601 7701 17635 7735
rect 19073 7701 19107 7735
rect 19533 7701 19567 7735
rect 20085 7701 20119 7735
rect 20361 7701 20395 7735
rect 20637 7701 20671 7735
rect 20913 7701 20947 7735
rect 21741 7701 21775 7735
rect 23397 7701 23431 7735
rect 23673 7701 23707 7735
rect 25053 7701 25087 7735
rect 25329 7701 25363 7735
rect 25605 7701 25639 7735
rect 26433 7701 26467 7735
rect 28181 7701 28215 7735
rect 28549 7701 28583 7735
rect 1593 7497 1627 7531
rect 2145 7497 2179 7531
rect 18889 7497 18923 7531
rect 19533 7497 19567 7531
rect 20361 7497 20395 7531
rect 21557 7497 21591 7531
rect 22017 7497 22051 7531
rect 22661 7497 22695 7531
rect 44097 7497 44131 7531
rect 45201 7497 45235 7531
rect 44741 7429 44775 7463
rect 1501 7361 1535 7395
rect 1961 7361 1995 7395
rect 19073 7361 19107 7395
rect 19349 7361 19383 7395
rect 19717 7361 19751 7395
rect 20085 7361 20119 7395
rect 20545 7361 20579 7395
rect 20821 7361 20855 7395
rect 21373 7361 21407 7395
rect 21833 7361 21867 7395
rect 22109 7361 22143 7395
rect 22385 7361 22419 7395
rect 22845 7361 22879 7395
rect 23121 7361 23155 7395
rect 23397 7361 23431 7395
rect 23673 7361 23707 7395
rect 23949 7361 23983 7395
rect 43913 7361 43947 7395
rect 44373 7361 44407 7395
rect 44925 7361 44959 7395
rect 19165 7225 19199 7259
rect 20637 7225 20671 7259
rect 19901 7157 19935 7191
rect 22293 7157 22327 7191
rect 22569 7157 22603 7191
rect 22937 7157 22971 7191
rect 23213 7157 23247 7191
rect 23857 7157 23891 7191
rect 24133 7157 24167 7191
rect 45385 6817 45419 6851
rect 23121 6749 23155 6783
rect 45109 6681 45143 6715
rect 22937 6613 22971 6647
rect 36093 4709 36127 4743
rect 23581 4573 23615 4607
rect 35909 4573 35943 4607
rect 23765 4437 23799 4471
rect 22661 4097 22695 4131
rect 23121 4097 23155 4131
rect 23673 4097 23707 4131
rect 27077 4097 27111 4131
rect 33701 4097 33735 4131
rect 35449 4097 35483 4131
rect 44557 4097 44591 4131
rect 22845 3961 22879 3995
rect 22937 3961 22971 3995
rect 35265 3961 35299 3995
rect 23857 3893 23891 3927
rect 27261 3893 27295 3927
rect 33885 3893 33919 3927
rect 44373 3893 44407 3927
rect 22017 3689 22051 3723
rect 33057 3689 33091 3723
rect 24041 3621 24075 3655
rect 22201 3485 22235 3519
rect 23857 3485 23891 3519
rect 33241 3485 33275 3519
rect 23029 3145 23063 3179
rect 23305 3145 23339 3179
rect 26433 3145 26467 3179
rect 39589 3145 39623 3179
rect 23213 3009 23247 3043
rect 23489 3009 23523 3043
rect 23581 3009 23615 3043
rect 26617 3009 26651 3043
rect 29285 3009 29319 3043
rect 39773 3009 39807 3043
rect 23765 2873 23799 2907
rect 29469 2873 29503 2907
rect 23213 2601 23247 2635
rect 28641 2601 28675 2635
rect 44649 2601 44683 2635
rect 45017 2601 45051 2635
rect 22753 2533 22787 2567
rect 24041 2533 24075 2567
rect 25053 2533 25087 2567
rect 45293 2533 45327 2567
rect 22937 2397 22971 2431
rect 23029 2397 23063 2431
rect 23397 2397 23431 2431
rect 23857 2397 23891 2431
rect 24869 2397 24903 2431
rect 28825 2397 28859 2431
rect 31493 2397 31527 2431
rect 38209 2397 38243 2431
rect 44833 2397 44867 2431
rect 45201 2397 45235 2431
rect 45477 2397 45511 2431
rect 20637 2329 20671 2363
rect 20821 2329 20855 2363
rect 23581 2261 23615 2295
rect 31677 2261 31711 2295
rect 38393 2261 38427 2295
rect 19625 2057 19659 2091
rect 22201 2057 22235 2091
rect 23305 2057 23339 2091
rect 24225 2057 24259 2091
rect 30849 2057 30883 2091
rect 37289 2057 37323 2091
rect 41797 2057 41831 2091
rect 43913 2057 43947 2091
rect 44649 2057 44683 2091
rect 22753 1989 22787 2023
rect 19809 1921 19843 1955
rect 22385 1921 22419 1955
rect 22569 1921 22603 1955
rect 23213 1921 23247 1955
rect 23489 1921 23523 1955
rect 24409 1921 24443 1955
rect 31033 1921 31067 1955
rect 37473 1921 37507 1955
rect 41981 1921 42015 1955
rect 44097 1921 44131 1955
rect 44833 1921 44867 1955
rect 23029 1785 23063 1819
rect 1685 1513 1719 1547
rect 19257 1513 19291 1547
rect 23581 1513 23615 1547
rect 27997 1513 28031 1547
rect 30205 1513 30239 1547
rect 41245 1513 41279 1547
rect 43453 1513 43487 1547
rect 45293 1513 45327 1547
rect 1501 1309 1535 1343
rect 3801 1309 3835 1343
rect 5917 1309 5951 1343
rect 8125 1309 8159 1343
rect 10333 1309 10367 1343
rect 12541 1309 12575 1343
rect 14749 1309 14783 1343
rect 17141 1309 17175 1343
rect 19441 1309 19475 1343
rect 21557 1309 21591 1343
rect 23765 1309 23799 1343
rect 25973 1309 26007 1343
rect 28181 1309 28215 1343
rect 30389 1309 30423 1343
rect 32597 1309 32631 1343
rect 34897 1309 34931 1343
rect 37013 1309 37047 1343
rect 39221 1309 39255 1343
rect 41429 1309 41463 1343
rect 43637 1309 43671 1343
rect 45477 1309 45511 1343
rect 3985 1173 4019 1207
rect 6101 1173 6135 1207
rect 8309 1173 8343 1207
rect 10517 1173 10551 1207
rect 12725 1173 12759 1207
rect 14933 1173 14967 1207
rect 16957 1173 16991 1207
rect 21373 1173 21407 1207
rect 25789 1173 25823 1207
rect 32413 1173 32447 1207
rect 34713 1173 34747 1207
rect 36829 1173 36863 1207
rect 39037 1173 39071 1207
<< metal1 >>
rect 9968 9948 17448 9976
rect 9968 9920 9996 9948
rect 17420 9920 17448 9948
rect 18138 9936 18144 9988
rect 18196 9976 18202 9988
rect 21818 9976 21824 9988
rect 18196 9948 21824 9976
rect 18196 9936 18202 9948
rect 21818 9936 21824 9948
rect 21876 9936 21882 9988
rect 22646 9936 22652 9988
rect 22704 9976 22710 9988
rect 32950 9976 32956 9988
rect 22704 9948 32956 9976
rect 22704 9936 22710 9948
rect 32950 9936 32956 9948
rect 33008 9936 33014 9988
rect 9950 9868 9956 9920
rect 10008 9868 10014 9920
rect 17402 9868 17408 9920
rect 17460 9868 17466 9920
rect 17494 9868 17500 9920
rect 17552 9908 17558 9920
rect 17552 9880 21864 9908
rect 17552 9868 17558 9880
rect 9398 9800 9404 9852
rect 9456 9840 9462 9852
rect 21450 9840 21456 9852
rect 9456 9812 21456 9840
rect 9456 9800 9462 9812
rect 21450 9800 21456 9812
rect 21508 9800 21514 9852
rect 21836 9840 21864 9880
rect 24486 9840 24492 9852
rect 21836 9812 24492 9840
rect 24486 9800 24492 9812
rect 24544 9800 24550 9852
rect 7190 9732 7196 9784
rect 7248 9772 7254 9784
rect 9674 9772 9680 9784
rect 7248 9744 9680 9772
rect 7248 9732 7254 9744
rect 9674 9732 9680 9744
rect 9732 9732 9738 9784
rect 13078 9732 13084 9784
rect 13136 9772 13142 9784
rect 21726 9772 21732 9784
rect 13136 9744 21732 9772
rect 13136 9732 13142 9744
rect 21726 9732 21732 9744
rect 21784 9732 21790 9784
rect 4430 9664 4436 9716
rect 4488 9704 4494 9716
rect 21542 9704 21548 9716
rect 4488 9676 21548 9704
rect 4488 9664 4494 9676
rect 21542 9664 21548 9676
rect 21600 9664 21606 9716
rect 9398 9636 9404 9648
rect 4080 9608 9404 9636
rect 4080 9512 4108 9608
rect 9398 9596 9404 9608
rect 9456 9596 9462 9648
rect 21726 9636 21732 9648
rect 12636 9608 21732 9636
rect 11606 9528 11612 9580
rect 11664 9568 11670 9580
rect 12636 9568 12664 9608
rect 21726 9596 21732 9608
rect 21784 9596 21790 9648
rect 11664 9540 12664 9568
rect 11664 9528 11670 9540
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 21358 9568 21364 9580
rect 12768 9540 21364 9568
rect 12768 9528 12774 9540
rect 21358 9528 21364 9540
rect 21416 9528 21422 9580
rect 38838 9568 38844 9580
rect 35866 9540 38844 9568
rect 4062 9460 4068 9512
rect 4120 9460 4126 9512
rect 9030 9460 9036 9512
rect 9088 9500 9094 9512
rect 21726 9500 21732 9512
rect 9088 9472 21732 9500
rect 9088 9460 9094 9472
rect 21726 9460 21732 9472
rect 21784 9460 21790 9512
rect 21818 9460 21824 9512
rect 21876 9500 21882 9512
rect 21876 9472 23888 9500
rect 21876 9460 21882 9472
rect 23860 9432 23888 9472
rect 23934 9460 23940 9512
rect 23992 9500 23998 9512
rect 35866 9500 35894 9540
rect 38838 9528 38844 9540
rect 38896 9528 38902 9580
rect 23992 9472 35894 9500
rect 23992 9460 23998 9472
rect 32858 9432 32864 9444
rect 12406 9404 16620 9432
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 12406 9364 12434 9404
rect 16592 9376 16620 9404
rect 16684 9404 23796 9432
rect 23860 9404 32864 9432
rect 8352 9336 12434 9364
rect 8352 9324 8358 9336
rect 16574 9324 16580 9376
rect 16632 9324 16638 9376
rect 16684 9296 16712 9404
rect 17402 9324 17408 9376
rect 17460 9364 17466 9376
rect 23658 9364 23664 9376
rect 17460 9336 23664 9364
rect 17460 9324 17466 9336
rect 23658 9324 23664 9336
rect 23716 9324 23722 9376
rect 23768 9364 23796 9404
rect 32858 9392 32864 9404
rect 32916 9392 32922 9444
rect 26142 9364 26148 9376
rect 23768 9336 26148 9364
rect 26142 9324 26148 9336
rect 26200 9324 26206 9376
rect 26234 9324 26240 9376
rect 26292 9364 26298 9376
rect 35158 9364 35164 9376
rect 26292 9336 35164 9364
rect 26292 9324 26298 9336
rect 35158 9324 35164 9336
rect 35216 9324 35222 9376
rect 2746 9268 16712 9296
rect 1486 9188 1492 9240
rect 1544 9228 1550 9240
rect 2746 9228 2774 9268
rect 16758 9256 16764 9308
rect 16816 9296 16822 9308
rect 27798 9296 27804 9308
rect 16816 9268 27804 9296
rect 16816 9256 16822 9268
rect 27798 9256 27804 9268
rect 27856 9256 27862 9308
rect 17494 9228 17500 9240
rect 1544 9200 2774 9228
rect 10428 9200 17500 9228
rect 1544 9188 1550 9200
rect 10428 9172 10456 9200
rect 17494 9188 17500 9200
rect 17552 9188 17558 9240
rect 19610 9228 19616 9240
rect 17604 9200 19616 9228
rect 10410 9120 10416 9172
rect 10468 9120 10474 9172
rect 17126 9160 17132 9172
rect 12406 9132 17132 9160
rect 7558 9052 7564 9104
rect 7616 9092 7622 9104
rect 12406 9092 12434 9132
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 7616 9064 12434 9092
rect 7616 9052 7622 9064
rect 12618 9052 12624 9104
rect 12676 9092 12682 9104
rect 17604 9092 17632 9200
rect 19610 9188 19616 9200
rect 19668 9188 19674 9240
rect 22094 9188 22100 9240
rect 22152 9228 22158 9240
rect 24394 9228 24400 9240
rect 22152 9200 24400 9228
rect 22152 9188 22158 9200
rect 24394 9188 24400 9200
rect 24452 9188 24458 9240
rect 24762 9188 24768 9240
rect 24820 9228 24826 9240
rect 31018 9228 31024 9240
rect 24820 9200 31024 9228
rect 24820 9188 24826 9200
rect 31018 9188 31024 9200
rect 31076 9188 31082 9240
rect 32214 9188 32220 9240
rect 32272 9228 32278 9240
rect 40954 9228 40960 9240
rect 32272 9200 40960 9228
rect 32272 9188 32278 9200
rect 40954 9188 40960 9200
rect 41012 9188 41018 9240
rect 20806 9160 20812 9172
rect 18064 9132 20812 9160
rect 18064 9104 18092 9132
rect 20806 9120 20812 9132
rect 20864 9120 20870 9172
rect 21008 9132 21312 9160
rect 12676 9064 17632 9092
rect 12676 9052 12682 9064
rect 18046 9052 18052 9104
rect 18104 9052 18110 9104
rect 18230 9052 18236 9104
rect 18288 9092 18294 9104
rect 21008 9092 21036 9132
rect 18288 9064 21036 9092
rect 21284 9092 21312 9132
rect 21726 9120 21732 9172
rect 21784 9160 21790 9172
rect 35894 9160 35900 9172
rect 21784 9132 35900 9160
rect 21784 9120 21790 9132
rect 35894 9120 35900 9132
rect 35952 9120 35958 9172
rect 37366 9120 37372 9172
rect 37424 9160 37430 9172
rect 43438 9160 43444 9172
rect 37424 9132 43444 9160
rect 37424 9120 37430 9132
rect 43438 9120 43444 9132
rect 43496 9120 43502 9172
rect 32766 9092 32772 9104
rect 21284 9064 32772 9092
rect 18288 9052 18294 9064
rect 32766 9052 32772 9064
rect 32824 9052 32830 9104
rect 35526 9052 35532 9104
rect 35584 9092 35590 9104
rect 35584 9064 42472 9092
rect 35584 9052 35590 9064
rect 13722 9024 13728 9036
rect 7116 8996 13728 9024
rect 7116 8832 7144 8996
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 16666 9024 16672 9036
rect 14016 8996 16672 9024
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 14016 8956 14044 8996
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 16942 8984 16948 9036
rect 17000 9024 17006 9036
rect 21082 9024 21088 9036
rect 17000 8996 21088 9024
rect 17000 8984 17006 8996
rect 21082 8984 21088 8996
rect 21140 8984 21146 9036
rect 21450 8984 21456 9036
rect 21508 9024 21514 9036
rect 24118 9024 24124 9036
rect 21508 8996 24124 9024
rect 21508 8984 21514 8996
rect 24118 8984 24124 8996
rect 24176 8984 24182 9036
rect 33962 8984 33968 9036
rect 34020 9024 34026 9036
rect 40678 9024 40684 9036
rect 34020 8996 40684 9024
rect 34020 8984 34026 8996
rect 40678 8984 40684 8996
rect 40736 8984 40742 9036
rect 10560 8928 14044 8956
rect 10560 8916 10566 8928
rect 14090 8916 14096 8968
rect 14148 8956 14154 8968
rect 23014 8956 23020 8968
rect 14148 8928 23020 8956
rect 14148 8916 14154 8928
rect 23014 8916 23020 8928
rect 23072 8916 23078 8968
rect 30282 8956 30288 8968
rect 24320 8928 30288 8956
rect 24320 8900 24348 8928
rect 30282 8916 30288 8928
rect 30340 8916 30346 8968
rect 33594 8916 33600 8968
rect 33652 8956 33658 8968
rect 38102 8956 38108 8968
rect 33652 8928 38108 8956
rect 33652 8916 33658 8928
rect 38102 8916 38108 8928
rect 38160 8916 38166 8968
rect 24026 8888 24032 8900
rect 9784 8860 24032 8888
rect 9784 8832 9812 8860
rect 24026 8848 24032 8860
rect 24084 8848 24090 8900
rect 24302 8848 24308 8900
rect 24360 8848 24366 8900
rect 27246 8848 27252 8900
rect 27304 8888 27310 8900
rect 30926 8888 30932 8900
rect 27304 8860 30932 8888
rect 27304 8848 27310 8860
rect 30926 8848 30932 8860
rect 30984 8848 30990 8900
rect 37182 8888 37188 8900
rect 31726 8860 37188 8888
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 7006 8820 7012 8832
rect 3384 8792 7012 8820
rect 3384 8780 3390 8792
rect 7006 8780 7012 8792
rect 7064 8780 7070 8832
rect 7098 8780 7104 8832
rect 7156 8780 7162 8832
rect 9766 8780 9772 8832
rect 9824 8780 9830 8832
rect 11514 8780 11520 8832
rect 11572 8820 11578 8832
rect 15102 8820 15108 8832
rect 11572 8792 15108 8820
rect 11572 8780 11578 8792
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 17034 8780 17040 8832
rect 17092 8820 17098 8832
rect 22094 8820 22100 8832
rect 17092 8792 22100 8820
rect 17092 8780 17098 8792
rect 22094 8780 22100 8792
rect 22152 8780 22158 8832
rect 22646 8780 22652 8832
rect 22704 8820 22710 8832
rect 31726 8820 31754 8860
rect 37182 8848 37188 8860
rect 37240 8848 37246 8900
rect 42444 8832 42472 9064
rect 22704 8792 31754 8820
rect 22704 8780 22710 8792
rect 31846 8780 31852 8832
rect 31904 8820 31910 8832
rect 37734 8820 37740 8832
rect 31904 8792 37740 8820
rect 31904 8780 31910 8792
rect 37734 8780 37740 8792
rect 37792 8780 37798 8832
rect 42426 8780 42432 8832
rect 42484 8780 42490 8832
rect 1104 8730 45976 8752
rect 1104 8678 12128 8730
rect 12180 8678 12192 8730
rect 12244 8678 12256 8730
rect 12308 8678 12320 8730
rect 12372 8678 12384 8730
rect 12436 8678 23306 8730
rect 23358 8678 23370 8730
rect 23422 8678 23434 8730
rect 23486 8678 23498 8730
rect 23550 8678 23562 8730
rect 23614 8678 34484 8730
rect 34536 8678 34548 8730
rect 34600 8678 34612 8730
rect 34664 8678 34676 8730
rect 34728 8678 34740 8730
rect 34792 8678 45662 8730
rect 45714 8678 45726 8730
rect 45778 8678 45790 8730
rect 45842 8678 45854 8730
rect 45906 8678 45918 8730
rect 45970 8678 45976 8730
rect 1104 8656 45976 8678
rect 1673 8619 1731 8625
rect 1673 8585 1685 8619
rect 1719 8616 1731 8619
rect 2498 8616 2504 8628
rect 1719 8588 2504 8616
rect 1719 8585 1731 8588
rect 1673 8579 1731 8585
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8616 2835 8619
rect 2866 8616 2872 8628
rect 2823 8588 2872 8616
rect 2823 8585 2835 8588
rect 2777 8579 2835 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 3145 8619 3203 8625
rect 3145 8585 3157 8619
rect 3191 8616 3203 8619
rect 3234 8616 3240 8628
rect 3191 8588 3240 8616
rect 3191 8585 3203 8588
rect 3145 8579 3203 8585
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 3513 8619 3571 8625
rect 3513 8585 3525 8619
rect 3559 8616 3571 8619
rect 3602 8616 3608 8628
rect 3559 8588 3608 8616
rect 3559 8585 3571 8588
rect 3513 8579 3571 8585
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 4338 8616 4344 8628
rect 4295 8588 4344 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4617 8619 4675 8625
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 5074 8616 5080 8628
rect 4663 8588 5080 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 5074 8576 5080 8588
rect 5132 8576 5138 8628
rect 5169 8619 5227 8625
rect 5169 8585 5181 8619
rect 5215 8616 5227 8619
rect 5442 8616 5448 8628
rect 5215 8588 5448 8616
rect 5215 8585 5227 8588
rect 5169 8579 5227 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 6089 8619 6147 8625
rect 6089 8585 6101 8619
rect 6135 8616 6147 8619
rect 6178 8616 6184 8628
rect 6135 8588 6184 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 6822 8576 6828 8628
rect 6880 8576 6886 8628
rect 7377 8619 7435 8625
rect 7377 8585 7389 8619
rect 7423 8616 7435 8619
rect 7650 8616 7656 8628
rect 7423 8588 7656 8616
rect 7423 8585 7435 8588
rect 7377 8579 7435 8585
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 8018 8616 8024 8628
rect 7791 8588 8024 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8616 8355 8619
rect 8386 8616 8392 8628
rect 8343 8588 8392 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 8665 8619 8723 8625
rect 8665 8585 8677 8619
rect 8711 8616 8723 8619
rect 8754 8616 8760 8628
rect 8711 8588 8760 8616
rect 8711 8585 8723 8588
rect 8665 8579 8723 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9217 8619 9275 8625
rect 9217 8585 9229 8619
rect 9263 8616 9275 8619
rect 9490 8616 9496 8628
rect 9263 8588 9496 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 9769 8619 9827 8625
rect 9769 8585 9781 8619
rect 9815 8616 9827 8619
rect 9858 8616 9864 8628
rect 9815 8588 9864 8616
rect 9815 8585 9827 8588
rect 9769 8579 9827 8585
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 10137 8619 10195 8625
rect 10137 8585 10149 8619
rect 10183 8616 10195 8619
rect 10594 8616 10600 8628
rect 10183 8588 10600 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 10689 8619 10747 8625
rect 10689 8585 10701 8619
rect 10735 8616 10747 8619
rect 10962 8616 10968 8628
rect 10735 8588 10968 8616
rect 10735 8585 10747 8588
rect 10689 8579 10747 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11241 8619 11299 8625
rect 11241 8585 11253 8619
rect 11287 8616 11299 8619
rect 11330 8616 11336 8628
rect 11287 8588 11336 8616
rect 11287 8585 11299 8588
rect 11241 8579 11299 8585
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 11793 8619 11851 8625
rect 11793 8585 11805 8619
rect 11839 8616 11851 8619
rect 11974 8616 11980 8628
rect 11839 8588 11980 8616
rect 11839 8585 11851 8588
rect 11793 8579 11851 8585
rect 11974 8576 11980 8588
rect 12032 8576 12038 8628
rect 12345 8619 12403 8625
rect 12345 8585 12357 8619
rect 12391 8616 12403 8619
rect 12434 8616 12440 8628
rect 12391 8588 12440 8616
rect 12391 8585 12403 8588
rect 12345 8579 12403 8585
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 12618 8616 12624 8628
rect 12544 8588 12624 8616
rect 2682 8508 2688 8560
rect 2740 8508 2746 8560
rect 3973 8551 4031 8557
rect 3973 8517 3985 8551
rect 4019 8548 4031 8551
rect 4062 8548 4068 8560
rect 4019 8520 4068 8548
rect 4019 8517 4031 8520
rect 3973 8511 4031 8517
rect 4062 8508 4068 8520
rect 4120 8508 4126 8560
rect 4893 8551 4951 8557
rect 4893 8517 4905 8551
rect 4939 8548 4951 8551
rect 4939 8520 10364 8548
rect 4939 8517 4951 8520
rect 4893 8511 4951 8517
rect 1486 8440 1492 8492
rect 1544 8440 1550 8492
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 2501 8483 2559 8489
rect 2501 8480 2513 8483
rect 2179 8452 2513 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 2501 8449 2513 8452
rect 2547 8480 2559 8483
rect 2700 8480 2728 8508
rect 2547 8452 2728 8480
rect 2547 8449 2559 8452
rect 2501 8443 2559 8449
rect 2958 8440 2964 8492
rect 3016 8440 3022 8492
rect 3326 8440 3332 8492
rect 3384 8440 3390 8492
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8449 4491 8483
rect 4433 8443 4491 8449
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 7098 8480 7104 8492
rect 6595 8452 7104 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 4448 8344 4476 8443
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8412 5687 8415
rect 5920 8412 5948 8443
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7190 8440 7196 8492
rect 7248 8440 7254 8492
rect 7558 8440 7564 8492
rect 7616 8440 7622 8492
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8480 8079 8483
rect 8294 8480 8300 8492
rect 8067 8452 8300 8480
rect 8067 8449 8079 8452
rect 8021 8443 8079 8449
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 8496 8412 8524 8443
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 9766 8480 9772 8492
rect 9539 8452 9772 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 9950 8440 9956 8492
rect 10008 8440 10014 8492
rect 10336 8480 10364 8520
rect 10410 8508 10416 8560
rect 10468 8508 10474 8560
rect 12544 8548 12572 8588
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 12897 8619 12955 8625
rect 12897 8585 12909 8619
rect 12943 8616 12955 8619
rect 13170 8616 13176 8628
rect 12943 8588 13176 8616
rect 12943 8585 12955 8588
rect 12897 8579 12955 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13265 8619 13323 8625
rect 13265 8585 13277 8619
rect 13311 8616 13323 8619
rect 13538 8616 13544 8628
rect 13311 8588 13544 8616
rect 13311 8585 13323 8588
rect 13265 8579 13323 8585
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 13817 8619 13875 8625
rect 13817 8585 13829 8619
rect 13863 8616 13875 8619
rect 13906 8616 13912 8628
rect 13863 8588 13912 8616
rect 13863 8585 13875 8588
rect 13817 8579 13875 8585
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 14369 8619 14427 8625
rect 14369 8585 14381 8619
rect 14415 8616 14427 8619
rect 14642 8616 14648 8628
rect 14415 8588 14648 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 14642 8576 14648 8588
rect 14700 8576 14706 8628
rect 14737 8619 14795 8625
rect 14737 8585 14749 8619
rect 14783 8616 14795 8619
rect 15010 8616 15016 8628
rect 14783 8588 15016 8616
rect 14783 8585 14795 8588
rect 14737 8579 14795 8585
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 15378 8616 15384 8628
rect 15335 8588 15384 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15841 8619 15899 8625
rect 15841 8585 15853 8619
rect 15887 8616 15899 8619
rect 16114 8616 16120 8628
rect 15887 8588 16120 8616
rect 15887 8585 15899 8588
rect 15841 8579 15899 8585
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16393 8619 16451 8625
rect 16393 8585 16405 8619
rect 16439 8616 16451 8619
rect 16482 8616 16488 8628
rect 16439 8588 16488 8616
rect 16439 8585 16451 8588
rect 16393 8579 16451 8585
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 16758 8576 16764 8628
rect 16816 8576 16822 8628
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 17129 8619 17187 8625
rect 17129 8616 17141 8619
rect 16908 8588 17141 8616
rect 16908 8576 16914 8588
rect 17129 8585 17141 8588
rect 17175 8585 17187 8619
rect 17129 8579 17187 8585
rect 17218 8576 17224 8628
rect 17276 8616 17282 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 17276 8588 17509 8616
rect 17276 8576 17282 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 17497 8579 17555 8585
rect 17586 8576 17592 8628
rect 17644 8616 17650 8628
rect 17865 8619 17923 8625
rect 17865 8616 17877 8619
rect 17644 8588 17877 8616
rect 17644 8576 17650 8588
rect 17865 8585 17877 8588
rect 17911 8585 17923 8619
rect 17865 8579 17923 8585
rect 17954 8576 17960 8628
rect 18012 8616 18018 8628
rect 18233 8619 18291 8625
rect 18233 8616 18245 8619
rect 18012 8588 18245 8616
rect 18012 8576 18018 8588
rect 18233 8585 18245 8588
rect 18279 8585 18291 8619
rect 18233 8579 18291 8585
rect 18690 8576 18696 8628
rect 18748 8616 18754 8628
rect 18969 8619 19027 8625
rect 18969 8616 18981 8619
rect 18748 8588 18981 8616
rect 18748 8576 18754 8588
rect 18969 8585 18981 8588
rect 19015 8585 19027 8619
rect 18969 8579 19027 8585
rect 19518 8576 19524 8628
rect 19576 8576 19582 8628
rect 20073 8619 20131 8625
rect 20073 8585 20085 8619
rect 20119 8585 20131 8619
rect 20073 8579 20131 8585
rect 16776 8548 16804 8576
rect 18506 8548 18512 8560
rect 10520 8520 12572 8548
rect 12636 8520 16804 8548
rect 17328 8520 18512 8548
rect 10520 8480 10548 8520
rect 10336 8452 10548 8480
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8480 11023 8483
rect 11514 8480 11520 8492
rect 11011 8452 11520 8480
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 11606 8440 11612 8492
rect 11664 8440 11670 8492
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8480 12127 8483
rect 12636 8480 12664 8520
rect 12115 8452 12664 8480
rect 12115 8449 12127 8452
rect 12069 8443 12127 8449
rect 12710 8440 12716 8492
rect 12768 8440 12774 8492
rect 13078 8440 13084 8492
rect 13136 8440 13142 8492
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8480 13599 8483
rect 14090 8480 14096 8492
rect 13587 8452 14096 8480
rect 13587 8449 13599 8452
rect 13541 8443 13599 8449
rect 14090 8440 14096 8452
rect 14148 8440 14154 8492
rect 14185 8483 14243 8489
rect 14185 8449 14197 8483
rect 14231 8480 14243 8483
rect 14458 8480 14464 8492
rect 14231 8452 14464 8480
rect 14231 8449 14243 8452
rect 14185 8443 14243 8449
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8480 14611 8483
rect 14918 8480 14924 8492
rect 14599 8452 14924 8480
rect 14599 8449 14611 8452
rect 14553 8443 14611 8449
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8480 15071 8483
rect 15562 8480 15568 8492
rect 15059 8452 15568 8480
rect 15059 8449 15071 8452
rect 15013 8443 15071 8449
rect 15562 8440 15568 8452
rect 15620 8440 15626 8492
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8480 15715 8483
rect 16022 8480 16028 8492
rect 15703 8452 16028 8480
rect 15703 8449 15715 8452
rect 15657 8443 15715 8449
rect 16022 8440 16028 8452
rect 16080 8440 16086 8492
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8480 16175 8483
rect 16850 8480 16856 8492
rect 16163 8452 16856 8480
rect 16163 8449 16175 8452
rect 16117 8443 16175 8449
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 16942 8440 16948 8492
rect 17000 8440 17006 8492
rect 17328 8489 17356 8520
rect 18506 8508 18512 8520
rect 18564 8508 18570 8560
rect 19334 8508 19340 8560
rect 19392 8548 19398 8560
rect 20088 8548 20116 8579
rect 21818 8576 21824 8628
rect 21876 8616 21882 8628
rect 22189 8619 22247 8625
rect 22189 8616 22201 8619
rect 21876 8588 22201 8616
rect 21876 8576 21882 8588
rect 22189 8585 22201 8588
rect 22235 8585 22247 8619
rect 22189 8579 22247 8585
rect 22462 8576 22468 8628
rect 22520 8576 22526 8628
rect 23014 8576 23020 8628
rect 23072 8576 23078 8628
rect 23934 8616 23940 8628
rect 23400 8588 23940 8616
rect 21266 8548 21272 8560
rect 19392 8520 20116 8548
rect 20824 8520 21272 8548
rect 19392 8508 19398 8520
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 17586 8440 17592 8492
rect 17644 8480 17650 8492
rect 17681 8483 17739 8489
rect 17681 8480 17693 8483
rect 17644 8452 17693 8480
rect 17644 8440 17650 8452
rect 17681 8449 17693 8452
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 10502 8412 10508 8424
rect 5675 8384 8340 8412
rect 8496 8384 10508 8412
rect 5675 8381 5687 8384
rect 5629 8375 5687 8381
rect 8202 8344 8208 8356
rect 4448 8316 8208 8344
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 8312 8276 8340 8384
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 10612 8384 17264 8412
rect 8386 8304 8392 8356
rect 8444 8344 8450 8356
rect 10612 8344 10640 8384
rect 17034 8344 17040 8356
rect 8444 8316 10640 8344
rect 10704 8316 17040 8344
rect 8444 8304 8450 8316
rect 10704 8276 10732 8316
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 17236 8344 17264 8384
rect 17494 8372 17500 8424
rect 17552 8412 17558 8424
rect 18156 8412 18184 8443
rect 18782 8440 18788 8492
rect 18840 8440 18846 8492
rect 19426 8440 19432 8492
rect 19484 8440 19490 8492
rect 19978 8440 19984 8492
rect 20036 8440 20042 8492
rect 20824 8489 20852 8520
rect 21266 8508 21272 8520
rect 21324 8508 21330 8560
rect 22002 8548 22008 8560
rect 21376 8520 22008 8548
rect 21376 8489 21404 8520
rect 22002 8508 22008 8520
rect 22060 8508 22066 8560
rect 22738 8548 22744 8560
rect 22112 8520 22744 8548
rect 22112 8489 22140 8520
rect 22738 8508 22744 8520
rect 22796 8508 22802 8560
rect 23290 8548 23296 8560
rect 22940 8520 23296 8548
rect 20809 8483 20867 8489
rect 20809 8449 20821 8483
rect 20855 8449 20867 8483
rect 20809 8443 20867 8449
rect 21085 8483 21143 8489
rect 21085 8449 21097 8483
rect 21131 8449 21143 8483
rect 21085 8443 21143 8449
rect 21361 8483 21419 8489
rect 21361 8449 21373 8483
rect 21407 8449 21419 8483
rect 21361 8443 21419 8449
rect 21637 8483 21695 8489
rect 21637 8449 21649 8483
rect 21683 8449 21695 8483
rect 21637 8443 21695 8449
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8449 22155 8483
rect 22097 8443 22155 8449
rect 22373 8483 22431 8489
rect 22373 8449 22385 8483
rect 22419 8449 22431 8483
rect 22373 8443 22431 8449
rect 17552 8384 18184 8412
rect 17552 8372 17558 8384
rect 19334 8372 19340 8424
rect 19392 8372 19398 8424
rect 21100 8412 21128 8443
rect 21450 8412 21456 8424
rect 21100 8384 21456 8412
rect 21450 8372 21456 8384
rect 21508 8372 21514 8424
rect 21652 8412 21680 8443
rect 22186 8412 22192 8424
rect 21652 8384 22192 8412
rect 22186 8372 22192 8384
rect 22244 8372 22250 8424
rect 22388 8412 22416 8443
rect 22646 8440 22652 8492
rect 22704 8440 22710 8492
rect 22940 8489 22968 8520
rect 23290 8508 23296 8520
rect 23348 8508 23354 8560
rect 22925 8483 22983 8489
rect 22925 8449 22937 8483
rect 22971 8449 22983 8483
rect 22925 8443 22983 8449
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8480 23259 8483
rect 23400 8480 23428 8588
rect 23934 8576 23940 8588
rect 23992 8576 23998 8628
rect 24026 8576 24032 8628
rect 24084 8576 24090 8628
rect 27246 8616 27252 8628
rect 24136 8588 27252 8616
rect 23247 8452 23428 8480
rect 23247 8449 23259 8452
rect 23201 8443 23259 8449
rect 23474 8440 23480 8492
rect 23532 8440 23538 8492
rect 23569 8483 23627 8489
rect 23569 8449 23581 8483
rect 23615 8449 23627 8483
rect 23569 8443 23627 8449
rect 23845 8483 23903 8489
rect 23845 8449 23857 8483
rect 23891 8480 23903 8483
rect 24136 8480 24164 8588
rect 27246 8576 27252 8588
rect 27304 8576 27310 8628
rect 27338 8576 27344 8628
rect 27396 8616 27402 8628
rect 27985 8619 28043 8625
rect 27985 8616 27997 8619
rect 27396 8588 27997 8616
rect 27396 8576 27402 8588
rect 27985 8585 27997 8588
rect 28031 8585 28043 8619
rect 27985 8579 28043 8585
rect 30193 8619 30251 8625
rect 30193 8585 30205 8619
rect 30239 8585 30251 8619
rect 30193 8579 30251 8585
rect 25130 8508 25136 8560
rect 25188 8548 25194 8560
rect 30208 8548 30236 8579
rect 30282 8576 30288 8628
rect 30340 8576 30346 8628
rect 30926 8576 30932 8628
rect 30984 8576 30990 8628
rect 31018 8576 31024 8628
rect 31076 8616 31082 8628
rect 32309 8619 32367 8625
rect 32309 8616 32321 8619
rect 31076 8588 32321 8616
rect 31076 8576 31082 8588
rect 32309 8585 32321 8588
rect 32355 8585 32367 8619
rect 32309 8579 32367 8585
rect 32585 8619 32643 8625
rect 32585 8585 32597 8619
rect 32631 8585 32643 8619
rect 32585 8579 32643 8585
rect 25188 8520 30236 8548
rect 30300 8548 30328 8576
rect 32600 8548 32628 8579
rect 32766 8576 32772 8628
rect 32824 8616 32830 8628
rect 34425 8619 34483 8625
rect 34425 8616 34437 8619
rect 32824 8588 34437 8616
rect 32824 8576 32830 8588
rect 34425 8585 34437 8588
rect 34471 8585 34483 8619
rect 34425 8579 34483 8585
rect 34885 8619 34943 8625
rect 34885 8585 34897 8619
rect 34931 8585 34943 8619
rect 34885 8579 34943 8585
rect 30300 8520 32628 8548
rect 25188 8508 25194 8520
rect 32858 8508 32864 8560
rect 32916 8548 32922 8560
rect 34900 8548 34928 8579
rect 35158 8576 35164 8628
rect 35216 8576 35222 8628
rect 36265 8619 36323 8625
rect 36265 8616 36277 8619
rect 35268 8588 36277 8616
rect 32916 8520 34928 8548
rect 32916 8508 32922 8520
rect 23891 8452 24164 8480
rect 23891 8449 23903 8452
rect 23845 8443 23903 8449
rect 23106 8412 23112 8424
rect 22388 8384 23112 8412
rect 23106 8372 23112 8384
rect 23164 8372 23170 8424
rect 23584 8412 23612 8443
rect 24210 8440 24216 8492
rect 24268 8480 24274 8492
rect 24581 8483 24639 8489
rect 24581 8480 24593 8483
rect 24268 8452 24593 8480
rect 24268 8440 24274 8452
rect 24581 8449 24593 8452
rect 24627 8449 24639 8483
rect 24581 8443 24639 8449
rect 24854 8440 24860 8492
rect 24912 8440 24918 8492
rect 24946 8440 24952 8492
rect 25004 8480 25010 8492
rect 25225 8483 25283 8489
rect 25225 8480 25237 8483
rect 25004 8452 25237 8480
rect 25004 8440 25010 8452
rect 25225 8449 25237 8452
rect 25271 8449 25283 8483
rect 25225 8443 25283 8449
rect 25314 8440 25320 8492
rect 25372 8480 25378 8492
rect 25593 8483 25651 8489
rect 25593 8480 25605 8483
rect 25372 8452 25605 8480
rect 25372 8440 25378 8452
rect 25593 8449 25605 8452
rect 25639 8449 25651 8483
rect 25593 8443 25651 8449
rect 25682 8440 25688 8492
rect 25740 8480 25746 8492
rect 25961 8483 26019 8489
rect 25961 8480 25973 8483
rect 25740 8452 25973 8480
rect 25740 8440 25746 8452
rect 25961 8449 25973 8452
rect 26007 8449 26019 8483
rect 25961 8443 26019 8449
rect 26050 8440 26056 8492
rect 26108 8480 26114 8492
rect 26329 8483 26387 8489
rect 26329 8480 26341 8483
rect 26108 8452 26341 8480
rect 26108 8440 26114 8452
rect 26329 8449 26341 8452
rect 26375 8449 26387 8483
rect 26329 8443 26387 8449
rect 26418 8440 26424 8492
rect 26476 8480 26482 8492
rect 26697 8483 26755 8489
rect 26697 8480 26709 8483
rect 26476 8452 26709 8480
rect 26476 8440 26482 8452
rect 26697 8449 26709 8452
rect 26743 8449 26755 8483
rect 26697 8443 26755 8449
rect 26786 8440 26792 8492
rect 26844 8480 26850 8492
rect 27157 8483 27215 8489
rect 27157 8480 27169 8483
rect 26844 8452 27169 8480
rect 26844 8440 26850 8452
rect 27157 8449 27169 8452
rect 27203 8449 27215 8483
rect 27157 8443 27215 8449
rect 27430 8440 27436 8492
rect 27488 8440 27494 8492
rect 27522 8440 27528 8492
rect 27580 8480 27586 8492
rect 27801 8483 27859 8489
rect 27801 8480 27813 8483
rect 27580 8452 27813 8480
rect 27580 8440 27586 8452
rect 27801 8449 27813 8452
rect 27847 8449 27859 8483
rect 27801 8443 27859 8449
rect 27890 8440 27896 8492
rect 27948 8480 27954 8492
rect 28169 8483 28227 8489
rect 28169 8480 28181 8483
rect 27948 8452 28181 8480
rect 27948 8440 27954 8452
rect 28169 8449 28181 8452
rect 28215 8449 28227 8483
rect 28169 8443 28227 8449
rect 28258 8440 28264 8492
rect 28316 8480 28322 8492
rect 28537 8483 28595 8489
rect 28537 8480 28549 8483
rect 28316 8452 28549 8480
rect 28316 8440 28322 8452
rect 28537 8449 28549 8452
rect 28583 8449 28595 8483
rect 28537 8443 28595 8449
rect 28626 8440 28632 8492
rect 28684 8480 28690 8492
rect 28905 8483 28963 8489
rect 28905 8480 28917 8483
rect 28684 8452 28917 8480
rect 28684 8440 28690 8452
rect 28905 8449 28917 8452
rect 28951 8449 28963 8483
rect 28905 8443 28963 8449
rect 28994 8440 29000 8492
rect 29052 8480 29058 8492
rect 29273 8483 29331 8489
rect 29273 8480 29285 8483
rect 29052 8452 29285 8480
rect 29052 8440 29058 8452
rect 29273 8449 29285 8452
rect 29319 8449 29331 8483
rect 29273 8443 29331 8449
rect 29362 8440 29368 8492
rect 29420 8480 29426 8492
rect 29733 8483 29791 8489
rect 29733 8480 29745 8483
rect 29420 8452 29745 8480
rect 29420 8440 29426 8452
rect 29733 8449 29745 8452
rect 29779 8449 29791 8483
rect 29733 8443 29791 8449
rect 30006 8440 30012 8492
rect 30064 8440 30070 8492
rect 30098 8440 30104 8492
rect 30156 8480 30162 8492
rect 30377 8483 30435 8489
rect 30377 8480 30389 8483
rect 30156 8452 30389 8480
rect 30156 8440 30162 8452
rect 30377 8449 30389 8452
rect 30423 8449 30435 8483
rect 30377 8443 30435 8449
rect 30466 8440 30472 8492
rect 30524 8480 30530 8492
rect 30745 8483 30803 8489
rect 30745 8480 30757 8483
rect 30524 8452 30757 8480
rect 30524 8440 30530 8452
rect 30745 8449 30757 8452
rect 30791 8449 30803 8483
rect 30745 8443 30803 8449
rect 30834 8440 30840 8492
rect 30892 8480 30898 8492
rect 31113 8483 31171 8489
rect 31113 8480 31125 8483
rect 30892 8452 31125 8480
rect 30892 8440 30898 8452
rect 31113 8449 31125 8452
rect 31159 8449 31171 8483
rect 31113 8443 31171 8449
rect 31202 8440 31208 8492
rect 31260 8480 31266 8492
rect 31481 8483 31539 8489
rect 31481 8480 31493 8483
rect 31260 8452 31493 8480
rect 31260 8440 31266 8452
rect 31481 8449 31493 8452
rect 31527 8449 31539 8483
rect 31481 8443 31539 8449
rect 31662 8440 31668 8492
rect 31720 8440 31726 8492
rect 32122 8440 32128 8492
rect 32180 8440 32186 8492
rect 32398 8440 32404 8492
rect 32456 8440 32462 8492
rect 32766 8440 32772 8492
rect 32824 8440 32830 8492
rect 33042 8440 33048 8492
rect 33100 8480 33106 8492
rect 33137 8483 33195 8489
rect 33137 8480 33149 8483
rect 33100 8452 33149 8480
rect 33100 8440 33106 8452
rect 33137 8449 33149 8452
rect 33183 8449 33195 8483
rect 33137 8443 33195 8449
rect 33502 8440 33508 8492
rect 33560 8440 33566 8492
rect 33870 8440 33876 8492
rect 33928 8440 33934 8492
rect 34238 8440 34244 8492
rect 34296 8440 34302 8492
rect 34330 8440 34336 8492
rect 34388 8480 34394 8492
rect 34701 8483 34759 8489
rect 34701 8480 34713 8483
rect 34388 8452 34713 8480
rect 34388 8440 34394 8452
rect 34701 8449 34713 8452
rect 34747 8449 34759 8483
rect 34701 8443 34759 8449
rect 34974 8440 34980 8492
rect 35032 8440 35038 8492
rect 23584 8384 24440 8412
rect 19352 8344 19380 8372
rect 17236 8316 19380 8344
rect 19610 8304 19616 8356
rect 19668 8344 19674 8356
rect 21913 8347 21971 8353
rect 19668 8316 21588 8344
rect 19668 8304 19674 8316
rect 8312 8248 10732 8276
rect 14274 8236 14280 8288
rect 14332 8276 14338 8288
rect 18690 8276 18696 8288
rect 14332 8248 18696 8276
rect 14332 8236 14338 8248
rect 18690 8236 18696 8248
rect 18748 8236 18754 8288
rect 19058 8236 19064 8288
rect 19116 8276 19122 8288
rect 19886 8276 19892 8288
rect 19116 8248 19892 8276
rect 19116 8236 19122 8248
rect 19886 8236 19892 8248
rect 19944 8236 19950 8288
rect 20622 8236 20628 8288
rect 20680 8236 20686 8288
rect 20898 8236 20904 8288
rect 20956 8236 20962 8288
rect 21174 8236 21180 8288
rect 21232 8236 21238 8288
rect 21450 8236 21456 8288
rect 21508 8236 21514 8288
rect 21560 8276 21588 8316
rect 21913 8313 21925 8347
rect 21959 8344 21971 8347
rect 22278 8344 22284 8356
rect 21959 8316 22284 8344
rect 21959 8313 21971 8316
rect 21913 8307 21971 8313
rect 22278 8304 22284 8316
rect 22336 8304 22342 8356
rect 23750 8304 23756 8356
rect 23808 8304 23814 8356
rect 24302 8344 24308 8356
rect 23860 8316 24308 8344
rect 22370 8276 22376 8288
rect 21560 8248 22376 8276
rect 22370 8236 22376 8248
rect 22428 8236 22434 8288
rect 22738 8236 22744 8288
rect 22796 8236 22802 8288
rect 23014 8236 23020 8288
rect 23072 8276 23078 8288
rect 23293 8279 23351 8285
rect 23293 8276 23305 8279
rect 23072 8248 23305 8276
rect 23072 8236 23078 8248
rect 23293 8245 23305 8248
rect 23339 8245 23351 8279
rect 23293 8239 23351 8245
rect 23382 8236 23388 8288
rect 23440 8276 23446 8288
rect 23860 8276 23888 8316
rect 24302 8304 24308 8316
rect 24360 8304 24366 8356
rect 24412 8353 24440 8384
rect 24486 8372 24492 8424
rect 24544 8412 24550 8424
rect 24544 8384 30604 8412
rect 24544 8372 24550 8384
rect 24397 8347 24455 8353
rect 24397 8313 24409 8347
rect 24443 8313 24455 8347
rect 24762 8344 24768 8356
rect 24397 8307 24455 8313
rect 24596 8316 24768 8344
rect 23440 8248 23888 8276
rect 23440 8236 23446 8248
rect 23934 8236 23940 8288
rect 23992 8276 23998 8288
rect 24596 8276 24624 8316
rect 24762 8304 24768 8316
rect 24820 8304 24826 8356
rect 26050 8304 26056 8356
rect 26108 8344 26114 8356
rect 26513 8347 26571 8353
rect 26513 8344 26525 8347
rect 26108 8316 26525 8344
rect 26108 8304 26114 8316
rect 26513 8313 26525 8316
rect 26559 8313 26571 8347
rect 26513 8307 26571 8313
rect 26786 8304 26792 8356
rect 26844 8344 26850 8356
rect 26844 8316 27108 8344
rect 26844 8304 26850 8316
rect 23992 8248 24624 8276
rect 23992 8236 23998 8248
rect 24670 8236 24676 8288
rect 24728 8236 24734 8288
rect 25038 8236 25044 8288
rect 25096 8236 25102 8288
rect 25406 8236 25412 8288
rect 25464 8236 25470 8288
rect 25590 8236 25596 8288
rect 25648 8276 25654 8288
rect 25777 8279 25835 8285
rect 25777 8276 25789 8279
rect 25648 8248 25789 8276
rect 25648 8236 25654 8248
rect 25777 8245 25789 8248
rect 25823 8245 25835 8279
rect 25777 8239 25835 8245
rect 25866 8236 25872 8288
rect 25924 8276 25930 8288
rect 26145 8279 26203 8285
rect 26145 8276 26157 8279
rect 25924 8248 26157 8276
rect 25924 8236 25930 8248
rect 26145 8245 26157 8248
rect 26191 8245 26203 8279
rect 26145 8239 26203 8245
rect 26418 8236 26424 8288
rect 26476 8276 26482 8288
rect 26973 8279 27031 8285
rect 26973 8276 26985 8279
rect 26476 8248 26985 8276
rect 26476 8236 26482 8248
rect 26973 8245 26985 8248
rect 27019 8245 27031 8279
rect 27080 8276 27108 8316
rect 27154 8304 27160 8356
rect 27212 8344 27218 8356
rect 30576 8353 30604 8384
rect 31754 8372 31760 8424
rect 31812 8412 31818 8424
rect 35268 8412 35296 8588
rect 36265 8585 36277 8588
rect 36311 8585 36323 8619
rect 36265 8579 36323 8585
rect 37001 8619 37059 8625
rect 37001 8585 37013 8619
rect 37047 8585 37059 8619
rect 37001 8579 37059 8585
rect 37016 8548 37044 8579
rect 37182 8576 37188 8628
rect 37240 8616 37246 8628
rect 37461 8619 37519 8625
rect 37461 8616 37473 8619
rect 37240 8588 37473 8616
rect 37240 8576 37246 8588
rect 37461 8585 37473 8588
rect 37507 8585 37519 8619
rect 37461 8579 37519 8585
rect 37734 8576 37740 8628
rect 37792 8576 37798 8628
rect 38102 8576 38108 8628
rect 38160 8576 38166 8628
rect 38838 8576 38844 8628
rect 38896 8576 38902 8628
rect 38930 8576 38936 8628
rect 38988 8616 38994 8628
rect 39209 8619 39267 8625
rect 39209 8616 39221 8619
rect 38988 8588 39221 8616
rect 38988 8576 38994 8588
rect 39209 8585 39221 8588
rect 39255 8585 39267 8619
rect 39209 8579 39267 8585
rect 39298 8576 39304 8628
rect 39356 8616 39362 8628
rect 39577 8619 39635 8625
rect 39577 8616 39589 8619
rect 39356 8588 39589 8616
rect 39356 8576 39362 8588
rect 39577 8585 39589 8588
rect 39623 8585 39635 8619
rect 39577 8579 39635 8585
rect 39666 8576 39672 8628
rect 39724 8616 39730 8628
rect 40037 8619 40095 8625
rect 40037 8616 40049 8619
rect 39724 8588 40049 8616
rect 39724 8576 39730 8588
rect 40037 8585 40049 8588
rect 40083 8585 40095 8619
rect 40037 8579 40095 8585
rect 40126 8576 40132 8628
rect 40184 8616 40190 8628
rect 40589 8619 40647 8625
rect 40589 8616 40601 8619
rect 40184 8588 40601 8616
rect 40184 8576 40190 8588
rect 40589 8585 40601 8588
rect 40635 8585 40647 8619
rect 40589 8579 40647 8585
rect 40678 8576 40684 8628
rect 40736 8576 40742 8628
rect 41138 8576 41144 8628
rect 41196 8616 41202 8628
rect 41509 8619 41567 8625
rect 41509 8616 41521 8619
rect 41196 8588 41521 8616
rect 41196 8576 41202 8588
rect 41509 8585 41521 8588
rect 41555 8585 41567 8619
rect 41509 8579 41567 8585
rect 41874 8576 41880 8628
rect 41932 8616 41938 8628
rect 42613 8619 42671 8625
rect 42613 8616 42625 8619
rect 41932 8588 42625 8616
rect 41932 8576 41938 8588
rect 42613 8585 42625 8588
rect 42659 8585 42671 8619
rect 42613 8579 42671 8585
rect 42981 8619 43039 8625
rect 42981 8585 42993 8619
rect 43027 8585 43039 8619
rect 42981 8579 43039 8585
rect 35636 8520 37044 8548
rect 38120 8548 38148 8576
rect 40497 8551 40555 8557
rect 40497 8548 40509 8551
rect 38120 8520 40509 8548
rect 35342 8440 35348 8492
rect 35400 8440 35406 8492
rect 31812 8384 35296 8412
rect 31812 8372 31818 8384
rect 27617 8347 27675 8353
rect 27617 8344 27629 8347
rect 27212 8316 27629 8344
rect 27212 8304 27218 8316
rect 27617 8313 27629 8316
rect 27663 8313 27675 8347
rect 30561 8347 30619 8353
rect 27617 8307 27675 8313
rect 27724 8316 30512 8344
rect 27249 8279 27307 8285
rect 27249 8276 27261 8279
rect 27080 8248 27261 8276
rect 26973 8239 27031 8245
rect 27249 8245 27261 8248
rect 27295 8245 27307 8279
rect 27249 8239 27307 8245
rect 27522 8236 27528 8288
rect 27580 8276 27586 8288
rect 27724 8276 27752 8316
rect 27580 8248 27752 8276
rect 27580 8236 27586 8248
rect 27890 8236 27896 8288
rect 27948 8276 27954 8288
rect 28353 8279 28411 8285
rect 28353 8276 28365 8279
rect 27948 8248 28365 8276
rect 27948 8236 27954 8248
rect 28353 8245 28365 8248
rect 28399 8245 28411 8279
rect 28353 8239 28411 8245
rect 28718 8236 28724 8288
rect 28776 8236 28782 8288
rect 29089 8279 29147 8285
rect 29089 8245 29101 8279
rect 29135 8276 29147 8279
rect 29270 8276 29276 8288
rect 29135 8248 29276 8276
rect 29135 8245 29147 8248
rect 29089 8239 29147 8245
rect 29270 8236 29276 8248
rect 29328 8236 29334 8288
rect 29546 8236 29552 8288
rect 29604 8236 29610 8288
rect 29822 8236 29828 8288
rect 29880 8236 29886 8288
rect 30484 8276 30512 8316
rect 30561 8313 30573 8347
rect 30607 8313 30619 8347
rect 30561 8307 30619 8313
rect 30650 8304 30656 8356
rect 30708 8344 30714 8356
rect 31849 8347 31907 8353
rect 31849 8344 31861 8347
rect 30708 8316 31861 8344
rect 30708 8304 30714 8316
rect 31849 8313 31861 8316
rect 31895 8313 31907 8347
rect 31849 8307 31907 8313
rect 31938 8304 31944 8356
rect 31996 8344 32002 8356
rect 34057 8347 34115 8353
rect 34057 8344 34069 8347
rect 31996 8316 34069 8344
rect 31996 8304 32002 8316
rect 34057 8313 34069 8316
rect 34103 8313 34115 8347
rect 34057 8307 34115 8313
rect 34146 8304 34152 8356
rect 34204 8344 34210 8356
rect 35529 8347 35587 8353
rect 35529 8344 35541 8347
rect 34204 8316 35541 8344
rect 34204 8304 34210 8316
rect 35529 8313 35541 8316
rect 35575 8313 35587 8347
rect 35529 8307 35587 8313
rect 31297 8279 31355 8285
rect 31297 8276 31309 8279
rect 30484 8248 31309 8276
rect 31297 8245 31309 8248
rect 31343 8245 31355 8279
rect 31297 8239 31355 8245
rect 32950 8236 32956 8288
rect 33008 8236 33014 8288
rect 33318 8236 33324 8288
rect 33376 8236 33382 8288
rect 33686 8236 33692 8288
rect 33744 8236 33750 8288
rect 33778 8236 33784 8288
rect 33836 8276 33842 8288
rect 35636 8276 35664 8520
rect 40497 8517 40509 8520
rect 40543 8517 40555 8551
rect 40696 8548 40724 8576
rect 41417 8551 41475 8557
rect 41417 8548 41429 8551
rect 40696 8520 41429 8548
rect 40497 8511 40555 8517
rect 41417 8517 41429 8520
rect 41463 8517 41475 8551
rect 41417 8511 41475 8517
rect 42242 8508 42248 8560
rect 42300 8548 42306 8560
rect 42996 8548 43024 8579
rect 43714 8576 43720 8628
rect 43772 8616 43778 8628
rect 44453 8619 44511 8625
rect 44453 8616 44465 8619
rect 43772 8588 44465 8616
rect 43772 8576 43778 8588
rect 44453 8585 44465 8588
rect 44499 8585 44511 8619
rect 44453 8579 44511 8585
rect 44818 8576 44824 8628
rect 44876 8616 44882 8628
rect 45189 8619 45247 8625
rect 45189 8616 45201 8619
rect 44876 8588 45201 8616
rect 44876 8576 44882 8588
rect 45189 8585 45201 8588
rect 45235 8585 45247 8619
rect 45189 8579 45247 8585
rect 42300 8520 43024 8548
rect 43364 8520 44128 8548
rect 42300 8508 42306 8520
rect 35710 8440 35716 8492
rect 35768 8440 35774 8492
rect 35894 8440 35900 8492
rect 35952 8440 35958 8492
rect 36078 8440 36084 8492
rect 36136 8440 36142 8492
rect 36446 8440 36452 8492
rect 36504 8440 36510 8492
rect 36814 8440 36820 8492
rect 36872 8440 36878 8492
rect 37090 8440 37096 8492
rect 37148 8480 37154 8492
rect 37277 8483 37335 8489
rect 37277 8480 37289 8483
rect 37148 8452 37289 8480
rect 37148 8440 37154 8452
rect 37277 8449 37289 8452
rect 37323 8449 37335 8483
rect 37277 8443 37335 8449
rect 37550 8440 37556 8492
rect 37608 8440 37614 8492
rect 37918 8440 37924 8492
rect 37976 8440 37982 8492
rect 38286 8440 38292 8492
rect 38344 8440 38350 8492
rect 38562 8440 38568 8492
rect 38620 8480 38626 8492
rect 38657 8483 38715 8489
rect 38657 8480 38669 8483
rect 38620 8452 38669 8480
rect 38620 8440 38626 8452
rect 38657 8449 38669 8452
rect 38703 8449 38715 8483
rect 38657 8443 38715 8449
rect 39025 8483 39083 8489
rect 39025 8449 39037 8483
rect 39071 8449 39083 8483
rect 39025 8443 39083 8449
rect 35912 8353 35940 8440
rect 36004 8384 38240 8412
rect 35897 8347 35955 8353
rect 35897 8313 35909 8347
rect 35943 8313 35955 8347
rect 35897 8307 35955 8313
rect 33836 8248 35664 8276
rect 33836 8236 33842 8248
rect 35802 8236 35808 8288
rect 35860 8276 35866 8288
rect 36004 8276 36032 8384
rect 36630 8304 36636 8356
rect 36688 8304 36694 8356
rect 38102 8304 38108 8356
rect 38160 8304 38166 8356
rect 38212 8344 38240 8384
rect 38378 8372 38384 8424
rect 38436 8412 38442 8424
rect 39040 8412 39068 8443
rect 39390 8440 39396 8492
rect 39448 8440 39454 8492
rect 39942 8440 39948 8492
rect 40000 8440 40006 8492
rect 40954 8440 40960 8492
rect 41012 8440 41018 8492
rect 41874 8440 41880 8492
rect 41932 8440 41938 8492
rect 42426 8440 42432 8492
rect 42484 8440 42490 8492
rect 42889 8483 42947 8489
rect 42889 8449 42901 8483
rect 42935 8449 42947 8483
rect 42889 8443 42947 8449
rect 42904 8412 42932 8443
rect 42978 8440 42984 8492
rect 43036 8480 43042 8492
rect 43364 8480 43392 8520
rect 43036 8452 43392 8480
rect 43036 8440 43042 8452
rect 43438 8440 43444 8492
rect 43496 8440 43502 8492
rect 43901 8483 43959 8489
rect 43901 8449 43913 8483
rect 43947 8449 43959 8483
rect 43901 8443 43959 8449
rect 38436 8384 39068 8412
rect 39132 8384 42932 8412
rect 38436 8372 38442 8384
rect 38212 8316 38424 8344
rect 35860 8248 36032 8276
rect 38396 8276 38424 8316
rect 38470 8304 38476 8356
rect 38528 8304 38534 8356
rect 39132 8344 39160 8384
rect 43070 8372 43076 8424
rect 43128 8412 43134 8424
rect 43916 8412 43944 8443
rect 43128 8384 43944 8412
rect 43128 8372 43134 8384
rect 38580 8316 39160 8344
rect 38580 8276 38608 8316
rect 40402 8304 40408 8356
rect 40460 8344 40466 8356
rect 41141 8347 41199 8353
rect 41141 8344 41153 8347
rect 40460 8316 41153 8344
rect 40460 8304 40466 8316
rect 41141 8313 41153 8316
rect 41187 8313 41199 8347
rect 41141 8307 41199 8313
rect 41506 8304 41512 8356
rect 41564 8344 41570 8356
rect 42061 8347 42119 8353
rect 42061 8344 42073 8347
rect 41564 8316 42073 8344
rect 41564 8304 41570 8316
rect 42061 8313 42073 8316
rect 42107 8313 42119 8347
rect 42061 8307 42119 8313
rect 42610 8304 42616 8356
rect 42668 8344 42674 8356
rect 44100 8353 44128 8520
rect 44358 8440 44364 8492
rect 44416 8440 44422 8492
rect 45094 8440 45100 8492
rect 45152 8440 45158 8492
rect 43625 8347 43683 8353
rect 43625 8344 43637 8347
rect 42668 8316 43637 8344
rect 42668 8304 42674 8316
rect 43625 8313 43637 8316
rect 43671 8313 43683 8347
rect 43625 8307 43683 8313
rect 44085 8347 44143 8353
rect 44085 8313 44097 8347
rect 44131 8313 44143 8347
rect 44085 8307 44143 8313
rect 38396 8248 38608 8276
rect 35860 8236 35866 8248
rect 1104 8186 45816 8208
rect 1104 8134 6539 8186
rect 6591 8134 6603 8186
rect 6655 8134 6667 8186
rect 6719 8134 6731 8186
rect 6783 8134 6795 8186
rect 6847 8134 17717 8186
rect 17769 8134 17781 8186
rect 17833 8134 17845 8186
rect 17897 8134 17909 8186
rect 17961 8134 17973 8186
rect 18025 8134 28895 8186
rect 28947 8134 28959 8186
rect 29011 8134 29023 8186
rect 29075 8134 29087 8186
rect 29139 8134 29151 8186
rect 29203 8134 40073 8186
rect 40125 8134 40137 8186
rect 40189 8134 40201 8186
rect 40253 8134 40265 8186
rect 40317 8134 40329 8186
rect 40381 8134 45816 8186
rect 1104 8112 45816 8134
rect 658 8032 664 8084
rect 716 8072 722 8084
rect 1857 8075 1915 8081
rect 1857 8072 1869 8075
rect 716 8044 1869 8072
rect 716 8032 722 8044
rect 1857 8041 1869 8044
rect 1903 8041 1915 8075
rect 1857 8035 1915 8041
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2188 8044 2973 8072
rect 2188 8032 2194 8044
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 2961 8035 3019 8041
rect 4617 8075 4675 8081
rect 4617 8041 4629 8075
rect 4663 8072 4675 8075
rect 4706 8072 4712 8084
rect 4663 8044 4712 8072
rect 4663 8041 4675 8044
rect 4617 8035 4675 8041
rect 4706 8032 4712 8044
rect 4764 8032 4770 8084
rect 5721 8075 5779 8081
rect 5721 8041 5733 8075
rect 5767 8072 5779 8075
rect 5810 8072 5816 8084
rect 5767 8044 5816 8072
rect 5767 8041 5779 8044
rect 5721 8035 5779 8041
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 6638 8032 6644 8084
rect 6696 8032 6702 8084
rect 7193 8075 7251 8081
rect 7193 8041 7205 8075
rect 7239 8072 7251 8075
rect 7282 8072 7288 8084
rect 7239 8044 7288 8072
rect 7239 8041 7251 8044
rect 7193 8035 7251 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 9214 8032 9220 8084
rect 9272 8032 9278 8084
rect 10137 8075 10195 8081
rect 10137 8041 10149 8075
rect 10183 8072 10195 8075
rect 10226 8072 10232 8084
rect 10183 8044 10232 8072
rect 10183 8041 10195 8044
rect 10137 8035 10195 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 11790 8032 11796 8084
rect 11848 8032 11854 8084
rect 12618 8072 12624 8084
rect 12406 8044 12624 8072
rect 1394 7964 1400 8016
rect 1452 8004 1458 8016
rect 2501 8007 2559 8013
rect 2501 8004 2513 8007
rect 1452 7976 2513 8004
rect 1452 7964 1458 7976
rect 2501 7973 2513 7976
rect 2547 7973 2559 8007
rect 2501 7967 2559 7973
rect 4154 7964 4160 8016
rect 4212 7964 4218 8016
rect 12406 8004 12434 8044
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 12713 8075 12771 8081
rect 12713 8041 12725 8075
rect 12759 8072 12771 8075
rect 12802 8072 12808 8084
rect 12759 8044 12808 8072
rect 12759 8041 12771 8044
rect 12713 8035 12771 8041
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 14366 8032 14372 8084
rect 14424 8032 14430 8084
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 15746 8072 15752 8084
rect 15703 8044 15752 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 15746 8032 15752 8044
rect 15804 8032 15810 8084
rect 17586 8032 17592 8084
rect 17644 8072 17650 8084
rect 17865 8075 17923 8081
rect 17865 8072 17877 8075
rect 17644 8044 17877 8072
rect 17644 8032 17650 8044
rect 17865 8041 17877 8044
rect 17911 8041 17923 8075
rect 17865 8035 17923 8041
rect 17972 8044 18276 8072
rect 6564 7976 12434 8004
rect 1780 7908 6500 7936
rect 1780 7877 1808 7908
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 4338 7868 4344 7880
rect 2823 7840 4344 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4430 7828 4436 7880
rect 4488 7828 4494 7880
rect 2314 7760 2320 7812
rect 2372 7760 2378 7812
rect 3970 7760 3976 7812
rect 4028 7760 4034 7812
rect 5445 7803 5503 7809
rect 5445 7769 5457 7803
rect 5491 7769 5503 7803
rect 6472 7800 6500 7908
rect 6564 7877 6592 7976
rect 17972 7936 18000 8044
rect 18141 8007 18199 8013
rect 18141 7973 18153 8007
rect 18187 7973 18199 8007
rect 18248 8004 18276 8044
rect 18322 8032 18328 8084
rect 18380 8072 18386 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 18380 8044 18613 8072
rect 18380 8032 18386 8044
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 18601 8035 18659 8041
rect 18690 8032 18696 8084
rect 18748 8032 18754 8084
rect 19426 8032 19432 8084
rect 19484 8072 19490 8084
rect 19613 8075 19671 8081
rect 19613 8072 19625 8075
rect 19484 8044 19625 8072
rect 19484 8032 19490 8044
rect 19613 8041 19625 8044
rect 19659 8041 19671 8075
rect 19613 8035 19671 8041
rect 19702 8032 19708 8084
rect 19760 8072 19766 8084
rect 20993 8075 21051 8081
rect 20993 8072 21005 8075
rect 19760 8044 21005 8072
rect 19760 8032 19766 8044
rect 20993 8041 21005 8044
rect 21039 8041 21051 8075
rect 20993 8035 21051 8041
rect 21082 8032 21088 8084
rect 21140 8072 21146 8084
rect 21269 8075 21327 8081
rect 21269 8072 21281 8075
rect 21140 8044 21281 8072
rect 21140 8032 21146 8044
rect 21269 8041 21281 8044
rect 21315 8041 21327 8075
rect 21269 8035 21327 8041
rect 21358 8032 21364 8084
rect 21416 8072 21422 8084
rect 21821 8075 21879 8081
rect 21821 8072 21833 8075
rect 21416 8044 21833 8072
rect 21416 8032 21422 8044
rect 21821 8041 21833 8044
rect 21867 8041 21879 8075
rect 21821 8035 21879 8041
rect 22554 8032 22560 8084
rect 22612 8032 22618 8084
rect 22830 8032 22836 8084
rect 22888 8032 22894 8084
rect 22922 8032 22928 8084
rect 22980 8072 22986 8084
rect 23109 8075 23167 8081
rect 23109 8072 23121 8075
rect 22980 8044 23121 8072
rect 22980 8032 22986 8044
rect 23109 8041 23121 8044
rect 23155 8041 23167 8075
rect 23109 8035 23167 8041
rect 23658 8032 23664 8084
rect 23716 8072 23722 8084
rect 23937 8075 23995 8081
rect 23937 8072 23949 8075
rect 23716 8044 23949 8072
rect 23716 8032 23722 8044
rect 23937 8041 23949 8044
rect 23983 8041 23995 8075
rect 23937 8035 23995 8041
rect 24210 8032 24216 8084
rect 24268 8032 24274 8084
rect 24578 8032 24584 8084
rect 24636 8072 24642 8084
rect 24765 8075 24823 8081
rect 24765 8072 24777 8075
rect 24636 8044 24777 8072
rect 24636 8032 24642 8044
rect 24765 8041 24777 8044
rect 24811 8041 24823 8075
rect 24765 8035 24823 8041
rect 25130 8032 25136 8084
rect 25188 8032 25194 8084
rect 25406 8032 25412 8084
rect 25464 8032 25470 8084
rect 25682 8032 25688 8084
rect 25740 8072 25746 8084
rect 25869 8075 25927 8081
rect 25869 8072 25881 8075
rect 25740 8044 25881 8072
rect 25740 8032 25746 8044
rect 25869 8041 25881 8044
rect 25915 8041 25927 8075
rect 25869 8035 25927 8041
rect 26142 8032 26148 8084
rect 26200 8032 26206 8084
rect 26694 8032 26700 8084
rect 26752 8032 26758 8084
rect 27062 8032 27068 8084
rect 27120 8032 27126 8084
rect 27798 8032 27804 8084
rect 27856 8032 27862 8084
rect 28905 8075 28963 8081
rect 28905 8072 28917 8075
rect 27908 8044 28917 8072
rect 18414 8004 18420 8016
rect 18248 7976 18420 8004
rect 18141 7967 18199 7973
rect 12084 7908 18000 7936
rect 18156 7936 18184 7967
rect 18414 7964 18420 7976
rect 18472 7964 18478 8016
rect 18506 7964 18512 8016
rect 18564 7964 18570 8016
rect 18708 8004 18736 8032
rect 22097 8007 22155 8013
rect 22097 8004 22109 8007
rect 18708 7976 22109 8004
rect 22097 7973 22109 7976
rect 22143 7973 22155 8007
rect 23566 8004 23572 8016
rect 22097 7967 22155 7973
rect 22296 7976 23572 8004
rect 18524 7936 18552 7964
rect 19702 7936 19708 7948
rect 18156 7908 18460 7936
rect 18524 7908 19708 7936
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 9674 7868 9680 7880
rect 7055 7840 9680 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7868 10011 7871
rect 12084 7868 12112 7908
rect 9999 7840 12112 7868
rect 9999 7837 10011 7840
rect 9953 7831 10011 7837
rect 12526 7828 12532 7880
rect 12584 7828 12590 7880
rect 15470 7828 15476 7880
rect 15528 7828 15534 7880
rect 17494 7828 17500 7880
rect 17552 7828 17558 7880
rect 17773 7871 17831 7877
rect 17773 7837 17785 7871
rect 17819 7868 17831 7871
rect 17954 7868 17960 7880
rect 17819 7840 17960 7868
rect 17819 7837 17831 7840
rect 17773 7831 17831 7837
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 18046 7828 18052 7880
rect 18104 7828 18110 7880
rect 18230 7828 18236 7880
rect 18288 7868 18294 7880
rect 18432 7877 18460 7908
rect 19702 7896 19708 7908
rect 19760 7896 19766 7948
rect 21726 7936 21732 7948
rect 19812 7908 21128 7936
rect 18325 7871 18383 7877
rect 18325 7868 18337 7871
rect 18288 7840 18337 7868
rect 18288 7828 18294 7840
rect 18325 7837 18337 7840
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7837 18475 7871
rect 18417 7831 18475 7837
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19242 7868 19248 7880
rect 18923 7840 19248 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 19334 7828 19340 7880
rect 19392 7828 19398 7880
rect 19812 7877 19840 7908
rect 19797 7871 19855 7877
rect 19797 7837 19809 7871
rect 19843 7837 19855 7871
rect 19797 7831 19855 7837
rect 19886 7828 19892 7880
rect 19944 7828 19950 7880
rect 20162 7828 20168 7880
rect 20220 7828 20226 7880
rect 20441 7871 20499 7877
rect 20441 7837 20453 7871
rect 20487 7868 20499 7871
rect 20622 7868 20628 7880
rect 20487 7840 20628 7868
rect 20487 7837 20499 7840
rect 20441 7831 20499 7837
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7868 20775 7871
rect 20898 7868 20904 7880
rect 20763 7840 20904 7868
rect 20763 7837 20775 7840
rect 20717 7831 20775 7837
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 6472 7772 9076 7800
rect 5445 7763 5503 7769
rect 5460 7732 5488 7763
rect 8938 7732 8944 7744
rect 5460 7704 8944 7732
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 9048 7732 9076 7772
rect 9122 7760 9128 7812
rect 9180 7760 9186 7812
rect 11698 7760 11704 7812
rect 11756 7760 11762 7812
rect 14274 7760 14280 7812
rect 14332 7760 14338 7812
rect 11790 7732 11796 7744
rect 9048 7704 11796 7732
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 17512 7732 17540 7828
rect 17862 7760 17868 7812
rect 17920 7800 17926 7812
rect 21100 7800 21128 7908
rect 21468 7908 21732 7936
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7868 21235 7871
rect 21358 7868 21364 7880
rect 21223 7840 21364 7868
rect 21223 7837 21235 7840
rect 21177 7831 21235 7837
rect 21358 7828 21364 7840
rect 21416 7828 21422 7880
rect 21468 7877 21496 7908
rect 21726 7896 21732 7908
rect 21784 7896 21790 7948
rect 21453 7871 21511 7877
rect 21453 7837 21465 7871
rect 21499 7837 21511 7871
rect 21453 7831 21511 7837
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7868 21603 7871
rect 21818 7868 21824 7880
rect 21591 7840 21824 7868
rect 21591 7837 21603 7840
rect 21545 7831 21603 7837
rect 21818 7828 21824 7840
rect 21876 7828 21882 7880
rect 22002 7828 22008 7880
rect 22060 7828 22066 7880
rect 22296 7877 22324 7976
rect 23566 7964 23572 7976
rect 23624 7964 23630 8016
rect 25148 8004 25176 8032
rect 23768 7976 25176 8004
rect 23014 7936 23020 7948
rect 22388 7908 23020 7936
rect 22388 7877 22416 7908
rect 23014 7896 23020 7908
rect 23072 7896 23078 7948
rect 22281 7871 22339 7877
rect 22281 7837 22293 7871
rect 22327 7837 22339 7871
rect 22281 7831 22339 7837
rect 22373 7871 22431 7877
rect 22373 7837 22385 7871
rect 22419 7837 22431 7871
rect 22373 7831 22431 7837
rect 22646 7828 22652 7880
rect 22704 7828 22710 7880
rect 22925 7871 22983 7877
rect 22925 7837 22937 7871
rect 22971 7868 22983 7871
rect 23106 7868 23112 7880
rect 22971 7840 23112 7868
rect 22971 7837 22983 7840
rect 22925 7831 22983 7837
rect 23106 7828 23112 7840
rect 23164 7828 23170 7880
rect 23198 7828 23204 7880
rect 23256 7828 23262 7880
rect 23768 7877 23796 7976
rect 25424 7936 25452 8032
rect 25498 7964 25504 8016
rect 25556 8004 25562 8016
rect 27433 8007 27491 8013
rect 27433 8004 27445 8007
rect 25556 7976 27445 8004
rect 25556 7964 25562 7976
rect 27433 7973 27445 7976
rect 27479 7973 27491 8007
rect 27433 7967 27491 7973
rect 24596 7908 24808 7936
rect 23477 7871 23535 7877
rect 23477 7837 23489 7871
rect 23523 7837 23535 7871
rect 23477 7831 23535 7837
rect 23753 7871 23811 7877
rect 23753 7837 23765 7871
rect 23799 7837 23811 7871
rect 23753 7831 23811 7837
rect 24029 7871 24087 7877
rect 24029 7837 24041 7871
rect 24075 7868 24087 7871
rect 24486 7868 24492 7880
rect 24075 7840 24492 7868
rect 24075 7837 24087 7840
rect 24029 7831 24087 7837
rect 21910 7800 21916 7812
rect 17920 7772 20944 7800
rect 21100 7772 21916 7800
rect 17920 7760 17926 7772
rect 17589 7735 17647 7741
rect 17589 7732 17601 7735
rect 17512 7704 17601 7732
rect 17589 7701 17601 7704
rect 17635 7701 17647 7735
rect 17589 7695 17647 7701
rect 17678 7692 17684 7744
rect 17736 7732 17742 7744
rect 19061 7735 19119 7741
rect 19061 7732 19073 7735
rect 17736 7704 19073 7732
rect 17736 7692 17742 7704
rect 19061 7701 19073 7704
rect 19107 7701 19119 7735
rect 19061 7695 19119 7701
rect 19518 7692 19524 7744
rect 19576 7692 19582 7744
rect 20070 7692 20076 7744
rect 20128 7692 20134 7744
rect 20346 7692 20352 7744
rect 20404 7692 20410 7744
rect 20438 7692 20444 7744
rect 20496 7732 20502 7744
rect 20916 7741 20944 7772
rect 21910 7760 21916 7772
rect 21968 7760 21974 7812
rect 23492 7800 23520 7831
rect 24486 7828 24492 7840
rect 24544 7828 24550 7880
rect 24596 7877 24624 7908
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 24670 7828 24676 7880
rect 24728 7828 24734 7880
rect 24688 7800 24716 7828
rect 22066 7772 23428 7800
rect 23492 7772 24716 7800
rect 24780 7800 24808 7908
rect 24872 7908 25452 7936
rect 24872 7877 24900 7908
rect 26786 7896 26792 7948
rect 26844 7896 26850 7948
rect 27338 7896 27344 7948
rect 27396 7896 27402 7948
rect 27908 7936 27936 8044
rect 28905 8041 28917 8044
rect 28951 8041 28963 8075
rect 28905 8035 28963 8041
rect 29270 8032 29276 8084
rect 29328 8032 29334 8084
rect 40770 8032 40776 8084
rect 40828 8072 40834 8084
rect 41141 8075 41199 8081
rect 41141 8072 41153 8075
rect 40828 8044 41153 8072
rect 40828 8032 40834 8044
rect 41141 8041 41153 8044
rect 41187 8041 41199 8075
rect 41141 8035 41199 8041
rect 44450 8032 44456 8084
rect 44508 8072 44514 8084
rect 45189 8075 45247 8081
rect 45189 8072 45201 8075
rect 44508 8044 45201 8072
rect 44508 8032 44514 8044
rect 45189 8041 45201 8044
rect 45235 8041 45247 8075
rect 45189 8035 45247 8041
rect 28718 8004 28724 8016
rect 27448 7908 27936 7936
rect 28000 7976 28724 8004
rect 24857 7871 24915 7877
rect 24857 7837 24869 7871
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 25038 7828 25044 7880
rect 25096 7868 25102 7880
rect 25133 7871 25191 7877
rect 25133 7868 25145 7871
rect 25096 7840 25145 7868
rect 25096 7828 25102 7840
rect 25133 7837 25145 7840
rect 25179 7837 25191 7871
rect 25133 7831 25191 7837
rect 25409 7871 25467 7877
rect 25409 7837 25421 7871
rect 25455 7868 25467 7871
rect 25590 7868 25596 7880
rect 25455 7840 25596 7868
rect 25455 7837 25467 7840
rect 25409 7831 25467 7837
rect 25590 7828 25596 7840
rect 25648 7828 25654 7880
rect 25685 7871 25743 7877
rect 25685 7837 25697 7871
rect 25731 7868 25743 7871
rect 25866 7868 25872 7880
rect 25731 7840 25872 7868
rect 25731 7837 25743 7840
rect 25685 7831 25743 7837
rect 25866 7828 25872 7840
rect 25924 7828 25930 7880
rect 25961 7871 26019 7877
rect 25961 7837 25973 7871
rect 26007 7868 26019 7871
rect 26050 7868 26056 7880
rect 26007 7840 26056 7868
rect 26007 7837 26019 7840
rect 25961 7831 26019 7837
rect 26050 7828 26056 7840
rect 26108 7828 26114 7880
rect 26237 7871 26295 7877
rect 26237 7837 26249 7871
rect 26283 7868 26295 7871
rect 26418 7868 26424 7880
rect 26283 7840 26424 7868
rect 26283 7837 26295 7840
rect 26237 7831 26295 7837
rect 26418 7828 26424 7840
rect 26476 7828 26482 7880
rect 26513 7871 26571 7877
rect 26513 7837 26525 7871
rect 26559 7868 26571 7871
rect 26804 7868 26832 7896
rect 26559 7840 26832 7868
rect 26881 7871 26939 7877
rect 26559 7837 26571 7840
rect 26513 7831 26571 7837
rect 26881 7837 26893 7871
rect 26927 7868 26939 7871
rect 27154 7868 27160 7880
rect 26927 7840 27160 7868
rect 26927 7837 26939 7840
rect 26881 7831 26939 7837
rect 27154 7828 27160 7840
rect 27212 7828 27218 7880
rect 27249 7871 27307 7877
rect 27249 7837 27261 7871
rect 27295 7868 27307 7871
rect 27356 7868 27384 7896
rect 27448 7880 27476 7908
rect 27295 7840 27384 7868
rect 27295 7837 27307 7840
rect 27249 7831 27307 7837
rect 27430 7828 27436 7880
rect 27488 7828 27494 7880
rect 27617 7871 27675 7877
rect 27617 7837 27629 7871
rect 27663 7868 27675 7871
rect 27890 7868 27896 7880
rect 27663 7840 27896 7868
rect 27663 7837 27675 7840
rect 27617 7831 27675 7837
rect 27890 7828 27896 7840
rect 27948 7828 27954 7880
rect 28000 7877 28028 7976
rect 28718 7964 28724 7976
rect 28776 7964 28782 8016
rect 29288 7936 29316 8032
rect 44545 8007 44603 8013
rect 44545 7973 44557 8007
rect 44591 8004 44603 8007
rect 45922 8004 45928 8016
rect 44591 7976 45928 8004
rect 44591 7973 44603 7976
rect 44545 7967 44603 7973
rect 45922 7964 45928 7976
rect 45980 7964 45986 8016
rect 28368 7908 29316 7936
rect 28368 7877 28396 7908
rect 27985 7871 28043 7877
rect 27985 7837 27997 7871
rect 28031 7837 28043 7871
rect 27985 7831 28043 7837
rect 28353 7871 28411 7877
rect 28353 7837 28365 7871
rect 28399 7837 28411 7871
rect 28353 7831 28411 7837
rect 28721 7871 28779 7877
rect 28721 7837 28733 7871
rect 28767 7868 28779 7871
rect 29546 7868 29552 7880
rect 28767 7840 29552 7868
rect 28767 7837 28779 7840
rect 28721 7831 28779 7837
rect 29546 7828 29552 7840
rect 29604 7828 29610 7880
rect 29822 7828 29828 7880
rect 29880 7828 29886 7880
rect 40954 7828 40960 7880
rect 41012 7828 41018 7880
rect 44085 7871 44143 7877
rect 44085 7837 44097 7871
rect 44131 7868 44143 7871
rect 46290 7868 46296 7880
rect 44131 7840 46296 7868
rect 44131 7837 44143 7840
rect 44085 7831 44143 7837
rect 46290 7828 46296 7840
rect 46348 7828 46354 7880
rect 29840 7800 29868 7828
rect 24780 7772 29868 7800
rect 43717 7803 43775 7809
rect 22066 7744 22094 7772
rect 20625 7735 20683 7741
rect 20625 7732 20637 7735
rect 20496 7704 20637 7732
rect 20496 7692 20502 7704
rect 20625 7701 20637 7704
rect 20671 7701 20683 7735
rect 20625 7695 20683 7701
rect 20901 7735 20959 7741
rect 20901 7701 20913 7735
rect 20947 7701 20959 7735
rect 20901 7695 20959 7701
rect 21726 7692 21732 7744
rect 21784 7692 21790 7744
rect 22002 7692 22008 7744
rect 22060 7704 22094 7744
rect 23400 7741 23428 7772
rect 43717 7769 43729 7803
rect 43763 7800 43775 7803
rect 44174 7800 44180 7812
rect 43763 7772 44180 7800
rect 43763 7769 43775 7772
rect 43717 7763 43775 7769
rect 44174 7760 44180 7772
rect 44232 7760 44238 7812
rect 44269 7803 44327 7809
rect 44269 7769 44281 7803
rect 44315 7800 44327 7803
rect 45002 7800 45008 7812
rect 44315 7772 45008 7800
rect 44315 7769 44327 7772
rect 44269 7763 44327 7769
rect 45002 7760 45008 7772
rect 45060 7760 45066 7812
rect 45097 7803 45155 7809
rect 45097 7769 45109 7803
rect 45143 7769 45155 7803
rect 45097 7763 45155 7769
rect 23385 7735 23443 7741
rect 22060 7692 22066 7704
rect 23385 7701 23397 7735
rect 23431 7701 23443 7735
rect 23385 7695 23443 7701
rect 23661 7735 23719 7741
rect 23661 7701 23673 7735
rect 23707 7732 23719 7735
rect 24118 7732 24124 7744
rect 23707 7704 24124 7732
rect 23707 7701 23719 7704
rect 23661 7695 23719 7701
rect 24118 7692 24124 7704
rect 24176 7692 24182 7744
rect 25038 7692 25044 7744
rect 25096 7692 25102 7744
rect 25314 7692 25320 7744
rect 25372 7692 25378 7744
rect 25590 7692 25596 7744
rect 25648 7692 25654 7744
rect 26418 7692 26424 7744
rect 26476 7692 26482 7744
rect 28166 7692 28172 7744
rect 28224 7692 28230 7744
rect 28534 7692 28540 7744
rect 28592 7692 28598 7744
rect 43898 7692 43904 7744
rect 43956 7732 43962 7744
rect 45112 7732 45140 7763
rect 43956 7704 45140 7732
rect 43956 7692 43962 7704
rect 1104 7642 45976 7664
rect 1104 7590 12128 7642
rect 12180 7590 12192 7642
rect 12244 7590 12256 7642
rect 12308 7590 12320 7642
rect 12372 7590 12384 7642
rect 12436 7590 23306 7642
rect 23358 7590 23370 7642
rect 23422 7590 23434 7642
rect 23486 7590 23498 7642
rect 23550 7590 23562 7642
rect 23614 7590 34484 7642
rect 34536 7590 34548 7642
rect 34600 7590 34612 7642
rect 34664 7590 34676 7642
rect 34728 7590 34740 7642
rect 34792 7590 45662 7642
rect 45714 7590 45726 7642
rect 45778 7590 45790 7642
rect 45842 7590 45854 7642
rect 45906 7590 45918 7642
rect 45970 7590 45976 7642
rect 1104 7568 45976 7590
rect 1026 7488 1032 7540
rect 1084 7528 1090 7540
rect 1581 7531 1639 7537
rect 1581 7528 1593 7531
rect 1084 7500 1593 7528
rect 1084 7488 1090 7500
rect 1581 7497 1593 7500
rect 1627 7497 1639 7531
rect 1581 7491 1639 7497
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 2133 7531 2191 7537
rect 2133 7528 2145 7531
rect 1820 7500 2145 7528
rect 1820 7488 1826 7500
rect 2133 7497 2145 7500
rect 2179 7497 2191 7531
rect 17678 7528 17684 7540
rect 2133 7491 2191 7497
rect 2746 7500 17684 7528
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7361 1547 7395
rect 1489 7355 1547 7361
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7392 2007 7395
rect 2746 7392 2774 7500
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 17862 7488 17868 7540
rect 17920 7488 17926 7540
rect 18877 7531 18935 7537
rect 18877 7497 18889 7531
rect 18923 7528 18935 7531
rect 19334 7528 19340 7540
rect 18923 7500 19340 7528
rect 18923 7497 18935 7500
rect 18877 7491 18935 7497
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 19521 7531 19579 7537
rect 19521 7497 19533 7531
rect 19567 7528 19579 7531
rect 19978 7528 19984 7540
rect 19567 7500 19984 7528
rect 19567 7497 19579 7500
rect 19521 7491 19579 7497
rect 19978 7488 19984 7500
rect 20036 7488 20042 7540
rect 20162 7488 20168 7540
rect 20220 7528 20226 7540
rect 20349 7531 20407 7537
rect 20349 7528 20361 7531
rect 20220 7500 20361 7528
rect 20220 7488 20226 7500
rect 20349 7497 20361 7500
rect 20395 7497 20407 7531
rect 20622 7528 20628 7540
rect 20349 7491 20407 7497
rect 20548 7500 20628 7528
rect 4338 7420 4344 7472
rect 4396 7460 4402 7472
rect 8294 7460 8300 7472
rect 4396 7432 8300 7460
rect 4396 7420 4402 7432
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 9122 7420 9128 7472
rect 9180 7420 9186 7472
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 17880 7460 17908 7488
rect 9732 7432 17908 7460
rect 18800 7432 20484 7460
rect 9732 7420 9738 7432
rect 1995 7364 2774 7392
rect 9140 7392 9168 7420
rect 9140 7364 15424 7392
rect 1995 7361 2007 7364
rect 1949 7355 2007 7361
rect 1504 7324 1532 7355
rect 15102 7324 15108 7336
rect 1504 7296 15108 7324
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 15396 7324 15424 7364
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 18800 7392 18828 7432
rect 15528 7364 18828 7392
rect 15528 7352 15534 7364
rect 19058 7352 19064 7404
rect 19116 7352 19122 7404
rect 19334 7352 19340 7404
rect 19392 7352 19398 7404
rect 19702 7352 19708 7404
rect 19760 7352 19766 7404
rect 19794 7352 19800 7404
rect 19852 7392 19858 7404
rect 20073 7395 20131 7401
rect 20073 7392 20085 7395
rect 19852 7364 20085 7392
rect 19852 7352 19858 7364
rect 20073 7361 20085 7364
rect 20119 7361 20131 7395
rect 20073 7355 20131 7361
rect 17218 7324 17224 7336
rect 15396 7296 17224 7324
rect 17218 7284 17224 7296
rect 17276 7284 17282 7336
rect 18782 7284 18788 7336
rect 18840 7284 18846 7336
rect 19886 7284 19892 7336
rect 19944 7284 19950 7336
rect 20456 7324 20484 7432
rect 20548 7401 20576 7500
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 21174 7488 21180 7540
rect 21232 7488 21238 7540
rect 21450 7488 21456 7540
rect 21508 7488 21514 7540
rect 21542 7488 21548 7540
rect 21600 7488 21606 7540
rect 21634 7488 21640 7540
rect 21692 7528 21698 7540
rect 22005 7531 22063 7537
rect 22005 7528 22017 7531
rect 21692 7500 22017 7528
rect 21692 7488 21698 7500
rect 22005 7497 22017 7500
rect 22051 7497 22063 7531
rect 22005 7491 22063 7497
rect 22649 7531 22707 7537
rect 22649 7497 22661 7531
rect 22695 7497 22707 7531
rect 22649 7491 22707 7497
rect 22848 7500 23336 7528
rect 20533 7395 20591 7401
rect 20533 7361 20545 7395
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 20806 7352 20812 7404
rect 20864 7352 20870 7404
rect 21192 7392 21220 7488
rect 21468 7460 21496 7488
rect 22664 7460 22692 7491
rect 21468 7432 21864 7460
rect 21836 7401 21864 7432
rect 21928 7432 22692 7460
rect 21361 7395 21419 7401
rect 21361 7392 21373 7395
rect 21192 7364 21373 7392
rect 21361 7361 21373 7364
rect 21407 7361 21419 7395
rect 21361 7355 21419 7361
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 21928 7324 21956 7432
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7392 22155 7395
rect 22278 7392 22284 7404
rect 22143 7364 22284 7392
rect 22143 7361 22155 7364
rect 22097 7355 22155 7361
rect 22278 7352 22284 7364
rect 22336 7352 22342 7404
rect 22373 7395 22431 7401
rect 22373 7361 22385 7395
rect 22419 7392 22431 7395
rect 22738 7392 22744 7404
rect 22419 7364 22744 7392
rect 22419 7361 22431 7364
rect 22373 7355 22431 7361
rect 22738 7352 22744 7364
rect 22796 7352 22802 7404
rect 22848 7401 22876 7500
rect 23308 7460 23336 7500
rect 23382 7488 23388 7540
rect 23440 7528 23446 7540
rect 31846 7528 31852 7540
rect 23440 7500 31852 7528
rect 23440 7488 23446 7500
rect 31846 7488 31852 7500
rect 31904 7488 31910 7540
rect 43346 7488 43352 7540
rect 43404 7528 43410 7540
rect 44085 7531 44143 7537
rect 44085 7528 44097 7531
rect 43404 7500 44097 7528
rect 43404 7488 43410 7500
rect 44085 7497 44097 7500
rect 44131 7497 44143 7531
rect 44085 7491 44143 7497
rect 45189 7531 45247 7537
rect 45189 7497 45201 7531
rect 45235 7528 45247 7531
rect 45554 7528 45560 7540
rect 45235 7500 45560 7528
rect 45235 7497 45247 7500
rect 45189 7491 45247 7497
rect 45554 7488 45560 7500
rect 45612 7488 45618 7540
rect 33778 7460 33784 7472
rect 23308 7432 33784 7460
rect 33778 7420 33784 7432
rect 33836 7420 33842 7472
rect 44729 7463 44787 7469
rect 44729 7429 44741 7463
rect 44775 7460 44787 7463
rect 44775 7432 45232 7460
rect 44775 7429 44787 7432
rect 44729 7423 44787 7429
rect 45204 7404 45232 7432
rect 22833 7395 22891 7401
rect 22833 7361 22845 7395
rect 22879 7361 22891 7395
rect 22833 7355 22891 7361
rect 23109 7395 23167 7401
rect 23109 7361 23121 7395
rect 23155 7392 23167 7395
rect 23198 7392 23204 7404
rect 23155 7364 23204 7392
rect 23155 7361 23167 7364
rect 23109 7355 23167 7361
rect 23198 7352 23204 7364
rect 23256 7352 23262 7404
rect 23290 7352 23296 7404
rect 23348 7352 23354 7404
rect 23385 7395 23443 7401
rect 23385 7361 23397 7395
rect 23431 7392 23443 7395
rect 23566 7392 23572 7404
rect 23431 7364 23572 7392
rect 23431 7361 23443 7364
rect 23385 7355 23443 7361
rect 23566 7352 23572 7364
rect 23624 7352 23630 7404
rect 23661 7395 23719 7401
rect 23661 7361 23673 7395
rect 23707 7392 23719 7395
rect 23842 7392 23848 7404
rect 23707 7364 23848 7392
rect 23707 7361 23719 7364
rect 23661 7355 23719 7361
rect 23842 7352 23848 7364
rect 23900 7352 23906 7404
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7392 23995 7395
rect 27522 7392 27528 7404
rect 23983 7364 27528 7392
rect 23983 7361 23995 7364
rect 23937 7355 23995 7361
rect 27522 7352 27528 7364
rect 27580 7352 27586 7404
rect 41414 7352 41420 7404
rect 41472 7392 41478 7404
rect 43901 7395 43959 7401
rect 43901 7392 43913 7395
rect 41472 7364 43913 7392
rect 41472 7352 41478 7364
rect 43901 7361 43913 7364
rect 43947 7361 43959 7395
rect 43901 7355 43959 7361
rect 44358 7352 44364 7404
rect 44416 7352 44422 7404
rect 44910 7352 44916 7404
rect 44968 7352 44974 7404
rect 45186 7352 45192 7404
rect 45244 7352 45250 7404
rect 20456 7296 21956 7324
rect 23308 7324 23336 7352
rect 30650 7324 30656 7336
rect 23308 7296 30656 7324
rect 30650 7284 30656 7296
rect 30708 7284 30714 7336
rect 2314 7216 2320 7268
rect 2372 7256 2378 7268
rect 9674 7256 9680 7268
rect 2372 7228 9680 7256
rect 2372 7216 2378 7228
rect 9674 7216 9680 7228
rect 9732 7216 9738 7268
rect 16666 7216 16672 7268
rect 16724 7256 16730 7268
rect 18506 7256 18512 7268
rect 16724 7228 18512 7256
rect 16724 7216 16730 7228
rect 18506 7216 18512 7228
rect 18564 7216 18570 7268
rect 18800 7256 18828 7284
rect 19153 7259 19211 7265
rect 19153 7256 19165 7259
rect 18800 7228 19165 7256
rect 19153 7225 19165 7228
rect 19199 7225 19211 7259
rect 19153 7219 19211 7225
rect 19242 7216 19248 7268
rect 19300 7216 19306 7268
rect 19904 7256 19932 7284
rect 20625 7259 20683 7265
rect 20625 7256 20637 7259
rect 19904 7228 20637 7256
rect 20625 7225 20637 7228
rect 20671 7225 20683 7259
rect 21634 7256 21640 7268
rect 20625 7219 20683 7225
rect 20732 7228 21640 7256
rect 14458 7148 14464 7200
rect 14516 7188 14522 7200
rect 19058 7188 19064 7200
rect 14516 7160 19064 7188
rect 14516 7148 14522 7160
rect 19058 7148 19064 7160
rect 19116 7148 19122 7200
rect 19260 7188 19288 7216
rect 20732 7200 20760 7228
rect 21634 7216 21640 7228
rect 21692 7216 21698 7268
rect 22204 7228 22968 7256
rect 19889 7191 19947 7197
rect 19889 7188 19901 7191
rect 19260 7160 19901 7188
rect 19889 7157 19901 7160
rect 19935 7157 19947 7191
rect 19889 7151 19947 7157
rect 20714 7148 20720 7200
rect 20772 7148 20778 7200
rect 21082 7148 21088 7200
rect 21140 7188 21146 7200
rect 22204 7188 22232 7228
rect 21140 7160 22232 7188
rect 21140 7148 21146 7160
rect 22278 7148 22284 7200
rect 22336 7148 22342 7200
rect 22370 7148 22376 7200
rect 22428 7188 22434 7200
rect 22940 7197 22968 7228
rect 23474 7216 23480 7268
rect 23532 7256 23538 7268
rect 33318 7256 33324 7268
rect 23532 7228 33324 7256
rect 23532 7216 23538 7228
rect 33318 7216 33324 7228
rect 33376 7216 33382 7268
rect 22557 7191 22615 7197
rect 22557 7188 22569 7191
rect 22428 7160 22569 7188
rect 22428 7148 22434 7160
rect 22557 7157 22569 7160
rect 22603 7157 22615 7191
rect 22557 7151 22615 7157
rect 22925 7191 22983 7197
rect 22925 7157 22937 7191
rect 22971 7157 22983 7191
rect 22925 7151 22983 7157
rect 23198 7148 23204 7200
rect 23256 7148 23262 7200
rect 23842 7148 23848 7200
rect 23900 7148 23906 7200
rect 24121 7191 24179 7197
rect 24121 7157 24133 7191
rect 24167 7188 24179 7191
rect 24394 7188 24400 7200
rect 24167 7160 24400 7188
rect 24167 7157 24179 7160
rect 24121 7151 24179 7157
rect 24394 7148 24400 7160
rect 24452 7148 24458 7200
rect 1104 7098 45816 7120
rect 1104 7046 6539 7098
rect 6591 7046 6603 7098
rect 6655 7046 6667 7098
rect 6719 7046 6731 7098
rect 6783 7046 6795 7098
rect 6847 7046 17717 7098
rect 17769 7046 17781 7098
rect 17833 7046 17845 7098
rect 17897 7046 17909 7098
rect 17961 7046 17973 7098
rect 18025 7046 28895 7098
rect 28947 7046 28959 7098
rect 29011 7046 29023 7098
rect 29075 7046 29087 7098
rect 29139 7046 29151 7098
rect 29203 7046 40073 7098
rect 40125 7046 40137 7098
rect 40189 7046 40201 7098
rect 40253 7046 40265 7098
rect 40317 7046 40329 7098
rect 40381 7046 45816 7098
rect 1104 7024 45816 7046
rect 12618 6944 12624 6996
rect 12676 6944 12682 6996
rect 15194 6944 15200 6996
rect 15252 6984 15258 6996
rect 21082 6984 21088 6996
rect 15252 6956 21088 6984
rect 15252 6944 15258 6956
rect 21082 6944 21088 6956
rect 21140 6944 21146 6996
rect 21358 6944 21364 6996
rect 21416 6984 21422 6996
rect 34146 6984 34152 6996
rect 21416 6956 34152 6984
rect 21416 6944 21422 6956
rect 34146 6944 34152 6956
rect 34204 6944 34210 6996
rect 12636 6916 12664 6944
rect 12636 6888 19380 6916
rect 19352 6848 19380 6888
rect 19702 6876 19708 6928
rect 19760 6916 19766 6928
rect 33686 6916 33692 6928
rect 19760 6888 33692 6916
rect 19760 6876 19766 6888
rect 33686 6876 33692 6888
rect 33744 6876 33750 6928
rect 20714 6848 20720 6860
rect 19352 6820 20720 6848
rect 20714 6808 20720 6820
rect 20772 6808 20778 6860
rect 44082 6808 44088 6860
rect 44140 6848 44146 6860
rect 45373 6851 45431 6857
rect 45373 6848 45385 6851
rect 44140 6820 45385 6848
rect 44140 6808 44146 6820
rect 45373 6817 45385 6820
rect 45419 6817 45431 6851
rect 45373 6811 45431 6817
rect 23109 6783 23167 6789
rect 23109 6749 23121 6783
rect 23155 6780 23167 6783
rect 36630 6780 36636 6792
rect 23155 6752 36636 6780
rect 23155 6749 23167 6752
rect 23109 6743 23167 6749
rect 36630 6740 36636 6752
rect 36688 6740 36694 6792
rect 3970 6672 3976 6724
rect 4028 6712 4034 6724
rect 25314 6712 25320 6724
rect 4028 6684 25320 6712
rect 4028 6672 4034 6684
rect 25314 6672 25320 6684
rect 25372 6672 25378 6724
rect 42794 6672 42800 6724
rect 42852 6712 42858 6724
rect 45097 6715 45155 6721
rect 45097 6712 45109 6715
rect 42852 6684 45109 6712
rect 42852 6672 42858 6684
rect 45097 6681 45109 6684
rect 45143 6681 45155 6715
rect 45097 6675 45155 6681
rect 16574 6604 16580 6656
rect 16632 6644 16638 6656
rect 22925 6647 22983 6653
rect 22925 6644 22937 6647
rect 16632 6616 22937 6644
rect 16632 6604 16638 6616
rect 22925 6613 22937 6616
rect 22971 6613 22983 6647
rect 22925 6607 22983 6613
rect 1104 6554 45976 6576
rect 1104 6502 12128 6554
rect 12180 6502 12192 6554
rect 12244 6502 12256 6554
rect 12308 6502 12320 6554
rect 12372 6502 12384 6554
rect 12436 6502 23306 6554
rect 23358 6502 23370 6554
rect 23422 6502 23434 6554
rect 23486 6502 23498 6554
rect 23550 6502 23562 6554
rect 23614 6502 34484 6554
rect 34536 6502 34548 6554
rect 34600 6502 34612 6554
rect 34664 6502 34676 6554
rect 34728 6502 34740 6554
rect 34792 6502 45662 6554
rect 45714 6502 45726 6554
rect 45778 6502 45790 6554
rect 45842 6502 45854 6554
rect 45906 6502 45918 6554
rect 45970 6502 45976 6554
rect 1104 6480 45976 6502
rect 24946 6196 24952 6248
rect 25004 6236 25010 6248
rect 39390 6236 39396 6248
rect 25004 6208 39396 6236
rect 25004 6196 25010 6208
rect 39390 6196 39396 6208
rect 39448 6196 39454 6248
rect 27246 6128 27252 6180
rect 27304 6168 27310 6180
rect 43070 6168 43076 6180
rect 27304 6140 43076 6168
rect 27304 6128 27310 6140
rect 43070 6128 43076 6140
rect 43128 6128 43134 6180
rect 1104 6010 45816 6032
rect 1104 5958 6539 6010
rect 6591 5958 6603 6010
rect 6655 5958 6667 6010
rect 6719 5958 6731 6010
rect 6783 5958 6795 6010
rect 6847 5958 17717 6010
rect 17769 5958 17781 6010
rect 17833 5958 17845 6010
rect 17897 5958 17909 6010
rect 17961 5958 17973 6010
rect 18025 5958 28895 6010
rect 28947 5958 28959 6010
rect 29011 5958 29023 6010
rect 29075 5958 29087 6010
rect 29139 5958 29151 6010
rect 29203 5958 40073 6010
rect 40125 5958 40137 6010
rect 40189 5958 40201 6010
rect 40253 5958 40265 6010
rect 40317 5958 40329 6010
rect 40381 5958 45816 6010
rect 1104 5936 45816 5958
rect 1104 5466 45976 5488
rect 1104 5414 12128 5466
rect 12180 5414 12192 5466
rect 12244 5414 12256 5466
rect 12308 5414 12320 5466
rect 12372 5414 12384 5466
rect 12436 5414 23306 5466
rect 23358 5414 23370 5466
rect 23422 5414 23434 5466
rect 23486 5414 23498 5466
rect 23550 5414 23562 5466
rect 23614 5414 34484 5466
rect 34536 5414 34548 5466
rect 34600 5414 34612 5466
rect 34664 5414 34676 5466
rect 34728 5414 34740 5466
rect 34792 5414 45662 5466
rect 45714 5414 45726 5466
rect 45778 5414 45790 5466
rect 45842 5414 45854 5466
rect 45906 5414 45918 5466
rect 45970 5414 45976 5466
rect 1104 5392 45976 5414
rect 1104 4922 45816 4944
rect 1104 4870 6539 4922
rect 6591 4870 6603 4922
rect 6655 4870 6667 4922
rect 6719 4870 6731 4922
rect 6783 4870 6795 4922
rect 6847 4870 17717 4922
rect 17769 4870 17781 4922
rect 17833 4870 17845 4922
rect 17897 4870 17909 4922
rect 17961 4870 17973 4922
rect 18025 4870 28895 4922
rect 28947 4870 28959 4922
rect 29011 4870 29023 4922
rect 29075 4870 29087 4922
rect 29139 4870 29151 4922
rect 29203 4870 40073 4922
rect 40125 4870 40137 4922
rect 40189 4870 40201 4922
rect 40253 4870 40265 4922
rect 40317 4870 40329 4922
rect 40381 4870 45816 4922
rect 1104 4848 45816 4870
rect 23106 4768 23112 4820
rect 23164 4808 23170 4820
rect 38378 4808 38384 4820
rect 23164 4780 38384 4808
rect 23164 4768 23170 4780
rect 38378 4768 38384 4780
rect 38436 4768 38442 4820
rect 43898 4768 43904 4820
rect 43956 4768 43962 4820
rect 36081 4743 36139 4749
rect 36081 4709 36093 4743
rect 36127 4740 36139 4743
rect 43916 4740 43944 4768
rect 36127 4712 43944 4740
rect 36127 4709 36139 4712
rect 36081 4703 36139 4709
rect 23569 4607 23627 4613
rect 23569 4573 23581 4607
rect 23615 4604 23627 4607
rect 23658 4604 23664 4616
rect 23615 4576 23664 4604
rect 23615 4573 23627 4576
rect 23569 4567 23627 4573
rect 23658 4564 23664 4576
rect 23716 4564 23722 4616
rect 35894 4564 35900 4616
rect 35952 4564 35958 4616
rect 39942 4536 39948 4548
rect 31726 4508 39948 4536
rect 23753 4471 23811 4477
rect 23753 4437 23765 4471
rect 23799 4468 23811 4471
rect 31726 4468 31754 4508
rect 39942 4496 39948 4508
rect 40000 4496 40006 4548
rect 23799 4440 31754 4468
rect 23799 4437 23811 4440
rect 23753 4431 23811 4437
rect 1104 4378 45976 4400
rect 1104 4326 12128 4378
rect 12180 4326 12192 4378
rect 12244 4326 12256 4378
rect 12308 4326 12320 4378
rect 12372 4326 12384 4378
rect 12436 4326 23306 4378
rect 23358 4326 23370 4378
rect 23422 4326 23434 4378
rect 23486 4326 23498 4378
rect 23550 4326 23562 4378
rect 23614 4326 34484 4378
rect 34536 4326 34548 4378
rect 34600 4326 34612 4378
rect 34664 4326 34676 4378
rect 34728 4326 34740 4378
rect 34792 4326 45662 4378
rect 45714 4326 45726 4378
rect 45778 4326 45790 4378
rect 45842 4326 45854 4378
rect 45906 4326 45918 4378
rect 45970 4326 45976 4378
rect 1104 4304 45976 4326
rect 22646 4088 22652 4140
rect 22704 4088 22710 4140
rect 23109 4131 23167 4137
rect 23109 4097 23121 4131
rect 23155 4097 23167 4131
rect 23109 4091 23167 4097
rect 20806 4020 20812 4072
rect 20864 4060 20870 4072
rect 23124 4060 23152 4091
rect 23198 4088 23204 4140
rect 23256 4128 23262 4140
rect 23661 4131 23719 4137
rect 23661 4128 23673 4131
rect 23256 4100 23673 4128
rect 23256 4088 23262 4100
rect 23661 4097 23673 4100
rect 23707 4097 23719 4131
rect 23661 4091 23719 4097
rect 27062 4088 27068 4140
rect 27120 4088 27126 4140
rect 33686 4088 33692 4140
rect 33744 4088 33750 4140
rect 35434 4088 35440 4140
rect 35492 4088 35498 4140
rect 44542 4088 44548 4140
rect 44600 4088 44606 4140
rect 35802 4060 35808 4072
rect 20864 4032 23152 4060
rect 23768 4032 35808 4060
rect 20864 4020 20870 4032
rect 22833 3995 22891 4001
rect 22833 3961 22845 3995
rect 22879 3961 22891 3995
rect 22833 3955 22891 3961
rect 22925 3995 22983 4001
rect 22925 3961 22937 3995
rect 22971 3992 22983 3995
rect 23658 3992 23664 4004
rect 22971 3964 23664 3992
rect 22971 3961 22983 3964
rect 22925 3955 22983 3961
rect 22848 3924 22876 3955
rect 23658 3952 23664 3964
rect 23716 3952 23722 4004
rect 23768 3924 23796 4032
rect 35802 4020 35808 4032
rect 35860 4020 35866 4072
rect 23860 3964 31754 3992
rect 23860 3933 23888 3964
rect 22848 3896 23796 3924
rect 23845 3927 23903 3933
rect 23845 3893 23857 3927
rect 23891 3893 23903 3927
rect 23845 3887 23903 3893
rect 27246 3884 27252 3936
rect 27304 3884 27310 3936
rect 31726 3924 31754 3964
rect 33594 3952 33600 4004
rect 33652 3952 33658 4004
rect 35253 3995 35311 4001
rect 35253 3961 35265 3995
rect 35299 3992 35311 3995
rect 35894 3992 35900 4004
rect 35299 3964 35900 3992
rect 35299 3961 35311 3964
rect 35253 3955 35311 3961
rect 35894 3952 35900 3964
rect 35952 3952 35958 4004
rect 33612 3924 33640 3952
rect 31726 3896 33640 3924
rect 33870 3884 33876 3936
rect 33928 3884 33934 3936
rect 44358 3884 44364 3936
rect 44416 3884 44422 3936
rect 1104 3834 45816 3856
rect 1104 3782 6539 3834
rect 6591 3782 6603 3834
rect 6655 3782 6667 3834
rect 6719 3782 6731 3834
rect 6783 3782 6795 3834
rect 6847 3782 17717 3834
rect 17769 3782 17781 3834
rect 17833 3782 17845 3834
rect 17897 3782 17909 3834
rect 17961 3782 17973 3834
rect 18025 3782 28895 3834
rect 28947 3782 28959 3834
rect 29011 3782 29023 3834
rect 29075 3782 29087 3834
rect 29139 3782 29151 3834
rect 29203 3782 40073 3834
rect 40125 3782 40137 3834
rect 40189 3782 40201 3834
rect 40253 3782 40265 3834
rect 40317 3782 40329 3834
rect 40381 3782 45816 3834
rect 1104 3760 45816 3782
rect 22005 3723 22063 3729
rect 22005 3689 22017 3723
rect 22051 3720 22063 3723
rect 22646 3720 22652 3732
rect 22051 3692 22652 3720
rect 22051 3689 22063 3692
rect 22005 3683 22063 3689
rect 22646 3680 22652 3692
rect 22704 3680 22710 3732
rect 33045 3723 33103 3729
rect 33045 3689 33057 3723
rect 33091 3720 33103 3723
rect 33686 3720 33692 3732
rect 33091 3692 33692 3720
rect 33091 3689 33103 3692
rect 33045 3683 33103 3689
rect 33686 3680 33692 3692
rect 33744 3680 33750 3732
rect 33870 3680 33876 3732
rect 33928 3720 33934 3732
rect 42794 3720 42800 3732
rect 33928 3692 42800 3720
rect 33928 3680 33934 3692
rect 42794 3680 42800 3692
rect 42852 3680 42858 3732
rect 24029 3655 24087 3661
rect 24029 3621 24041 3655
rect 24075 3652 24087 3655
rect 32214 3652 32220 3664
rect 24075 3624 32220 3652
rect 24075 3621 24087 3624
rect 24029 3615 24087 3621
rect 32214 3612 32220 3624
rect 32272 3612 32278 3664
rect 21358 3476 21364 3528
rect 21416 3516 21422 3528
rect 22189 3519 22247 3525
rect 22189 3516 22201 3519
rect 21416 3488 22201 3516
rect 21416 3476 21422 3488
rect 22189 3485 22201 3488
rect 22235 3485 22247 3519
rect 22189 3479 22247 3485
rect 23014 3476 23020 3528
rect 23072 3516 23078 3528
rect 23845 3519 23903 3525
rect 23845 3516 23857 3519
rect 23072 3488 23857 3516
rect 23072 3476 23078 3488
rect 23845 3485 23857 3488
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33229 3519 33287 3525
rect 33229 3516 33241 3519
rect 32456 3488 33241 3516
rect 32456 3476 32462 3488
rect 33229 3485 33241 3488
rect 33275 3485 33287 3519
rect 33229 3479 33287 3485
rect 23934 3408 23940 3460
rect 23992 3448 23998 3460
rect 33962 3448 33968 3460
rect 23992 3420 33968 3448
rect 23992 3408 23998 3420
rect 33962 3408 33968 3420
rect 34020 3408 34026 3460
rect 1104 3290 45976 3312
rect 1104 3238 12128 3290
rect 12180 3238 12192 3290
rect 12244 3238 12256 3290
rect 12308 3238 12320 3290
rect 12372 3238 12384 3290
rect 12436 3238 23306 3290
rect 23358 3238 23370 3290
rect 23422 3238 23434 3290
rect 23486 3238 23498 3290
rect 23550 3238 23562 3290
rect 23614 3238 34484 3290
rect 34536 3238 34548 3290
rect 34600 3238 34612 3290
rect 34664 3238 34676 3290
rect 34728 3238 34740 3290
rect 34792 3238 45662 3290
rect 45714 3238 45726 3290
rect 45778 3238 45790 3290
rect 45842 3238 45854 3290
rect 45906 3238 45918 3290
rect 45970 3238 45976 3290
rect 1104 3216 45976 3238
rect 23014 3136 23020 3188
rect 23072 3136 23078 3188
rect 23198 3136 23204 3188
rect 23256 3176 23262 3188
rect 23293 3179 23351 3185
rect 23293 3176 23305 3179
rect 23256 3148 23305 3176
rect 23256 3136 23262 3148
rect 23293 3145 23305 3148
rect 23339 3145 23351 3179
rect 23293 3139 23351 3145
rect 26421 3179 26479 3185
rect 26421 3145 26433 3179
rect 26467 3176 26479 3179
rect 27062 3176 27068 3188
rect 26467 3148 27068 3176
rect 26467 3145 26479 3148
rect 26421 3139 26479 3145
rect 27062 3136 27068 3148
rect 27120 3136 27126 3188
rect 39577 3179 39635 3185
rect 39577 3145 39589 3179
rect 39623 3176 39635 3179
rect 44542 3176 44548 3188
rect 39623 3148 44548 3176
rect 39623 3145 39635 3148
rect 39577 3139 39635 3145
rect 44542 3136 44548 3148
rect 44600 3136 44606 3188
rect 19242 3000 19248 3052
rect 19300 3040 19306 3052
rect 23201 3043 23259 3049
rect 23201 3040 23213 3043
rect 19300 3012 23213 3040
rect 19300 3000 19306 3012
rect 23201 3009 23213 3012
rect 23247 3009 23259 3043
rect 23201 3003 23259 3009
rect 23477 3043 23535 3049
rect 23477 3009 23489 3043
rect 23523 3009 23535 3043
rect 23477 3003 23535 3009
rect 23492 2972 23520 3003
rect 23566 3000 23572 3052
rect 23624 3000 23630 3052
rect 25774 3000 25780 3052
rect 25832 3040 25838 3052
rect 26605 3043 26663 3049
rect 26605 3040 26617 3043
rect 25832 3012 26617 3040
rect 25832 3000 25838 3012
rect 26605 3009 26617 3012
rect 26651 3009 26663 3043
rect 26605 3003 26663 3009
rect 29270 3000 29276 3052
rect 29328 3000 29334 3052
rect 39022 3000 39028 3052
rect 39080 3040 39086 3052
rect 39761 3043 39819 3049
rect 39761 3040 39773 3043
rect 39080 3012 39773 3040
rect 39080 3000 39086 3012
rect 39761 3009 39773 3012
rect 39807 3009 39819 3043
rect 39761 3003 39819 3009
rect 23658 2972 23664 2984
rect 23492 2944 23664 2972
rect 23658 2932 23664 2944
rect 23716 2932 23722 2984
rect 40954 2972 40960 2984
rect 23768 2944 40960 2972
rect 23768 2913 23796 2944
rect 40954 2932 40960 2944
rect 41012 2932 41018 2984
rect 23753 2907 23811 2913
rect 23753 2873 23765 2907
rect 23799 2873 23811 2907
rect 23753 2867 23811 2873
rect 29457 2907 29515 2913
rect 29457 2873 29469 2907
rect 29503 2904 29515 2907
rect 41414 2904 41420 2916
rect 29503 2876 41420 2904
rect 29503 2873 29515 2876
rect 29457 2867 29515 2873
rect 41414 2864 41420 2876
rect 41472 2864 41478 2916
rect 1104 2746 45816 2768
rect 1104 2694 6539 2746
rect 6591 2694 6603 2746
rect 6655 2694 6667 2746
rect 6719 2694 6731 2746
rect 6783 2694 6795 2746
rect 6847 2694 17717 2746
rect 17769 2694 17781 2746
rect 17833 2694 17845 2746
rect 17897 2694 17909 2746
rect 17961 2694 17973 2746
rect 18025 2694 28895 2746
rect 28947 2694 28959 2746
rect 29011 2694 29023 2746
rect 29075 2694 29087 2746
rect 29139 2694 29151 2746
rect 29203 2694 40073 2746
rect 40125 2694 40137 2746
rect 40189 2694 40201 2746
rect 40253 2694 40265 2746
rect 40317 2694 40329 2746
rect 40381 2694 45816 2746
rect 1104 2672 45816 2694
rect 23201 2635 23259 2641
rect 23201 2601 23213 2635
rect 23247 2632 23259 2635
rect 28629 2635 28687 2641
rect 23247 2604 28580 2632
rect 23247 2601 23259 2604
rect 23201 2595 23259 2601
rect 22741 2567 22799 2573
rect 22741 2533 22753 2567
rect 22787 2564 22799 2567
rect 23566 2564 23572 2576
rect 22787 2536 23572 2564
rect 22787 2533 22799 2536
rect 22741 2527 22799 2533
rect 23566 2524 23572 2536
rect 23624 2524 23630 2576
rect 24029 2567 24087 2573
rect 24029 2533 24041 2567
rect 24075 2564 24087 2567
rect 24946 2564 24952 2576
rect 24075 2536 24952 2564
rect 24075 2533 24087 2536
rect 24029 2527 24087 2533
rect 24946 2524 24952 2536
rect 25004 2524 25010 2576
rect 25041 2567 25099 2573
rect 25041 2533 25053 2567
rect 25087 2564 25099 2567
rect 28552 2564 28580 2604
rect 28629 2601 28641 2635
rect 28675 2632 28687 2635
rect 29270 2632 29276 2644
rect 28675 2604 29276 2632
rect 28675 2601 28687 2604
rect 28629 2595 28687 2601
rect 29270 2592 29276 2604
rect 29328 2592 29334 2644
rect 44174 2592 44180 2644
rect 44232 2592 44238 2644
rect 44637 2635 44695 2641
rect 44637 2601 44649 2635
rect 44683 2632 44695 2635
rect 44910 2632 44916 2644
rect 44683 2604 44916 2632
rect 44683 2601 44695 2604
rect 44637 2595 44695 2601
rect 44910 2592 44916 2604
rect 44968 2592 44974 2644
rect 45002 2592 45008 2644
rect 45060 2592 45066 2644
rect 41874 2564 41880 2576
rect 25087 2536 26234 2564
rect 28552 2536 41880 2564
rect 25087 2533 25099 2536
rect 25041 2527 25099 2533
rect 26206 2496 26234 2536
rect 41874 2524 41880 2536
rect 41932 2524 41938 2576
rect 44192 2564 44220 2592
rect 45281 2567 45339 2573
rect 45281 2564 45293 2567
rect 44192 2536 45293 2564
rect 45281 2533 45293 2536
rect 45327 2533 45339 2567
rect 45281 2527 45339 2533
rect 37366 2496 37372 2508
rect 26206 2468 37372 2496
rect 37366 2456 37372 2468
rect 37424 2456 37430 2508
rect 44266 2496 44272 2508
rect 40052 2468 44272 2496
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 22925 2431 22983 2437
rect 22925 2428 22937 2431
rect 20772 2400 22937 2428
rect 20772 2388 20778 2400
rect 22925 2397 22937 2400
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 23014 2388 23020 2440
rect 23072 2388 23078 2440
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23385 2431 23443 2437
rect 23385 2428 23397 2431
rect 23256 2400 23397 2428
rect 23256 2388 23262 2400
rect 23385 2397 23397 2400
rect 23431 2397 23443 2431
rect 23385 2391 23443 2397
rect 23842 2388 23848 2440
rect 23900 2388 23906 2440
rect 24854 2388 24860 2440
rect 24912 2388 24918 2440
rect 28810 2388 28816 2440
rect 28868 2388 28874 2440
rect 31478 2388 31484 2440
rect 31536 2388 31542 2440
rect 38194 2388 38200 2440
rect 38252 2388 38258 2440
rect 20622 2320 20628 2372
rect 20680 2320 20686 2372
rect 20809 2363 20867 2369
rect 20809 2329 20821 2363
rect 20855 2360 20867 2363
rect 35526 2360 35532 2372
rect 20855 2332 35532 2360
rect 20855 2329 20867 2332
rect 20809 2323 20867 2329
rect 35526 2320 35532 2332
rect 35584 2320 35590 2372
rect 40052 2360 40080 2468
rect 44266 2456 44272 2468
rect 44324 2456 44330 2508
rect 41782 2388 41788 2440
rect 41840 2428 41846 2440
rect 44821 2431 44879 2437
rect 44821 2428 44833 2431
rect 41840 2400 44833 2428
rect 41840 2388 41846 2400
rect 44821 2397 44833 2400
rect 44867 2397 44879 2431
rect 44821 2391 44879 2397
rect 45189 2431 45247 2437
rect 45189 2397 45201 2431
rect 45235 2397 45247 2431
rect 45189 2391 45247 2397
rect 35866 2332 40080 2360
rect 23569 2295 23627 2301
rect 23569 2261 23581 2295
rect 23615 2292 23627 2295
rect 23934 2292 23940 2304
rect 23615 2264 23940 2292
rect 23615 2261 23627 2264
rect 23569 2255 23627 2261
rect 23934 2252 23940 2264
rect 23992 2252 23998 2304
rect 31665 2295 31723 2301
rect 31665 2261 31677 2295
rect 31711 2292 31723 2295
rect 35866 2292 35894 2332
rect 43898 2320 43904 2372
rect 43956 2360 43962 2372
rect 45204 2360 45232 2391
rect 45462 2388 45468 2440
rect 45520 2388 45526 2440
rect 43956 2332 45232 2360
rect 43956 2320 43962 2332
rect 31711 2264 35894 2292
rect 38381 2295 38439 2301
rect 31711 2261 31723 2264
rect 31665 2255 31723 2261
rect 38381 2261 38393 2295
rect 38427 2292 38439 2295
rect 45094 2292 45100 2304
rect 38427 2264 45100 2292
rect 38427 2261 38439 2264
rect 38381 2255 38439 2261
rect 45094 2252 45100 2264
rect 45152 2252 45158 2304
rect 1104 2202 45976 2224
rect 1104 2150 12128 2202
rect 12180 2150 12192 2202
rect 12244 2150 12256 2202
rect 12308 2150 12320 2202
rect 12372 2150 12384 2202
rect 12436 2150 23306 2202
rect 23358 2150 23370 2202
rect 23422 2150 23434 2202
rect 23486 2150 23498 2202
rect 23550 2150 23562 2202
rect 23614 2150 34484 2202
rect 34536 2150 34548 2202
rect 34600 2150 34612 2202
rect 34664 2150 34676 2202
rect 34728 2150 34740 2202
rect 34792 2150 45662 2202
rect 45714 2150 45726 2202
rect 45778 2150 45790 2202
rect 45842 2150 45854 2202
rect 45906 2150 45918 2202
rect 45970 2150 45976 2202
rect 1104 2128 45976 2150
rect 19613 2091 19671 2097
rect 19613 2057 19625 2091
rect 19659 2088 19671 2091
rect 20622 2088 20628 2100
rect 19659 2060 20628 2088
rect 19659 2057 19671 2060
rect 19613 2051 19671 2057
rect 20622 2048 20628 2060
rect 20680 2048 20686 2100
rect 22189 2091 22247 2097
rect 22189 2057 22201 2091
rect 22235 2088 22247 2091
rect 23014 2088 23020 2100
rect 22235 2060 23020 2088
rect 22235 2057 22247 2060
rect 22189 2051 22247 2057
rect 23014 2048 23020 2060
rect 23072 2048 23078 2100
rect 23106 2048 23112 2100
rect 23164 2048 23170 2100
rect 23198 2048 23204 2100
rect 23256 2088 23262 2100
rect 23293 2091 23351 2097
rect 23293 2088 23305 2091
rect 23256 2060 23305 2088
rect 23256 2048 23262 2060
rect 23293 2057 23305 2060
rect 23339 2057 23351 2091
rect 23293 2051 23351 2057
rect 23842 2048 23848 2100
rect 23900 2048 23906 2100
rect 24213 2091 24271 2097
rect 24213 2057 24225 2091
rect 24259 2088 24271 2091
rect 24854 2088 24860 2100
rect 24259 2060 24860 2088
rect 24259 2057 24271 2060
rect 24213 2051 24271 2057
rect 24854 2048 24860 2060
rect 24912 2048 24918 2100
rect 30837 2091 30895 2097
rect 30837 2057 30849 2091
rect 30883 2088 30895 2091
rect 31478 2088 31484 2100
rect 30883 2060 31484 2088
rect 30883 2057 30895 2060
rect 30837 2051 30895 2057
rect 31478 2048 31484 2060
rect 31536 2048 31542 2100
rect 37277 2091 37335 2097
rect 37277 2057 37289 2091
rect 37323 2088 37335 2091
rect 38194 2088 38200 2100
rect 37323 2060 38200 2088
rect 37323 2057 37335 2060
rect 37277 2051 37335 2057
rect 38194 2048 38200 2060
rect 38252 2048 38258 2100
rect 41782 2048 41788 2100
rect 41840 2048 41846 2100
rect 43898 2048 43904 2100
rect 43956 2048 43962 2100
rect 44637 2091 44695 2097
rect 44637 2057 44649 2091
rect 44683 2088 44695 2091
rect 45462 2088 45468 2100
rect 44683 2060 45468 2088
rect 44683 2057 44695 2060
rect 44637 2051 44695 2057
rect 45462 2048 45468 2060
rect 45520 2048 45526 2100
rect 22741 2023 22799 2029
rect 22741 1989 22753 2023
rect 22787 2020 22799 2023
rect 23124 2020 23152 2048
rect 22787 1992 23152 2020
rect 22787 1989 22799 1992
rect 22741 1983 22799 1989
rect 19794 1912 19800 1964
rect 19852 1912 19858 1964
rect 20898 1912 20904 1964
rect 20956 1952 20962 1964
rect 22373 1955 22431 1961
rect 22373 1952 22385 1955
rect 20956 1924 22385 1952
rect 20956 1912 20962 1924
rect 22373 1921 22385 1924
rect 22419 1921 22431 1955
rect 22373 1915 22431 1921
rect 22557 1955 22615 1961
rect 22557 1921 22569 1955
rect 22603 1921 22615 1955
rect 22557 1915 22615 1921
rect 1670 1844 1676 1896
rect 1728 1884 1734 1896
rect 22572 1884 22600 1915
rect 23198 1912 23204 1964
rect 23256 1912 23262 1964
rect 23477 1955 23535 1961
rect 23477 1921 23489 1955
rect 23523 1921 23535 1955
rect 23477 1915 23535 1921
rect 1728 1856 22600 1884
rect 1728 1844 1734 1856
rect 22646 1844 22652 1896
rect 22704 1884 22710 1896
rect 23492 1884 23520 1915
rect 22704 1856 23520 1884
rect 22704 1844 22710 1856
rect 23017 1819 23075 1825
rect 23017 1785 23029 1819
rect 23063 1816 23075 1819
rect 23860 1816 23888 2048
rect 24394 1912 24400 1964
rect 24452 1912 24458 1964
rect 31018 1912 31024 1964
rect 31076 1912 31082 1964
rect 37458 1912 37464 1964
rect 37516 1912 37522 1964
rect 41966 1912 41972 1964
rect 42024 1912 42030 1964
rect 44082 1912 44088 1964
rect 44140 1912 44146 1964
rect 44818 1912 44824 1964
rect 44876 1912 44882 1964
rect 23063 1788 23888 1816
rect 23063 1785 23075 1788
rect 23017 1779 23075 1785
rect 1104 1658 45816 1680
rect 1104 1606 6539 1658
rect 6591 1606 6603 1658
rect 6655 1606 6667 1658
rect 6719 1606 6731 1658
rect 6783 1606 6795 1658
rect 6847 1606 17717 1658
rect 17769 1606 17781 1658
rect 17833 1606 17845 1658
rect 17897 1606 17909 1658
rect 17961 1606 17973 1658
rect 18025 1606 28895 1658
rect 28947 1606 28959 1658
rect 29011 1606 29023 1658
rect 29075 1606 29087 1658
rect 29139 1606 29151 1658
rect 29203 1606 40073 1658
rect 40125 1606 40137 1658
rect 40189 1606 40201 1658
rect 40253 1606 40265 1658
rect 40317 1606 40329 1658
rect 40381 1606 45816 1658
rect 1104 1584 45816 1606
rect 1670 1504 1676 1556
rect 1728 1504 1734 1556
rect 19245 1547 19303 1553
rect 19245 1513 19257 1547
rect 19291 1544 19303 1547
rect 19794 1544 19800 1556
rect 19291 1516 19800 1544
rect 19291 1513 19303 1516
rect 19245 1507 19303 1513
rect 19794 1504 19800 1516
rect 19852 1504 19858 1556
rect 23569 1547 23627 1553
rect 23569 1513 23581 1547
rect 23615 1544 23627 1547
rect 24394 1544 24400 1556
rect 23615 1516 24400 1544
rect 23615 1513 23627 1516
rect 23569 1507 23627 1513
rect 24394 1504 24400 1516
rect 24452 1504 24458 1556
rect 27985 1547 28043 1553
rect 27985 1513 27997 1547
rect 28031 1544 28043 1547
rect 28810 1544 28816 1556
rect 28031 1516 28816 1544
rect 28031 1513 28043 1516
rect 27985 1507 28043 1513
rect 28810 1504 28816 1516
rect 28868 1504 28874 1556
rect 30193 1547 30251 1553
rect 30193 1513 30205 1547
rect 30239 1544 30251 1547
rect 31018 1544 31024 1556
rect 30239 1516 31024 1544
rect 30239 1513 30251 1516
rect 30193 1507 30251 1513
rect 31018 1504 31024 1516
rect 31076 1504 31082 1556
rect 41233 1547 41291 1553
rect 41233 1513 41245 1547
rect 41279 1544 41291 1547
rect 41966 1544 41972 1556
rect 41279 1516 41972 1544
rect 41279 1513 41291 1516
rect 41233 1507 41291 1513
rect 41966 1504 41972 1516
rect 42024 1504 42030 1556
rect 43441 1547 43499 1553
rect 43441 1513 43453 1547
rect 43487 1544 43499 1547
rect 44082 1544 44088 1556
rect 43487 1516 44088 1544
rect 43487 1513 43499 1516
rect 43441 1507 43499 1513
rect 44082 1504 44088 1516
rect 44140 1504 44146 1556
rect 44818 1504 44824 1556
rect 44876 1544 44882 1556
rect 45281 1547 45339 1553
rect 45281 1544 45293 1547
rect 44876 1516 45293 1544
rect 44876 1504 44882 1516
rect 45281 1513 45293 1516
rect 45327 1513 45339 1547
rect 45281 1507 45339 1513
rect 1486 1300 1492 1352
rect 1544 1300 1550 1352
rect 3786 1300 3792 1352
rect 3844 1300 3850 1352
rect 5902 1300 5908 1352
rect 5960 1300 5966 1352
rect 8110 1300 8116 1352
rect 8168 1300 8174 1352
rect 10318 1300 10324 1352
rect 10376 1300 10382 1352
rect 12526 1300 12532 1352
rect 12584 1300 12590 1352
rect 14734 1300 14740 1352
rect 14792 1300 14798 1352
rect 16546 1312 17080 1340
rect 16546 1272 16574 1312
rect 3988 1244 11744 1272
rect 3988 1213 4016 1244
rect 11716 1216 11744 1244
rect 12728 1244 16574 1272
rect 17052 1272 17080 1312
rect 17126 1300 17132 1352
rect 17184 1300 17190 1352
rect 19426 1300 19432 1352
rect 19484 1300 19490 1352
rect 20714 1300 20720 1352
rect 20772 1300 20778 1352
rect 21542 1300 21548 1352
rect 21600 1300 21606 1352
rect 23750 1300 23756 1352
rect 23808 1300 23814 1352
rect 25958 1300 25964 1352
rect 26016 1300 26022 1352
rect 28166 1300 28172 1352
rect 28224 1300 28230 1352
rect 30374 1300 30380 1352
rect 30432 1300 30438 1352
rect 32582 1300 32588 1352
rect 32640 1300 32646 1352
rect 34882 1300 34888 1352
rect 34940 1300 34946 1352
rect 35434 1300 35440 1352
rect 35492 1300 35498 1352
rect 36998 1300 37004 1352
rect 37056 1300 37062 1352
rect 37458 1300 37464 1352
rect 37516 1300 37522 1352
rect 39206 1300 39212 1352
rect 39264 1300 39270 1352
rect 41414 1300 41420 1352
rect 41472 1300 41478 1352
rect 43622 1300 43628 1352
rect 43680 1300 43686 1352
rect 45465 1343 45523 1349
rect 45465 1309 45477 1343
rect 45511 1340 45523 1343
rect 45554 1340 45560 1352
rect 45511 1312 45560 1340
rect 45511 1309 45523 1312
rect 45465 1303 45523 1309
rect 45554 1300 45560 1312
rect 45612 1300 45618 1352
rect 20732 1272 20760 1300
rect 17052 1244 20760 1272
rect 3973 1207 4031 1213
rect 3973 1173 3985 1207
rect 4019 1173 4031 1207
rect 3973 1167 4031 1173
rect 6086 1164 6092 1216
rect 6144 1164 6150 1216
rect 8294 1164 8300 1216
rect 8352 1164 8358 1216
rect 10502 1164 10508 1216
rect 10560 1164 10566 1216
rect 11698 1164 11704 1216
rect 11756 1164 11762 1216
rect 12728 1213 12756 1244
rect 20898 1232 20904 1284
rect 20956 1232 20962 1284
rect 12713 1207 12771 1213
rect 12713 1173 12725 1207
rect 12759 1173 12771 1207
rect 12713 1167 12771 1173
rect 14921 1207 14979 1213
rect 14921 1173 14933 1207
rect 14967 1204 14979 1207
rect 16850 1204 16856 1216
rect 14967 1176 16856 1204
rect 14967 1173 14979 1176
rect 14921 1167 14979 1173
rect 16850 1164 16856 1176
rect 16908 1164 16914 1216
rect 16945 1207 17003 1213
rect 16945 1173 16957 1207
rect 16991 1204 17003 1207
rect 20916 1204 20944 1232
rect 16991 1176 20944 1204
rect 16991 1173 17003 1176
rect 16945 1167 17003 1173
rect 21358 1164 21364 1216
rect 21416 1164 21422 1216
rect 25774 1164 25780 1216
rect 25832 1164 25838 1216
rect 32398 1164 32404 1216
rect 32456 1164 32462 1216
rect 34701 1207 34759 1213
rect 34701 1173 34713 1207
rect 34747 1204 34759 1207
rect 35452 1204 35480 1300
rect 34747 1176 35480 1204
rect 36817 1207 36875 1213
rect 34747 1173 34759 1176
rect 34701 1167 34759 1173
rect 36817 1173 36829 1207
rect 36863 1204 36875 1207
rect 37476 1204 37504 1300
rect 36863 1176 37504 1204
rect 36863 1173 36875 1176
rect 36817 1167 36875 1173
rect 39022 1164 39028 1216
rect 39080 1164 39086 1216
rect 1104 1114 45976 1136
rect 1104 1062 12128 1114
rect 12180 1062 12192 1114
rect 12244 1062 12256 1114
rect 12308 1062 12320 1114
rect 12372 1062 12384 1114
rect 12436 1062 23306 1114
rect 23358 1062 23370 1114
rect 23422 1062 23434 1114
rect 23486 1062 23498 1114
rect 23550 1062 23562 1114
rect 23614 1062 34484 1114
rect 34536 1062 34548 1114
rect 34600 1062 34612 1114
rect 34664 1062 34676 1114
rect 34728 1062 34740 1114
rect 34792 1062 45662 1114
rect 45714 1062 45726 1114
rect 45778 1062 45790 1114
rect 45842 1062 45854 1114
rect 45906 1062 45918 1114
rect 45970 1062 45976 1114
rect 1104 1040 45976 1062
rect 6086 960 6092 1012
rect 6144 1000 6150 1012
rect 6144 972 6914 1000
rect 6144 960 6150 972
rect 6886 796 6914 972
rect 10502 960 10508 1012
rect 10560 1000 10566 1012
rect 10560 972 16804 1000
rect 10560 960 10566 972
rect 11698 892 11704 944
rect 11756 932 11762 944
rect 16574 932 16580 944
rect 11756 904 16580 932
rect 11756 892 11762 904
rect 16574 892 16580 904
rect 16632 892 16638 944
rect 16776 932 16804 972
rect 16850 960 16856 1012
rect 16908 1000 16914 1012
rect 22646 1000 22652 1012
rect 16908 972 22652 1000
rect 16908 960 16914 972
rect 22646 960 22652 972
rect 22704 960 22710 1012
rect 19242 932 19248 944
rect 16776 904 19248 932
rect 19242 892 19248 904
rect 19300 892 19306 944
rect 20806 824 20812 876
rect 20864 824 20870 876
rect 20824 796 20852 824
rect 6886 768 20852 796
rect 8294 688 8300 740
rect 8352 688 8358 740
rect 16574 688 16580 740
rect 16632 728 16638 740
rect 23198 728 23204 740
rect 16632 700 23204 728
rect 16632 688 16638 700
rect 23198 688 23204 700
rect 23256 688 23262 740
rect 8312 660 8340 688
rect 23658 660 23664 672
rect 8312 632 23664 660
rect 23658 620 23664 632
rect 23716 620 23722 672
<< via1 >>
rect 18144 9936 18196 9988
rect 21824 9936 21876 9988
rect 22652 9936 22704 9988
rect 32956 9936 33008 9988
rect 9956 9868 10008 9920
rect 17408 9868 17460 9920
rect 17500 9868 17552 9920
rect 9404 9800 9456 9852
rect 21456 9800 21508 9852
rect 24492 9800 24544 9852
rect 7196 9732 7248 9784
rect 9680 9732 9732 9784
rect 13084 9732 13136 9784
rect 21732 9732 21784 9784
rect 4436 9664 4488 9716
rect 21548 9664 21600 9716
rect 9404 9596 9456 9648
rect 11612 9528 11664 9580
rect 21732 9596 21784 9648
rect 12716 9528 12768 9580
rect 21364 9528 21416 9580
rect 4068 9460 4120 9512
rect 9036 9460 9088 9512
rect 21732 9460 21784 9512
rect 21824 9460 21876 9512
rect 23940 9460 23992 9512
rect 38844 9528 38896 9580
rect 8300 9324 8352 9376
rect 16580 9324 16632 9376
rect 17408 9324 17460 9376
rect 23664 9324 23716 9376
rect 32864 9392 32916 9444
rect 26148 9324 26200 9376
rect 26240 9324 26292 9376
rect 35164 9324 35216 9376
rect 1492 9188 1544 9240
rect 16764 9256 16816 9308
rect 27804 9256 27856 9308
rect 17500 9188 17552 9240
rect 10416 9120 10468 9172
rect 7564 9052 7616 9104
rect 17132 9120 17184 9172
rect 12624 9052 12676 9104
rect 19616 9188 19668 9240
rect 22100 9188 22152 9240
rect 24400 9188 24452 9240
rect 24768 9188 24820 9240
rect 31024 9188 31076 9240
rect 32220 9188 32272 9240
rect 40960 9188 41012 9240
rect 20812 9120 20864 9172
rect 18052 9052 18104 9104
rect 18236 9052 18288 9104
rect 21732 9120 21784 9172
rect 35900 9120 35952 9172
rect 37372 9120 37424 9172
rect 43444 9120 43496 9172
rect 32772 9052 32824 9104
rect 35532 9052 35584 9104
rect 13728 8984 13780 9036
rect 10508 8916 10560 8968
rect 16672 8984 16724 9036
rect 16948 8984 17000 9036
rect 21088 8984 21140 9036
rect 21456 8984 21508 9036
rect 24124 8984 24176 9036
rect 33968 8984 34020 9036
rect 40684 8984 40736 9036
rect 14096 8916 14148 8968
rect 23020 8916 23072 8968
rect 30288 8916 30340 8968
rect 33600 8916 33652 8968
rect 38108 8916 38160 8968
rect 24032 8848 24084 8900
rect 24308 8848 24360 8900
rect 27252 8848 27304 8900
rect 30932 8848 30984 8900
rect 3332 8780 3384 8832
rect 7012 8780 7064 8832
rect 7104 8780 7156 8832
rect 9772 8780 9824 8832
rect 11520 8780 11572 8832
rect 15108 8780 15160 8832
rect 17040 8780 17092 8832
rect 22100 8780 22152 8832
rect 22652 8780 22704 8832
rect 37188 8848 37240 8900
rect 31852 8780 31904 8832
rect 37740 8780 37792 8832
rect 42432 8780 42484 8832
rect 12128 8678 12180 8730
rect 12192 8678 12244 8730
rect 12256 8678 12308 8730
rect 12320 8678 12372 8730
rect 12384 8678 12436 8730
rect 23306 8678 23358 8730
rect 23370 8678 23422 8730
rect 23434 8678 23486 8730
rect 23498 8678 23550 8730
rect 23562 8678 23614 8730
rect 34484 8678 34536 8730
rect 34548 8678 34600 8730
rect 34612 8678 34664 8730
rect 34676 8678 34728 8730
rect 34740 8678 34792 8730
rect 45662 8678 45714 8730
rect 45726 8678 45778 8730
rect 45790 8678 45842 8730
rect 45854 8678 45906 8730
rect 45918 8678 45970 8730
rect 2504 8576 2556 8628
rect 2872 8576 2924 8628
rect 3240 8576 3292 8628
rect 3608 8576 3660 8628
rect 4344 8576 4396 8628
rect 5080 8576 5132 8628
rect 5448 8576 5500 8628
rect 6184 8576 6236 8628
rect 6828 8619 6880 8628
rect 6828 8585 6837 8619
rect 6837 8585 6871 8619
rect 6871 8585 6880 8619
rect 6828 8576 6880 8585
rect 7656 8576 7708 8628
rect 8024 8576 8076 8628
rect 8392 8576 8444 8628
rect 8760 8576 8812 8628
rect 9496 8576 9548 8628
rect 9864 8576 9916 8628
rect 10600 8576 10652 8628
rect 10968 8576 11020 8628
rect 11336 8576 11388 8628
rect 11980 8576 12032 8628
rect 12440 8576 12492 8628
rect 2688 8508 2740 8560
rect 4068 8508 4120 8560
rect 1492 8483 1544 8492
rect 1492 8449 1501 8483
rect 1501 8449 1535 8483
rect 1535 8449 1544 8483
rect 1492 8440 1544 8449
rect 2964 8483 3016 8492
rect 2964 8449 2973 8483
rect 2973 8449 3007 8483
rect 3007 8449 3016 8483
rect 2964 8440 3016 8449
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 7104 8440 7156 8492
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 8300 8440 8352 8492
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 9772 8440 9824 8492
rect 9956 8483 10008 8492
rect 9956 8449 9965 8483
rect 9965 8449 9999 8483
rect 9999 8449 10008 8483
rect 9956 8440 10008 8449
rect 10416 8551 10468 8560
rect 10416 8517 10425 8551
rect 10425 8517 10459 8551
rect 10459 8517 10468 8551
rect 10416 8508 10468 8517
rect 12624 8576 12676 8628
rect 13176 8576 13228 8628
rect 13544 8576 13596 8628
rect 13912 8576 13964 8628
rect 14648 8576 14700 8628
rect 15016 8576 15068 8628
rect 15384 8576 15436 8628
rect 16120 8576 16172 8628
rect 16488 8576 16540 8628
rect 16764 8576 16816 8628
rect 16856 8576 16908 8628
rect 17224 8576 17276 8628
rect 17592 8576 17644 8628
rect 17960 8576 18012 8628
rect 18696 8576 18748 8628
rect 19524 8619 19576 8628
rect 19524 8585 19533 8619
rect 19533 8585 19567 8619
rect 19567 8585 19576 8619
rect 19524 8576 19576 8585
rect 11520 8440 11572 8492
rect 11612 8483 11664 8492
rect 11612 8449 11621 8483
rect 11621 8449 11655 8483
rect 11655 8449 11664 8483
rect 11612 8440 11664 8449
rect 12716 8483 12768 8492
rect 12716 8449 12725 8483
rect 12725 8449 12759 8483
rect 12759 8449 12768 8483
rect 12716 8440 12768 8449
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 14096 8440 14148 8492
rect 14464 8440 14516 8492
rect 14924 8440 14976 8492
rect 15568 8440 15620 8492
rect 16028 8440 16080 8492
rect 16856 8440 16908 8492
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 18512 8508 18564 8560
rect 19340 8508 19392 8560
rect 21824 8576 21876 8628
rect 22468 8619 22520 8628
rect 22468 8585 22477 8619
rect 22477 8585 22511 8619
rect 22511 8585 22520 8619
rect 22468 8576 22520 8585
rect 23020 8619 23072 8628
rect 23020 8585 23029 8619
rect 23029 8585 23063 8619
rect 23063 8585 23072 8619
rect 23020 8576 23072 8585
rect 17592 8440 17644 8492
rect 8208 8304 8260 8356
rect 10508 8372 10560 8424
rect 8392 8304 8444 8356
rect 17040 8304 17092 8356
rect 17500 8372 17552 8424
rect 18788 8483 18840 8492
rect 18788 8449 18797 8483
rect 18797 8449 18831 8483
rect 18831 8449 18840 8483
rect 18788 8440 18840 8449
rect 19432 8483 19484 8492
rect 19432 8449 19441 8483
rect 19441 8449 19475 8483
rect 19475 8449 19484 8483
rect 19432 8440 19484 8449
rect 19984 8483 20036 8492
rect 19984 8449 19993 8483
rect 19993 8449 20027 8483
rect 20027 8449 20036 8483
rect 19984 8440 20036 8449
rect 21272 8508 21324 8560
rect 22008 8508 22060 8560
rect 22744 8508 22796 8560
rect 19340 8372 19392 8424
rect 21456 8372 21508 8424
rect 22192 8372 22244 8424
rect 22652 8483 22704 8492
rect 22652 8449 22661 8483
rect 22661 8449 22695 8483
rect 22695 8449 22704 8483
rect 22652 8440 22704 8449
rect 23296 8508 23348 8560
rect 23940 8576 23992 8628
rect 24032 8619 24084 8628
rect 24032 8585 24041 8619
rect 24041 8585 24075 8619
rect 24075 8585 24084 8619
rect 24032 8576 24084 8585
rect 23480 8483 23532 8492
rect 23480 8449 23489 8483
rect 23489 8449 23523 8483
rect 23523 8449 23532 8483
rect 23480 8440 23532 8449
rect 27252 8576 27304 8628
rect 27344 8576 27396 8628
rect 25136 8508 25188 8560
rect 30288 8576 30340 8628
rect 30932 8619 30984 8628
rect 30932 8585 30941 8619
rect 30941 8585 30975 8619
rect 30975 8585 30984 8619
rect 30932 8576 30984 8585
rect 31024 8576 31076 8628
rect 32772 8576 32824 8628
rect 32864 8508 32916 8560
rect 35164 8619 35216 8628
rect 35164 8585 35173 8619
rect 35173 8585 35207 8619
rect 35207 8585 35216 8619
rect 35164 8576 35216 8585
rect 23112 8372 23164 8424
rect 24216 8440 24268 8492
rect 24860 8483 24912 8492
rect 24860 8449 24869 8483
rect 24869 8449 24903 8483
rect 24903 8449 24912 8483
rect 24860 8440 24912 8449
rect 24952 8440 25004 8492
rect 25320 8440 25372 8492
rect 25688 8440 25740 8492
rect 26056 8440 26108 8492
rect 26424 8440 26476 8492
rect 26792 8440 26844 8492
rect 27436 8483 27488 8492
rect 27436 8449 27445 8483
rect 27445 8449 27479 8483
rect 27479 8449 27488 8483
rect 27436 8440 27488 8449
rect 27528 8440 27580 8492
rect 27896 8440 27948 8492
rect 28264 8440 28316 8492
rect 28632 8440 28684 8492
rect 29000 8440 29052 8492
rect 29368 8440 29420 8492
rect 30012 8483 30064 8492
rect 30012 8449 30021 8483
rect 30021 8449 30055 8483
rect 30055 8449 30064 8483
rect 30012 8440 30064 8449
rect 30104 8440 30156 8492
rect 30472 8440 30524 8492
rect 30840 8440 30892 8492
rect 31208 8440 31260 8492
rect 31668 8483 31720 8492
rect 31668 8449 31677 8483
rect 31677 8449 31711 8483
rect 31711 8449 31720 8483
rect 31668 8440 31720 8449
rect 32128 8483 32180 8492
rect 32128 8449 32137 8483
rect 32137 8449 32171 8483
rect 32171 8449 32180 8483
rect 32128 8440 32180 8449
rect 32404 8483 32456 8492
rect 32404 8449 32413 8483
rect 32413 8449 32447 8483
rect 32447 8449 32456 8483
rect 32404 8440 32456 8449
rect 32772 8483 32824 8492
rect 32772 8449 32781 8483
rect 32781 8449 32815 8483
rect 32815 8449 32824 8483
rect 32772 8440 32824 8449
rect 33048 8440 33100 8492
rect 33508 8483 33560 8492
rect 33508 8449 33517 8483
rect 33517 8449 33551 8483
rect 33551 8449 33560 8483
rect 33508 8440 33560 8449
rect 33876 8483 33928 8492
rect 33876 8449 33885 8483
rect 33885 8449 33919 8483
rect 33919 8449 33928 8483
rect 33876 8440 33928 8449
rect 34244 8483 34296 8492
rect 34244 8449 34253 8483
rect 34253 8449 34287 8483
rect 34287 8449 34296 8483
rect 34244 8440 34296 8449
rect 34336 8440 34388 8492
rect 34980 8483 35032 8492
rect 34980 8449 34989 8483
rect 34989 8449 35023 8483
rect 35023 8449 35032 8483
rect 34980 8440 35032 8449
rect 19616 8304 19668 8356
rect 14280 8236 14332 8288
rect 18696 8236 18748 8288
rect 19064 8236 19116 8288
rect 19892 8236 19944 8288
rect 20628 8279 20680 8288
rect 20628 8245 20637 8279
rect 20637 8245 20671 8279
rect 20671 8245 20680 8279
rect 20628 8236 20680 8245
rect 20904 8279 20956 8288
rect 20904 8245 20913 8279
rect 20913 8245 20947 8279
rect 20947 8245 20956 8279
rect 20904 8236 20956 8245
rect 21180 8279 21232 8288
rect 21180 8245 21189 8279
rect 21189 8245 21223 8279
rect 21223 8245 21232 8279
rect 21180 8236 21232 8245
rect 21456 8279 21508 8288
rect 21456 8245 21465 8279
rect 21465 8245 21499 8279
rect 21499 8245 21508 8279
rect 21456 8236 21508 8245
rect 22284 8304 22336 8356
rect 23756 8347 23808 8356
rect 23756 8313 23765 8347
rect 23765 8313 23799 8347
rect 23799 8313 23808 8347
rect 23756 8304 23808 8313
rect 22376 8236 22428 8288
rect 22744 8279 22796 8288
rect 22744 8245 22753 8279
rect 22753 8245 22787 8279
rect 22787 8245 22796 8279
rect 22744 8236 22796 8245
rect 23020 8236 23072 8288
rect 23388 8236 23440 8288
rect 24308 8304 24360 8356
rect 24492 8372 24544 8424
rect 23940 8236 23992 8288
rect 24768 8304 24820 8356
rect 26056 8304 26108 8356
rect 26792 8304 26844 8356
rect 24676 8279 24728 8288
rect 24676 8245 24685 8279
rect 24685 8245 24719 8279
rect 24719 8245 24728 8279
rect 24676 8236 24728 8245
rect 25044 8279 25096 8288
rect 25044 8245 25053 8279
rect 25053 8245 25087 8279
rect 25087 8245 25096 8279
rect 25044 8236 25096 8245
rect 25412 8279 25464 8288
rect 25412 8245 25421 8279
rect 25421 8245 25455 8279
rect 25455 8245 25464 8279
rect 25412 8236 25464 8245
rect 25596 8236 25648 8288
rect 25872 8236 25924 8288
rect 26424 8236 26476 8288
rect 27160 8304 27212 8356
rect 31760 8372 31812 8424
rect 37188 8576 37240 8628
rect 37740 8619 37792 8628
rect 37740 8585 37749 8619
rect 37749 8585 37783 8619
rect 37783 8585 37792 8619
rect 37740 8576 37792 8585
rect 38108 8576 38160 8628
rect 38844 8619 38896 8628
rect 38844 8585 38853 8619
rect 38853 8585 38887 8619
rect 38887 8585 38896 8619
rect 38844 8576 38896 8585
rect 38936 8576 38988 8628
rect 39304 8576 39356 8628
rect 39672 8576 39724 8628
rect 40132 8576 40184 8628
rect 40684 8576 40736 8628
rect 41144 8576 41196 8628
rect 41880 8576 41932 8628
rect 35348 8483 35400 8492
rect 35348 8449 35357 8483
rect 35357 8449 35391 8483
rect 35391 8449 35400 8483
rect 35348 8440 35400 8449
rect 27528 8236 27580 8288
rect 27896 8236 27948 8288
rect 28724 8279 28776 8288
rect 28724 8245 28733 8279
rect 28733 8245 28767 8279
rect 28767 8245 28776 8279
rect 28724 8236 28776 8245
rect 29276 8236 29328 8288
rect 29552 8279 29604 8288
rect 29552 8245 29561 8279
rect 29561 8245 29595 8279
rect 29595 8245 29604 8279
rect 29552 8236 29604 8245
rect 29828 8279 29880 8288
rect 29828 8245 29837 8279
rect 29837 8245 29871 8279
rect 29871 8245 29880 8279
rect 29828 8236 29880 8245
rect 30656 8304 30708 8356
rect 31944 8304 31996 8356
rect 34152 8304 34204 8356
rect 32956 8279 33008 8288
rect 32956 8245 32965 8279
rect 32965 8245 32999 8279
rect 32999 8245 33008 8279
rect 32956 8236 33008 8245
rect 33324 8279 33376 8288
rect 33324 8245 33333 8279
rect 33333 8245 33367 8279
rect 33367 8245 33376 8279
rect 33324 8236 33376 8245
rect 33692 8279 33744 8288
rect 33692 8245 33701 8279
rect 33701 8245 33735 8279
rect 33735 8245 33744 8279
rect 33692 8236 33744 8245
rect 33784 8236 33836 8288
rect 42248 8508 42300 8560
rect 43720 8576 43772 8628
rect 44824 8576 44876 8628
rect 35716 8483 35768 8492
rect 35716 8449 35725 8483
rect 35725 8449 35759 8483
rect 35759 8449 35768 8483
rect 35716 8440 35768 8449
rect 35900 8440 35952 8492
rect 36084 8483 36136 8492
rect 36084 8449 36093 8483
rect 36093 8449 36127 8483
rect 36127 8449 36136 8483
rect 36084 8440 36136 8449
rect 36452 8483 36504 8492
rect 36452 8449 36461 8483
rect 36461 8449 36495 8483
rect 36495 8449 36504 8483
rect 36452 8440 36504 8449
rect 36820 8483 36872 8492
rect 36820 8449 36829 8483
rect 36829 8449 36863 8483
rect 36863 8449 36872 8483
rect 36820 8440 36872 8449
rect 37096 8440 37148 8492
rect 37556 8483 37608 8492
rect 37556 8449 37565 8483
rect 37565 8449 37599 8483
rect 37599 8449 37608 8483
rect 37556 8440 37608 8449
rect 37924 8483 37976 8492
rect 37924 8449 37933 8483
rect 37933 8449 37967 8483
rect 37967 8449 37976 8483
rect 37924 8440 37976 8449
rect 38292 8483 38344 8492
rect 38292 8449 38301 8483
rect 38301 8449 38335 8483
rect 38335 8449 38344 8483
rect 38292 8440 38344 8449
rect 38568 8440 38620 8492
rect 35808 8236 35860 8288
rect 36636 8347 36688 8356
rect 36636 8313 36645 8347
rect 36645 8313 36679 8347
rect 36679 8313 36688 8347
rect 36636 8304 36688 8313
rect 38108 8347 38160 8356
rect 38108 8313 38117 8347
rect 38117 8313 38151 8347
rect 38151 8313 38160 8347
rect 38108 8304 38160 8313
rect 38384 8372 38436 8424
rect 39396 8483 39448 8492
rect 39396 8449 39405 8483
rect 39405 8449 39439 8483
rect 39439 8449 39448 8483
rect 39396 8440 39448 8449
rect 39948 8483 40000 8492
rect 39948 8449 39957 8483
rect 39957 8449 39991 8483
rect 39991 8449 40000 8483
rect 39948 8440 40000 8449
rect 40960 8483 41012 8492
rect 40960 8449 40969 8483
rect 40969 8449 41003 8483
rect 41003 8449 41012 8483
rect 40960 8440 41012 8449
rect 41880 8483 41932 8492
rect 41880 8449 41889 8483
rect 41889 8449 41923 8483
rect 41923 8449 41932 8483
rect 41880 8440 41932 8449
rect 42432 8483 42484 8492
rect 42432 8449 42441 8483
rect 42441 8449 42475 8483
rect 42475 8449 42484 8483
rect 42432 8440 42484 8449
rect 42984 8440 43036 8492
rect 43444 8483 43496 8492
rect 43444 8449 43453 8483
rect 43453 8449 43487 8483
rect 43487 8449 43496 8483
rect 43444 8440 43496 8449
rect 38476 8347 38528 8356
rect 38476 8313 38485 8347
rect 38485 8313 38519 8347
rect 38519 8313 38528 8347
rect 38476 8304 38528 8313
rect 43076 8372 43128 8424
rect 40408 8304 40460 8356
rect 41512 8304 41564 8356
rect 42616 8304 42668 8356
rect 44364 8483 44416 8492
rect 44364 8449 44373 8483
rect 44373 8449 44407 8483
rect 44407 8449 44416 8483
rect 44364 8440 44416 8449
rect 45100 8483 45152 8492
rect 45100 8449 45109 8483
rect 45109 8449 45143 8483
rect 45143 8449 45152 8483
rect 45100 8440 45152 8449
rect 6539 8134 6591 8186
rect 6603 8134 6655 8186
rect 6667 8134 6719 8186
rect 6731 8134 6783 8186
rect 6795 8134 6847 8186
rect 17717 8134 17769 8186
rect 17781 8134 17833 8186
rect 17845 8134 17897 8186
rect 17909 8134 17961 8186
rect 17973 8134 18025 8186
rect 28895 8134 28947 8186
rect 28959 8134 29011 8186
rect 29023 8134 29075 8186
rect 29087 8134 29139 8186
rect 29151 8134 29203 8186
rect 40073 8134 40125 8186
rect 40137 8134 40189 8186
rect 40201 8134 40253 8186
rect 40265 8134 40317 8186
rect 40329 8134 40381 8186
rect 664 8032 716 8084
rect 2136 8032 2188 8084
rect 4712 8032 4764 8084
rect 5816 8032 5868 8084
rect 6644 8075 6696 8084
rect 6644 8041 6653 8075
rect 6653 8041 6687 8075
rect 6687 8041 6696 8075
rect 6644 8032 6696 8041
rect 7288 8032 7340 8084
rect 9220 8075 9272 8084
rect 9220 8041 9229 8075
rect 9229 8041 9263 8075
rect 9263 8041 9272 8075
rect 9220 8032 9272 8041
rect 10232 8032 10284 8084
rect 11796 8075 11848 8084
rect 11796 8041 11805 8075
rect 11805 8041 11839 8075
rect 11839 8041 11848 8075
rect 11796 8032 11848 8041
rect 1400 7964 1452 8016
rect 4160 8007 4212 8016
rect 4160 7973 4169 8007
rect 4169 7973 4203 8007
rect 4203 7973 4212 8007
rect 4160 7964 4212 7973
rect 12624 8032 12676 8084
rect 12808 8032 12860 8084
rect 14372 8075 14424 8084
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 15752 8032 15804 8084
rect 17592 8032 17644 8084
rect 4344 7828 4396 7880
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 2320 7803 2372 7812
rect 2320 7769 2329 7803
rect 2329 7769 2363 7803
rect 2363 7769 2372 7803
rect 2320 7760 2372 7769
rect 3976 7803 4028 7812
rect 3976 7769 3985 7803
rect 3985 7769 4019 7803
rect 4019 7769 4028 7803
rect 3976 7760 4028 7769
rect 18328 8032 18380 8084
rect 18696 8032 18748 8084
rect 19432 8032 19484 8084
rect 19708 8032 19760 8084
rect 21088 8032 21140 8084
rect 21364 8032 21416 8084
rect 22560 8075 22612 8084
rect 22560 8041 22569 8075
rect 22569 8041 22603 8075
rect 22603 8041 22612 8075
rect 22560 8032 22612 8041
rect 22836 8075 22888 8084
rect 22836 8041 22845 8075
rect 22845 8041 22879 8075
rect 22879 8041 22888 8075
rect 22836 8032 22888 8041
rect 22928 8032 22980 8084
rect 23664 8032 23716 8084
rect 24216 8075 24268 8084
rect 24216 8041 24225 8075
rect 24225 8041 24259 8075
rect 24259 8041 24268 8075
rect 24216 8032 24268 8041
rect 24584 8032 24636 8084
rect 25136 8032 25188 8084
rect 25412 8032 25464 8084
rect 25688 8032 25740 8084
rect 26148 8075 26200 8084
rect 26148 8041 26157 8075
rect 26157 8041 26191 8075
rect 26191 8041 26200 8075
rect 26148 8032 26200 8041
rect 26700 8075 26752 8084
rect 26700 8041 26709 8075
rect 26709 8041 26743 8075
rect 26743 8041 26752 8075
rect 26700 8032 26752 8041
rect 27068 8075 27120 8084
rect 27068 8041 27077 8075
rect 27077 8041 27111 8075
rect 27111 8041 27120 8075
rect 27068 8032 27120 8041
rect 27804 8075 27856 8084
rect 27804 8041 27813 8075
rect 27813 8041 27847 8075
rect 27847 8041 27856 8075
rect 27804 8032 27856 8041
rect 18420 7964 18472 8016
rect 18512 7964 18564 8016
rect 9680 7828 9732 7880
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 17500 7828 17552 7880
rect 17960 7828 18012 7880
rect 18052 7871 18104 7880
rect 18052 7837 18061 7871
rect 18061 7837 18095 7871
rect 18095 7837 18104 7871
rect 18052 7828 18104 7837
rect 18236 7828 18288 7880
rect 19708 7896 19760 7948
rect 19248 7828 19300 7880
rect 19340 7871 19392 7880
rect 19340 7837 19349 7871
rect 19349 7837 19383 7871
rect 19383 7837 19392 7871
rect 19340 7828 19392 7837
rect 19892 7871 19944 7880
rect 19892 7837 19901 7871
rect 19901 7837 19935 7871
rect 19935 7837 19944 7871
rect 19892 7828 19944 7837
rect 20168 7871 20220 7880
rect 20168 7837 20177 7871
rect 20177 7837 20211 7871
rect 20211 7837 20220 7871
rect 20168 7828 20220 7837
rect 20628 7828 20680 7880
rect 20904 7828 20956 7880
rect 8944 7692 8996 7744
rect 9128 7803 9180 7812
rect 9128 7769 9137 7803
rect 9137 7769 9171 7803
rect 9171 7769 9180 7803
rect 9128 7760 9180 7769
rect 11704 7803 11756 7812
rect 11704 7769 11713 7803
rect 11713 7769 11747 7803
rect 11747 7769 11756 7803
rect 11704 7760 11756 7769
rect 14280 7803 14332 7812
rect 14280 7769 14289 7803
rect 14289 7769 14323 7803
rect 14323 7769 14332 7803
rect 14280 7760 14332 7769
rect 11796 7692 11848 7744
rect 17868 7760 17920 7812
rect 21364 7828 21416 7880
rect 21732 7896 21784 7948
rect 21824 7828 21876 7880
rect 22008 7871 22060 7880
rect 22008 7837 22017 7871
rect 22017 7837 22051 7871
rect 22051 7837 22060 7871
rect 22008 7828 22060 7837
rect 23572 7964 23624 8016
rect 23020 7896 23072 7948
rect 22652 7871 22704 7880
rect 22652 7837 22661 7871
rect 22661 7837 22695 7871
rect 22695 7837 22704 7871
rect 22652 7828 22704 7837
rect 23112 7828 23164 7880
rect 23204 7871 23256 7880
rect 23204 7837 23213 7871
rect 23213 7837 23247 7871
rect 23247 7837 23256 7871
rect 23204 7828 23256 7837
rect 25504 7964 25556 8016
rect 17684 7692 17736 7744
rect 19524 7735 19576 7744
rect 19524 7701 19533 7735
rect 19533 7701 19567 7735
rect 19567 7701 19576 7735
rect 19524 7692 19576 7701
rect 20076 7735 20128 7744
rect 20076 7701 20085 7735
rect 20085 7701 20119 7735
rect 20119 7701 20128 7735
rect 20076 7692 20128 7701
rect 20352 7735 20404 7744
rect 20352 7701 20361 7735
rect 20361 7701 20395 7735
rect 20395 7701 20404 7735
rect 20352 7692 20404 7701
rect 20444 7692 20496 7744
rect 21916 7760 21968 7812
rect 24492 7828 24544 7880
rect 24676 7828 24728 7880
rect 26792 7896 26844 7948
rect 27344 7896 27396 7948
rect 29276 8032 29328 8084
rect 40776 8032 40828 8084
rect 44456 8032 44508 8084
rect 25044 7828 25096 7880
rect 25596 7828 25648 7880
rect 25872 7828 25924 7880
rect 26056 7828 26108 7880
rect 26424 7828 26476 7880
rect 27160 7828 27212 7880
rect 27436 7828 27488 7880
rect 27896 7828 27948 7880
rect 28724 7964 28776 8016
rect 45928 7964 45980 8016
rect 29552 7828 29604 7880
rect 29828 7828 29880 7880
rect 40960 7871 41012 7880
rect 40960 7837 40969 7871
rect 40969 7837 41003 7871
rect 41003 7837 41012 7871
rect 40960 7828 41012 7837
rect 46296 7828 46348 7880
rect 21732 7735 21784 7744
rect 21732 7701 21741 7735
rect 21741 7701 21775 7735
rect 21775 7701 21784 7735
rect 21732 7692 21784 7701
rect 22008 7692 22060 7744
rect 44180 7760 44232 7812
rect 45008 7760 45060 7812
rect 24124 7692 24176 7744
rect 25044 7735 25096 7744
rect 25044 7701 25053 7735
rect 25053 7701 25087 7735
rect 25087 7701 25096 7735
rect 25044 7692 25096 7701
rect 25320 7735 25372 7744
rect 25320 7701 25329 7735
rect 25329 7701 25363 7735
rect 25363 7701 25372 7735
rect 25320 7692 25372 7701
rect 25596 7735 25648 7744
rect 25596 7701 25605 7735
rect 25605 7701 25639 7735
rect 25639 7701 25648 7735
rect 25596 7692 25648 7701
rect 26424 7735 26476 7744
rect 26424 7701 26433 7735
rect 26433 7701 26467 7735
rect 26467 7701 26476 7735
rect 26424 7692 26476 7701
rect 28172 7735 28224 7744
rect 28172 7701 28181 7735
rect 28181 7701 28215 7735
rect 28215 7701 28224 7735
rect 28172 7692 28224 7701
rect 28540 7735 28592 7744
rect 28540 7701 28549 7735
rect 28549 7701 28583 7735
rect 28583 7701 28592 7735
rect 28540 7692 28592 7701
rect 43904 7692 43956 7744
rect 12128 7590 12180 7642
rect 12192 7590 12244 7642
rect 12256 7590 12308 7642
rect 12320 7590 12372 7642
rect 12384 7590 12436 7642
rect 23306 7590 23358 7642
rect 23370 7590 23422 7642
rect 23434 7590 23486 7642
rect 23498 7590 23550 7642
rect 23562 7590 23614 7642
rect 34484 7590 34536 7642
rect 34548 7590 34600 7642
rect 34612 7590 34664 7642
rect 34676 7590 34728 7642
rect 34740 7590 34792 7642
rect 45662 7590 45714 7642
rect 45726 7590 45778 7642
rect 45790 7590 45842 7642
rect 45854 7590 45906 7642
rect 45918 7590 45970 7642
rect 1032 7488 1084 7540
rect 1768 7488 1820 7540
rect 17684 7488 17736 7540
rect 17868 7488 17920 7540
rect 19340 7488 19392 7540
rect 19984 7488 20036 7540
rect 20168 7488 20220 7540
rect 4344 7420 4396 7472
rect 8300 7420 8352 7472
rect 9128 7420 9180 7472
rect 9680 7420 9732 7472
rect 15108 7284 15160 7336
rect 15476 7352 15528 7404
rect 19064 7395 19116 7404
rect 19064 7361 19073 7395
rect 19073 7361 19107 7395
rect 19107 7361 19116 7395
rect 19064 7352 19116 7361
rect 19340 7395 19392 7404
rect 19340 7361 19349 7395
rect 19349 7361 19383 7395
rect 19383 7361 19392 7395
rect 19340 7352 19392 7361
rect 19708 7395 19760 7404
rect 19708 7361 19717 7395
rect 19717 7361 19751 7395
rect 19751 7361 19760 7395
rect 19708 7352 19760 7361
rect 19800 7352 19852 7404
rect 17224 7284 17276 7336
rect 18788 7284 18840 7336
rect 19892 7284 19944 7336
rect 20628 7488 20680 7540
rect 21180 7488 21232 7540
rect 21456 7488 21508 7540
rect 21548 7531 21600 7540
rect 21548 7497 21557 7531
rect 21557 7497 21591 7531
rect 21591 7497 21600 7531
rect 21548 7488 21600 7497
rect 21640 7488 21692 7540
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 22284 7352 22336 7404
rect 22744 7352 22796 7404
rect 23388 7488 23440 7540
rect 31852 7488 31904 7540
rect 43352 7488 43404 7540
rect 45560 7488 45612 7540
rect 33784 7420 33836 7472
rect 23204 7352 23256 7404
rect 23296 7352 23348 7404
rect 23572 7352 23624 7404
rect 23848 7352 23900 7404
rect 27528 7352 27580 7404
rect 41420 7352 41472 7404
rect 44364 7395 44416 7404
rect 44364 7361 44373 7395
rect 44373 7361 44407 7395
rect 44407 7361 44416 7395
rect 44364 7352 44416 7361
rect 44916 7395 44968 7404
rect 44916 7361 44925 7395
rect 44925 7361 44959 7395
rect 44959 7361 44968 7395
rect 44916 7352 44968 7361
rect 45192 7352 45244 7404
rect 30656 7284 30708 7336
rect 2320 7216 2372 7268
rect 9680 7216 9732 7268
rect 16672 7216 16724 7268
rect 18512 7216 18564 7268
rect 19248 7216 19300 7268
rect 14464 7148 14516 7200
rect 19064 7148 19116 7200
rect 21640 7216 21692 7268
rect 20720 7148 20772 7200
rect 21088 7148 21140 7200
rect 22284 7191 22336 7200
rect 22284 7157 22293 7191
rect 22293 7157 22327 7191
rect 22327 7157 22336 7191
rect 22284 7148 22336 7157
rect 22376 7148 22428 7200
rect 23480 7216 23532 7268
rect 33324 7216 33376 7268
rect 23204 7191 23256 7200
rect 23204 7157 23213 7191
rect 23213 7157 23247 7191
rect 23247 7157 23256 7191
rect 23204 7148 23256 7157
rect 23848 7191 23900 7200
rect 23848 7157 23857 7191
rect 23857 7157 23891 7191
rect 23891 7157 23900 7191
rect 23848 7148 23900 7157
rect 24400 7148 24452 7200
rect 6539 7046 6591 7098
rect 6603 7046 6655 7098
rect 6667 7046 6719 7098
rect 6731 7046 6783 7098
rect 6795 7046 6847 7098
rect 17717 7046 17769 7098
rect 17781 7046 17833 7098
rect 17845 7046 17897 7098
rect 17909 7046 17961 7098
rect 17973 7046 18025 7098
rect 28895 7046 28947 7098
rect 28959 7046 29011 7098
rect 29023 7046 29075 7098
rect 29087 7046 29139 7098
rect 29151 7046 29203 7098
rect 40073 7046 40125 7098
rect 40137 7046 40189 7098
rect 40201 7046 40253 7098
rect 40265 7046 40317 7098
rect 40329 7046 40381 7098
rect 12624 6944 12676 6996
rect 15200 6944 15252 6996
rect 21088 6944 21140 6996
rect 21364 6944 21416 6996
rect 34152 6944 34204 6996
rect 19708 6876 19760 6928
rect 33692 6876 33744 6928
rect 20720 6808 20772 6860
rect 44088 6808 44140 6860
rect 36636 6740 36688 6792
rect 3976 6672 4028 6724
rect 25320 6672 25372 6724
rect 42800 6672 42852 6724
rect 16580 6604 16632 6656
rect 12128 6502 12180 6554
rect 12192 6502 12244 6554
rect 12256 6502 12308 6554
rect 12320 6502 12372 6554
rect 12384 6502 12436 6554
rect 23306 6502 23358 6554
rect 23370 6502 23422 6554
rect 23434 6502 23486 6554
rect 23498 6502 23550 6554
rect 23562 6502 23614 6554
rect 34484 6502 34536 6554
rect 34548 6502 34600 6554
rect 34612 6502 34664 6554
rect 34676 6502 34728 6554
rect 34740 6502 34792 6554
rect 45662 6502 45714 6554
rect 45726 6502 45778 6554
rect 45790 6502 45842 6554
rect 45854 6502 45906 6554
rect 45918 6502 45970 6554
rect 24952 6196 25004 6248
rect 39396 6196 39448 6248
rect 27252 6128 27304 6180
rect 43076 6128 43128 6180
rect 6539 5958 6591 6010
rect 6603 5958 6655 6010
rect 6667 5958 6719 6010
rect 6731 5958 6783 6010
rect 6795 5958 6847 6010
rect 17717 5958 17769 6010
rect 17781 5958 17833 6010
rect 17845 5958 17897 6010
rect 17909 5958 17961 6010
rect 17973 5958 18025 6010
rect 28895 5958 28947 6010
rect 28959 5958 29011 6010
rect 29023 5958 29075 6010
rect 29087 5958 29139 6010
rect 29151 5958 29203 6010
rect 40073 5958 40125 6010
rect 40137 5958 40189 6010
rect 40201 5958 40253 6010
rect 40265 5958 40317 6010
rect 40329 5958 40381 6010
rect 12128 5414 12180 5466
rect 12192 5414 12244 5466
rect 12256 5414 12308 5466
rect 12320 5414 12372 5466
rect 12384 5414 12436 5466
rect 23306 5414 23358 5466
rect 23370 5414 23422 5466
rect 23434 5414 23486 5466
rect 23498 5414 23550 5466
rect 23562 5414 23614 5466
rect 34484 5414 34536 5466
rect 34548 5414 34600 5466
rect 34612 5414 34664 5466
rect 34676 5414 34728 5466
rect 34740 5414 34792 5466
rect 45662 5414 45714 5466
rect 45726 5414 45778 5466
rect 45790 5414 45842 5466
rect 45854 5414 45906 5466
rect 45918 5414 45970 5466
rect 6539 4870 6591 4922
rect 6603 4870 6655 4922
rect 6667 4870 6719 4922
rect 6731 4870 6783 4922
rect 6795 4870 6847 4922
rect 17717 4870 17769 4922
rect 17781 4870 17833 4922
rect 17845 4870 17897 4922
rect 17909 4870 17961 4922
rect 17973 4870 18025 4922
rect 28895 4870 28947 4922
rect 28959 4870 29011 4922
rect 29023 4870 29075 4922
rect 29087 4870 29139 4922
rect 29151 4870 29203 4922
rect 40073 4870 40125 4922
rect 40137 4870 40189 4922
rect 40201 4870 40253 4922
rect 40265 4870 40317 4922
rect 40329 4870 40381 4922
rect 23112 4768 23164 4820
rect 38384 4768 38436 4820
rect 43904 4768 43956 4820
rect 23664 4564 23716 4616
rect 35900 4607 35952 4616
rect 35900 4573 35909 4607
rect 35909 4573 35943 4607
rect 35943 4573 35952 4607
rect 35900 4564 35952 4573
rect 39948 4496 40000 4548
rect 12128 4326 12180 4378
rect 12192 4326 12244 4378
rect 12256 4326 12308 4378
rect 12320 4326 12372 4378
rect 12384 4326 12436 4378
rect 23306 4326 23358 4378
rect 23370 4326 23422 4378
rect 23434 4326 23486 4378
rect 23498 4326 23550 4378
rect 23562 4326 23614 4378
rect 34484 4326 34536 4378
rect 34548 4326 34600 4378
rect 34612 4326 34664 4378
rect 34676 4326 34728 4378
rect 34740 4326 34792 4378
rect 45662 4326 45714 4378
rect 45726 4326 45778 4378
rect 45790 4326 45842 4378
rect 45854 4326 45906 4378
rect 45918 4326 45970 4378
rect 22652 4131 22704 4140
rect 22652 4097 22661 4131
rect 22661 4097 22695 4131
rect 22695 4097 22704 4131
rect 22652 4088 22704 4097
rect 20812 4020 20864 4072
rect 23204 4088 23256 4140
rect 27068 4131 27120 4140
rect 27068 4097 27077 4131
rect 27077 4097 27111 4131
rect 27111 4097 27120 4131
rect 27068 4088 27120 4097
rect 33692 4131 33744 4140
rect 33692 4097 33701 4131
rect 33701 4097 33735 4131
rect 33735 4097 33744 4131
rect 33692 4088 33744 4097
rect 35440 4131 35492 4140
rect 35440 4097 35449 4131
rect 35449 4097 35483 4131
rect 35483 4097 35492 4131
rect 35440 4088 35492 4097
rect 44548 4131 44600 4140
rect 44548 4097 44557 4131
rect 44557 4097 44591 4131
rect 44591 4097 44600 4131
rect 44548 4088 44600 4097
rect 23664 3952 23716 4004
rect 35808 4020 35860 4072
rect 27252 3927 27304 3936
rect 27252 3893 27261 3927
rect 27261 3893 27295 3927
rect 27295 3893 27304 3927
rect 27252 3884 27304 3893
rect 33600 3952 33652 4004
rect 35900 3952 35952 4004
rect 33876 3927 33928 3936
rect 33876 3893 33885 3927
rect 33885 3893 33919 3927
rect 33919 3893 33928 3927
rect 33876 3884 33928 3893
rect 44364 3927 44416 3936
rect 44364 3893 44373 3927
rect 44373 3893 44407 3927
rect 44407 3893 44416 3927
rect 44364 3884 44416 3893
rect 6539 3782 6591 3834
rect 6603 3782 6655 3834
rect 6667 3782 6719 3834
rect 6731 3782 6783 3834
rect 6795 3782 6847 3834
rect 17717 3782 17769 3834
rect 17781 3782 17833 3834
rect 17845 3782 17897 3834
rect 17909 3782 17961 3834
rect 17973 3782 18025 3834
rect 28895 3782 28947 3834
rect 28959 3782 29011 3834
rect 29023 3782 29075 3834
rect 29087 3782 29139 3834
rect 29151 3782 29203 3834
rect 40073 3782 40125 3834
rect 40137 3782 40189 3834
rect 40201 3782 40253 3834
rect 40265 3782 40317 3834
rect 40329 3782 40381 3834
rect 22652 3680 22704 3732
rect 33692 3680 33744 3732
rect 33876 3680 33928 3732
rect 42800 3680 42852 3732
rect 32220 3612 32272 3664
rect 21364 3476 21416 3528
rect 23020 3476 23072 3528
rect 32404 3476 32456 3528
rect 23940 3408 23992 3460
rect 33968 3408 34020 3460
rect 12128 3238 12180 3290
rect 12192 3238 12244 3290
rect 12256 3238 12308 3290
rect 12320 3238 12372 3290
rect 12384 3238 12436 3290
rect 23306 3238 23358 3290
rect 23370 3238 23422 3290
rect 23434 3238 23486 3290
rect 23498 3238 23550 3290
rect 23562 3238 23614 3290
rect 34484 3238 34536 3290
rect 34548 3238 34600 3290
rect 34612 3238 34664 3290
rect 34676 3238 34728 3290
rect 34740 3238 34792 3290
rect 45662 3238 45714 3290
rect 45726 3238 45778 3290
rect 45790 3238 45842 3290
rect 45854 3238 45906 3290
rect 45918 3238 45970 3290
rect 23020 3179 23072 3188
rect 23020 3145 23029 3179
rect 23029 3145 23063 3179
rect 23063 3145 23072 3179
rect 23020 3136 23072 3145
rect 23204 3136 23256 3188
rect 27068 3136 27120 3188
rect 44548 3136 44600 3188
rect 19248 3000 19300 3052
rect 23572 3043 23624 3052
rect 23572 3009 23581 3043
rect 23581 3009 23615 3043
rect 23615 3009 23624 3043
rect 23572 3000 23624 3009
rect 25780 3000 25832 3052
rect 29276 3043 29328 3052
rect 29276 3009 29285 3043
rect 29285 3009 29319 3043
rect 29319 3009 29328 3043
rect 29276 3000 29328 3009
rect 39028 3000 39080 3052
rect 23664 2932 23716 2984
rect 40960 2932 41012 2984
rect 41420 2864 41472 2916
rect 6539 2694 6591 2746
rect 6603 2694 6655 2746
rect 6667 2694 6719 2746
rect 6731 2694 6783 2746
rect 6795 2694 6847 2746
rect 17717 2694 17769 2746
rect 17781 2694 17833 2746
rect 17845 2694 17897 2746
rect 17909 2694 17961 2746
rect 17973 2694 18025 2746
rect 28895 2694 28947 2746
rect 28959 2694 29011 2746
rect 29023 2694 29075 2746
rect 29087 2694 29139 2746
rect 29151 2694 29203 2746
rect 40073 2694 40125 2746
rect 40137 2694 40189 2746
rect 40201 2694 40253 2746
rect 40265 2694 40317 2746
rect 40329 2694 40381 2746
rect 23572 2524 23624 2576
rect 24952 2524 25004 2576
rect 29276 2592 29328 2644
rect 44180 2592 44232 2644
rect 44916 2592 44968 2644
rect 45008 2635 45060 2644
rect 45008 2601 45017 2635
rect 45017 2601 45051 2635
rect 45051 2601 45060 2635
rect 45008 2592 45060 2601
rect 41880 2524 41932 2576
rect 37372 2456 37424 2508
rect 20720 2388 20772 2440
rect 23020 2431 23072 2440
rect 23020 2397 23029 2431
rect 23029 2397 23063 2431
rect 23063 2397 23072 2431
rect 23020 2388 23072 2397
rect 23204 2388 23256 2440
rect 23848 2431 23900 2440
rect 23848 2397 23857 2431
rect 23857 2397 23891 2431
rect 23891 2397 23900 2431
rect 23848 2388 23900 2397
rect 24860 2431 24912 2440
rect 24860 2397 24869 2431
rect 24869 2397 24903 2431
rect 24903 2397 24912 2431
rect 24860 2388 24912 2397
rect 28816 2431 28868 2440
rect 28816 2397 28825 2431
rect 28825 2397 28859 2431
rect 28859 2397 28868 2431
rect 28816 2388 28868 2397
rect 31484 2431 31536 2440
rect 31484 2397 31493 2431
rect 31493 2397 31527 2431
rect 31527 2397 31536 2431
rect 31484 2388 31536 2397
rect 38200 2431 38252 2440
rect 38200 2397 38209 2431
rect 38209 2397 38243 2431
rect 38243 2397 38252 2431
rect 38200 2388 38252 2397
rect 20628 2363 20680 2372
rect 20628 2329 20637 2363
rect 20637 2329 20671 2363
rect 20671 2329 20680 2363
rect 20628 2320 20680 2329
rect 35532 2320 35584 2372
rect 44272 2456 44324 2508
rect 41788 2388 41840 2440
rect 23940 2252 23992 2304
rect 43904 2320 43956 2372
rect 45468 2431 45520 2440
rect 45468 2397 45477 2431
rect 45477 2397 45511 2431
rect 45511 2397 45520 2431
rect 45468 2388 45520 2397
rect 45100 2252 45152 2304
rect 12128 2150 12180 2202
rect 12192 2150 12244 2202
rect 12256 2150 12308 2202
rect 12320 2150 12372 2202
rect 12384 2150 12436 2202
rect 23306 2150 23358 2202
rect 23370 2150 23422 2202
rect 23434 2150 23486 2202
rect 23498 2150 23550 2202
rect 23562 2150 23614 2202
rect 34484 2150 34536 2202
rect 34548 2150 34600 2202
rect 34612 2150 34664 2202
rect 34676 2150 34728 2202
rect 34740 2150 34792 2202
rect 45662 2150 45714 2202
rect 45726 2150 45778 2202
rect 45790 2150 45842 2202
rect 45854 2150 45906 2202
rect 45918 2150 45970 2202
rect 20628 2048 20680 2100
rect 23020 2048 23072 2100
rect 23112 2048 23164 2100
rect 23204 2048 23256 2100
rect 23848 2048 23900 2100
rect 24860 2048 24912 2100
rect 31484 2048 31536 2100
rect 38200 2048 38252 2100
rect 41788 2091 41840 2100
rect 41788 2057 41797 2091
rect 41797 2057 41831 2091
rect 41831 2057 41840 2091
rect 41788 2048 41840 2057
rect 43904 2091 43956 2100
rect 43904 2057 43913 2091
rect 43913 2057 43947 2091
rect 43947 2057 43956 2091
rect 43904 2048 43956 2057
rect 45468 2048 45520 2100
rect 19800 1955 19852 1964
rect 19800 1921 19809 1955
rect 19809 1921 19843 1955
rect 19843 1921 19852 1955
rect 19800 1912 19852 1921
rect 20904 1912 20956 1964
rect 1676 1844 1728 1896
rect 23204 1955 23256 1964
rect 23204 1921 23213 1955
rect 23213 1921 23247 1955
rect 23247 1921 23256 1955
rect 23204 1912 23256 1921
rect 22652 1844 22704 1896
rect 24400 1955 24452 1964
rect 24400 1921 24409 1955
rect 24409 1921 24443 1955
rect 24443 1921 24452 1955
rect 24400 1912 24452 1921
rect 31024 1955 31076 1964
rect 31024 1921 31033 1955
rect 31033 1921 31067 1955
rect 31067 1921 31076 1955
rect 31024 1912 31076 1921
rect 37464 1955 37516 1964
rect 37464 1921 37473 1955
rect 37473 1921 37507 1955
rect 37507 1921 37516 1955
rect 37464 1912 37516 1921
rect 41972 1955 42024 1964
rect 41972 1921 41981 1955
rect 41981 1921 42015 1955
rect 42015 1921 42024 1955
rect 41972 1912 42024 1921
rect 44088 1955 44140 1964
rect 44088 1921 44097 1955
rect 44097 1921 44131 1955
rect 44131 1921 44140 1955
rect 44088 1912 44140 1921
rect 44824 1955 44876 1964
rect 44824 1921 44833 1955
rect 44833 1921 44867 1955
rect 44867 1921 44876 1955
rect 44824 1912 44876 1921
rect 6539 1606 6591 1658
rect 6603 1606 6655 1658
rect 6667 1606 6719 1658
rect 6731 1606 6783 1658
rect 6795 1606 6847 1658
rect 17717 1606 17769 1658
rect 17781 1606 17833 1658
rect 17845 1606 17897 1658
rect 17909 1606 17961 1658
rect 17973 1606 18025 1658
rect 28895 1606 28947 1658
rect 28959 1606 29011 1658
rect 29023 1606 29075 1658
rect 29087 1606 29139 1658
rect 29151 1606 29203 1658
rect 40073 1606 40125 1658
rect 40137 1606 40189 1658
rect 40201 1606 40253 1658
rect 40265 1606 40317 1658
rect 40329 1606 40381 1658
rect 1676 1547 1728 1556
rect 1676 1513 1685 1547
rect 1685 1513 1719 1547
rect 1719 1513 1728 1547
rect 1676 1504 1728 1513
rect 19800 1504 19852 1556
rect 24400 1504 24452 1556
rect 28816 1504 28868 1556
rect 31024 1504 31076 1556
rect 41972 1504 42024 1556
rect 44088 1504 44140 1556
rect 44824 1504 44876 1556
rect 1492 1343 1544 1352
rect 1492 1309 1501 1343
rect 1501 1309 1535 1343
rect 1535 1309 1544 1343
rect 1492 1300 1544 1309
rect 3792 1343 3844 1352
rect 3792 1309 3801 1343
rect 3801 1309 3835 1343
rect 3835 1309 3844 1343
rect 3792 1300 3844 1309
rect 5908 1343 5960 1352
rect 5908 1309 5917 1343
rect 5917 1309 5951 1343
rect 5951 1309 5960 1343
rect 5908 1300 5960 1309
rect 8116 1343 8168 1352
rect 8116 1309 8125 1343
rect 8125 1309 8159 1343
rect 8159 1309 8168 1343
rect 8116 1300 8168 1309
rect 10324 1343 10376 1352
rect 10324 1309 10333 1343
rect 10333 1309 10367 1343
rect 10367 1309 10376 1343
rect 10324 1300 10376 1309
rect 12532 1343 12584 1352
rect 12532 1309 12541 1343
rect 12541 1309 12575 1343
rect 12575 1309 12584 1343
rect 12532 1300 12584 1309
rect 14740 1343 14792 1352
rect 14740 1309 14749 1343
rect 14749 1309 14783 1343
rect 14783 1309 14792 1343
rect 14740 1300 14792 1309
rect 17132 1343 17184 1352
rect 17132 1309 17141 1343
rect 17141 1309 17175 1343
rect 17175 1309 17184 1343
rect 17132 1300 17184 1309
rect 19432 1343 19484 1352
rect 19432 1309 19441 1343
rect 19441 1309 19475 1343
rect 19475 1309 19484 1343
rect 19432 1300 19484 1309
rect 20720 1300 20772 1352
rect 21548 1343 21600 1352
rect 21548 1309 21557 1343
rect 21557 1309 21591 1343
rect 21591 1309 21600 1343
rect 21548 1300 21600 1309
rect 23756 1343 23808 1352
rect 23756 1309 23765 1343
rect 23765 1309 23799 1343
rect 23799 1309 23808 1343
rect 23756 1300 23808 1309
rect 25964 1343 26016 1352
rect 25964 1309 25973 1343
rect 25973 1309 26007 1343
rect 26007 1309 26016 1343
rect 25964 1300 26016 1309
rect 28172 1343 28224 1352
rect 28172 1309 28181 1343
rect 28181 1309 28215 1343
rect 28215 1309 28224 1343
rect 28172 1300 28224 1309
rect 30380 1343 30432 1352
rect 30380 1309 30389 1343
rect 30389 1309 30423 1343
rect 30423 1309 30432 1343
rect 30380 1300 30432 1309
rect 32588 1343 32640 1352
rect 32588 1309 32597 1343
rect 32597 1309 32631 1343
rect 32631 1309 32640 1343
rect 32588 1300 32640 1309
rect 34888 1343 34940 1352
rect 34888 1309 34897 1343
rect 34897 1309 34931 1343
rect 34931 1309 34940 1343
rect 34888 1300 34940 1309
rect 35440 1300 35492 1352
rect 37004 1343 37056 1352
rect 37004 1309 37013 1343
rect 37013 1309 37047 1343
rect 37047 1309 37056 1343
rect 37004 1300 37056 1309
rect 37464 1300 37516 1352
rect 39212 1343 39264 1352
rect 39212 1309 39221 1343
rect 39221 1309 39255 1343
rect 39255 1309 39264 1343
rect 39212 1300 39264 1309
rect 41420 1343 41472 1352
rect 41420 1309 41429 1343
rect 41429 1309 41463 1343
rect 41463 1309 41472 1343
rect 41420 1300 41472 1309
rect 43628 1343 43680 1352
rect 43628 1309 43637 1343
rect 43637 1309 43671 1343
rect 43671 1309 43680 1343
rect 43628 1300 43680 1309
rect 45560 1300 45612 1352
rect 6092 1207 6144 1216
rect 6092 1173 6101 1207
rect 6101 1173 6135 1207
rect 6135 1173 6144 1207
rect 6092 1164 6144 1173
rect 8300 1207 8352 1216
rect 8300 1173 8309 1207
rect 8309 1173 8343 1207
rect 8343 1173 8352 1207
rect 8300 1164 8352 1173
rect 10508 1207 10560 1216
rect 10508 1173 10517 1207
rect 10517 1173 10551 1207
rect 10551 1173 10560 1207
rect 10508 1164 10560 1173
rect 11704 1164 11756 1216
rect 20904 1232 20956 1284
rect 16856 1164 16908 1216
rect 21364 1207 21416 1216
rect 21364 1173 21373 1207
rect 21373 1173 21407 1207
rect 21407 1173 21416 1207
rect 21364 1164 21416 1173
rect 25780 1207 25832 1216
rect 25780 1173 25789 1207
rect 25789 1173 25823 1207
rect 25823 1173 25832 1207
rect 25780 1164 25832 1173
rect 32404 1207 32456 1216
rect 32404 1173 32413 1207
rect 32413 1173 32447 1207
rect 32447 1173 32456 1207
rect 32404 1164 32456 1173
rect 39028 1207 39080 1216
rect 39028 1173 39037 1207
rect 39037 1173 39071 1207
rect 39071 1173 39080 1207
rect 39028 1164 39080 1173
rect 12128 1062 12180 1114
rect 12192 1062 12244 1114
rect 12256 1062 12308 1114
rect 12320 1062 12372 1114
rect 12384 1062 12436 1114
rect 23306 1062 23358 1114
rect 23370 1062 23422 1114
rect 23434 1062 23486 1114
rect 23498 1062 23550 1114
rect 23562 1062 23614 1114
rect 34484 1062 34536 1114
rect 34548 1062 34600 1114
rect 34612 1062 34664 1114
rect 34676 1062 34728 1114
rect 34740 1062 34792 1114
rect 45662 1062 45714 1114
rect 45726 1062 45778 1114
rect 45790 1062 45842 1114
rect 45854 1062 45906 1114
rect 45918 1062 45970 1114
rect 6092 960 6144 1012
rect 10508 960 10560 1012
rect 11704 892 11756 944
rect 16580 892 16632 944
rect 16856 960 16908 1012
rect 22652 960 22704 1012
rect 19248 892 19300 944
rect 20812 824 20864 876
rect 8300 688 8352 740
rect 16580 688 16632 740
rect 23204 688 23256 740
rect 23664 620 23716 672
<< metal2 >>
rect 662 9840 718 10000
rect 1030 9840 1086 10000
rect 1398 9840 1454 10000
rect 1766 9840 1822 10000
rect 2134 9840 2190 10000
rect 2502 9840 2558 10000
rect 2870 9840 2926 10000
rect 3238 9840 3294 10000
rect 3606 9840 3662 10000
rect 3974 9840 4030 10000
rect 4342 9840 4398 10000
rect 4710 9840 4766 10000
rect 5078 9840 5134 10000
rect 5446 9840 5502 10000
rect 5814 9840 5870 10000
rect 6182 9840 6238 10000
rect 6550 9840 6606 10000
rect 6918 9840 6974 10000
rect 7286 9840 7342 10000
rect 7654 9840 7710 10000
rect 8022 9840 8078 10000
rect 8390 9840 8446 10000
rect 8758 9840 8814 10000
rect 9126 9840 9182 10000
rect 9404 9852 9456 9858
rect 676 8090 704 9840
rect 664 8084 716 8090
rect 664 8026 716 8032
rect 1044 7546 1072 9840
rect 1412 8022 1440 9840
rect 1492 9240 1544 9246
rect 1492 9182 1544 9188
rect 1504 8498 1532 9182
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1400 8016 1452 8022
rect 1400 7958 1452 7964
rect 1780 7546 1808 9840
rect 2148 8090 2176 9840
rect 2516 8634 2544 9840
rect 2686 8936 2742 8945
rect 2686 8871 2742 8880
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2700 8566 2728 8871
rect 2884 8634 2912 9840
rect 3252 8634 3280 9840
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 3344 8498 3372 8774
rect 3620 8634 3648 9840
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 1032 7540 1084 7546
rect 1032 7482 1084 7488
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 2332 7274 2360 7754
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2976 6905 3004 8434
rect 3988 8004 4016 9840
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4080 8566 4108 9454
rect 4356 8634 4384 9840
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 4160 8016 4212 8022
rect 3988 7976 4160 8004
rect 4160 7958 4212 7964
rect 4448 7886 4476 9658
rect 4724 8090 4752 9840
rect 5092 8634 5120 9840
rect 5460 8634 5488 9840
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5828 8090 5856 9840
rect 6196 8634 6224 9840
rect 6564 8786 6592 9840
rect 6932 9058 6960 9840
rect 7196 9784 7248 9790
rect 7196 9726 7248 9732
rect 6472 8758 6592 8786
rect 6840 9030 6960 9058
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 5816 8084 5868 8090
rect 6472 8072 6500 8758
rect 6840 8634 6868 9030
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6539 8188 6847 8197
rect 6539 8186 6545 8188
rect 6601 8186 6625 8188
rect 6681 8186 6705 8188
rect 6761 8186 6785 8188
rect 6841 8186 6847 8188
rect 6601 8134 6603 8186
rect 6783 8134 6785 8186
rect 6539 8132 6545 8134
rect 6601 8132 6625 8134
rect 6681 8132 6705 8134
rect 6761 8132 6785 8134
rect 6841 8132 6847 8134
rect 6539 8123 6847 8132
rect 6644 8084 6696 8090
rect 6472 8044 6644 8072
rect 5816 8026 5868 8032
rect 6644 8026 6696 8032
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 2962 6896 3018 6905
rect 2962 6831 3018 6840
rect 3988 6730 4016 7754
rect 4356 7478 4384 7822
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 6539 7100 6847 7109
rect 6539 7098 6545 7100
rect 6601 7098 6625 7100
rect 6681 7098 6705 7100
rect 6761 7098 6785 7100
rect 6841 7098 6847 7100
rect 6601 7046 6603 7098
rect 6783 7046 6785 7098
rect 6539 7044 6545 7046
rect 6601 7044 6625 7046
rect 6681 7044 6705 7046
rect 6761 7044 6785 7046
rect 6841 7044 6847 7046
rect 6539 7035 6847 7044
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 7024 6225 7052 8774
rect 7116 8498 7144 8774
rect 7208 8498 7236 9726
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7300 8090 7328 9840
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7576 8498 7604 9046
rect 7668 8634 7696 9840
rect 8036 8634 8064 9840
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8312 8498 8340 9318
rect 8404 8634 8432 9840
rect 8772 8634 8800 9840
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 9048 8498 9076 9454
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8220 8362 8432 8378
rect 8208 8356 8444 8362
rect 8260 8350 8392 8356
rect 8208 8298 8260 8304
rect 8392 8298 8444 8304
rect 7288 8084 7340 8090
rect 9140 8072 9168 9840
rect 9494 9840 9550 10000
rect 9862 9840 9918 10000
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9404 9794 9456 9800
rect 9416 9654 9444 9794
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9508 8634 9536 9840
rect 9680 9784 9732 9790
rect 9678 9752 9680 9761
rect 9732 9752 9734 9761
rect 9678 9687 9734 9696
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9784 8498 9812 8774
rect 9876 8634 9904 9840
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9968 8498 9996 9862
rect 10230 9840 10286 10000
rect 10598 9840 10654 10000
rect 10966 9840 11022 10000
rect 11334 9840 11390 10000
rect 11702 9840 11758 10000
rect 12070 9840 12126 10000
rect 12438 9840 12494 10000
rect 12806 9840 12862 10000
rect 13174 9840 13230 10000
rect 13542 9840 13598 10000
rect 13910 9840 13966 10000
rect 14278 9840 14334 10000
rect 14646 9840 14702 10000
rect 15014 9840 15070 10000
rect 15382 9840 15438 10000
rect 15750 9840 15806 10000
rect 16118 9840 16174 10000
rect 16486 9840 16542 10000
rect 16854 9840 16910 10000
rect 17222 9840 17278 10000
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 10244 8090 10272 9840
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10428 8566 10456 9114
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10520 8430 10548 8910
rect 10612 8634 10640 9840
rect 10980 8634 11008 9840
rect 11348 8634 11376 9840
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11532 8498 11560 8774
rect 11624 8498 11652 9522
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 9220 8084 9272 8090
rect 9140 8044 9220 8072
rect 7288 8026 7340 8032
rect 9220 8026 9272 8032
rect 10232 8084 10284 8090
rect 11716 8072 11744 9840
rect 12084 8922 12112 9840
rect 12452 9194 12480 9840
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12452 9166 12572 9194
rect 11992 8894 12112 8922
rect 11992 8634 12020 8894
rect 12128 8732 12436 8741
rect 12128 8730 12134 8732
rect 12190 8730 12214 8732
rect 12270 8730 12294 8732
rect 12350 8730 12374 8732
rect 12430 8730 12436 8732
rect 12190 8678 12192 8730
rect 12372 8678 12374 8730
rect 12128 8676 12134 8678
rect 12190 8676 12214 8678
rect 12270 8676 12294 8678
rect 12350 8676 12374 8678
rect 12430 8676 12436 8678
rect 12128 8667 12436 8676
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 12440 8628 12492 8634
rect 12544 8616 12572 9166
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12636 8634 12664 9046
rect 12492 8588 12572 8616
rect 12624 8628 12676 8634
rect 12440 8570 12492 8576
rect 12624 8570 12676 8576
rect 12728 8498 12756 9522
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12820 8090 12848 9840
rect 13084 9784 13136 9790
rect 13084 9726 13136 9732
rect 13096 8498 13124 9726
rect 13188 8634 13216 9840
rect 13556 8634 13584 9840
rect 13726 9208 13782 9217
rect 13726 9143 13782 9152
rect 13740 9042 13768 9143
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13924 8634 13952 9840
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 14108 8498 14136 8910
rect 14292 8820 14320 9840
rect 14292 8792 14412 8820
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 11796 8084 11848 8090
rect 11716 8044 11796 8072
rect 10232 8026 10284 8032
rect 11796 8026 11848 8032
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12530 7984 12586 7993
rect 12530 7919 12586 7928
rect 12544 7886 12572 7919
rect 9680 7880 9732 7886
rect 12532 7880 12584 7886
rect 9680 7822 9732 7828
rect 11794 7848 11850 7857
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8312 6361 8340 7414
rect 8298 6352 8354 6361
rect 8298 6287 8354 6296
rect 7010 6216 7066 6225
rect 7010 6151 7066 6160
rect 6539 6012 6847 6021
rect 6539 6010 6545 6012
rect 6601 6010 6625 6012
rect 6681 6010 6705 6012
rect 6761 6010 6785 6012
rect 6841 6010 6847 6012
rect 6601 5958 6603 6010
rect 6783 5958 6785 6010
rect 6539 5956 6545 5958
rect 6601 5956 6625 5958
rect 6681 5956 6705 5958
rect 6761 5956 6785 5958
rect 6841 5956 6847 5958
rect 6539 5947 6847 5956
rect 8956 5817 8984 7686
rect 9140 7478 9168 7754
rect 9692 7478 9720 7822
rect 11704 7812 11756 7818
rect 12532 7822 12584 7828
rect 11794 7783 11850 7792
rect 11704 7754 11756 7760
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9678 7304 9734 7313
rect 9678 7239 9680 7248
rect 9732 7239 9734 7248
rect 9680 7210 9732 7216
rect 11716 6769 11744 7754
rect 11808 7750 11836 7783
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 12128 7644 12436 7653
rect 12128 7642 12134 7644
rect 12190 7642 12214 7644
rect 12270 7642 12294 7644
rect 12350 7642 12374 7644
rect 12430 7642 12436 7644
rect 12190 7590 12192 7642
rect 12372 7590 12374 7642
rect 12128 7588 12134 7590
rect 12190 7588 12214 7590
rect 12270 7588 12294 7590
rect 12350 7588 12374 7590
rect 12430 7588 12436 7590
rect 12128 7579 12436 7588
rect 12636 7002 12664 8026
rect 14292 7818 14320 8230
rect 14384 8090 14412 8792
rect 14660 8634 14688 9840
rect 15028 8634 15056 9840
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15120 8537 15148 8774
rect 15396 8634 15424 9840
rect 15566 8664 15622 8673
rect 15384 8628 15436 8634
rect 15566 8599 15622 8608
rect 15384 8570 15436 8576
rect 15106 8528 15162 8537
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14924 8492 14976 8498
rect 14976 8452 15056 8480
rect 15580 8498 15608 8599
rect 15106 8463 15162 8472
rect 15568 8492 15620 8498
rect 14924 8434 14976 8440
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14476 7206 14504 8434
rect 15028 8378 15056 8452
rect 15568 8434 15620 8440
rect 15028 8350 15240 8378
rect 15106 7576 15162 7585
rect 15106 7511 15162 7520
rect 15120 7342 15148 7511
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 15212 7002 15240 8350
rect 15764 8090 15792 9840
rect 16132 8634 16160 9840
rect 16500 8634 16528 9840
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16592 8945 16620 9318
rect 16764 9308 16816 9314
rect 16764 9250 16816 9256
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16578 8936 16634 8945
rect 16578 8871 16634 8880
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16028 8492 16080 8498
rect 16080 8452 16620 8480
rect 16028 8434 16080 8440
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15488 7410 15516 7822
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 11702 6760 11758 6769
rect 11702 6695 11758 6704
rect 16592 6662 16620 8452
rect 16684 7274 16712 8978
rect 16776 8634 16804 9250
rect 16868 8634 16896 9840
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16960 8498 16988 8978
rect 17040 8832 17092 8838
rect 17144 8809 17172 9114
rect 17040 8774 17092 8780
rect 17130 8800 17186 8809
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16868 8401 16896 8434
rect 16854 8392 16910 8401
rect 17052 8362 17080 8774
rect 17130 8735 17186 8744
rect 17236 8634 17264 9840
rect 17420 9382 17448 9862
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17512 9246 17540 9862
rect 17590 9840 17646 10000
rect 17958 9840 18014 10000
rect 18144 9988 18196 9994
rect 18144 9930 18196 9936
rect 17500 9240 17552 9246
rect 17500 9182 17552 9188
rect 17604 8634 17632 9840
rect 17972 8634 18000 9840
rect 18052 9104 18104 9110
rect 18052 9046 18104 9052
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 16854 8327 16910 8336
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 17512 7886 17540 8366
rect 17604 8090 17632 8434
rect 17717 8188 18025 8197
rect 17717 8186 17723 8188
rect 17779 8186 17803 8188
rect 17859 8186 17883 8188
rect 17939 8186 17963 8188
rect 18019 8186 18025 8188
rect 17779 8134 17781 8186
rect 17961 8134 17963 8186
rect 17717 8132 17723 8134
rect 17779 8132 17803 8134
rect 17859 8132 17883 8134
rect 17939 8132 17963 8134
rect 18019 8132 18025 8134
rect 17717 8123 18025 8132
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 18064 7886 18092 9046
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17684 7744 17736 7750
rect 17222 7712 17278 7721
rect 17684 7686 17736 7692
rect 17222 7647 17278 7656
rect 17236 7342 17264 7647
rect 17696 7546 17724 7686
rect 17880 7546 17908 7754
rect 17972 7698 18000 7822
rect 18156 7698 18184 9930
rect 18326 9840 18382 10000
rect 18694 9840 18750 10000
rect 19062 9840 19118 10000
rect 19168 9846 19380 9874
rect 18236 9104 18288 9110
rect 18236 9046 18288 9052
rect 18248 7886 18276 9046
rect 18340 8090 18368 9840
rect 18708 8634 18736 9840
rect 19076 9738 19104 9840
rect 19168 9738 19196 9846
rect 19076 9710 19196 9738
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 19352 8566 19380 9846
rect 19430 9840 19486 10000
rect 19798 9840 19854 10000
rect 19904 9846 20116 9874
rect 19444 8616 19472 9840
rect 19616 9240 19668 9246
rect 19616 9182 19668 9188
rect 19524 8628 19576 8634
rect 19444 8588 19524 8616
rect 19524 8570 19576 8576
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 18418 8120 18474 8129
rect 18328 8084 18380 8090
rect 18418 8055 18474 8064
rect 18328 8026 18380 8032
rect 18432 8022 18460 8055
rect 18524 8022 18552 8502
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18708 8090 18736 8230
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 18512 8016 18564 8022
rect 18512 7958 18564 7964
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 17972 7670 18184 7698
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18800 7342 18828 8434
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19064 8288 19116 8294
rect 19352 8265 19380 8366
rect 19064 8230 19116 8236
rect 19338 8256 19394 8265
rect 19076 7410 19104 8230
rect 19338 8191 19394 8200
rect 19444 8090 19472 8434
rect 19628 8362 19656 9182
rect 19616 8356 19668 8362
rect 19616 8298 19668 8304
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 19720 7954 19748 8026
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 19260 7274 19288 7822
rect 19352 7546 19380 7822
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19338 7440 19394 7449
rect 19338 7375 19340 7384
rect 19392 7375 19394 7384
rect 19340 7346 19392 7352
rect 19536 7313 19564 7686
rect 19812 7410 19840 9840
rect 19904 8294 19932 9846
rect 20088 9738 20116 9846
rect 20166 9840 20222 10000
rect 20534 9840 20590 10000
rect 20902 9840 20958 10000
rect 21270 9840 21326 10000
rect 21456 9852 21508 9858
rect 20180 9738 20208 9840
rect 20088 9710 20208 9738
rect 20258 9752 20314 9761
rect 20314 9710 20484 9738
rect 20258 9687 20314 9696
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19522 7304 19578 7313
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 19248 7268 19300 7274
rect 19522 7239 19578 7248
rect 19248 7210 19300 7216
rect 17717 7100 18025 7109
rect 17717 7098 17723 7100
rect 17779 7098 17803 7100
rect 17859 7098 17883 7100
rect 17939 7098 17963 7100
rect 18019 7098 18025 7100
rect 17779 7046 17781 7098
rect 17961 7046 17963 7098
rect 17717 7044 17723 7046
rect 17779 7044 17803 7046
rect 17859 7044 17883 7046
rect 17939 7044 17963 7046
rect 18019 7044 18025 7046
rect 17717 7035 18025 7044
rect 18524 7041 18552 7210
rect 19064 7200 19116 7206
rect 19062 7168 19064 7177
rect 19116 7168 19118 7177
rect 19062 7103 19118 7112
rect 18510 7032 18566 7041
rect 18510 6967 18566 6976
rect 19720 6934 19748 7346
rect 19904 7342 19932 7822
rect 19996 7546 20024 8434
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20350 7848 20406 7857
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 20088 7585 20116 7686
rect 20074 7576 20130 7585
rect 19984 7540 20036 7546
rect 20180 7546 20208 7822
rect 20350 7783 20406 7792
rect 20364 7750 20392 7783
rect 20456 7750 20484 9710
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20074 7511 20130 7520
rect 20168 7540 20220 7546
rect 19984 7482 20036 7488
rect 20168 7482 20220 7488
rect 20548 7392 20576 9840
rect 20810 9208 20866 9217
rect 20810 9143 20812 9152
rect 20864 9143 20866 9152
rect 20812 9114 20864 9120
rect 20916 8650 20944 9840
rect 21088 9036 21140 9042
rect 21088 8978 21140 8984
rect 20824 8622 20944 8650
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 7886 20668 8230
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20628 7540 20680 7546
rect 20824 7528 20852 8622
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20916 7886 20944 8230
rect 21100 8090 21128 8978
rect 21284 8566 21312 9840
rect 21638 9840 21694 10000
rect 21824 9988 21876 9994
rect 21824 9930 21876 9936
rect 21730 9888 21786 9897
rect 21456 9794 21508 9800
rect 21362 9752 21418 9761
rect 21362 9687 21418 9696
rect 21376 9586 21404 9687
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21468 9042 21496 9794
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21560 9353 21588 9658
rect 21546 9344 21602 9353
rect 21546 9279 21602 9288
rect 21456 9036 21508 9042
rect 21456 8978 21508 8984
rect 21272 8560 21324 8566
rect 21272 8502 21324 8508
rect 21456 8424 21508 8430
rect 21178 8392 21234 8401
rect 21234 8350 21312 8378
rect 21652 8412 21680 9840
rect 21730 9823 21786 9832
rect 21744 9790 21772 9823
rect 21732 9784 21784 9790
rect 21732 9726 21784 9732
rect 21732 9648 21784 9654
rect 21730 9616 21732 9625
rect 21784 9616 21786 9625
rect 21730 9551 21786 9560
rect 21836 9518 21864 9930
rect 22006 9840 22062 10000
rect 22374 9840 22430 10000
rect 22652 9988 22704 9994
rect 22652 9930 22704 9936
rect 21732 9512 21784 9518
rect 21730 9480 21732 9489
rect 21824 9512 21876 9518
rect 21784 9480 21786 9489
rect 21824 9454 21876 9460
rect 21730 9415 21786 9424
rect 21732 9172 21784 9178
rect 21732 9114 21784 9120
rect 21508 8384 21680 8412
rect 21456 8366 21508 8372
rect 21178 8327 21234 8336
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 21192 7546 21220 8230
rect 21284 8106 21312 8350
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21284 8090 21404 8106
rect 21284 8084 21416 8090
rect 21284 8078 21364 8084
rect 21364 8026 21416 8032
rect 21364 7880 21416 7886
rect 21364 7822 21416 7828
rect 20680 7500 20852 7528
rect 21180 7540 21232 7546
rect 20628 7482 20680 7488
rect 21180 7482 21232 7488
rect 20812 7404 20864 7410
rect 20548 7364 20812 7392
rect 20812 7346 20864 7352
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 19708 6928 19760 6934
rect 19708 6870 19760 6876
rect 20732 6866 20760 7142
rect 21100 7002 21128 7142
rect 21376 7002 21404 7822
rect 21468 7546 21496 8230
rect 21744 7954 21772 9114
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21732 7948 21784 7954
rect 21732 7890 21784 7896
rect 21836 7886 21864 8570
rect 22020 8566 22048 9840
rect 22098 9480 22154 9489
rect 22098 9415 22154 9424
rect 22112 9246 22140 9415
rect 22100 9240 22152 9246
rect 22100 9182 22152 9188
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 21824 7880 21876 7886
rect 21546 7848 21602 7857
rect 22008 7880 22060 7886
rect 21824 7822 21876 7828
rect 22006 7848 22008 7857
rect 22060 7848 22062 7857
rect 21546 7783 21602 7792
rect 21916 7812 21968 7818
rect 21560 7546 21588 7783
rect 22006 7783 22062 7792
rect 21916 7754 21968 7760
rect 21732 7744 21784 7750
rect 21732 7686 21784 7692
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21548 7540 21600 7546
rect 21548 7482 21600 7488
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21652 7274 21680 7482
rect 21640 7268 21692 7274
rect 21640 7210 21692 7216
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 21364 6996 21416 7002
rect 21364 6938 21416 6944
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 12128 6556 12436 6565
rect 12128 6554 12134 6556
rect 12190 6554 12214 6556
rect 12270 6554 12294 6556
rect 12350 6554 12374 6556
rect 12430 6554 12436 6556
rect 12190 6502 12192 6554
rect 12372 6502 12374 6554
rect 12128 6500 12134 6502
rect 12190 6500 12214 6502
rect 12270 6500 12294 6502
rect 12350 6500 12374 6502
rect 12430 6500 12436 6502
rect 12128 6491 12436 6500
rect 17717 6012 18025 6021
rect 17717 6010 17723 6012
rect 17779 6010 17803 6012
rect 17859 6010 17883 6012
rect 17939 6010 17963 6012
rect 18019 6010 18025 6012
rect 17779 5958 17781 6010
rect 17961 5958 17963 6010
rect 17717 5956 17723 5958
rect 17779 5956 17803 5958
rect 17859 5956 17883 5958
rect 17939 5956 17963 5958
rect 18019 5956 18025 5958
rect 17717 5947 18025 5956
rect 21744 5817 21772 7686
rect 21928 7313 21956 7754
rect 22008 7744 22060 7750
rect 22006 7712 22008 7721
rect 22060 7712 22062 7721
rect 22006 7647 22062 7656
rect 21914 7304 21970 7313
rect 21914 7239 21970 7248
rect 22112 7154 22140 8774
rect 22388 8514 22416 9840
rect 22664 8922 22692 9930
rect 22742 9840 22798 10000
rect 23110 9840 23166 10000
rect 23216 9846 23428 9874
rect 22572 8894 22692 8922
rect 22466 8664 22522 8673
rect 22466 8599 22468 8608
rect 22520 8599 22522 8608
rect 22468 8570 22520 8576
rect 22204 8486 22416 8514
rect 22204 8430 22232 8486
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 22572 8378 22600 8894
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 22664 8498 22692 8774
rect 22756 8566 22784 9840
rect 23020 8968 23072 8974
rect 22834 8936 22890 8945
rect 22890 8894 22968 8922
rect 23020 8910 23072 8916
rect 22834 8871 22890 8880
rect 22834 8800 22890 8809
rect 22834 8735 22890 8744
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22284 8356 22336 8362
rect 22572 8350 22692 8378
rect 22284 8298 22336 8304
rect 22296 7410 22324 8298
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22558 8256 22614 8265
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 22388 7206 22416 8230
rect 22558 8191 22614 8200
rect 22572 8090 22600 8191
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 22664 7886 22692 8350
rect 22744 8288 22796 8294
rect 22744 8230 22796 8236
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 22756 7410 22784 8230
rect 22848 8090 22876 8735
rect 22940 8090 22968 8894
rect 23032 8634 23060 8910
rect 23020 8628 23072 8634
rect 23020 8570 23072 8576
rect 23124 8430 23152 9840
rect 23216 8548 23244 9846
rect 23400 9738 23428 9846
rect 23478 9840 23534 10000
rect 23846 9840 23902 10000
rect 24214 9840 24270 10000
rect 24492 9852 24544 9858
rect 23492 9738 23520 9840
rect 23400 9710 23520 9738
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 23754 9344 23810 9353
rect 23306 8732 23614 8741
rect 23306 8730 23312 8732
rect 23368 8730 23392 8732
rect 23448 8730 23472 8732
rect 23528 8730 23552 8732
rect 23608 8730 23614 8732
rect 23368 8678 23370 8730
rect 23550 8678 23552 8730
rect 23306 8676 23312 8678
rect 23368 8676 23392 8678
rect 23448 8676 23472 8678
rect 23528 8676 23552 8678
rect 23608 8676 23614 8678
rect 23306 8667 23614 8676
rect 23296 8560 23348 8566
rect 23216 8520 23296 8548
rect 23296 8502 23348 8508
rect 23478 8528 23534 8537
rect 23478 8463 23480 8472
rect 23532 8463 23534 8472
rect 23480 8434 23532 8440
rect 23112 8424 23164 8430
rect 23112 8366 23164 8372
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 22928 8084 22980 8090
rect 22928 8026 22980 8032
rect 23032 7954 23060 8230
rect 23400 7970 23428 8230
rect 23676 8090 23704 9318
rect 23754 9279 23810 9288
rect 23768 8362 23796 9279
rect 23860 8537 23888 9840
rect 23940 9512 23992 9518
rect 23940 9454 23992 9460
rect 23952 8634 23980 9454
rect 24124 9036 24176 9042
rect 24124 8978 24176 8984
rect 24032 8900 24084 8906
rect 24032 8842 24084 8848
rect 24044 8634 24072 8842
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 24032 8628 24084 8634
rect 24032 8570 24084 8576
rect 23846 8528 23902 8537
rect 23846 8463 23902 8472
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23940 8288 23992 8294
rect 23860 8236 23940 8242
rect 23860 8230 23992 8236
rect 23860 8214 23980 8230
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 23124 7942 23428 7970
rect 23572 8016 23624 8022
rect 23624 7964 23796 7970
rect 23572 7958 23796 7964
rect 23584 7942 23796 7958
rect 23124 7886 23152 7942
rect 23112 7880 23164 7886
rect 23112 7822 23164 7828
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23216 7528 23244 7822
rect 23306 7644 23614 7653
rect 23306 7642 23312 7644
rect 23368 7642 23392 7644
rect 23448 7642 23472 7644
rect 23528 7642 23552 7644
rect 23608 7642 23614 7644
rect 23368 7590 23370 7642
rect 23550 7590 23552 7642
rect 23306 7588 23312 7590
rect 23368 7588 23392 7590
rect 23448 7588 23472 7590
rect 23528 7588 23552 7590
rect 23608 7588 23614 7590
rect 23306 7579 23614 7588
rect 23388 7540 23440 7546
rect 23216 7500 23336 7528
rect 23308 7410 23336 7500
rect 23388 7482 23440 7488
rect 22744 7404 22796 7410
rect 22744 7346 22796 7352
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 23296 7404 23348 7410
rect 23296 7346 23348 7352
rect 23216 7290 23244 7346
rect 23400 7290 23428 7482
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 23216 7262 23428 7290
rect 23478 7304 23534 7313
rect 23478 7239 23480 7248
rect 23532 7239 23534 7248
rect 23480 7210 23532 7216
rect 22284 7200 22336 7206
rect 22112 7148 22284 7154
rect 22112 7142 22336 7148
rect 22376 7200 22428 7206
rect 23204 7200 23256 7206
rect 22376 7142 22428 7148
rect 23202 7168 23204 7177
rect 23584 7177 23612 7346
rect 23768 7313 23796 7942
rect 23860 7410 23888 8214
rect 24136 7750 24164 8978
rect 24228 8498 24256 9840
rect 24582 9840 24638 10000
rect 24688 9846 24900 9874
rect 24492 9794 24544 9800
rect 24400 9240 24452 9246
rect 24400 9182 24452 9188
rect 24308 8900 24360 8906
rect 24308 8842 24360 8848
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24320 8362 24348 8842
rect 24308 8356 24360 8362
rect 24308 8298 24360 8304
rect 24214 8120 24270 8129
rect 24214 8055 24216 8064
rect 24268 8055 24270 8064
rect 24216 8026 24268 8032
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 23754 7304 23810 7313
rect 23754 7239 23810 7248
rect 24412 7206 24440 9182
rect 24504 8514 24532 9794
rect 24596 9738 24624 9840
rect 24688 9738 24716 9846
rect 24596 9710 24716 9738
rect 24768 9240 24820 9246
rect 24768 9182 24820 9188
rect 24504 8486 24624 8514
rect 24492 8424 24544 8430
rect 24492 8366 24544 8372
rect 24504 7886 24532 8366
rect 24596 8090 24624 8486
rect 24780 8362 24808 9182
rect 24872 8498 24900 9846
rect 24950 9840 25006 10000
rect 25318 9840 25374 10000
rect 25686 9840 25742 10000
rect 26054 9840 26110 10000
rect 26422 9840 26478 10000
rect 26698 9888 26754 9897
rect 24964 8498 24992 9840
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 25044 8288 25096 8294
rect 25044 8230 25096 8236
rect 24584 8084 24636 8090
rect 24584 8026 24636 8032
rect 24688 7886 24716 8230
rect 25056 7886 25084 8230
rect 25148 8090 25176 8502
rect 25332 8498 25360 9840
rect 25594 9072 25650 9081
rect 25594 9007 25650 9016
rect 25320 8492 25372 8498
rect 25320 8434 25372 8440
rect 25608 8378 25636 9007
rect 25700 8498 25728 9840
rect 26068 8498 26096 9840
rect 26148 9376 26200 9382
rect 26148 9318 26200 9324
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 25688 8492 25740 8498
rect 25688 8434 25740 8440
rect 26056 8492 26108 8498
rect 26056 8434 26108 8440
rect 25608 8350 25728 8378
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25596 8288 25648 8294
rect 25596 8230 25648 8236
rect 25424 8090 25452 8230
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 25412 8084 25464 8090
rect 25412 8026 25464 8032
rect 25504 8016 25556 8022
rect 25502 7984 25504 7993
rect 25556 7984 25558 7993
rect 25502 7919 25558 7928
rect 25608 7886 25636 8230
rect 25700 8090 25728 8350
rect 26056 8356 26108 8362
rect 26056 8298 26108 8304
rect 25872 8288 25924 8294
rect 25872 8230 25924 8236
rect 25688 8084 25740 8090
rect 25688 8026 25740 8032
rect 25884 7886 25912 8230
rect 26068 7886 26096 8298
rect 26160 8090 26188 9318
rect 26252 9217 26280 9318
rect 26238 9208 26294 9217
rect 26238 9143 26294 9152
rect 26436 8498 26464 9840
rect 26790 9840 26846 10000
rect 27158 9840 27214 10000
rect 27264 9846 27476 9874
rect 26698 9823 26754 9832
rect 26424 8492 26476 8498
rect 26424 8434 26476 8440
rect 26424 8288 26476 8294
rect 26424 8230 26476 8236
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 26436 7886 26464 8230
rect 26712 8090 26740 9823
rect 26804 8498 26832 9840
rect 27066 9752 27122 9761
rect 27172 9738 27200 9840
rect 27264 9738 27292 9846
rect 27172 9710 27292 9738
rect 27066 9687 27122 9696
rect 26792 8492 26844 8498
rect 26792 8434 26844 8440
rect 26792 8356 26844 8362
rect 26792 8298 26844 8304
rect 26700 8084 26752 8090
rect 26700 8026 26752 8032
rect 26804 7954 26832 8298
rect 27080 8090 27108 9687
rect 27252 8900 27304 8906
rect 27252 8842 27304 8848
rect 27264 8634 27292 8842
rect 27252 8628 27304 8634
rect 27252 8570 27304 8576
rect 27344 8628 27396 8634
rect 27344 8570 27396 8576
rect 27160 8356 27212 8362
rect 27160 8298 27212 8304
rect 27068 8084 27120 8090
rect 27068 8026 27120 8032
rect 26792 7948 26844 7954
rect 26792 7890 26844 7896
rect 27172 7886 27200 8298
rect 27356 7954 27384 8570
rect 27448 8498 27476 9846
rect 27526 9840 27582 10000
rect 27894 9840 27950 10000
rect 28262 9840 28318 10000
rect 28630 9840 28686 10000
rect 28998 9840 29054 10000
rect 29366 9840 29422 10000
rect 29734 9840 29790 10000
rect 29840 9846 30052 9874
rect 27540 8498 27568 9840
rect 27804 9308 27856 9314
rect 27804 9250 27856 9256
rect 27436 8492 27488 8498
rect 27436 8434 27488 8440
rect 27528 8492 27580 8498
rect 27528 8434 27580 8440
rect 27434 8392 27490 8401
rect 27434 8327 27490 8336
rect 27344 7948 27396 7954
rect 27344 7890 27396 7896
rect 27448 7886 27476 8327
rect 27528 8288 27580 8294
rect 27528 8230 27580 8236
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 24676 7880 24728 7886
rect 25044 7880 25096 7886
rect 24676 7822 24728 7828
rect 24766 7848 24822 7857
rect 25044 7822 25096 7828
rect 25596 7880 25648 7886
rect 25596 7822 25648 7828
rect 25872 7880 25924 7886
rect 25872 7822 25924 7828
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 26424 7880 26476 7886
rect 26424 7822 26476 7828
rect 27160 7880 27212 7886
rect 27160 7822 27212 7828
rect 27436 7880 27488 7886
rect 27436 7822 27488 7828
rect 24766 7783 24822 7792
rect 23848 7200 23900 7206
rect 23256 7168 23258 7177
rect 22112 7126 22324 7142
rect 23202 7103 23258 7112
rect 23570 7168 23626 7177
rect 23848 7142 23900 7148
rect 24400 7200 24452 7206
rect 24780 7177 24808 7783
rect 25044 7744 25096 7750
rect 25044 7686 25096 7692
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25596 7744 25648 7750
rect 25596 7686 25648 7692
rect 26424 7744 26476 7750
rect 26424 7686 26476 7692
rect 24400 7142 24452 7148
rect 24766 7168 24822 7177
rect 23570 7103 23626 7112
rect 23860 7041 23888 7142
rect 24766 7103 24822 7112
rect 23846 7032 23902 7041
rect 23846 6967 23902 6976
rect 23306 6556 23614 6565
rect 23306 6554 23312 6556
rect 23368 6554 23392 6556
rect 23448 6554 23472 6556
rect 23528 6554 23552 6556
rect 23608 6554 23614 6556
rect 23368 6502 23370 6554
rect 23550 6502 23552 6554
rect 23306 6500 23312 6502
rect 23368 6500 23392 6502
rect 23448 6500 23472 6502
rect 23528 6500 23552 6502
rect 23608 6500 23614 6502
rect 23306 6491 23614 6500
rect 24952 6248 25004 6254
rect 25056 6225 25084 7686
rect 25332 6730 25360 7686
rect 25608 6905 25636 7686
rect 25594 6896 25650 6905
rect 25594 6831 25650 6840
rect 25320 6724 25372 6730
rect 25320 6666 25372 6672
rect 26436 6361 26464 7686
rect 27540 7410 27568 8230
rect 27816 8090 27844 9250
rect 27908 8498 27936 9840
rect 28170 9616 28226 9625
rect 28170 9551 28226 9560
rect 27896 8492 27948 8498
rect 27896 8434 27948 8440
rect 27896 8288 27948 8294
rect 27896 8230 27948 8236
rect 27804 8084 27856 8090
rect 27804 8026 27856 8032
rect 27908 7886 27936 8230
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 28184 7750 28212 9551
rect 28276 8498 28304 9840
rect 28644 8498 28672 9840
rect 29012 8498 29040 9840
rect 29380 8498 29408 9840
rect 29748 9738 29776 9840
rect 29840 9738 29868 9846
rect 29748 9710 29868 9738
rect 30024 8498 30052 9846
rect 30102 9840 30158 10000
rect 30470 9840 30526 10000
rect 30838 9840 30894 10000
rect 31206 9840 31262 10000
rect 31574 9840 31630 10000
rect 31942 9840 31998 10000
rect 32310 9840 32366 10000
rect 32678 9840 32734 10000
rect 32956 9988 33008 9994
rect 32956 9930 33008 9936
rect 30116 8498 30144 9840
rect 30288 8968 30340 8974
rect 30288 8910 30340 8916
rect 30300 8634 30328 8910
rect 30288 8628 30340 8634
rect 30288 8570 30340 8576
rect 30484 8498 30512 9840
rect 30852 8498 30880 9840
rect 31024 9240 31076 9246
rect 31024 9182 31076 9188
rect 30932 8900 30984 8906
rect 30932 8842 30984 8848
rect 30944 8634 30972 8842
rect 31036 8634 31064 9182
rect 30932 8628 30984 8634
rect 30932 8570 30984 8576
rect 31024 8628 31076 8634
rect 31024 8570 31076 8576
rect 31220 8498 31248 9840
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 28632 8492 28684 8498
rect 28632 8434 28684 8440
rect 29000 8492 29052 8498
rect 29000 8434 29052 8440
rect 29368 8492 29420 8498
rect 29368 8434 29420 8440
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 30104 8492 30156 8498
rect 30104 8434 30156 8440
rect 30472 8492 30524 8498
rect 30472 8434 30524 8440
rect 30840 8492 30892 8498
rect 30840 8434 30892 8440
rect 31208 8492 31260 8498
rect 31588 8480 31616 9840
rect 31852 8832 31904 8838
rect 31852 8774 31904 8780
rect 31668 8492 31720 8498
rect 31588 8452 31668 8480
rect 31208 8434 31260 8440
rect 31668 8434 31720 8440
rect 31760 8424 31812 8430
rect 31680 8372 31760 8378
rect 31680 8366 31812 8372
rect 30656 8356 30708 8362
rect 30656 8298 30708 8304
rect 31680 8350 31800 8366
rect 28724 8288 28776 8294
rect 28724 8230 28776 8236
rect 29276 8288 29328 8294
rect 29276 8230 29328 8236
rect 29552 8288 29604 8294
rect 29552 8230 29604 8236
rect 29828 8288 29880 8294
rect 29828 8230 29880 8236
rect 28736 8022 28764 8230
rect 28895 8188 29203 8197
rect 28895 8186 28901 8188
rect 28957 8186 28981 8188
rect 29037 8186 29061 8188
rect 29117 8186 29141 8188
rect 29197 8186 29203 8188
rect 28957 8134 28959 8186
rect 29139 8134 29141 8186
rect 28895 8132 28901 8134
rect 28957 8132 28981 8134
rect 29037 8132 29061 8134
rect 29117 8132 29141 8134
rect 29197 8132 29203 8134
rect 28895 8123 29203 8132
rect 29288 8090 29316 8230
rect 29276 8084 29328 8090
rect 29276 8026 29328 8032
rect 28724 8016 28776 8022
rect 28724 7958 28776 7964
rect 29564 7886 29592 8230
rect 29840 7886 29868 8230
rect 29552 7880 29604 7886
rect 29552 7822 29604 7828
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 28172 7744 28224 7750
rect 28172 7686 28224 7692
rect 28540 7744 28592 7750
rect 28540 7686 28592 7692
rect 27528 7404 27580 7410
rect 27528 7346 27580 7352
rect 28552 6769 28580 7686
rect 30668 7342 30696 8298
rect 31680 7721 31708 8350
rect 31666 7712 31722 7721
rect 31666 7647 31722 7656
rect 31864 7546 31892 8774
rect 31956 8480 31984 9840
rect 32220 9240 32272 9246
rect 32220 9182 32272 9188
rect 32128 8492 32180 8498
rect 31956 8452 32128 8480
rect 32128 8434 32180 8440
rect 31944 8356 31996 8362
rect 31944 8298 31996 8304
rect 31852 7540 31904 7546
rect 31852 7482 31904 7488
rect 31956 7449 31984 8298
rect 31942 7440 31998 7449
rect 31942 7375 31998 7384
rect 30656 7336 30708 7342
rect 30656 7278 30708 7284
rect 28895 7100 29203 7109
rect 28895 7098 28901 7100
rect 28957 7098 28981 7100
rect 29037 7098 29061 7100
rect 29117 7098 29141 7100
rect 29197 7098 29203 7100
rect 28957 7046 28959 7098
rect 29139 7046 29141 7098
rect 28895 7044 28901 7046
rect 28957 7044 28981 7046
rect 29037 7044 29061 7046
rect 29117 7044 29141 7046
rect 29197 7044 29203 7046
rect 28895 7035 29203 7044
rect 28538 6760 28594 6769
rect 28538 6695 28594 6704
rect 26422 6352 26478 6361
rect 26422 6287 26478 6296
rect 24952 6190 25004 6196
rect 25042 6216 25098 6225
rect 8942 5808 8998 5817
rect 8942 5743 8998 5752
rect 21730 5808 21786 5817
rect 21730 5743 21786 5752
rect 12128 5468 12436 5477
rect 12128 5466 12134 5468
rect 12190 5466 12214 5468
rect 12270 5466 12294 5468
rect 12350 5466 12374 5468
rect 12430 5466 12436 5468
rect 12190 5414 12192 5466
rect 12372 5414 12374 5466
rect 12128 5412 12134 5414
rect 12190 5412 12214 5414
rect 12270 5412 12294 5414
rect 12350 5412 12374 5414
rect 12430 5412 12436 5414
rect 12128 5403 12436 5412
rect 23306 5468 23614 5477
rect 23306 5466 23312 5468
rect 23368 5466 23392 5468
rect 23448 5466 23472 5468
rect 23528 5466 23552 5468
rect 23608 5466 23614 5468
rect 23368 5414 23370 5466
rect 23550 5414 23552 5466
rect 23306 5412 23312 5414
rect 23368 5412 23392 5414
rect 23448 5412 23472 5414
rect 23528 5412 23552 5414
rect 23608 5412 23614 5414
rect 23306 5403 23614 5412
rect 6539 4924 6847 4933
rect 6539 4922 6545 4924
rect 6601 4922 6625 4924
rect 6681 4922 6705 4924
rect 6761 4922 6785 4924
rect 6841 4922 6847 4924
rect 6601 4870 6603 4922
rect 6783 4870 6785 4922
rect 6539 4868 6545 4870
rect 6601 4868 6625 4870
rect 6681 4868 6705 4870
rect 6761 4868 6785 4870
rect 6841 4868 6847 4870
rect 6539 4859 6847 4868
rect 17717 4924 18025 4933
rect 17717 4922 17723 4924
rect 17779 4922 17803 4924
rect 17859 4922 17883 4924
rect 17939 4922 17963 4924
rect 18019 4922 18025 4924
rect 17779 4870 17781 4922
rect 17961 4870 17963 4922
rect 17717 4868 17723 4870
rect 17779 4868 17803 4870
rect 17859 4868 17883 4870
rect 17939 4868 17963 4870
rect 18019 4868 18025 4870
rect 17717 4859 18025 4868
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 12128 4380 12436 4389
rect 12128 4378 12134 4380
rect 12190 4378 12214 4380
rect 12270 4378 12294 4380
rect 12350 4378 12374 4380
rect 12430 4378 12436 4380
rect 12190 4326 12192 4378
rect 12372 4326 12374 4378
rect 12128 4324 12134 4326
rect 12190 4324 12214 4326
rect 12270 4324 12294 4326
rect 12350 4324 12374 4326
rect 12430 4324 12436 4326
rect 12128 4315 12436 4324
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 6539 3836 6847 3845
rect 6539 3834 6545 3836
rect 6601 3834 6625 3836
rect 6681 3834 6705 3836
rect 6761 3834 6785 3836
rect 6841 3834 6847 3836
rect 6601 3782 6603 3834
rect 6783 3782 6785 3834
rect 6539 3780 6545 3782
rect 6601 3780 6625 3782
rect 6681 3780 6705 3782
rect 6761 3780 6785 3782
rect 6841 3780 6847 3782
rect 6539 3771 6847 3780
rect 17717 3836 18025 3845
rect 17717 3834 17723 3836
rect 17779 3834 17803 3836
rect 17859 3834 17883 3836
rect 17939 3834 17963 3836
rect 18019 3834 18025 3836
rect 17779 3782 17781 3834
rect 17961 3782 17963 3834
rect 17717 3780 17723 3782
rect 17779 3780 17803 3782
rect 17859 3780 17883 3782
rect 17939 3780 17963 3782
rect 18019 3780 18025 3782
rect 17717 3771 18025 3780
rect 12128 3292 12436 3301
rect 12128 3290 12134 3292
rect 12190 3290 12214 3292
rect 12270 3290 12294 3292
rect 12350 3290 12374 3292
rect 12430 3290 12436 3292
rect 12190 3238 12192 3290
rect 12372 3238 12374 3290
rect 12128 3236 12134 3238
rect 12190 3236 12214 3238
rect 12270 3236 12294 3238
rect 12350 3236 12374 3238
rect 12430 3236 12436 3238
rect 12128 3227 12436 3236
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 6539 2748 6847 2757
rect 6539 2746 6545 2748
rect 6601 2746 6625 2748
rect 6681 2746 6705 2748
rect 6761 2746 6785 2748
rect 6841 2746 6847 2748
rect 6601 2694 6603 2746
rect 6783 2694 6785 2746
rect 6539 2692 6545 2694
rect 6601 2692 6625 2694
rect 6681 2692 6705 2694
rect 6761 2692 6785 2694
rect 6841 2692 6847 2694
rect 6539 2683 6847 2692
rect 17717 2748 18025 2757
rect 17717 2746 17723 2748
rect 17779 2746 17803 2748
rect 17859 2746 17883 2748
rect 17939 2746 17963 2748
rect 18019 2746 18025 2748
rect 17779 2694 17781 2746
rect 17961 2694 17963 2746
rect 17717 2692 17723 2694
rect 17779 2692 17803 2694
rect 17859 2692 17883 2694
rect 17939 2692 17963 2694
rect 18019 2692 18025 2694
rect 17717 2683 18025 2692
rect 12128 2204 12436 2213
rect 12128 2202 12134 2204
rect 12190 2202 12214 2204
rect 12270 2202 12294 2204
rect 12350 2202 12374 2204
rect 12430 2202 12436 2204
rect 12190 2150 12192 2202
rect 12372 2150 12374 2202
rect 12128 2148 12134 2150
rect 12190 2148 12214 2150
rect 12270 2148 12294 2150
rect 12350 2148 12374 2150
rect 12430 2148 12436 2150
rect 12128 2139 12436 2148
rect 1676 1896 1728 1902
rect 1676 1838 1728 1844
rect 1688 1562 1716 1838
rect 6539 1660 6847 1669
rect 6539 1658 6545 1660
rect 6601 1658 6625 1660
rect 6681 1658 6705 1660
rect 6761 1658 6785 1660
rect 6841 1658 6847 1660
rect 6601 1606 6603 1658
rect 6783 1606 6785 1658
rect 6539 1604 6545 1606
rect 6601 1604 6625 1606
rect 6681 1604 6705 1606
rect 6761 1604 6785 1606
rect 6841 1604 6847 1606
rect 6539 1595 6847 1604
rect 17717 1660 18025 1669
rect 17717 1658 17723 1660
rect 17779 1658 17803 1660
rect 17859 1658 17883 1660
rect 17939 1658 17963 1660
rect 18019 1658 18025 1660
rect 17779 1606 17781 1658
rect 17961 1606 17963 1658
rect 17717 1604 17723 1606
rect 17779 1604 17803 1606
rect 17859 1604 17883 1606
rect 17939 1604 17963 1606
rect 18019 1604 18025 1606
rect 17717 1595 18025 1604
rect 1676 1556 1728 1562
rect 1676 1498 1728 1504
rect 1492 1352 1544 1358
rect 1492 1294 1544 1300
rect 3792 1352 3844 1358
rect 3792 1294 3844 1300
rect 5908 1352 5960 1358
rect 5908 1294 5960 1300
rect 8116 1352 8168 1358
rect 8116 1294 8168 1300
rect 10324 1352 10376 1358
rect 10324 1294 10376 1300
rect 12532 1352 12584 1358
rect 12532 1294 12584 1300
rect 14740 1352 14792 1358
rect 14740 1294 14792 1300
rect 17132 1352 17184 1358
rect 17132 1294 17184 1300
rect 1398 82 1454 160
rect 1504 82 1532 1294
rect 1398 54 1532 82
rect 3606 82 3662 160
rect 3804 82 3832 1294
rect 3606 54 3832 82
rect 5814 82 5870 160
rect 5920 82 5948 1294
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 6104 1018 6132 1158
rect 6092 1012 6144 1018
rect 6092 954 6144 960
rect 5814 54 5948 82
rect 8022 82 8078 160
rect 8128 82 8156 1294
rect 8300 1216 8352 1222
rect 8300 1158 8352 1164
rect 8312 746 8340 1158
rect 8300 740 8352 746
rect 8300 682 8352 688
rect 8022 54 8156 82
rect 10230 82 10286 160
rect 10336 82 10364 1294
rect 10508 1216 10560 1222
rect 10508 1158 10560 1164
rect 11704 1216 11756 1222
rect 11704 1158 11756 1164
rect 10520 1018 10548 1158
rect 10508 1012 10560 1018
rect 10508 954 10560 960
rect 11716 950 11744 1158
rect 12128 1116 12436 1125
rect 12128 1114 12134 1116
rect 12190 1114 12214 1116
rect 12270 1114 12294 1116
rect 12350 1114 12374 1116
rect 12430 1114 12436 1116
rect 12190 1062 12192 1114
rect 12372 1062 12374 1114
rect 12128 1060 12134 1062
rect 12190 1060 12214 1062
rect 12270 1060 12294 1062
rect 12350 1060 12374 1062
rect 12430 1060 12436 1062
rect 12128 1051 12436 1060
rect 11704 944 11756 950
rect 11704 886 11756 892
rect 10230 54 10364 82
rect 12438 82 12494 160
rect 12544 82 12572 1294
rect 12438 54 12572 82
rect 14646 82 14702 160
rect 14752 82 14780 1294
rect 16856 1216 16908 1222
rect 16856 1158 16908 1164
rect 16868 1018 16896 1158
rect 16856 1012 16908 1018
rect 16856 954 16908 960
rect 16580 944 16632 950
rect 16580 886 16632 892
rect 16592 746 16620 886
rect 16580 740 16632 746
rect 16580 682 16632 688
rect 14646 54 14780 82
rect 16854 82 16910 160
rect 17144 82 17172 1294
rect 19260 950 19288 2994
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 20640 2106 20668 2314
rect 20628 2100 20680 2106
rect 20628 2042 20680 2048
rect 19800 1964 19852 1970
rect 19800 1906 19852 1912
rect 19812 1562 19840 1906
rect 19800 1556 19852 1562
rect 19800 1498 19852 1504
rect 20732 1358 20760 2382
rect 19432 1352 19484 1358
rect 19432 1294 19484 1300
rect 20720 1352 20772 1358
rect 20720 1294 20772 1300
rect 19248 944 19300 950
rect 19248 886 19300 892
rect 16854 54 17172 82
rect 19062 82 19118 160
rect 19444 82 19472 1294
rect 20824 882 20852 4014
rect 22664 3738 22692 4082
rect 22652 3732 22704 3738
rect 22652 3674 22704 3680
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 20904 1964 20956 1970
rect 20904 1906 20956 1912
rect 20916 1290 20944 1906
rect 20904 1284 20956 1290
rect 20904 1226 20956 1232
rect 21376 1222 21404 3470
rect 23032 3194 23060 3470
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 23032 2106 23060 2382
rect 23124 2106 23152 4762
rect 23664 4616 23716 4622
rect 23664 4558 23716 4564
rect 23306 4380 23614 4389
rect 23306 4378 23312 4380
rect 23368 4378 23392 4380
rect 23448 4378 23472 4380
rect 23528 4378 23552 4380
rect 23608 4378 23614 4380
rect 23368 4326 23370 4378
rect 23550 4326 23552 4378
rect 23306 4324 23312 4326
rect 23368 4324 23392 4326
rect 23448 4324 23472 4326
rect 23528 4324 23552 4326
rect 23608 4324 23614 4326
rect 23306 4315 23614 4324
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23216 3194 23244 4082
rect 23676 4010 23704 4558
rect 23664 4004 23716 4010
rect 23664 3946 23716 3952
rect 23940 3460 23992 3466
rect 23940 3402 23992 3408
rect 23306 3292 23614 3301
rect 23306 3290 23312 3292
rect 23368 3290 23392 3292
rect 23448 3290 23472 3292
rect 23528 3290 23552 3292
rect 23608 3290 23614 3292
rect 23368 3238 23370 3290
rect 23550 3238 23552 3290
rect 23306 3236 23312 3238
rect 23368 3236 23392 3238
rect 23448 3236 23472 3238
rect 23528 3236 23552 3238
rect 23608 3236 23614 3238
rect 23306 3227 23614 3236
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 23584 2582 23612 2994
rect 23664 2984 23716 2990
rect 23664 2926 23716 2932
rect 23572 2576 23624 2582
rect 23572 2518 23624 2524
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23216 2106 23244 2382
rect 23306 2204 23614 2213
rect 23306 2202 23312 2204
rect 23368 2202 23392 2204
rect 23448 2202 23472 2204
rect 23528 2202 23552 2204
rect 23608 2202 23614 2204
rect 23368 2150 23370 2202
rect 23550 2150 23552 2202
rect 23306 2148 23312 2150
rect 23368 2148 23392 2150
rect 23448 2148 23472 2150
rect 23528 2148 23552 2150
rect 23608 2148 23614 2150
rect 23306 2139 23614 2148
rect 23020 2100 23072 2106
rect 23020 2042 23072 2048
rect 23112 2100 23164 2106
rect 23112 2042 23164 2048
rect 23204 2100 23256 2106
rect 23204 2042 23256 2048
rect 23204 1964 23256 1970
rect 23204 1906 23256 1912
rect 22652 1896 22704 1902
rect 22652 1838 22704 1844
rect 21548 1352 21600 1358
rect 21548 1294 21600 1300
rect 21364 1216 21416 1222
rect 21364 1158 21416 1164
rect 20812 876 20864 882
rect 20812 818 20864 824
rect 19062 54 19472 82
rect 21270 82 21326 160
rect 21560 82 21588 1294
rect 22664 1018 22692 1838
rect 22652 1012 22704 1018
rect 22652 954 22704 960
rect 23216 746 23244 1906
rect 23306 1116 23614 1125
rect 23306 1114 23312 1116
rect 23368 1114 23392 1116
rect 23448 1114 23472 1116
rect 23528 1114 23552 1116
rect 23608 1114 23614 1116
rect 23368 1062 23370 1114
rect 23550 1062 23552 1114
rect 23306 1060 23312 1062
rect 23368 1060 23392 1062
rect 23448 1060 23472 1062
rect 23528 1060 23552 1062
rect 23608 1060 23614 1062
rect 23306 1051 23614 1060
rect 23204 740 23256 746
rect 23204 682 23256 688
rect 23676 678 23704 2926
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 23860 2106 23888 2382
rect 23952 2310 23980 3402
rect 24964 2582 24992 6190
rect 25042 6151 25098 6160
rect 27252 6180 27304 6186
rect 27252 6122 27304 6128
rect 27068 4140 27120 4146
rect 27068 4082 27120 4088
rect 27080 3194 27108 4082
rect 27264 3942 27292 6122
rect 28895 6012 29203 6021
rect 28895 6010 28901 6012
rect 28957 6010 28981 6012
rect 29037 6010 29061 6012
rect 29117 6010 29141 6012
rect 29197 6010 29203 6012
rect 28957 5958 28959 6010
rect 29139 5958 29141 6010
rect 28895 5956 28901 5958
rect 28957 5956 28981 5958
rect 29037 5956 29061 5958
rect 29117 5956 29141 5958
rect 29197 5956 29203 5958
rect 28895 5947 29203 5956
rect 28895 4924 29203 4933
rect 28895 4922 28901 4924
rect 28957 4922 28981 4924
rect 29037 4922 29061 4924
rect 29117 4922 29141 4924
rect 29197 4922 29203 4924
rect 28957 4870 28959 4922
rect 29139 4870 29141 4922
rect 28895 4868 28901 4870
rect 28957 4868 28981 4870
rect 29037 4868 29061 4870
rect 29117 4868 29141 4870
rect 29197 4868 29203 4870
rect 28895 4859 29203 4868
rect 27252 3936 27304 3942
rect 27252 3878 27304 3884
rect 28895 3836 29203 3845
rect 28895 3834 28901 3836
rect 28957 3834 28981 3836
rect 29037 3834 29061 3836
rect 29117 3834 29141 3836
rect 29197 3834 29203 3836
rect 28957 3782 28959 3834
rect 29139 3782 29141 3834
rect 28895 3780 28901 3782
rect 28957 3780 28981 3782
rect 29037 3780 29061 3782
rect 29117 3780 29141 3782
rect 29197 3780 29203 3782
rect 28895 3771 29203 3780
rect 32232 3670 32260 9182
rect 32324 8480 32352 9840
rect 32404 8492 32456 8498
rect 32324 8452 32404 8480
rect 32692 8480 32720 9840
rect 32864 9444 32916 9450
rect 32864 9386 32916 9392
rect 32772 9104 32824 9110
rect 32772 9046 32824 9052
rect 32784 8634 32812 9046
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 32876 8566 32904 9386
rect 32864 8560 32916 8566
rect 32864 8502 32916 8508
rect 32772 8492 32824 8498
rect 32692 8452 32772 8480
rect 32404 8434 32456 8440
rect 32772 8434 32824 8440
rect 32968 8294 32996 9930
rect 33046 9840 33102 10000
rect 33414 9840 33470 10000
rect 33782 9840 33838 10000
rect 34150 9840 34206 10000
rect 34518 9840 34574 10000
rect 34886 9840 34942 10000
rect 35254 9840 35310 10000
rect 35622 9840 35678 10000
rect 35990 9840 36046 10000
rect 36358 9840 36414 10000
rect 36726 9840 36782 10000
rect 37094 9840 37150 10000
rect 37462 9840 37518 10000
rect 37830 9840 37886 10000
rect 38198 9840 38254 10000
rect 38566 9840 38622 10000
rect 38934 9840 38990 10000
rect 39302 9840 39358 10000
rect 39670 9840 39726 10000
rect 40038 9840 40094 10000
rect 40406 9840 40462 10000
rect 40774 9840 40830 10000
rect 41142 9840 41198 10000
rect 41510 9840 41566 10000
rect 41878 9840 41934 10000
rect 42246 9840 42302 10000
rect 42614 9840 42670 10000
rect 42982 9840 43038 10000
rect 43350 9840 43406 10000
rect 43718 9840 43774 10000
rect 44086 9840 44142 10000
rect 44454 9840 44510 10000
rect 44822 9840 44878 10000
rect 45190 9840 45246 10000
rect 45558 9840 45614 10000
rect 45926 9840 45982 10000
rect 46294 9840 46350 10000
rect 33060 8498 33088 9840
rect 33048 8492 33100 8498
rect 33428 8480 33456 9840
rect 33600 8968 33652 8974
rect 33600 8910 33652 8916
rect 33508 8492 33560 8498
rect 33428 8452 33508 8480
rect 33048 8434 33100 8440
rect 33508 8434 33560 8440
rect 32956 8288 33008 8294
rect 32956 8230 33008 8236
rect 33324 8288 33376 8294
rect 33324 8230 33376 8236
rect 33336 7274 33364 8230
rect 33324 7268 33376 7274
rect 33324 7210 33376 7216
rect 33612 4010 33640 8910
rect 33796 8480 33824 9840
rect 33968 9036 34020 9042
rect 33968 8978 34020 8984
rect 33876 8492 33928 8498
rect 33796 8452 33876 8480
rect 33876 8434 33928 8440
rect 33692 8288 33744 8294
rect 33692 8230 33744 8236
rect 33784 8288 33836 8294
rect 33784 8230 33836 8236
rect 33704 6934 33732 8230
rect 33796 7478 33824 8230
rect 33784 7472 33836 7478
rect 33784 7414 33836 7420
rect 33692 6928 33744 6934
rect 33692 6870 33744 6876
rect 33692 4140 33744 4146
rect 33692 4082 33744 4088
rect 33600 4004 33652 4010
rect 33600 3946 33652 3952
rect 33704 3738 33732 4082
rect 33876 3936 33928 3942
rect 33876 3878 33928 3884
rect 33888 3738 33916 3878
rect 33692 3732 33744 3738
rect 33692 3674 33744 3680
rect 33876 3732 33928 3738
rect 33876 3674 33928 3680
rect 32220 3664 32272 3670
rect 32220 3606 32272 3612
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 25780 3052 25832 3058
rect 25780 2994 25832 3000
rect 29276 3052 29328 3058
rect 29276 2994 29328 3000
rect 24952 2576 25004 2582
rect 24952 2518 25004 2524
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 23940 2304 23992 2310
rect 23940 2246 23992 2252
rect 24872 2106 24900 2382
rect 23848 2100 23900 2106
rect 23848 2042 23900 2048
rect 24860 2100 24912 2106
rect 24860 2042 24912 2048
rect 24400 1964 24452 1970
rect 24400 1906 24452 1912
rect 24412 1562 24440 1906
rect 24400 1556 24452 1562
rect 24400 1498 24452 1504
rect 23756 1352 23808 1358
rect 23756 1294 23808 1300
rect 23664 672 23716 678
rect 23664 614 23716 620
rect 23492 190 23612 218
rect 23492 160 23520 190
rect 21270 54 21588 82
rect 1398 0 1454 54
rect 3606 0 3662 54
rect 5814 0 5870 54
rect 8022 0 8078 54
rect 10230 0 10286 54
rect 12438 0 12494 54
rect 14646 0 14702 54
rect 16854 0 16910 54
rect 19062 0 19118 54
rect 21270 0 21326 54
rect 23478 0 23534 160
rect 23584 82 23612 190
rect 23768 82 23796 1294
rect 25792 1222 25820 2994
rect 28895 2748 29203 2757
rect 28895 2746 28901 2748
rect 28957 2746 28981 2748
rect 29037 2746 29061 2748
rect 29117 2746 29141 2748
rect 29197 2746 29203 2748
rect 28957 2694 28959 2746
rect 29139 2694 29141 2746
rect 28895 2692 28901 2694
rect 28957 2692 28981 2694
rect 29037 2692 29061 2694
rect 29117 2692 29141 2694
rect 29197 2692 29203 2694
rect 28895 2683 29203 2692
rect 29288 2650 29316 2994
rect 29276 2644 29328 2650
rect 29276 2586 29328 2592
rect 28816 2440 28868 2446
rect 28816 2382 28868 2388
rect 31484 2440 31536 2446
rect 31484 2382 31536 2388
rect 28828 1562 28856 2382
rect 31496 2106 31524 2382
rect 31484 2100 31536 2106
rect 31484 2042 31536 2048
rect 31024 1964 31076 1970
rect 31024 1906 31076 1912
rect 28895 1660 29203 1669
rect 28895 1658 28901 1660
rect 28957 1658 28981 1660
rect 29037 1658 29061 1660
rect 29117 1658 29141 1660
rect 29197 1658 29203 1660
rect 28957 1606 28959 1658
rect 29139 1606 29141 1658
rect 28895 1604 28901 1606
rect 28957 1604 28981 1606
rect 29037 1604 29061 1606
rect 29117 1604 29141 1606
rect 29197 1604 29203 1606
rect 28895 1595 29203 1604
rect 31036 1562 31064 1906
rect 28816 1556 28868 1562
rect 28816 1498 28868 1504
rect 31024 1556 31076 1562
rect 31024 1498 31076 1504
rect 25964 1352 26016 1358
rect 25964 1294 26016 1300
rect 28172 1352 28224 1358
rect 28172 1294 28224 1300
rect 30380 1352 30432 1358
rect 30380 1294 30432 1300
rect 25780 1216 25832 1222
rect 25780 1158 25832 1164
rect 23584 54 23796 82
rect 25686 82 25742 160
rect 25976 82 26004 1294
rect 25686 54 26004 82
rect 27894 82 27950 160
rect 28184 82 28212 1294
rect 27894 54 28212 82
rect 30102 82 30158 160
rect 30392 82 30420 1294
rect 32416 1222 32444 3470
rect 33980 3466 34008 8978
rect 34164 8480 34192 9840
rect 34532 8922 34560 9840
rect 34348 8894 34560 8922
rect 34348 8498 34376 8894
rect 34484 8732 34792 8741
rect 34484 8730 34490 8732
rect 34546 8730 34570 8732
rect 34626 8730 34650 8732
rect 34706 8730 34730 8732
rect 34786 8730 34792 8732
rect 34546 8678 34548 8730
rect 34728 8678 34730 8730
rect 34484 8676 34490 8678
rect 34546 8676 34570 8678
rect 34626 8676 34650 8678
rect 34706 8676 34730 8678
rect 34786 8676 34792 8678
rect 34484 8667 34792 8676
rect 34244 8492 34296 8498
rect 34164 8452 34244 8480
rect 34244 8434 34296 8440
rect 34336 8492 34388 8498
rect 34900 8480 34928 9840
rect 35164 9376 35216 9382
rect 35164 9318 35216 9324
rect 35176 8634 35204 9318
rect 35164 8628 35216 8634
rect 35164 8570 35216 8576
rect 34980 8492 35032 8498
rect 34900 8452 34980 8480
rect 34336 8434 34388 8440
rect 35268 8480 35296 9840
rect 35532 9104 35584 9110
rect 35532 9046 35584 9052
rect 35348 8492 35400 8498
rect 35268 8452 35348 8480
rect 34980 8434 35032 8440
rect 35348 8434 35400 8440
rect 34152 8356 34204 8362
rect 34152 8298 34204 8304
rect 34164 7002 34192 8298
rect 34484 7644 34792 7653
rect 34484 7642 34490 7644
rect 34546 7642 34570 7644
rect 34626 7642 34650 7644
rect 34706 7642 34730 7644
rect 34786 7642 34792 7644
rect 34546 7590 34548 7642
rect 34728 7590 34730 7642
rect 34484 7588 34490 7590
rect 34546 7588 34570 7590
rect 34626 7588 34650 7590
rect 34706 7588 34730 7590
rect 34786 7588 34792 7590
rect 34484 7579 34792 7588
rect 34152 6996 34204 7002
rect 34152 6938 34204 6944
rect 34484 6556 34792 6565
rect 34484 6554 34490 6556
rect 34546 6554 34570 6556
rect 34626 6554 34650 6556
rect 34706 6554 34730 6556
rect 34786 6554 34792 6556
rect 34546 6502 34548 6554
rect 34728 6502 34730 6554
rect 34484 6500 34490 6502
rect 34546 6500 34570 6502
rect 34626 6500 34650 6502
rect 34706 6500 34730 6502
rect 34786 6500 34792 6502
rect 34484 6491 34792 6500
rect 34484 5468 34792 5477
rect 34484 5466 34490 5468
rect 34546 5466 34570 5468
rect 34626 5466 34650 5468
rect 34706 5466 34730 5468
rect 34786 5466 34792 5468
rect 34546 5414 34548 5466
rect 34728 5414 34730 5466
rect 34484 5412 34490 5414
rect 34546 5412 34570 5414
rect 34626 5412 34650 5414
rect 34706 5412 34730 5414
rect 34786 5412 34792 5414
rect 34484 5403 34792 5412
rect 34484 4380 34792 4389
rect 34484 4378 34490 4380
rect 34546 4378 34570 4380
rect 34626 4378 34650 4380
rect 34706 4378 34730 4380
rect 34786 4378 34792 4380
rect 34546 4326 34548 4378
rect 34728 4326 34730 4378
rect 34484 4324 34490 4326
rect 34546 4324 34570 4326
rect 34626 4324 34650 4326
rect 34706 4324 34730 4326
rect 34786 4324 34792 4326
rect 34484 4315 34792 4324
rect 35440 4140 35492 4146
rect 35440 4082 35492 4088
rect 33968 3460 34020 3466
rect 33968 3402 34020 3408
rect 34484 3292 34792 3301
rect 34484 3290 34490 3292
rect 34546 3290 34570 3292
rect 34626 3290 34650 3292
rect 34706 3290 34730 3292
rect 34786 3290 34792 3292
rect 34546 3238 34548 3290
rect 34728 3238 34730 3290
rect 34484 3236 34490 3238
rect 34546 3236 34570 3238
rect 34626 3236 34650 3238
rect 34706 3236 34730 3238
rect 34786 3236 34792 3238
rect 34484 3227 34792 3236
rect 34484 2204 34792 2213
rect 34484 2202 34490 2204
rect 34546 2202 34570 2204
rect 34626 2202 34650 2204
rect 34706 2202 34730 2204
rect 34786 2202 34792 2204
rect 34546 2150 34548 2202
rect 34728 2150 34730 2202
rect 34484 2148 34490 2150
rect 34546 2148 34570 2150
rect 34626 2148 34650 2150
rect 34706 2148 34730 2150
rect 34786 2148 34792 2150
rect 34484 2139 34792 2148
rect 35452 1358 35480 4082
rect 35544 2378 35572 9046
rect 35636 8480 35664 9840
rect 35900 9172 35952 9178
rect 35900 9114 35952 9120
rect 35912 8498 35940 9114
rect 35716 8492 35768 8498
rect 35636 8452 35716 8480
rect 35716 8434 35768 8440
rect 35900 8492 35952 8498
rect 36004 8480 36032 9840
rect 36084 8492 36136 8498
rect 36004 8452 36084 8480
rect 35900 8434 35952 8440
rect 36372 8480 36400 9840
rect 36452 8492 36504 8498
rect 36372 8452 36452 8480
rect 36084 8434 36136 8440
rect 36740 8480 36768 9840
rect 37108 8498 37136 9840
rect 37372 9172 37424 9178
rect 37372 9114 37424 9120
rect 37188 8900 37240 8906
rect 37188 8842 37240 8848
rect 37200 8634 37228 8842
rect 37188 8628 37240 8634
rect 37188 8570 37240 8576
rect 36820 8492 36872 8498
rect 36740 8452 36820 8480
rect 36452 8434 36504 8440
rect 36820 8434 36872 8440
rect 37096 8492 37148 8498
rect 37096 8434 37148 8440
rect 36636 8356 36688 8362
rect 36636 8298 36688 8304
rect 35808 8288 35860 8294
rect 35808 8230 35860 8236
rect 35820 4078 35848 8230
rect 36648 6798 36676 8298
rect 36636 6792 36688 6798
rect 36636 6734 36688 6740
rect 35900 4616 35952 4622
rect 35900 4558 35952 4564
rect 35808 4072 35860 4078
rect 35808 4014 35860 4020
rect 35912 4010 35940 4558
rect 35900 4004 35952 4010
rect 35900 3946 35952 3952
rect 37384 2514 37412 9114
rect 37476 8480 37504 9840
rect 37740 8832 37792 8838
rect 37740 8774 37792 8780
rect 37752 8634 37780 8774
rect 37740 8628 37792 8634
rect 37740 8570 37792 8576
rect 37556 8492 37608 8498
rect 37476 8452 37556 8480
rect 37844 8480 37872 9840
rect 38108 8968 38160 8974
rect 38108 8910 38160 8916
rect 38120 8634 38148 8910
rect 38108 8628 38160 8634
rect 38108 8570 38160 8576
rect 37924 8492 37976 8498
rect 37844 8452 37924 8480
rect 37556 8434 37608 8440
rect 38212 8480 38240 9840
rect 38580 8498 38608 9840
rect 38844 9580 38896 9586
rect 38844 9522 38896 9528
rect 38856 8634 38884 9522
rect 38948 8634 38976 9840
rect 39316 8634 39344 9840
rect 39684 8634 39712 9840
rect 40052 9092 40080 9840
rect 40052 9064 40172 9092
rect 40144 8634 40172 9064
rect 38844 8628 38896 8634
rect 38844 8570 38896 8576
rect 38936 8628 38988 8634
rect 38936 8570 38988 8576
rect 39304 8628 39356 8634
rect 39304 8570 39356 8576
rect 39672 8628 39724 8634
rect 39672 8570 39724 8576
rect 40132 8628 40184 8634
rect 40132 8570 40184 8576
rect 38292 8492 38344 8498
rect 38212 8452 38292 8480
rect 37924 8434 37976 8440
rect 38292 8434 38344 8440
rect 38568 8492 38620 8498
rect 38568 8434 38620 8440
rect 39396 8492 39448 8498
rect 39396 8434 39448 8440
rect 39948 8492 40000 8498
rect 39948 8434 40000 8440
rect 38384 8424 38436 8430
rect 38384 8366 38436 8372
rect 38108 8356 38160 8362
rect 38108 8298 38160 8304
rect 38120 7857 38148 8298
rect 38106 7848 38162 7857
rect 38106 7783 38162 7792
rect 38396 4826 38424 8366
rect 38476 8356 38528 8362
rect 38476 8298 38528 8304
rect 38488 7313 38516 8298
rect 38474 7304 38530 7313
rect 38474 7239 38530 7248
rect 39408 6254 39436 8434
rect 39396 6248 39448 6254
rect 39396 6190 39448 6196
rect 38384 4820 38436 4826
rect 38384 4762 38436 4768
rect 39960 4554 39988 8434
rect 40420 8362 40448 9840
rect 40684 9036 40736 9042
rect 40684 8978 40736 8984
rect 40696 8634 40724 8978
rect 40684 8628 40736 8634
rect 40684 8570 40736 8576
rect 40408 8356 40460 8362
rect 40408 8298 40460 8304
rect 40073 8188 40381 8197
rect 40073 8186 40079 8188
rect 40135 8186 40159 8188
rect 40215 8186 40239 8188
rect 40295 8186 40319 8188
rect 40375 8186 40381 8188
rect 40135 8134 40137 8186
rect 40317 8134 40319 8186
rect 40073 8132 40079 8134
rect 40135 8132 40159 8134
rect 40215 8132 40239 8134
rect 40295 8132 40319 8134
rect 40375 8132 40381 8134
rect 40073 8123 40381 8132
rect 40788 8090 40816 9840
rect 40960 9240 41012 9246
rect 40960 9182 41012 9188
rect 40972 8498 41000 9182
rect 41156 8634 41184 9840
rect 41144 8628 41196 8634
rect 41144 8570 41196 8576
rect 40960 8492 41012 8498
rect 40960 8434 41012 8440
rect 41524 8362 41552 9840
rect 41892 8634 41920 9840
rect 41880 8628 41932 8634
rect 41880 8570 41932 8576
rect 42260 8566 42288 9840
rect 42432 8832 42484 8838
rect 42432 8774 42484 8780
rect 42248 8560 42300 8566
rect 42248 8502 42300 8508
rect 42444 8498 42472 8774
rect 41880 8492 41932 8498
rect 41880 8434 41932 8440
rect 42432 8492 42484 8498
rect 42432 8434 42484 8440
rect 41512 8356 41564 8362
rect 41512 8298 41564 8304
rect 40776 8084 40828 8090
rect 40776 8026 40828 8032
rect 40960 7880 41012 7886
rect 40960 7822 41012 7828
rect 40073 7100 40381 7109
rect 40073 7098 40079 7100
rect 40135 7098 40159 7100
rect 40215 7098 40239 7100
rect 40295 7098 40319 7100
rect 40375 7098 40381 7100
rect 40135 7046 40137 7098
rect 40317 7046 40319 7098
rect 40073 7044 40079 7046
rect 40135 7044 40159 7046
rect 40215 7044 40239 7046
rect 40295 7044 40319 7046
rect 40375 7044 40381 7046
rect 40073 7035 40381 7044
rect 40073 6012 40381 6021
rect 40073 6010 40079 6012
rect 40135 6010 40159 6012
rect 40215 6010 40239 6012
rect 40295 6010 40319 6012
rect 40375 6010 40381 6012
rect 40135 5958 40137 6010
rect 40317 5958 40319 6010
rect 40073 5956 40079 5958
rect 40135 5956 40159 5958
rect 40215 5956 40239 5958
rect 40295 5956 40319 5958
rect 40375 5956 40381 5958
rect 40073 5947 40381 5956
rect 40073 4924 40381 4933
rect 40073 4922 40079 4924
rect 40135 4922 40159 4924
rect 40215 4922 40239 4924
rect 40295 4922 40319 4924
rect 40375 4922 40381 4924
rect 40135 4870 40137 4922
rect 40317 4870 40319 4922
rect 40073 4868 40079 4870
rect 40135 4868 40159 4870
rect 40215 4868 40239 4870
rect 40295 4868 40319 4870
rect 40375 4868 40381 4870
rect 40073 4859 40381 4868
rect 39948 4548 40000 4554
rect 39948 4490 40000 4496
rect 40073 3836 40381 3845
rect 40073 3834 40079 3836
rect 40135 3834 40159 3836
rect 40215 3834 40239 3836
rect 40295 3834 40319 3836
rect 40375 3834 40381 3836
rect 40135 3782 40137 3834
rect 40317 3782 40319 3834
rect 40073 3780 40079 3782
rect 40135 3780 40159 3782
rect 40215 3780 40239 3782
rect 40295 3780 40319 3782
rect 40375 3780 40381 3782
rect 40073 3771 40381 3780
rect 39028 3052 39080 3058
rect 39028 2994 39080 3000
rect 37372 2508 37424 2514
rect 37372 2450 37424 2456
rect 38200 2440 38252 2446
rect 38200 2382 38252 2388
rect 35532 2372 35584 2378
rect 35532 2314 35584 2320
rect 38212 2106 38240 2382
rect 38200 2100 38252 2106
rect 38200 2042 38252 2048
rect 37464 1964 37516 1970
rect 37464 1906 37516 1912
rect 37476 1358 37504 1906
rect 32588 1352 32640 1358
rect 32588 1294 32640 1300
rect 34888 1352 34940 1358
rect 34888 1294 34940 1300
rect 35440 1352 35492 1358
rect 35440 1294 35492 1300
rect 37004 1352 37056 1358
rect 37004 1294 37056 1300
rect 37464 1352 37516 1358
rect 37464 1294 37516 1300
rect 32404 1216 32456 1222
rect 32404 1158 32456 1164
rect 30102 54 30420 82
rect 32310 82 32366 160
rect 32600 82 32628 1294
rect 34484 1116 34792 1125
rect 34484 1114 34490 1116
rect 34546 1114 34570 1116
rect 34626 1114 34650 1116
rect 34706 1114 34730 1116
rect 34786 1114 34792 1116
rect 34546 1062 34548 1114
rect 34728 1062 34730 1114
rect 34484 1060 34490 1062
rect 34546 1060 34570 1062
rect 34626 1060 34650 1062
rect 34706 1060 34730 1062
rect 34786 1060 34792 1062
rect 34484 1051 34792 1060
rect 32310 54 32628 82
rect 34518 82 34574 160
rect 34900 82 34928 1294
rect 34518 54 34928 82
rect 36726 82 36782 160
rect 37016 82 37044 1294
rect 39040 1222 39068 2994
rect 40972 2990 41000 7822
rect 41420 7404 41472 7410
rect 41420 7346 41472 7352
rect 40960 2984 41012 2990
rect 40960 2926 41012 2932
rect 41432 2922 41460 7346
rect 41420 2916 41472 2922
rect 41420 2858 41472 2864
rect 40073 2748 40381 2757
rect 40073 2746 40079 2748
rect 40135 2746 40159 2748
rect 40215 2746 40239 2748
rect 40295 2746 40319 2748
rect 40375 2746 40381 2748
rect 40135 2694 40137 2746
rect 40317 2694 40319 2746
rect 40073 2692 40079 2694
rect 40135 2692 40159 2694
rect 40215 2692 40239 2694
rect 40295 2692 40319 2694
rect 40375 2692 40381 2694
rect 40073 2683 40381 2692
rect 41892 2582 41920 8434
rect 42628 8362 42656 9840
rect 42996 8498 43024 9840
rect 42984 8492 43036 8498
rect 42984 8434 43036 8440
rect 43076 8424 43128 8430
rect 43076 8366 43128 8372
rect 42616 8356 42668 8362
rect 42616 8298 42668 8304
rect 42800 6724 42852 6730
rect 42800 6666 42852 6672
rect 42812 3738 42840 6666
rect 43088 6186 43116 8366
rect 43364 7546 43392 9840
rect 43444 9172 43496 9178
rect 43444 9114 43496 9120
rect 43456 8498 43484 9114
rect 43732 8634 43760 9840
rect 43720 8628 43772 8634
rect 43720 8570 43772 8576
rect 43444 8492 43496 8498
rect 43444 8434 43496 8440
rect 43904 7744 43956 7750
rect 43904 7686 43956 7692
rect 43352 7540 43404 7546
rect 43352 7482 43404 7488
rect 43076 6180 43128 6186
rect 43076 6122 43128 6128
rect 43916 4826 43944 7686
rect 44100 6866 44128 9840
rect 44364 8492 44416 8498
rect 44284 8452 44364 8480
rect 44180 7812 44232 7818
rect 44180 7754 44232 7760
rect 44088 6860 44140 6866
rect 44088 6802 44140 6808
rect 43904 4820 43956 4826
rect 43904 4762 43956 4768
rect 42800 3732 42852 3738
rect 42800 3674 42852 3680
rect 44192 2650 44220 7754
rect 44180 2644 44232 2650
rect 44180 2586 44232 2592
rect 41880 2576 41932 2582
rect 41880 2518 41932 2524
rect 44284 2514 44312 8452
rect 44364 8434 44416 8440
rect 44468 8090 44496 9840
rect 44836 8634 44864 9840
rect 44824 8628 44876 8634
rect 44824 8570 44876 8576
rect 45100 8492 45152 8498
rect 45100 8434 45152 8440
rect 44456 8084 44508 8090
rect 44456 8026 44508 8032
rect 45008 7812 45060 7818
rect 45008 7754 45060 7760
rect 44364 7404 44416 7410
rect 44364 7346 44416 7352
rect 44916 7404 44968 7410
rect 44916 7346 44968 7352
rect 44376 3942 44404 7346
rect 44548 4140 44600 4146
rect 44548 4082 44600 4088
rect 44364 3936 44416 3942
rect 44364 3878 44416 3884
rect 44560 3194 44588 4082
rect 44548 3188 44600 3194
rect 44548 3130 44600 3136
rect 44928 2650 44956 7346
rect 45020 2650 45048 7754
rect 44916 2644 44968 2650
rect 44916 2586 44968 2592
rect 45008 2644 45060 2650
rect 45008 2586 45060 2592
rect 44272 2508 44324 2514
rect 44272 2450 44324 2456
rect 41788 2440 41840 2446
rect 41788 2382 41840 2388
rect 41800 2106 41828 2382
rect 43904 2372 43956 2378
rect 43904 2314 43956 2320
rect 43916 2106 43944 2314
rect 45112 2310 45140 8434
rect 45204 7410 45232 9840
rect 45572 7546 45600 9840
rect 45940 8922 45968 9840
rect 45940 8894 46060 8922
rect 45662 8732 45970 8741
rect 45662 8730 45668 8732
rect 45724 8730 45748 8732
rect 45804 8730 45828 8732
rect 45884 8730 45908 8732
rect 45964 8730 45970 8732
rect 45724 8678 45726 8730
rect 45906 8678 45908 8730
rect 45662 8676 45668 8678
rect 45724 8676 45748 8678
rect 45804 8676 45828 8678
rect 45884 8676 45908 8678
rect 45964 8676 45970 8678
rect 45662 8667 45970 8676
rect 46032 8514 46060 8894
rect 45940 8486 46060 8514
rect 45940 8022 45968 8486
rect 45928 8016 45980 8022
rect 45928 7958 45980 7964
rect 46308 7886 46336 9840
rect 46296 7880 46348 7886
rect 46296 7822 46348 7828
rect 45662 7644 45970 7653
rect 45662 7642 45668 7644
rect 45724 7642 45748 7644
rect 45804 7642 45828 7644
rect 45884 7642 45908 7644
rect 45964 7642 45970 7644
rect 45724 7590 45726 7642
rect 45906 7590 45908 7642
rect 45662 7588 45668 7590
rect 45724 7588 45748 7590
rect 45804 7588 45828 7590
rect 45884 7588 45908 7590
rect 45964 7588 45970 7590
rect 45662 7579 45970 7588
rect 45560 7540 45612 7546
rect 45560 7482 45612 7488
rect 45192 7404 45244 7410
rect 45192 7346 45244 7352
rect 45662 6556 45970 6565
rect 45662 6554 45668 6556
rect 45724 6554 45748 6556
rect 45804 6554 45828 6556
rect 45884 6554 45908 6556
rect 45964 6554 45970 6556
rect 45724 6502 45726 6554
rect 45906 6502 45908 6554
rect 45662 6500 45668 6502
rect 45724 6500 45748 6502
rect 45804 6500 45828 6502
rect 45884 6500 45908 6502
rect 45964 6500 45970 6502
rect 45662 6491 45970 6500
rect 45662 5468 45970 5477
rect 45662 5466 45668 5468
rect 45724 5466 45748 5468
rect 45804 5466 45828 5468
rect 45884 5466 45908 5468
rect 45964 5466 45970 5468
rect 45724 5414 45726 5466
rect 45906 5414 45908 5466
rect 45662 5412 45668 5414
rect 45724 5412 45748 5414
rect 45804 5412 45828 5414
rect 45884 5412 45908 5414
rect 45964 5412 45970 5414
rect 45662 5403 45970 5412
rect 45662 4380 45970 4389
rect 45662 4378 45668 4380
rect 45724 4378 45748 4380
rect 45804 4378 45828 4380
rect 45884 4378 45908 4380
rect 45964 4378 45970 4380
rect 45724 4326 45726 4378
rect 45906 4326 45908 4378
rect 45662 4324 45668 4326
rect 45724 4324 45748 4326
rect 45804 4324 45828 4326
rect 45884 4324 45908 4326
rect 45964 4324 45970 4326
rect 45662 4315 45970 4324
rect 45662 3292 45970 3301
rect 45662 3290 45668 3292
rect 45724 3290 45748 3292
rect 45804 3290 45828 3292
rect 45884 3290 45908 3292
rect 45964 3290 45970 3292
rect 45724 3238 45726 3290
rect 45906 3238 45908 3290
rect 45662 3236 45668 3238
rect 45724 3236 45748 3238
rect 45804 3236 45828 3238
rect 45884 3236 45908 3238
rect 45964 3236 45970 3238
rect 45662 3227 45970 3236
rect 45468 2440 45520 2446
rect 45468 2382 45520 2388
rect 45100 2304 45152 2310
rect 45100 2246 45152 2252
rect 45480 2106 45508 2382
rect 45662 2204 45970 2213
rect 45662 2202 45668 2204
rect 45724 2202 45748 2204
rect 45804 2202 45828 2204
rect 45884 2202 45908 2204
rect 45964 2202 45970 2204
rect 45724 2150 45726 2202
rect 45906 2150 45908 2202
rect 45662 2148 45668 2150
rect 45724 2148 45748 2150
rect 45804 2148 45828 2150
rect 45884 2148 45908 2150
rect 45964 2148 45970 2150
rect 45662 2139 45970 2148
rect 41788 2100 41840 2106
rect 41788 2042 41840 2048
rect 43904 2100 43956 2106
rect 43904 2042 43956 2048
rect 45468 2100 45520 2106
rect 45468 2042 45520 2048
rect 41972 1964 42024 1970
rect 41972 1906 42024 1912
rect 44088 1964 44140 1970
rect 44088 1906 44140 1912
rect 44824 1964 44876 1970
rect 44824 1906 44876 1912
rect 40073 1660 40381 1669
rect 40073 1658 40079 1660
rect 40135 1658 40159 1660
rect 40215 1658 40239 1660
rect 40295 1658 40319 1660
rect 40375 1658 40381 1660
rect 40135 1606 40137 1658
rect 40317 1606 40319 1658
rect 40073 1604 40079 1606
rect 40135 1604 40159 1606
rect 40215 1604 40239 1606
rect 40295 1604 40319 1606
rect 40375 1604 40381 1606
rect 40073 1595 40381 1604
rect 41984 1562 42012 1906
rect 44100 1562 44128 1906
rect 44836 1562 44864 1906
rect 41972 1556 42024 1562
rect 41972 1498 42024 1504
rect 44088 1556 44140 1562
rect 44088 1498 44140 1504
rect 44824 1556 44876 1562
rect 44824 1498 44876 1504
rect 39212 1352 39264 1358
rect 39212 1294 39264 1300
rect 41420 1352 41472 1358
rect 41420 1294 41472 1300
rect 43628 1352 43680 1358
rect 43628 1294 43680 1300
rect 45560 1352 45612 1358
rect 45560 1294 45612 1300
rect 39028 1216 39080 1222
rect 39028 1158 39080 1164
rect 36726 54 37044 82
rect 38934 82 38990 160
rect 39224 82 39252 1294
rect 38934 54 39252 82
rect 41142 82 41198 160
rect 41432 82 41460 1294
rect 41142 54 41460 82
rect 43350 82 43406 160
rect 43640 82 43668 1294
rect 45572 160 45600 1294
rect 45662 1116 45970 1125
rect 45662 1114 45668 1116
rect 45724 1114 45748 1116
rect 45804 1114 45828 1116
rect 45884 1114 45908 1116
rect 45964 1114 45970 1116
rect 45724 1062 45726 1114
rect 45906 1062 45908 1114
rect 45662 1060 45668 1062
rect 45724 1060 45748 1062
rect 45804 1060 45828 1062
rect 45884 1060 45908 1062
rect 45964 1060 45970 1062
rect 45662 1051 45970 1060
rect 43350 54 43668 82
rect 25686 0 25742 54
rect 27894 0 27950 54
rect 30102 0 30158 54
rect 32310 0 32366 54
rect 34518 0 34574 54
rect 36726 0 36782 54
rect 38934 0 38990 54
rect 41142 0 41198 54
rect 43350 0 43406 54
rect 45558 0 45614 160
<< via2 >>
rect 2686 8880 2742 8936
rect 6545 8186 6601 8188
rect 6625 8186 6681 8188
rect 6705 8186 6761 8188
rect 6785 8186 6841 8188
rect 6545 8134 6591 8186
rect 6591 8134 6601 8186
rect 6625 8134 6655 8186
rect 6655 8134 6667 8186
rect 6667 8134 6681 8186
rect 6705 8134 6719 8186
rect 6719 8134 6731 8186
rect 6731 8134 6761 8186
rect 6785 8134 6795 8186
rect 6795 8134 6841 8186
rect 6545 8132 6601 8134
rect 6625 8132 6681 8134
rect 6705 8132 6761 8134
rect 6785 8132 6841 8134
rect 2962 6840 3018 6896
rect 6545 7098 6601 7100
rect 6625 7098 6681 7100
rect 6705 7098 6761 7100
rect 6785 7098 6841 7100
rect 6545 7046 6591 7098
rect 6591 7046 6601 7098
rect 6625 7046 6655 7098
rect 6655 7046 6667 7098
rect 6667 7046 6681 7098
rect 6705 7046 6719 7098
rect 6719 7046 6731 7098
rect 6731 7046 6761 7098
rect 6785 7046 6795 7098
rect 6795 7046 6841 7098
rect 6545 7044 6601 7046
rect 6625 7044 6681 7046
rect 6705 7044 6761 7046
rect 6785 7044 6841 7046
rect 9678 9732 9680 9752
rect 9680 9732 9732 9752
rect 9732 9732 9734 9752
rect 9678 9696 9734 9732
rect 12134 8730 12190 8732
rect 12214 8730 12270 8732
rect 12294 8730 12350 8732
rect 12374 8730 12430 8732
rect 12134 8678 12180 8730
rect 12180 8678 12190 8730
rect 12214 8678 12244 8730
rect 12244 8678 12256 8730
rect 12256 8678 12270 8730
rect 12294 8678 12308 8730
rect 12308 8678 12320 8730
rect 12320 8678 12350 8730
rect 12374 8678 12384 8730
rect 12384 8678 12430 8730
rect 12134 8676 12190 8678
rect 12214 8676 12270 8678
rect 12294 8676 12350 8678
rect 12374 8676 12430 8678
rect 13726 9152 13782 9208
rect 12530 7928 12586 7984
rect 8298 6296 8354 6352
rect 7010 6160 7066 6216
rect 6545 6010 6601 6012
rect 6625 6010 6681 6012
rect 6705 6010 6761 6012
rect 6785 6010 6841 6012
rect 6545 5958 6591 6010
rect 6591 5958 6601 6010
rect 6625 5958 6655 6010
rect 6655 5958 6667 6010
rect 6667 5958 6681 6010
rect 6705 5958 6719 6010
rect 6719 5958 6731 6010
rect 6731 5958 6761 6010
rect 6785 5958 6795 6010
rect 6795 5958 6841 6010
rect 6545 5956 6601 5958
rect 6625 5956 6681 5958
rect 6705 5956 6761 5958
rect 6785 5956 6841 5958
rect 11794 7792 11850 7848
rect 9678 7268 9734 7304
rect 9678 7248 9680 7268
rect 9680 7248 9732 7268
rect 9732 7248 9734 7268
rect 12134 7642 12190 7644
rect 12214 7642 12270 7644
rect 12294 7642 12350 7644
rect 12374 7642 12430 7644
rect 12134 7590 12180 7642
rect 12180 7590 12190 7642
rect 12214 7590 12244 7642
rect 12244 7590 12256 7642
rect 12256 7590 12270 7642
rect 12294 7590 12308 7642
rect 12308 7590 12320 7642
rect 12320 7590 12350 7642
rect 12374 7590 12384 7642
rect 12384 7590 12430 7642
rect 12134 7588 12190 7590
rect 12214 7588 12270 7590
rect 12294 7588 12350 7590
rect 12374 7588 12430 7590
rect 15566 8608 15622 8664
rect 15106 8472 15162 8528
rect 15106 7520 15162 7576
rect 16578 8880 16634 8936
rect 11702 6704 11758 6760
rect 16854 8336 16910 8392
rect 17130 8744 17186 8800
rect 17723 8186 17779 8188
rect 17803 8186 17859 8188
rect 17883 8186 17939 8188
rect 17963 8186 18019 8188
rect 17723 8134 17769 8186
rect 17769 8134 17779 8186
rect 17803 8134 17833 8186
rect 17833 8134 17845 8186
rect 17845 8134 17859 8186
rect 17883 8134 17897 8186
rect 17897 8134 17909 8186
rect 17909 8134 17939 8186
rect 17963 8134 17973 8186
rect 17973 8134 18019 8186
rect 17723 8132 17779 8134
rect 17803 8132 17859 8134
rect 17883 8132 17939 8134
rect 17963 8132 18019 8134
rect 17222 7656 17278 7712
rect 18418 8064 18474 8120
rect 19338 8200 19394 8256
rect 19338 7404 19394 7440
rect 19338 7384 19340 7404
rect 19340 7384 19392 7404
rect 19392 7384 19394 7404
rect 20258 9696 20314 9752
rect 19522 7248 19578 7304
rect 17723 7098 17779 7100
rect 17803 7098 17859 7100
rect 17883 7098 17939 7100
rect 17963 7098 18019 7100
rect 17723 7046 17769 7098
rect 17769 7046 17779 7098
rect 17803 7046 17833 7098
rect 17833 7046 17845 7098
rect 17845 7046 17859 7098
rect 17883 7046 17897 7098
rect 17897 7046 17909 7098
rect 17909 7046 17939 7098
rect 17963 7046 17973 7098
rect 17973 7046 18019 7098
rect 17723 7044 17779 7046
rect 17803 7044 17859 7046
rect 17883 7044 17939 7046
rect 17963 7044 18019 7046
rect 19062 7148 19064 7168
rect 19064 7148 19116 7168
rect 19116 7148 19118 7168
rect 19062 7112 19118 7148
rect 18510 6976 18566 7032
rect 20074 7520 20130 7576
rect 20350 7792 20406 7848
rect 20810 9172 20866 9208
rect 20810 9152 20812 9172
rect 20812 9152 20864 9172
rect 20864 9152 20866 9172
rect 21362 9696 21418 9752
rect 21546 9288 21602 9344
rect 21178 8336 21234 8392
rect 21730 9832 21786 9888
rect 21730 9596 21732 9616
rect 21732 9596 21784 9616
rect 21784 9596 21786 9616
rect 21730 9560 21786 9596
rect 21730 9460 21732 9480
rect 21732 9460 21784 9480
rect 21784 9460 21786 9480
rect 21730 9424 21786 9460
rect 22098 9424 22154 9480
rect 21546 7792 21602 7848
rect 22006 7828 22008 7848
rect 22008 7828 22060 7848
rect 22060 7828 22062 7848
rect 22006 7792 22062 7828
rect 12134 6554 12190 6556
rect 12214 6554 12270 6556
rect 12294 6554 12350 6556
rect 12374 6554 12430 6556
rect 12134 6502 12180 6554
rect 12180 6502 12190 6554
rect 12214 6502 12244 6554
rect 12244 6502 12256 6554
rect 12256 6502 12270 6554
rect 12294 6502 12308 6554
rect 12308 6502 12320 6554
rect 12320 6502 12350 6554
rect 12374 6502 12384 6554
rect 12384 6502 12430 6554
rect 12134 6500 12190 6502
rect 12214 6500 12270 6502
rect 12294 6500 12350 6502
rect 12374 6500 12430 6502
rect 17723 6010 17779 6012
rect 17803 6010 17859 6012
rect 17883 6010 17939 6012
rect 17963 6010 18019 6012
rect 17723 5958 17769 6010
rect 17769 5958 17779 6010
rect 17803 5958 17833 6010
rect 17833 5958 17845 6010
rect 17845 5958 17859 6010
rect 17883 5958 17897 6010
rect 17897 5958 17909 6010
rect 17909 5958 17939 6010
rect 17963 5958 17973 6010
rect 17973 5958 18019 6010
rect 17723 5956 17779 5958
rect 17803 5956 17859 5958
rect 17883 5956 17939 5958
rect 17963 5956 18019 5958
rect 22006 7692 22008 7712
rect 22008 7692 22060 7712
rect 22060 7692 22062 7712
rect 22006 7656 22062 7692
rect 21914 7248 21970 7304
rect 22466 8628 22522 8664
rect 22466 8608 22468 8628
rect 22468 8608 22520 8628
rect 22520 8608 22522 8628
rect 22834 8880 22890 8936
rect 22834 8744 22890 8800
rect 22558 8200 22614 8256
rect 23312 8730 23368 8732
rect 23392 8730 23448 8732
rect 23472 8730 23528 8732
rect 23552 8730 23608 8732
rect 23312 8678 23358 8730
rect 23358 8678 23368 8730
rect 23392 8678 23422 8730
rect 23422 8678 23434 8730
rect 23434 8678 23448 8730
rect 23472 8678 23486 8730
rect 23486 8678 23498 8730
rect 23498 8678 23528 8730
rect 23552 8678 23562 8730
rect 23562 8678 23608 8730
rect 23312 8676 23368 8678
rect 23392 8676 23448 8678
rect 23472 8676 23528 8678
rect 23552 8676 23608 8678
rect 23478 8492 23534 8528
rect 23478 8472 23480 8492
rect 23480 8472 23532 8492
rect 23532 8472 23534 8492
rect 23754 9288 23810 9344
rect 23846 8472 23902 8528
rect 23312 7642 23368 7644
rect 23392 7642 23448 7644
rect 23472 7642 23528 7644
rect 23552 7642 23608 7644
rect 23312 7590 23358 7642
rect 23358 7590 23368 7642
rect 23392 7590 23422 7642
rect 23422 7590 23434 7642
rect 23434 7590 23448 7642
rect 23472 7590 23486 7642
rect 23486 7590 23498 7642
rect 23498 7590 23528 7642
rect 23552 7590 23562 7642
rect 23562 7590 23608 7642
rect 23312 7588 23368 7590
rect 23392 7588 23448 7590
rect 23472 7588 23528 7590
rect 23552 7588 23608 7590
rect 23478 7268 23534 7304
rect 23478 7248 23480 7268
rect 23480 7248 23532 7268
rect 23532 7248 23534 7268
rect 24214 8084 24270 8120
rect 24214 8064 24216 8084
rect 24216 8064 24268 8084
rect 24268 8064 24270 8084
rect 23754 7248 23810 7304
rect 25594 9016 25650 9072
rect 25502 7964 25504 7984
rect 25504 7964 25556 7984
rect 25556 7964 25558 7984
rect 25502 7928 25558 7964
rect 26238 9152 26294 9208
rect 26698 9832 26754 9888
rect 27066 9696 27122 9752
rect 27434 8336 27490 8392
rect 24766 7792 24822 7848
rect 23202 7148 23204 7168
rect 23204 7148 23256 7168
rect 23256 7148 23258 7168
rect 23202 7112 23258 7148
rect 23570 7112 23626 7168
rect 24766 7112 24822 7168
rect 23846 6976 23902 7032
rect 23312 6554 23368 6556
rect 23392 6554 23448 6556
rect 23472 6554 23528 6556
rect 23552 6554 23608 6556
rect 23312 6502 23358 6554
rect 23358 6502 23368 6554
rect 23392 6502 23422 6554
rect 23422 6502 23434 6554
rect 23434 6502 23448 6554
rect 23472 6502 23486 6554
rect 23486 6502 23498 6554
rect 23498 6502 23528 6554
rect 23552 6502 23562 6554
rect 23562 6502 23608 6554
rect 23312 6500 23368 6502
rect 23392 6500 23448 6502
rect 23472 6500 23528 6502
rect 23552 6500 23608 6502
rect 25594 6840 25650 6896
rect 28170 9560 28226 9616
rect 28901 8186 28957 8188
rect 28981 8186 29037 8188
rect 29061 8186 29117 8188
rect 29141 8186 29197 8188
rect 28901 8134 28947 8186
rect 28947 8134 28957 8186
rect 28981 8134 29011 8186
rect 29011 8134 29023 8186
rect 29023 8134 29037 8186
rect 29061 8134 29075 8186
rect 29075 8134 29087 8186
rect 29087 8134 29117 8186
rect 29141 8134 29151 8186
rect 29151 8134 29197 8186
rect 28901 8132 28957 8134
rect 28981 8132 29037 8134
rect 29061 8132 29117 8134
rect 29141 8132 29197 8134
rect 31666 7656 31722 7712
rect 31942 7384 31998 7440
rect 28901 7098 28957 7100
rect 28981 7098 29037 7100
rect 29061 7098 29117 7100
rect 29141 7098 29197 7100
rect 28901 7046 28947 7098
rect 28947 7046 28957 7098
rect 28981 7046 29011 7098
rect 29011 7046 29023 7098
rect 29023 7046 29037 7098
rect 29061 7046 29075 7098
rect 29075 7046 29087 7098
rect 29087 7046 29117 7098
rect 29141 7046 29151 7098
rect 29151 7046 29197 7098
rect 28901 7044 28957 7046
rect 28981 7044 29037 7046
rect 29061 7044 29117 7046
rect 29141 7044 29197 7046
rect 28538 6704 28594 6760
rect 26422 6296 26478 6352
rect 8942 5752 8998 5808
rect 21730 5752 21786 5808
rect 12134 5466 12190 5468
rect 12214 5466 12270 5468
rect 12294 5466 12350 5468
rect 12374 5466 12430 5468
rect 12134 5414 12180 5466
rect 12180 5414 12190 5466
rect 12214 5414 12244 5466
rect 12244 5414 12256 5466
rect 12256 5414 12270 5466
rect 12294 5414 12308 5466
rect 12308 5414 12320 5466
rect 12320 5414 12350 5466
rect 12374 5414 12384 5466
rect 12384 5414 12430 5466
rect 12134 5412 12190 5414
rect 12214 5412 12270 5414
rect 12294 5412 12350 5414
rect 12374 5412 12430 5414
rect 23312 5466 23368 5468
rect 23392 5466 23448 5468
rect 23472 5466 23528 5468
rect 23552 5466 23608 5468
rect 23312 5414 23358 5466
rect 23358 5414 23368 5466
rect 23392 5414 23422 5466
rect 23422 5414 23434 5466
rect 23434 5414 23448 5466
rect 23472 5414 23486 5466
rect 23486 5414 23498 5466
rect 23498 5414 23528 5466
rect 23552 5414 23562 5466
rect 23562 5414 23608 5466
rect 23312 5412 23368 5414
rect 23392 5412 23448 5414
rect 23472 5412 23528 5414
rect 23552 5412 23608 5414
rect 6545 4922 6601 4924
rect 6625 4922 6681 4924
rect 6705 4922 6761 4924
rect 6785 4922 6841 4924
rect 6545 4870 6591 4922
rect 6591 4870 6601 4922
rect 6625 4870 6655 4922
rect 6655 4870 6667 4922
rect 6667 4870 6681 4922
rect 6705 4870 6719 4922
rect 6719 4870 6731 4922
rect 6731 4870 6761 4922
rect 6785 4870 6795 4922
rect 6795 4870 6841 4922
rect 6545 4868 6601 4870
rect 6625 4868 6681 4870
rect 6705 4868 6761 4870
rect 6785 4868 6841 4870
rect 17723 4922 17779 4924
rect 17803 4922 17859 4924
rect 17883 4922 17939 4924
rect 17963 4922 18019 4924
rect 17723 4870 17769 4922
rect 17769 4870 17779 4922
rect 17803 4870 17833 4922
rect 17833 4870 17845 4922
rect 17845 4870 17859 4922
rect 17883 4870 17897 4922
rect 17897 4870 17909 4922
rect 17909 4870 17939 4922
rect 17963 4870 17973 4922
rect 17973 4870 18019 4922
rect 17723 4868 17779 4870
rect 17803 4868 17859 4870
rect 17883 4868 17939 4870
rect 17963 4868 18019 4870
rect 12134 4378 12190 4380
rect 12214 4378 12270 4380
rect 12294 4378 12350 4380
rect 12374 4378 12430 4380
rect 12134 4326 12180 4378
rect 12180 4326 12190 4378
rect 12214 4326 12244 4378
rect 12244 4326 12256 4378
rect 12256 4326 12270 4378
rect 12294 4326 12308 4378
rect 12308 4326 12320 4378
rect 12320 4326 12350 4378
rect 12374 4326 12384 4378
rect 12384 4326 12430 4378
rect 12134 4324 12190 4326
rect 12214 4324 12270 4326
rect 12294 4324 12350 4326
rect 12374 4324 12430 4326
rect 6545 3834 6601 3836
rect 6625 3834 6681 3836
rect 6705 3834 6761 3836
rect 6785 3834 6841 3836
rect 6545 3782 6591 3834
rect 6591 3782 6601 3834
rect 6625 3782 6655 3834
rect 6655 3782 6667 3834
rect 6667 3782 6681 3834
rect 6705 3782 6719 3834
rect 6719 3782 6731 3834
rect 6731 3782 6761 3834
rect 6785 3782 6795 3834
rect 6795 3782 6841 3834
rect 6545 3780 6601 3782
rect 6625 3780 6681 3782
rect 6705 3780 6761 3782
rect 6785 3780 6841 3782
rect 17723 3834 17779 3836
rect 17803 3834 17859 3836
rect 17883 3834 17939 3836
rect 17963 3834 18019 3836
rect 17723 3782 17769 3834
rect 17769 3782 17779 3834
rect 17803 3782 17833 3834
rect 17833 3782 17845 3834
rect 17845 3782 17859 3834
rect 17883 3782 17897 3834
rect 17897 3782 17909 3834
rect 17909 3782 17939 3834
rect 17963 3782 17973 3834
rect 17973 3782 18019 3834
rect 17723 3780 17779 3782
rect 17803 3780 17859 3782
rect 17883 3780 17939 3782
rect 17963 3780 18019 3782
rect 12134 3290 12190 3292
rect 12214 3290 12270 3292
rect 12294 3290 12350 3292
rect 12374 3290 12430 3292
rect 12134 3238 12180 3290
rect 12180 3238 12190 3290
rect 12214 3238 12244 3290
rect 12244 3238 12256 3290
rect 12256 3238 12270 3290
rect 12294 3238 12308 3290
rect 12308 3238 12320 3290
rect 12320 3238 12350 3290
rect 12374 3238 12384 3290
rect 12384 3238 12430 3290
rect 12134 3236 12190 3238
rect 12214 3236 12270 3238
rect 12294 3236 12350 3238
rect 12374 3236 12430 3238
rect 6545 2746 6601 2748
rect 6625 2746 6681 2748
rect 6705 2746 6761 2748
rect 6785 2746 6841 2748
rect 6545 2694 6591 2746
rect 6591 2694 6601 2746
rect 6625 2694 6655 2746
rect 6655 2694 6667 2746
rect 6667 2694 6681 2746
rect 6705 2694 6719 2746
rect 6719 2694 6731 2746
rect 6731 2694 6761 2746
rect 6785 2694 6795 2746
rect 6795 2694 6841 2746
rect 6545 2692 6601 2694
rect 6625 2692 6681 2694
rect 6705 2692 6761 2694
rect 6785 2692 6841 2694
rect 17723 2746 17779 2748
rect 17803 2746 17859 2748
rect 17883 2746 17939 2748
rect 17963 2746 18019 2748
rect 17723 2694 17769 2746
rect 17769 2694 17779 2746
rect 17803 2694 17833 2746
rect 17833 2694 17845 2746
rect 17845 2694 17859 2746
rect 17883 2694 17897 2746
rect 17897 2694 17909 2746
rect 17909 2694 17939 2746
rect 17963 2694 17973 2746
rect 17973 2694 18019 2746
rect 17723 2692 17779 2694
rect 17803 2692 17859 2694
rect 17883 2692 17939 2694
rect 17963 2692 18019 2694
rect 12134 2202 12190 2204
rect 12214 2202 12270 2204
rect 12294 2202 12350 2204
rect 12374 2202 12430 2204
rect 12134 2150 12180 2202
rect 12180 2150 12190 2202
rect 12214 2150 12244 2202
rect 12244 2150 12256 2202
rect 12256 2150 12270 2202
rect 12294 2150 12308 2202
rect 12308 2150 12320 2202
rect 12320 2150 12350 2202
rect 12374 2150 12384 2202
rect 12384 2150 12430 2202
rect 12134 2148 12190 2150
rect 12214 2148 12270 2150
rect 12294 2148 12350 2150
rect 12374 2148 12430 2150
rect 6545 1658 6601 1660
rect 6625 1658 6681 1660
rect 6705 1658 6761 1660
rect 6785 1658 6841 1660
rect 6545 1606 6591 1658
rect 6591 1606 6601 1658
rect 6625 1606 6655 1658
rect 6655 1606 6667 1658
rect 6667 1606 6681 1658
rect 6705 1606 6719 1658
rect 6719 1606 6731 1658
rect 6731 1606 6761 1658
rect 6785 1606 6795 1658
rect 6795 1606 6841 1658
rect 6545 1604 6601 1606
rect 6625 1604 6681 1606
rect 6705 1604 6761 1606
rect 6785 1604 6841 1606
rect 17723 1658 17779 1660
rect 17803 1658 17859 1660
rect 17883 1658 17939 1660
rect 17963 1658 18019 1660
rect 17723 1606 17769 1658
rect 17769 1606 17779 1658
rect 17803 1606 17833 1658
rect 17833 1606 17845 1658
rect 17845 1606 17859 1658
rect 17883 1606 17897 1658
rect 17897 1606 17909 1658
rect 17909 1606 17939 1658
rect 17963 1606 17973 1658
rect 17973 1606 18019 1658
rect 17723 1604 17779 1606
rect 17803 1604 17859 1606
rect 17883 1604 17939 1606
rect 17963 1604 18019 1606
rect 12134 1114 12190 1116
rect 12214 1114 12270 1116
rect 12294 1114 12350 1116
rect 12374 1114 12430 1116
rect 12134 1062 12180 1114
rect 12180 1062 12190 1114
rect 12214 1062 12244 1114
rect 12244 1062 12256 1114
rect 12256 1062 12270 1114
rect 12294 1062 12308 1114
rect 12308 1062 12320 1114
rect 12320 1062 12350 1114
rect 12374 1062 12384 1114
rect 12384 1062 12430 1114
rect 12134 1060 12190 1062
rect 12214 1060 12270 1062
rect 12294 1060 12350 1062
rect 12374 1060 12430 1062
rect 23312 4378 23368 4380
rect 23392 4378 23448 4380
rect 23472 4378 23528 4380
rect 23552 4378 23608 4380
rect 23312 4326 23358 4378
rect 23358 4326 23368 4378
rect 23392 4326 23422 4378
rect 23422 4326 23434 4378
rect 23434 4326 23448 4378
rect 23472 4326 23486 4378
rect 23486 4326 23498 4378
rect 23498 4326 23528 4378
rect 23552 4326 23562 4378
rect 23562 4326 23608 4378
rect 23312 4324 23368 4326
rect 23392 4324 23448 4326
rect 23472 4324 23528 4326
rect 23552 4324 23608 4326
rect 23312 3290 23368 3292
rect 23392 3290 23448 3292
rect 23472 3290 23528 3292
rect 23552 3290 23608 3292
rect 23312 3238 23358 3290
rect 23358 3238 23368 3290
rect 23392 3238 23422 3290
rect 23422 3238 23434 3290
rect 23434 3238 23448 3290
rect 23472 3238 23486 3290
rect 23486 3238 23498 3290
rect 23498 3238 23528 3290
rect 23552 3238 23562 3290
rect 23562 3238 23608 3290
rect 23312 3236 23368 3238
rect 23392 3236 23448 3238
rect 23472 3236 23528 3238
rect 23552 3236 23608 3238
rect 23312 2202 23368 2204
rect 23392 2202 23448 2204
rect 23472 2202 23528 2204
rect 23552 2202 23608 2204
rect 23312 2150 23358 2202
rect 23358 2150 23368 2202
rect 23392 2150 23422 2202
rect 23422 2150 23434 2202
rect 23434 2150 23448 2202
rect 23472 2150 23486 2202
rect 23486 2150 23498 2202
rect 23498 2150 23528 2202
rect 23552 2150 23562 2202
rect 23562 2150 23608 2202
rect 23312 2148 23368 2150
rect 23392 2148 23448 2150
rect 23472 2148 23528 2150
rect 23552 2148 23608 2150
rect 23312 1114 23368 1116
rect 23392 1114 23448 1116
rect 23472 1114 23528 1116
rect 23552 1114 23608 1116
rect 23312 1062 23358 1114
rect 23358 1062 23368 1114
rect 23392 1062 23422 1114
rect 23422 1062 23434 1114
rect 23434 1062 23448 1114
rect 23472 1062 23486 1114
rect 23486 1062 23498 1114
rect 23498 1062 23528 1114
rect 23552 1062 23562 1114
rect 23562 1062 23608 1114
rect 23312 1060 23368 1062
rect 23392 1060 23448 1062
rect 23472 1060 23528 1062
rect 23552 1060 23608 1062
rect 25042 6160 25098 6216
rect 28901 6010 28957 6012
rect 28981 6010 29037 6012
rect 29061 6010 29117 6012
rect 29141 6010 29197 6012
rect 28901 5958 28947 6010
rect 28947 5958 28957 6010
rect 28981 5958 29011 6010
rect 29011 5958 29023 6010
rect 29023 5958 29037 6010
rect 29061 5958 29075 6010
rect 29075 5958 29087 6010
rect 29087 5958 29117 6010
rect 29141 5958 29151 6010
rect 29151 5958 29197 6010
rect 28901 5956 28957 5958
rect 28981 5956 29037 5958
rect 29061 5956 29117 5958
rect 29141 5956 29197 5958
rect 28901 4922 28957 4924
rect 28981 4922 29037 4924
rect 29061 4922 29117 4924
rect 29141 4922 29197 4924
rect 28901 4870 28947 4922
rect 28947 4870 28957 4922
rect 28981 4870 29011 4922
rect 29011 4870 29023 4922
rect 29023 4870 29037 4922
rect 29061 4870 29075 4922
rect 29075 4870 29087 4922
rect 29087 4870 29117 4922
rect 29141 4870 29151 4922
rect 29151 4870 29197 4922
rect 28901 4868 28957 4870
rect 28981 4868 29037 4870
rect 29061 4868 29117 4870
rect 29141 4868 29197 4870
rect 28901 3834 28957 3836
rect 28981 3834 29037 3836
rect 29061 3834 29117 3836
rect 29141 3834 29197 3836
rect 28901 3782 28947 3834
rect 28947 3782 28957 3834
rect 28981 3782 29011 3834
rect 29011 3782 29023 3834
rect 29023 3782 29037 3834
rect 29061 3782 29075 3834
rect 29075 3782 29087 3834
rect 29087 3782 29117 3834
rect 29141 3782 29151 3834
rect 29151 3782 29197 3834
rect 28901 3780 28957 3782
rect 28981 3780 29037 3782
rect 29061 3780 29117 3782
rect 29141 3780 29197 3782
rect 28901 2746 28957 2748
rect 28981 2746 29037 2748
rect 29061 2746 29117 2748
rect 29141 2746 29197 2748
rect 28901 2694 28947 2746
rect 28947 2694 28957 2746
rect 28981 2694 29011 2746
rect 29011 2694 29023 2746
rect 29023 2694 29037 2746
rect 29061 2694 29075 2746
rect 29075 2694 29087 2746
rect 29087 2694 29117 2746
rect 29141 2694 29151 2746
rect 29151 2694 29197 2746
rect 28901 2692 28957 2694
rect 28981 2692 29037 2694
rect 29061 2692 29117 2694
rect 29141 2692 29197 2694
rect 28901 1658 28957 1660
rect 28981 1658 29037 1660
rect 29061 1658 29117 1660
rect 29141 1658 29197 1660
rect 28901 1606 28947 1658
rect 28947 1606 28957 1658
rect 28981 1606 29011 1658
rect 29011 1606 29023 1658
rect 29023 1606 29037 1658
rect 29061 1606 29075 1658
rect 29075 1606 29087 1658
rect 29087 1606 29117 1658
rect 29141 1606 29151 1658
rect 29151 1606 29197 1658
rect 28901 1604 28957 1606
rect 28981 1604 29037 1606
rect 29061 1604 29117 1606
rect 29141 1604 29197 1606
rect 34490 8730 34546 8732
rect 34570 8730 34626 8732
rect 34650 8730 34706 8732
rect 34730 8730 34786 8732
rect 34490 8678 34536 8730
rect 34536 8678 34546 8730
rect 34570 8678 34600 8730
rect 34600 8678 34612 8730
rect 34612 8678 34626 8730
rect 34650 8678 34664 8730
rect 34664 8678 34676 8730
rect 34676 8678 34706 8730
rect 34730 8678 34740 8730
rect 34740 8678 34786 8730
rect 34490 8676 34546 8678
rect 34570 8676 34626 8678
rect 34650 8676 34706 8678
rect 34730 8676 34786 8678
rect 34490 7642 34546 7644
rect 34570 7642 34626 7644
rect 34650 7642 34706 7644
rect 34730 7642 34786 7644
rect 34490 7590 34536 7642
rect 34536 7590 34546 7642
rect 34570 7590 34600 7642
rect 34600 7590 34612 7642
rect 34612 7590 34626 7642
rect 34650 7590 34664 7642
rect 34664 7590 34676 7642
rect 34676 7590 34706 7642
rect 34730 7590 34740 7642
rect 34740 7590 34786 7642
rect 34490 7588 34546 7590
rect 34570 7588 34626 7590
rect 34650 7588 34706 7590
rect 34730 7588 34786 7590
rect 34490 6554 34546 6556
rect 34570 6554 34626 6556
rect 34650 6554 34706 6556
rect 34730 6554 34786 6556
rect 34490 6502 34536 6554
rect 34536 6502 34546 6554
rect 34570 6502 34600 6554
rect 34600 6502 34612 6554
rect 34612 6502 34626 6554
rect 34650 6502 34664 6554
rect 34664 6502 34676 6554
rect 34676 6502 34706 6554
rect 34730 6502 34740 6554
rect 34740 6502 34786 6554
rect 34490 6500 34546 6502
rect 34570 6500 34626 6502
rect 34650 6500 34706 6502
rect 34730 6500 34786 6502
rect 34490 5466 34546 5468
rect 34570 5466 34626 5468
rect 34650 5466 34706 5468
rect 34730 5466 34786 5468
rect 34490 5414 34536 5466
rect 34536 5414 34546 5466
rect 34570 5414 34600 5466
rect 34600 5414 34612 5466
rect 34612 5414 34626 5466
rect 34650 5414 34664 5466
rect 34664 5414 34676 5466
rect 34676 5414 34706 5466
rect 34730 5414 34740 5466
rect 34740 5414 34786 5466
rect 34490 5412 34546 5414
rect 34570 5412 34626 5414
rect 34650 5412 34706 5414
rect 34730 5412 34786 5414
rect 34490 4378 34546 4380
rect 34570 4378 34626 4380
rect 34650 4378 34706 4380
rect 34730 4378 34786 4380
rect 34490 4326 34536 4378
rect 34536 4326 34546 4378
rect 34570 4326 34600 4378
rect 34600 4326 34612 4378
rect 34612 4326 34626 4378
rect 34650 4326 34664 4378
rect 34664 4326 34676 4378
rect 34676 4326 34706 4378
rect 34730 4326 34740 4378
rect 34740 4326 34786 4378
rect 34490 4324 34546 4326
rect 34570 4324 34626 4326
rect 34650 4324 34706 4326
rect 34730 4324 34786 4326
rect 34490 3290 34546 3292
rect 34570 3290 34626 3292
rect 34650 3290 34706 3292
rect 34730 3290 34786 3292
rect 34490 3238 34536 3290
rect 34536 3238 34546 3290
rect 34570 3238 34600 3290
rect 34600 3238 34612 3290
rect 34612 3238 34626 3290
rect 34650 3238 34664 3290
rect 34664 3238 34676 3290
rect 34676 3238 34706 3290
rect 34730 3238 34740 3290
rect 34740 3238 34786 3290
rect 34490 3236 34546 3238
rect 34570 3236 34626 3238
rect 34650 3236 34706 3238
rect 34730 3236 34786 3238
rect 34490 2202 34546 2204
rect 34570 2202 34626 2204
rect 34650 2202 34706 2204
rect 34730 2202 34786 2204
rect 34490 2150 34536 2202
rect 34536 2150 34546 2202
rect 34570 2150 34600 2202
rect 34600 2150 34612 2202
rect 34612 2150 34626 2202
rect 34650 2150 34664 2202
rect 34664 2150 34676 2202
rect 34676 2150 34706 2202
rect 34730 2150 34740 2202
rect 34740 2150 34786 2202
rect 34490 2148 34546 2150
rect 34570 2148 34626 2150
rect 34650 2148 34706 2150
rect 34730 2148 34786 2150
rect 38106 7792 38162 7848
rect 38474 7248 38530 7304
rect 40079 8186 40135 8188
rect 40159 8186 40215 8188
rect 40239 8186 40295 8188
rect 40319 8186 40375 8188
rect 40079 8134 40125 8186
rect 40125 8134 40135 8186
rect 40159 8134 40189 8186
rect 40189 8134 40201 8186
rect 40201 8134 40215 8186
rect 40239 8134 40253 8186
rect 40253 8134 40265 8186
rect 40265 8134 40295 8186
rect 40319 8134 40329 8186
rect 40329 8134 40375 8186
rect 40079 8132 40135 8134
rect 40159 8132 40215 8134
rect 40239 8132 40295 8134
rect 40319 8132 40375 8134
rect 40079 7098 40135 7100
rect 40159 7098 40215 7100
rect 40239 7098 40295 7100
rect 40319 7098 40375 7100
rect 40079 7046 40125 7098
rect 40125 7046 40135 7098
rect 40159 7046 40189 7098
rect 40189 7046 40201 7098
rect 40201 7046 40215 7098
rect 40239 7046 40253 7098
rect 40253 7046 40265 7098
rect 40265 7046 40295 7098
rect 40319 7046 40329 7098
rect 40329 7046 40375 7098
rect 40079 7044 40135 7046
rect 40159 7044 40215 7046
rect 40239 7044 40295 7046
rect 40319 7044 40375 7046
rect 40079 6010 40135 6012
rect 40159 6010 40215 6012
rect 40239 6010 40295 6012
rect 40319 6010 40375 6012
rect 40079 5958 40125 6010
rect 40125 5958 40135 6010
rect 40159 5958 40189 6010
rect 40189 5958 40201 6010
rect 40201 5958 40215 6010
rect 40239 5958 40253 6010
rect 40253 5958 40265 6010
rect 40265 5958 40295 6010
rect 40319 5958 40329 6010
rect 40329 5958 40375 6010
rect 40079 5956 40135 5958
rect 40159 5956 40215 5958
rect 40239 5956 40295 5958
rect 40319 5956 40375 5958
rect 40079 4922 40135 4924
rect 40159 4922 40215 4924
rect 40239 4922 40295 4924
rect 40319 4922 40375 4924
rect 40079 4870 40125 4922
rect 40125 4870 40135 4922
rect 40159 4870 40189 4922
rect 40189 4870 40201 4922
rect 40201 4870 40215 4922
rect 40239 4870 40253 4922
rect 40253 4870 40265 4922
rect 40265 4870 40295 4922
rect 40319 4870 40329 4922
rect 40329 4870 40375 4922
rect 40079 4868 40135 4870
rect 40159 4868 40215 4870
rect 40239 4868 40295 4870
rect 40319 4868 40375 4870
rect 40079 3834 40135 3836
rect 40159 3834 40215 3836
rect 40239 3834 40295 3836
rect 40319 3834 40375 3836
rect 40079 3782 40125 3834
rect 40125 3782 40135 3834
rect 40159 3782 40189 3834
rect 40189 3782 40201 3834
rect 40201 3782 40215 3834
rect 40239 3782 40253 3834
rect 40253 3782 40265 3834
rect 40265 3782 40295 3834
rect 40319 3782 40329 3834
rect 40329 3782 40375 3834
rect 40079 3780 40135 3782
rect 40159 3780 40215 3782
rect 40239 3780 40295 3782
rect 40319 3780 40375 3782
rect 34490 1114 34546 1116
rect 34570 1114 34626 1116
rect 34650 1114 34706 1116
rect 34730 1114 34786 1116
rect 34490 1062 34536 1114
rect 34536 1062 34546 1114
rect 34570 1062 34600 1114
rect 34600 1062 34612 1114
rect 34612 1062 34626 1114
rect 34650 1062 34664 1114
rect 34664 1062 34676 1114
rect 34676 1062 34706 1114
rect 34730 1062 34740 1114
rect 34740 1062 34786 1114
rect 34490 1060 34546 1062
rect 34570 1060 34626 1062
rect 34650 1060 34706 1062
rect 34730 1060 34786 1062
rect 40079 2746 40135 2748
rect 40159 2746 40215 2748
rect 40239 2746 40295 2748
rect 40319 2746 40375 2748
rect 40079 2694 40125 2746
rect 40125 2694 40135 2746
rect 40159 2694 40189 2746
rect 40189 2694 40201 2746
rect 40201 2694 40215 2746
rect 40239 2694 40253 2746
rect 40253 2694 40265 2746
rect 40265 2694 40295 2746
rect 40319 2694 40329 2746
rect 40329 2694 40375 2746
rect 40079 2692 40135 2694
rect 40159 2692 40215 2694
rect 40239 2692 40295 2694
rect 40319 2692 40375 2694
rect 45668 8730 45724 8732
rect 45748 8730 45804 8732
rect 45828 8730 45884 8732
rect 45908 8730 45964 8732
rect 45668 8678 45714 8730
rect 45714 8678 45724 8730
rect 45748 8678 45778 8730
rect 45778 8678 45790 8730
rect 45790 8678 45804 8730
rect 45828 8678 45842 8730
rect 45842 8678 45854 8730
rect 45854 8678 45884 8730
rect 45908 8678 45918 8730
rect 45918 8678 45964 8730
rect 45668 8676 45724 8678
rect 45748 8676 45804 8678
rect 45828 8676 45884 8678
rect 45908 8676 45964 8678
rect 45668 7642 45724 7644
rect 45748 7642 45804 7644
rect 45828 7642 45884 7644
rect 45908 7642 45964 7644
rect 45668 7590 45714 7642
rect 45714 7590 45724 7642
rect 45748 7590 45778 7642
rect 45778 7590 45790 7642
rect 45790 7590 45804 7642
rect 45828 7590 45842 7642
rect 45842 7590 45854 7642
rect 45854 7590 45884 7642
rect 45908 7590 45918 7642
rect 45918 7590 45964 7642
rect 45668 7588 45724 7590
rect 45748 7588 45804 7590
rect 45828 7588 45884 7590
rect 45908 7588 45964 7590
rect 45668 6554 45724 6556
rect 45748 6554 45804 6556
rect 45828 6554 45884 6556
rect 45908 6554 45964 6556
rect 45668 6502 45714 6554
rect 45714 6502 45724 6554
rect 45748 6502 45778 6554
rect 45778 6502 45790 6554
rect 45790 6502 45804 6554
rect 45828 6502 45842 6554
rect 45842 6502 45854 6554
rect 45854 6502 45884 6554
rect 45908 6502 45918 6554
rect 45918 6502 45964 6554
rect 45668 6500 45724 6502
rect 45748 6500 45804 6502
rect 45828 6500 45884 6502
rect 45908 6500 45964 6502
rect 45668 5466 45724 5468
rect 45748 5466 45804 5468
rect 45828 5466 45884 5468
rect 45908 5466 45964 5468
rect 45668 5414 45714 5466
rect 45714 5414 45724 5466
rect 45748 5414 45778 5466
rect 45778 5414 45790 5466
rect 45790 5414 45804 5466
rect 45828 5414 45842 5466
rect 45842 5414 45854 5466
rect 45854 5414 45884 5466
rect 45908 5414 45918 5466
rect 45918 5414 45964 5466
rect 45668 5412 45724 5414
rect 45748 5412 45804 5414
rect 45828 5412 45884 5414
rect 45908 5412 45964 5414
rect 45668 4378 45724 4380
rect 45748 4378 45804 4380
rect 45828 4378 45884 4380
rect 45908 4378 45964 4380
rect 45668 4326 45714 4378
rect 45714 4326 45724 4378
rect 45748 4326 45778 4378
rect 45778 4326 45790 4378
rect 45790 4326 45804 4378
rect 45828 4326 45842 4378
rect 45842 4326 45854 4378
rect 45854 4326 45884 4378
rect 45908 4326 45918 4378
rect 45918 4326 45964 4378
rect 45668 4324 45724 4326
rect 45748 4324 45804 4326
rect 45828 4324 45884 4326
rect 45908 4324 45964 4326
rect 45668 3290 45724 3292
rect 45748 3290 45804 3292
rect 45828 3290 45884 3292
rect 45908 3290 45964 3292
rect 45668 3238 45714 3290
rect 45714 3238 45724 3290
rect 45748 3238 45778 3290
rect 45778 3238 45790 3290
rect 45790 3238 45804 3290
rect 45828 3238 45842 3290
rect 45842 3238 45854 3290
rect 45854 3238 45884 3290
rect 45908 3238 45918 3290
rect 45918 3238 45964 3290
rect 45668 3236 45724 3238
rect 45748 3236 45804 3238
rect 45828 3236 45884 3238
rect 45908 3236 45964 3238
rect 45668 2202 45724 2204
rect 45748 2202 45804 2204
rect 45828 2202 45884 2204
rect 45908 2202 45964 2204
rect 45668 2150 45714 2202
rect 45714 2150 45724 2202
rect 45748 2150 45778 2202
rect 45778 2150 45790 2202
rect 45790 2150 45804 2202
rect 45828 2150 45842 2202
rect 45842 2150 45854 2202
rect 45854 2150 45884 2202
rect 45908 2150 45918 2202
rect 45918 2150 45964 2202
rect 45668 2148 45724 2150
rect 45748 2148 45804 2150
rect 45828 2148 45884 2150
rect 45908 2148 45964 2150
rect 40079 1658 40135 1660
rect 40159 1658 40215 1660
rect 40239 1658 40295 1660
rect 40319 1658 40375 1660
rect 40079 1606 40125 1658
rect 40125 1606 40135 1658
rect 40159 1606 40189 1658
rect 40189 1606 40201 1658
rect 40201 1606 40215 1658
rect 40239 1606 40253 1658
rect 40253 1606 40265 1658
rect 40265 1606 40295 1658
rect 40319 1606 40329 1658
rect 40329 1606 40375 1658
rect 40079 1604 40135 1606
rect 40159 1604 40215 1606
rect 40239 1604 40295 1606
rect 40319 1604 40375 1606
rect 45668 1114 45724 1116
rect 45748 1114 45804 1116
rect 45828 1114 45884 1116
rect 45908 1114 45964 1116
rect 45668 1062 45714 1114
rect 45714 1062 45724 1114
rect 45748 1062 45778 1114
rect 45778 1062 45790 1114
rect 45790 1062 45804 1114
rect 45828 1062 45842 1114
rect 45842 1062 45854 1114
rect 45854 1062 45884 1114
rect 45908 1062 45918 1114
rect 45918 1062 45964 1114
rect 45668 1060 45724 1062
rect 45748 1060 45804 1062
rect 45828 1060 45884 1062
rect 45908 1060 45964 1062
<< metal3 >>
rect 21725 9890 21791 9893
rect 26693 9890 26759 9893
rect 21725 9888 26759 9890
rect 21725 9832 21730 9888
rect 21786 9832 26698 9888
rect 26754 9832 26759 9888
rect 21725 9830 26759 9832
rect 21725 9827 21791 9830
rect 26693 9827 26759 9830
rect 9673 9754 9739 9757
rect 20253 9754 20319 9757
rect 9673 9752 20319 9754
rect 9673 9696 9678 9752
rect 9734 9696 20258 9752
rect 20314 9696 20319 9752
rect 9673 9694 20319 9696
rect 9673 9691 9739 9694
rect 20253 9691 20319 9694
rect 21357 9754 21423 9757
rect 27061 9754 27127 9757
rect 21357 9752 27127 9754
rect 21357 9696 21362 9752
rect 21418 9696 27066 9752
rect 27122 9696 27127 9752
rect 21357 9694 27127 9696
rect 21357 9691 21423 9694
rect 27061 9691 27127 9694
rect 21725 9618 21791 9621
rect 28165 9618 28231 9621
rect 21725 9616 28231 9618
rect 21725 9560 21730 9616
rect 21786 9560 28170 9616
rect 28226 9560 28231 9616
rect 21725 9558 28231 9560
rect 21725 9555 21791 9558
rect 28165 9555 28231 9558
rect 21725 9482 21791 9485
rect 22093 9482 22159 9485
rect 21725 9480 22159 9482
rect 21725 9424 21730 9480
rect 21786 9424 22098 9480
rect 22154 9424 22159 9480
rect 21725 9422 22159 9424
rect 21725 9419 21791 9422
rect 22093 9419 22159 9422
rect 21541 9346 21607 9349
rect 23749 9346 23815 9349
rect 21541 9344 23815 9346
rect 21541 9288 21546 9344
rect 21602 9288 23754 9344
rect 23810 9288 23815 9344
rect 21541 9286 23815 9288
rect 21541 9283 21607 9286
rect 23749 9283 23815 9286
rect 13721 9210 13787 9213
rect 20662 9210 20668 9212
rect 13721 9208 20668 9210
rect 13721 9152 13726 9208
rect 13782 9152 20668 9208
rect 13721 9150 20668 9152
rect 13721 9147 13787 9150
rect 20662 9148 20668 9150
rect 20732 9148 20738 9212
rect 20805 9210 20871 9213
rect 26233 9210 26299 9213
rect 20805 9208 26299 9210
rect 20805 9152 20810 9208
rect 20866 9152 26238 9208
rect 26294 9152 26299 9208
rect 20805 9150 26299 9152
rect 20805 9147 20871 9150
rect 26233 9147 26299 9150
rect 25589 9074 25655 9077
rect 2730 9072 25655 9074
rect 2730 9016 25594 9072
rect 25650 9016 25655 9072
rect 2730 9014 25655 9016
rect 2730 8941 2790 9014
rect 25589 9011 25655 9014
rect 2681 8936 2790 8941
rect 2681 8880 2686 8936
rect 2742 8880 2790 8936
rect 2681 8878 2790 8880
rect 16573 8938 16639 8941
rect 22829 8938 22895 8941
rect 16573 8936 22895 8938
rect 16573 8880 16578 8936
rect 16634 8880 22834 8936
rect 22890 8880 22895 8936
rect 16573 8878 22895 8880
rect 2681 8875 2747 8878
rect 16573 8875 16639 8878
rect 22829 8875 22895 8878
rect 17125 8802 17191 8805
rect 22829 8802 22895 8805
rect 17125 8800 22895 8802
rect 17125 8744 17130 8800
rect 17186 8744 22834 8800
rect 22890 8744 22895 8800
rect 17125 8742 22895 8744
rect 17125 8739 17191 8742
rect 22829 8739 22895 8742
rect 12124 8736 12440 8737
rect 12124 8672 12130 8736
rect 12194 8672 12210 8736
rect 12274 8672 12290 8736
rect 12354 8672 12370 8736
rect 12434 8672 12440 8736
rect 12124 8671 12440 8672
rect 23302 8736 23618 8737
rect 23302 8672 23308 8736
rect 23372 8672 23388 8736
rect 23452 8672 23468 8736
rect 23532 8672 23548 8736
rect 23612 8672 23618 8736
rect 23302 8671 23618 8672
rect 34480 8736 34796 8737
rect 34480 8672 34486 8736
rect 34550 8672 34566 8736
rect 34630 8672 34646 8736
rect 34710 8672 34726 8736
rect 34790 8672 34796 8736
rect 34480 8671 34796 8672
rect 45658 8736 45974 8737
rect 45658 8672 45664 8736
rect 45728 8672 45744 8736
rect 45808 8672 45824 8736
rect 45888 8672 45904 8736
rect 45968 8672 45974 8736
rect 45658 8671 45974 8672
rect 15561 8666 15627 8669
rect 22461 8666 22527 8669
rect 15561 8664 22527 8666
rect 15561 8608 15566 8664
rect 15622 8608 22466 8664
rect 22522 8608 22527 8664
rect 15561 8606 22527 8608
rect 15561 8603 15627 8606
rect 22461 8603 22527 8606
rect 15101 8530 15167 8533
rect 23473 8530 23539 8533
rect 23841 8530 23907 8533
rect 15101 8528 22110 8530
rect 15101 8472 15106 8528
rect 15162 8472 22110 8528
rect 15101 8470 22110 8472
rect 15101 8467 15167 8470
rect 16849 8394 16915 8397
rect 21173 8394 21239 8397
rect 16849 8392 21239 8394
rect 16849 8336 16854 8392
rect 16910 8336 21178 8392
rect 21234 8336 21239 8392
rect 16849 8334 21239 8336
rect 22050 8394 22110 8470
rect 23473 8528 23907 8530
rect 23473 8472 23478 8528
rect 23534 8472 23846 8528
rect 23902 8472 23907 8528
rect 23473 8470 23907 8472
rect 23473 8467 23539 8470
rect 23841 8467 23907 8470
rect 27429 8394 27495 8397
rect 22050 8392 27495 8394
rect 22050 8336 27434 8392
rect 27490 8336 27495 8392
rect 22050 8334 27495 8336
rect 16849 8331 16915 8334
rect 21173 8331 21239 8334
rect 27429 8331 27495 8334
rect 19333 8258 19399 8261
rect 22553 8258 22619 8261
rect 19333 8256 22619 8258
rect 19333 8200 19338 8256
rect 19394 8200 22558 8256
rect 22614 8200 22619 8256
rect 19333 8198 22619 8200
rect 19333 8195 19399 8198
rect 22553 8195 22619 8198
rect 6535 8192 6851 8193
rect 6535 8128 6541 8192
rect 6605 8128 6621 8192
rect 6685 8128 6701 8192
rect 6765 8128 6781 8192
rect 6845 8128 6851 8192
rect 6535 8127 6851 8128
rect 17713 8192 18029 8193
rect 17713 8128 17719 8192
rect 17783 8128 17799 8192
rect 17863 8128 17879 8192
rect 17943 8128 17959 8192
rect 18023 8128 18029 8192
rect 17713 8127 18029 8128
rect 28891 8192 29207 8193
rect 28891 8128 28897 8192
rect 28961 8128 28977 8192
rect 29041 8128 29057 8192
rect 29121 8128 29137 8192
rect 29201 8128 29207 8192
rect 28891 8127 29207 8128
rect 40069 8192 40385 8193
rect 40069 8128 40075 8192
rect 40139 8128 40155 8192
rect 40219 8128 40235 8192
rect 40299 8128 40315 8192
rect 40379 8128 40385 8192
rect 40069 8127 40385 8128
rect 18413 8122 18479 8125
rect 24209 8122 24275 8125
rect 18413 8120 24275 8122
rect 18413 8064 18418 8120
rect 18474 8064 24214 8120
rect 24270 8064 24275 8120
rect 18413 8062 24275 8064
rect 18413 8059 18479 8062
rect 24209 8059 24275 8062
rect 12525 7986 12591 7989
rect 25497 7986 25563 7989
rect 12525 7984 25563 7986
rect 12525 7928 12530 7984
rect 12586 7928 25502 7984
rect 25558 7928 25563 7984
rect 12525 7926 25563 7928
rect 12525 7923 12591 7926
rect 25497 7923 25563 7926
rect 11789 7850 11855 7853
rect 20345 7850 20411 7853
rect 11789 7848 20411 7850
rect 11789 7792 11794 7848
rect 11850 7792 20350 7848
rect 20406 7792 20411 7848
rect 11789 7790 20411 7792
rect 11789 7787 11855 7790
rect 20345 7787 20411 7790
rect 20662 7788 20668 7852
rect 20732 7850 20738 7852
rect 21541 7850 21607 7853
rect 20732 7848 21607 7850
rect 20732 7792 21546 7848
rect 21602 7792 21607 7848
rect 20732 7790 21607 7792
rect 20732 7788 20738 7790
rect 21541 7787 21607 7790
rect 22001 7850 22067 7853
rect 24761 7850 24827 7853
rect 38101 7850 38167 7853
rect 22001 7848 24594 7850
rect 22001 7792 22006 7848
rect 22062 7792 24594 7848
rect 22001 7790 24594 7792
rect 22001 7787 22067 7790
rect 17217 7714 17283 7717
rect 22001 7714 22067 7717
rect 17217 7712 22067 7714
rect 17217 7656 17222 7712
rect 17278 7656 22006 7712
rect 22062 7656 22067 7712
rect 17217 7654 22067 7656
rect 24534 7714 24594 7790
rect 24761 7848 38167 7850
rect 24761 7792 24766 7848
rect 24822 7792 38106 7848
rect 38162 7792 38167 7848
rect 24761 7790 38167 7792
rect 24761 7787 24827 7790
rect 38101 7787 38167 7790
rect 31661 7714 31727 7717
rect 24534 7712 31727 7714
rect 24534 7656 31666 7712
rect 31722 7656 31727 7712
rect 24534 7654 31727 7656
rect 17217 7651 17283 7654
rect 22001 7651 22067 7654
rect 31661 7651 31727 7654
rect 12124 7648 12440 7649
rect 12124 7584 12130 7648
rect 12194 7584 12210 7648
rect 12274 7584 12290 7648
rect 12354 7584 12370 7648
rect 12434 7584 12440 7648
rect 12124 7583 12440 7584
rect 23302 7648 23618 7649
rect 23302 7584 23308 7648
rect 23372 7584 23388 7648
rect 23452 7584 23468 7648
rect 23532 7584 23548 7648
rect 23612 7584 23618 7648
rect 23302 7583 23618 7584
rect 34480 7648 34796 7649
rect 34480 7584 34486 7648
rect 34550 7584 34566 7648
rect 34630 7584 34646 7648
rect 34710 7584 34726 7648
rect 34790 7584 34796 7648
rect 34480 7583 34796 7584
rect 45658 7648 45974 7649
rect 45658 7584 45664 7648
rect 45728 7584 45744 7648
rect 45808 7584 45824 7648
rect 45888 7584 45904 7648
rect 45968 7584 45974 7648
rect 45658 7583 45974 7584
rect 15101 7578 15167 7581
rect 20069 7578 20135 7581
rect 15101 7576 20135 7578
rect 15101 7520 15106 7576
rect 15162 7520 20074 7576
rect 20130 7520 20135 7576
rect 15101 7518 20135 7520
rect 15101 7515 15167 7518
rect 20069 7515 20135 7518
rect 19333 7442 19399 7445
rect 31937 7442 32003 7445
rect 19333 7440 32003 7442
rect 19333 7384 19338 7440
rect 19394 7384 31942 7440
rect 31998 7384 32003 7440
rect 19333 7382 32003 7384
rect 19333 7379 19399 7382
rect 31937 7379 32003 7382
rect 9673 7306 9739 7309
rect 19517 7306 19583 7309
rect 9673 7304 19583 7306
rect 9673 7248 9678 7304
rect 9734 7248 19522 7304
rect 19578 7248 19583 7304
rect 9673 7246 19583 7248
rect 9673 7243 9739 7246
rect 19517 7243 19583 7246
rect 21909 7306 21975 7309
rect 23473 7306 23539 7309
rect 21909 7304 23539 7306
rect 21909 7248 21914 7304
rect 21970 7248 23478 7304
rect 23534 7248 23539 7304
rect 21909 7246 23539 7248
rect 21909 7243 21975 7246
rect 23473 7243 23539 7246
rect 23749 7306 23815 7309
rect 38469 7306 38535 7309
rect 23749 7304 38535 7306
rect 23749 7248 23754 7304
rect 23810 7248 38474 7304
rect 38530 7248 38535 7304
rect 23749 7246 38535 7248
rect 23749 7243 23815 7246
rect 38469 7243 38535 7246
rect 19057 7170 19123 7173
rect 23197 7170 23263 7173
rect 19057 7168 23263 7170
rect 19057 7112 19062 7168
rect 19118 7112 23202 7168
rect 23258 7112 23263 7168
rect 19057 7110 23263 7112
rect 19057 7107 19123 7110
rect 23197 7107 23263 7110
rect 23565 7170 23631 7173
rect 24761 7170 24827 7173
rect 23565 7168 24827 7170
rect 23565 7112 23570 7168
rect 23626 7112 24766 7168
rect 24822 7112 24827 7168
rect 23565 7110 24827 7112
rect 23565 7107 23631 7110
rect 24761 7107 24827 7110
rect 6535 7104 6851 7105
rect 6535 7040 6541 7104
rect 6605 7040 6621 7104
rect 6685 7040 6701 7104
rect 6765 7040 6781 7104
rect 6845 7040 6851 7104
rect 6535 7039 6851 7040
rect 17713 7104 18029 7105
rect 17713 7040 17719 7104
rect 17783 7040 17799 7104
rect 17863 7040 17879 7104
rect 17943 7040 17959 7104
rect 18023 7040 18029 7104
rect 17713 7039 18029 7040
rect 28891 7104 29207 7105
rect 28891 7040 28897 7104
rect 28961 7040 28977 7104
rect 29041 7040 29057 7104
rect 29121 7040 29137 7104
rect 29201 7040 29207 7104
rect 28891 7039 29207 7040
rect 40069 7104 40385 7105
rect 40069 7040 40075 7104
rect 40139 7040 40155 7104
rect 40219 7040 40235 7104
rect 40299 7040 40315 7104
rect 40379 7040 40385 7104
rect 40069 7039 40385 7040
rect 18505 7034 18571 7037
rect 23841 7034 23907 7037
rect 18505 7032 23907 7034
rect 18505 6976 18510 7032
rect 18566 6976 23846 7032
rect 23902 6976 23907 7032
rect 18505 6974 23907 6976
rect 18505 6971 18571 6974
rect 23841 6971 23907 6974
rect 2957 6898 3023 6901
rect 25589 6898 25655 6901
rect 2957 6896 25655 6898
rect 2957 6840 2962 6896
rect 3018 6840 25594 6896
rect 25650 6840 25655 6896
rect 2957 6838 25655 6840
rect 2957 6835 3023 6838
rect 25589 6835 25655 6838
rect 11697 6762 11763 6765
rect 28533 6762 28599 6765
rect 11697 6760 28599 6762
rect 11697 6704 11702 6760
rect 11758 6704 28538 6760
rect 28594 6704 28599 6760
rect 11697 6702 28599 6704
rect 11697 6699 11763 6702
rect 28533 6699 28599 6702
rect 12124 6560 12440 6561
rect 12124 6496 12130 6560
rect 12194 6496 12210 6560
rect 12274 6496 12290 6560
rect 12354 6496 12370 6560
rect 12434 6496 12440 6560
rect 12124 6495 12440 6496
rect 23302 6560 23618 6561
rect 23302 6496 23308 6560
rect 23372 6496 23388 6560
rect 23452 6496 23468 6560
rect 23532 6496 23548 6560
rect 23612 6496 23618 6560
rect 23302 6495 23618 6496
rect 34480 6560 34796 6561
rect 34480 6496 34486 6560
rect 34550 6496 34566 6560
rect 34630 6496 34646 6560
rect 34710 6496 34726 6560
rect 34790 6496 34796 6560
rect 34480 6495 34796 6496
rect 45658 6560 45974 6561
rect 45658 6496 45664 6560
rect 45728 6496 45744 6560
rect 45808 6496 45824 6560
rect 45888 6496 45904 6560
rect 45968 6496 45974 6560
rect 45658 6495 45974 6496
rect 8293 6354 8359 6357
rect 26417 6354 26483 6357
rect 8293 6352 26483 6354
rect 8293 6296 8298 6352
rect 8354 6296 26422 6352
rect 26478 6296 26483 6352
rect 8293 6294 26483 6296
rect 8293 6291 8359 6294
rect 26417 6291 26483 6294
rect 7005 6218 7071 6221
rect 25037 6218 25103 6221
rect 7005 6216 25103 6218
rect 7005 6160 7010 6216
rect 7066 6160 25042 6216
rect 25098 6160 25103 6216
rect 7005 6158 25103 6160
rect 7005 6155 7071 6158
rect 25037 6155 25103 6158
rect 6535 6016 6851 6017
rect 6535 5952 6541 6016
rect 6605 5952 6621 6016
rect 6685 5952 6701 6016
rect 6765 5952 6781 6016
rect 6845 5952 6851 6016
rect 6535 5951 6851 5952
rect 17713 6016 18029 6017
rect 17713 5952 17719 6016
rect 17783 5952 17799 6016
rect 17863 5952 17879 6016
rect 17943 5952 17959 6016
rect 18023 5952 18029 6016
rect 17713 5951 18029 5952
rect 28891 6016 29207 6017
rect 28891 5952 28897 6016
rect 28961 5952 28977 6016
rect 29041 5952 29057 6016
rect 29121 5952 29137 6016
rect 29201 5952 29207 6016
rect 28891 5951 29207 5952
rect 40069 6016 40385 6017
rect 40069 5952 40075 6016
rect 40139 5952 40155 6016
rect 40219 5952 40235 6016
rect 40299 5952 40315 6016
rect 40379 5952 40385 6016
rect 40069 5951 40385 5952
rect 8937 5810 9003 5813
rect 21725 5810 21791 5813
rect 8937 5808 21791 5810
rect 8937 5752 8942 5808
rect 8998 5752 21730 5808
rect 21786 5752 21791 5808
rect 8937 5750 21791 5752
rect 8937 5747 9003 5750
rect 21725 5747 21791 5750
rect 12124 5472 12440 5473
rect 12124 5408 12130 5472
rect 12194 5408 12210 5472
rect 12274 5408 12290 5472
rect 12354 5408 12370 5472
rect 12434 5408 12440 5472
rect 12124 5407 12440 5408
rect 23302 5472 23618 5473
rect 23302 5408 23308 5472
rect 23372 5408 23388 5472
rect 23452 5408 23468 5472
rect 23532 5408 23548 5472
rect 23612 5408 23618 5472
rect 23302 5407 23618 5408
rect 34480 5472 34796 5473
rect 34480 5408 34486 5472
rect 34550 5408 34566 5472
rect 34630 5408 34646 5472
rect 34710 5408 34726 5472
rect 34790 5408 34796 5472
rect 34480 5407 34796 5408
rect 45658 5472 45974 5473
rect 45658 5408 45664 5472
rect 45728 5408 45744 5472
rect 45808 5408 45824 5472
rect 45888 5408 45904 5472
rect 45968 5408 45974 5472
rect 45658 5407 45974 5408
rect 6535 4928 6851 4929
rect 6535 4864 6541 4928
rect 6605 4864 6621 4928
rect 6685 4864 6701 4928
rect 6765 4864 6781 4928
rect 6845 4864 6851 4928
rect 6535 4863 6851 4864
rect 17713 4928 18029 4929
rect 17713 4864 17719 4928
rect 17783 4864 17799 4928
rect 17863 4864 17879 4928
rect 17943 4864 17959 4928
rect 18023 4864 18029 4928
rect 17713 4863 18029 4864
rect 28891 4928 29207 4929
rect 28891 4864 28897 4928
rect 28961 4864 28977 4928
rect 29041 4864 29057 4928
rect 29121 4864 29137 4928
rect 29201 4864 29207 4928
rect 28891 4863 29207 4864
rect 40069 4928 40385 4929
rect 40069 4864 40075 4928
rect 40139 4864 40155 4928
rect 40219 4864 40235 4928
rect 40299 4864 40315 4928
rect 40379 4864 40385 4928
rect 40069 4863 40385 4864
rect 12124 4384 12440 4385
rect 12124 4320 12130 4384
rect 12194 4320 12210 4384
rect 12274 4320 12290 4384
rect 12354 4320 12370 4384
rect 12434 4320 12440 4384
rect 12124 4319 12440 4320
rect 23302 4384 23618 4385
rect 23302 4320 23308 4384
rect 23372 4320 23388 4384
rect 23452 4320 23468 4384
rect 23532 4320 23548 4384
rect 23612 4320 23618 4384
rect 23302 4319 23618 4320
rect 34480 4384 34796 4385
rect 34480 4320 34486 4384
rect 34550 4320 34566 4384
rect 34630 4320 34646 4384
rect 34710 4320 34726 4384
rect 34790 4320 34796 4384
rect 34480 4319 34796 4320
rect 45658 4384 45974 4385
rect 45658 4320 45664 4384
rect 45728 4320 45744 4384
rect 45808 4320 45824 4384
rect 45888 4320 45904 4384
rect 45968 4320 45974 4384
rect 45658 4319 45974 4320
rect 6535 3840 6851 3841
rect 6535 3776 6541 3840
rect 6605 3776 6621 3840
rect 6685 3776 6701 3840
rect 6765 3776 6781 3840
rect 6845 3776 6851 3840
rect 6535 3775 6851 3776
rect 17713 3840 18029 3841
rect 17713 3776 17719 3840
rect 17783 3776 17799 3840
rect 17863 3776 17879 3840
rect 17943 3776 17959 3840
rect 18023 3776 18029 3840
rect 17713 3775 18029 3776
rect 28891 3840 29207 3841
rect 28891 3776 28897 3840
rect 28961 3776 28977 3840
rect 29041 3776 29057 3840
rect 29121 3776 29137 3840
rect 29201 3776 29207 3840
rect 28891 3775 29207 3776
rect 40069 3840 40385 3841
rect 40069 3776 40075 3840
rect 40139 3776 40155 3840
rect 40219 3776 40235 3840
rect 40299 3776 40315 3840
rect 40379 3776 40385 3840
rect 40069 3775 40385 3776
rect 12124 3296 12440 3297
rect 12124 3232 12130 3296
rect 12194 3232 12210 3296
rect 12274 3232 12290 3296
rect 12354 3232 12370 3296
rect 12434 3232 12440 3296
rect 12124 3231 12440 3232
rect 23302 3296 23618 3297
rect 23302 3232 23308 3296
rect 23372 3232 23388 3296
rect 23452 3232 23468 3296
rect 23532 3232 23548 3296
rect 23612 3232 23618 3296
rect 23302 3231 23618 3232
rect 34480 3296 34796 3297
rect 34480 3232 34486 3296
rect 34550 3232 34566 3296
rect 34630 3232 34646 3296
rect 34710 3232 34726 3296
rect 34790 3232 34796 3296
rect 34480 3231 34796 3232
rect 45658 3296 45974 3297
rect 45658 3232 45664 3296
rect 45728 3232 45744 3296
rect 45808 3232 45824 3296
rect 45888 3232 45904 3296
rect 45968 3232 45974 3296
rect 45658 3231 45974 3232
rect 6535 2752 6851 2753
rect 6535 2688 6541 2752
rect 6605 2688 6621 2752
rect 6685 2688 6701 2752
rect 6765 2688 6781 2752
rect 6845 2688 6851 2752
rect 6535 2687 6851 2688
rect 17713 2752 18029 2753
rect 17713 2688 17719 2752
rect 17783 2688 17799 2752
rect 17863 2688 17879 2752
rect 17943 2688 17959 2752
rect 18023 2688 18029 2752
rect 17713 2687 18029 2688
rect 28891 2752 29207 2753
rect 28891 2688 28897 2752
rect 28961 2688 28977 2752
rect 29041 2688 29057 2752
rect 29121 2688 29137 2752
rect 29201 2688 29207 2752
rect 28891 2687 29207 2688
rect 40069 2752 40385 2753
rect 40069 2688 40075 2752
rect 40139 2688 40155 2752
rect 40219 2688 40235 2752
rect 40299 2688 40315 2752
rect 40379 2688 40385 2752
rect 40069 2687 40385 2688
rect 12124 2208 12440 2209
rect 12124 2144 12130 2208
rect 12194 2144 12210 2208
rect 12274 2144 12290 2208
rect 12354 2144 12370 2208
rect 12434 2144 12440 2208
rect 12124 2143 12440 2144
rect 23302 2208 23618 2209
rect 23302 2144 23308 2208
rect 23372 2144 23388 2208
rect 23452 2144 23468 2208
rect 23532 2144 23548 2208
rect 23612 2144 23618 2208
rect 23302 2143 23618 2144
rect 34480 2208 34796 2209
rect 34480 2144 34486 2208
rect 34550 2144 34566 2208
rect 34630 2144 34646 2208
rect 34710 2144 34726 2208
rect 34790 2144 34796 2208
rect 34480 2143 34796 2144
rect 45658 2208 45974 2209
rect 45658 2144 45664 2208
rect 45728 2144 45744 2208
rect 45808 2144 45824 2208
rect 45888 2144 45904 2208
rect 45968 2144 45974 2208
rect 45658 2143 45974 2144
rect 6535 1664 6851 1665
rect 6535 1600 6541 1664
rect 6605 1600 6621 1664
rect 6685 1600 6701 1664
rect 6765 1600 6781 1664
rect 6845 1600 6851 1664
rect 6535 1599 6851 1600
rect 17713 1664 18029 1665
rect 17713 1600 17719 1664
rect 17783 1600 17799 1664
rect 17863 1600 17879 1664
rect 17943 1600 17959 1664
rect 18023 1600 18029 1664
rect 17713 1599 18029 1600
rect 28891 1664 29207 1665
rect 28891 1600 28897 1664
rect 28961 1600 28977 1664
rect 29041 1600 29057 1664
rect 29121 1600 29137 1664
rect 29201 1600 29207 1664
rect 28891 1599 29207 1600
rect 40069 1664 40385 1665
rect 40069 1600 40075 1664
rect 40139 1600 40155 1664
rect 40219 1600 40235 1664
rect 40299 1600 40315 1664
rect 40379 1600 40385 1664
rect 40069 1599 40385 1600
rect 12124 1120 12440 1121
rect 12124 1056 12130 1120
rect 12194 1056 12210 1120
rect 12274 1056 12290 1120
rect 12354 1056 12370 1120
rect 12434 1056 12440 1120
rect 12124 1055 12440 1056
rect 23302 1120 23618 1121
rect 23302 1056 23308 1120
rect 23372 1056 23388 1120
rect 23452 1056 23468 1120
rect 23532 1056 23548 1120
rect 23612 1056 23618 1120
rect 23302 1055 23618 1056
rect 34480 1120 34796 1121
rect 34480 1056 34486 1120
rect 34550 1056 34566 1120
rect 34630 1056 34646 1120
rect 34710 1056 34726 1120
rect 34790 1056 34796 1120
rect 34480 1055 34796 1056
rect 45658 1120 45974 1121
rect 45658 1056 45664 1120
rect 45728 1056 45744 1120
rect 45808 1056 45824 1120
rect 45888 1056 45904 1120
rect 45968 1056 45974 1120
rect 45658 1055 45974 1056
<< via3 >>
rect 20668 9148 20732 9212
rect 12130 8732 12194 8736
rect 12130 8676 12134 8732
rect 12134 8676 12190 8732
rect 12190 8676 12194 8732
rect 12130 8672 12194 8676
rect 12210 8732 12274 8736
rect 12210 8676 12214 8732
rect 12214 8676 12270 8732
rect 12270 8676 12274 8732
rect 12210 8672 12274 8676
rect 12290 8732 12354 8736
rect 12290 8676 12294 8732
rect 12294 8676 12350 8732
rect 12350 8676 12354 8732
rect 12290 8672 12354 8676
rect 12370 8732 12434 8736
rect 12370 8676 12374 8732
rect 12374 8676 12430 8732
rect 12430 8676 12434 8732
rect 12370 8672 12434 8676
rect 23308 8732 23372 8736
rect 23308 8676 23312 8732
rect 23312 8676 23368 8732
rect 23368 8676 23372 8732
rect 23308 8672 23372 8676
rect 23388 8732 23452 8736
rect 23388 8676 23392 8732
rect 23392 8676 23448 8732
rect 23448 8676 23452 8732
rect 23388 8672 23452 8676
rect 23468 8732 23532 8736
rect 23468 8676 23472 8732
rect 23472 8676 23528 8732
rect 23528 8676 23532 8732
rect 23468 8672 23532 8676
rect 23548 8732 23612 8736
rect 23548 8676 23552 8732
rect 23552 8676 23608 8732
rect 23608 8676 23612 8732
rect 23548 8672 23612 8676
rect 34486 8732 34550 8736
rect 34486 8676 34490 8732
rect 34490 8676 34546 8732
rect 34546 8676 34550 8732
rect 34486 8672 34550 8676
rect 34566 8732 34630 8736
rect 34566 8676 34570 8732
rect 34570 8676 34626 8732
rect 34626 8676 34630 8732
rect 34566 8672 34630 8676
rect 34646 8732 34710 8736
rect 34646 8676 34650 8732
rect 34650 8676 34706 8732
rect 34706 8676 34710 8732
rect 34646 8672 34710 8676
rect 34726 8732 34790 8736
rect 34726 8676 34730 8732
rect 34730 8676 34786 8732
rect 34786 8676 34790 8732
rect 34726 8672 34790 8676
rect 45664 8732 45728 8736
rect 45664 8676 45668 8732
rect 45668 8676 45724 8732
rect 45724 8676 45728 8732
rect 45664 8672 45728 8676
rect 45744 8732 45808 8736
rect 45744 8676 45748 8732
rect 45748 8676 45804 8732
rect 45804 8676 45808 8732
rect 45744 8672 45808 8676
rect 45824 8732 45888 8736
rect 45824 8676 45828 8732
rect 45828 8676 45884 8732
rect 45884 8676 45888 8732
rect 45824 8672 45888 8676
rect 45904 8732 45968 8736
rect 45904 8676 45908 8732
rect 45908 8676 45964 8732
rect 45964 8676 45968 8732
rect 45904 8672 45968 8676
rect 6541 8188 6605 8192
rect 6541 8132 6545 8188
rect 6545 8132 6601 8188
rect 6601 8132 6605 8188
rect 6541 8128 6605 8132
rect 6621 8188 6685 8192
rect 6621 8132 6625 8188
rect 6625 8132 6681 8188
rect 6681 8132 6685 8188
rect 6621 8128 6685 8132
rect 6701 8188 6765 8192
rect 6701 8132 6705 8188
rect 6705 8132 6761 8188
rect 6761 8132 6765 8188
rect 6701 8128 6765 8132
rect 6781 8188 6845 8192
rect 6781 8132 6785 8188
rect 6785 8132 6841 8188
rect 6841 8132 6845 8188
rect 6781 8128 6845 8132
rect 17719 8188 17783 8192
rect 17719 8132 17723 8188
rect 17723 8132 17779 8188
rect 17779 8132 17783 8188
rect 17719 8128 17783 8132
rect 17799 8188 17863 8192
rect 17799 8132 17803 8188
rect 17803 8132 17859 8188
rect 17859 8132 17863 8188
rect 17799 8128 17863 8132
rect 17879 8188 17943 8192
rect 17879 8132 17883 8188
rect 17883 8132 17939 8188
rect 17939 8132 17943 8188
rect 17879 8128 17943 8132
rect 17959 8188 18023 8192
rect 17959 8132 17963 8188
rect 17963 8132 18019 8188
rect 18019 8132 18023 8188
rect 17959 8128 18023 8132
rect 28897 8188 28961 8192
rect 28897 8132 28901 8188
rect 28901 8132 28957 8188
rect 28957 8132 28961 8188
rect 28897 8128 28961 8132
rect 28977 8188 29041 8192
rect 28977 8132 28981 8188
rect 28981 8132 29037 8188
rect 29037 8132 29041 8188
rect 28977 8128 29041 8132
rect 29057 8188 29121 8192
rect 29057 8132 29061 8188
rect 29061 8132 29117 8188
rect 29117 8132 29121 8188
rect 29057 8128 29121 8132
rect 29137 8188 29201 8192
rect 29137 8132 29141 8188
rect 29141 8132 29197 8188
rect 29197 8132 29201 8188
rect 29137 8128 29201 8132
rect 40075 8188 40139 8192
rect 40075 8132 40079 8188
rect 40079 8132 40135 8188
rect 40135 8132 40139 8188
rect 40075 8128 40139 8132
rect 40155 8188 40219 8192
rect 40155 8132 40159 8188
rect 40159 8132 40215 8188
rect 40215 8132 40219 8188
rect 40155 8128 40219 8132
rect 40235 8188 40299 8192
rect 40235 8132 40239 8188
rect 40239 8132 40295 8188
rect 40295 8132 40299 8188
rect 40235 8128 40299 8132
rect 40315 8188 40379 8192
rect 40315 8132 40319 8188
rect 40319 8132 40375 8188
rect 40375 8132 40379 8188
rect 40315 8128 40379 8132
rect 20668 7788 20732 7852
rect 12130 7644 12194 7648
rect 12130 7588 12134 7644
rect 12134 7588 12190 7644
rect 12190 7588 12194 7644
rect 12130 7584 12194 7588
rect 12210 7644 12274 7648
rect 12210 7588 12214 7644
rect 12214 7588 12270 7644
rect 12270 7588 12274 7644
rect 12210 7584 12274 7588
rect 12290 7644 12354 7648
rect 12290 7588 12294 7644
rect 12294 7588 12350 7644
rect 12350 7588 12354 7644
rect 12290 7584 12354 7588
rect 12370 7644 12434 7648
rect 12370 7588 12374 7644
rect 12374 7588 12430 7644
rect 12430 7588 12434 7644
rect 12370 7584 12434 7588
rect 23308 7644 23372 7648
rect 23308 7588 23312 7644
rect 23312 7588 23368 7644
rect 23368 7588 23372 7644
rect 23308 7584 23372 7588
rect 23388 7644 23452 7648
rect 23388 7588 23392 7644
rect 23392 7588 23448 7644
rect 23448 7588 23452 7644
rect 23388 7584 23452 7588
rect 23468 7644 23532 7648
rect 23468 7588 23472 7644
rect 23472 7588 23528 7644
rect 23528 7588 23532 7644
rect 23468 7584 23532 7588
rect 23548 7644 23612 7648
rect 23548 7588 23552 7644
rect 23552 7588 23608 7644
rect 23608 7588 23612 7644
rect 23548 7584 23612 7588
rect 34486 7644 34550 7648
rect 34486 7588 34490 7644
rect 34490 7588 34546 7644
rect 34546 7588 34550 7644
rect 34486 7584 34550 7588
rect 34566 7644 34630 7648
rect 34566 7588 34570 7644
rect 34570 7588 34626 7644
rect 34626 7588 34630 7644
rect 34566 7584 34630 7588
rect 34646 7644 34710 7648
rect 34646 7588 34650 7644
rect 34650 7588 34706 7644
rect 34706 7588 34710 7644
rect 34646 7584 34710 7588
rect 34726 7644 34790 7648
rect 34726 7588 34730 7644
rect 34730 7588 34786 7644
rect 34786 7588 34790 7644
rect 34726 7584 34790 7588
rect 45664 7644 45728 7648
rect 45664 7588 45668 7644
rect 45668 7588 45724 7644
rect 45724 7588 45728 7644
rect 45664 7584 45728 7588
rect 45744 7644 45808 7648
rect 45744 7588 45748 7644
rect 45748 7588 45804 7644
rect 45804 7588 45808 7644
rect 45744 7584 45808 7588
rect 45824 7644 45888 7648
rect 45824 7588 45828 7644
rect 45828 7588 45884 7644
rect 45884 7588 45888 7644
rect 45824 7584 45888 7588
rect 45904 7644 45968 7648
rect 45904 7588 45908 7644
rect 45908 7588 45964 7644
rect 45964 7588 45968 7644
rect 45904 7584 45968 7588
rect 6541 7100 6605 7104
rect 6541 7044 6545 7100
rect 6545 7044 6601 7100
rect 6601 7044 6605 7100
rect 6541 7040 6605 7044
rect 6621 7100 6685 7104
rect 6621 7044 6625 7100
rect 6625 7044 6681 7100
rect 6681 7044 6685 7100
rect 6621 7040 6685 7044
rect 6701 7100 6765 7104
rect 6701 7044 6705 7100
rect 6705 7044 6761 7100
rect 6761 7044 6765 7100
rect 6701 7040 6765 7044
rect 6781 7100 6845 7104
rect 6781 7044 6785 7100
rect 6785 7044 6841 7100
rect 6841 7044 6845 7100
rect 6781 7040 6845 7044
rect 17719 7100 17783 7104
rect 17719 7044 17723 7100
rect 17723 7044 17779 7100
rect 17779 7044 17783 7100
rect 17719 7040 17783 7044
rect 17799 7100 17863 7104
rect 17799 7044 17803 7100
rect 17803 7044 17859 7100
rect 17859 7044 17863 7100
rect 17799 7040 17863 7044
rect 17879 7100 17943 7104
rect 17879 7044 17883 7100
rect 17883 7044 17939 7100
rect 17939 7044 17943 7100
rect 17879 7040 17943 7044
rect 17959 7100 18023 7104
rect 17959 7044 17963 7100
rect 17963 7044 18019 7100
rect 18019 7044 18023 7100
rect 17959 7040 18023 7044
rect 28897 7100 28961 7104
rect 28897 7044 28901 7100
rect 28901 7044 28957 7100
rect 28957 7044 28961 7100
rect 28897 7040 28961 7044
rect 28977 7100 29041 7104
rect 28977 7044 28981 7100
rect 28981 7044 29037 7100
rect 29037 7044 29041 7100
rect 28977 7040 29041 7044
rect 29057 7100 29121 7104
rect 29057 7044 29061 7100
rect 29061 7044 29117 7100
rect 29117 7044 29121 7100
rect 29057 7040 29121 7044
rect 29137 7100 29201 7104
rect 29137 7044 29141 7100
rect 29141 7044 29197 7100
rect 29197 7044 29201 7100
rect 29137 7040 29201 7044
rect 40075 7100 40139 7104
rect 40075 7044 40079 7100
rect 40079 7044 40135 7100
rect 40135 7044 40139 7100
rect 40075 7040 40139 7044
rect 40155 7100 40219 7104
rect 40155 7044 40159 7100
rect 40159 7044 40215 7100
rect 40215 7044 40219 7100
rect 40155 7040 40219 7044
rect 40235 7100 40299 7104
rect 40235 7044 40239 7100
rect 40239 7044 40295 7100
rect 40295 7044 40299 7100
rect 40235 7040 40299 7044
rect 40315 7100 40379 7104
rect 40315 7044 40319 7100
rect 40319 7044 40375 7100
rect 40375 7044 40379 7100
rect 40315 7040 40379 7044
rect 12130 6556 12194 6560
rect 12130 6500 12134 6556
rect 12134 6500 12190 6556
rect 12190 6500 12194 6556
rect 12130 6496 12194 6500
rect 12210 6556 12274 6560
rect 12210 6500 12214 6556
rect 12214 6500 12270 6556
rect 12270 6500 12274 6556
rect 12210 6496 12274 6500
rect 12290 6556 12354 6560
rect 12290 6500 12294 6556
rect 12294 6500 12350 6556
rect 12350 6500 12354 6556
rect 12290 6496 12354 6500
rect 12370 6556 12434 6560
rect 12370 6500 12374 6556
rect 12374 6500 12430 6556
rect 12430 6500 12434 6556
rect 12370 6496 12434 6500
rect 23308 6556 23372 6560
rect 23308 6500 23312 6556
rect 23312 6500 23368 6556
rect 23368 6500 23372 6556
rect 23308 6496 23372 6500
rect 23388 6556 23452 6560
rect 23388 6500 23392 6556
rect 23392 6500 23448 6556
rect 23448 6500 23452 6556
rect 23388 6496 23452 6500
rect 23468 6556 23532 6560
rect 23468 6500 23472 6556
rect 23472 6500 23528 6556
rect 23528 6500 23532 6556
rect 23468 6496 23532 6500
rect 23548 6556 23612 6560
rect 23548 6500 23552 6556
rect 23552 6500 23608 6556
rect 23608 6500 23612 6556
rect 23548 6496 23612 6500
rect 34486 6556 34550 6560
rect 34486 6500 34490 6556
rect 34490 6500 34546 6556
rect 34546 6500 34550 6556
rect 34486 6496 34550 6500
rect 34566 6556 34630 6560
rect 34566 6500 34570 6556
rect 34570 6500 34626 6556
rect 34626 6500 34630 6556
rect 34566 6496 34630 6500
rect 34646 6556 34710 6560
rect 34646 6500 34650 6556
rect 34650 6500 34706 6556
rect 34706 6500 34710 6556
rect 34646 6496 34710 6500
rect 34726 6556 34790 6560
rect 34726 6500 34730 6556
rect 34730 6500 34786 6556
rect 34786 6500 34790 6556
rect 34726 6496 34790 6500
rect 45664 6556 45728 6560
rect 45664 6500 45668 6556
rect 45668 6500 45724 6556
rect 45724 6500 45728 6556
rect 45664 6496 45728 6500
rect 45744 6556 45808 6560
rect 45744 6500 45748 6556
rect 45748 6500 45804 6556
rect 45804 6500 45808 6556
rect 45744 6496 45808 6500
rect 45824 6556 45888 6560
rect 45824 6500 45828 6556
rect 45828 6500 45884 6556
rect 45884 6500 45888 6556
rect 45824 6496 45888 6500
rect 45904 6556 45968 6560
rect 45904 6500 45908 6556
rect 45908 6500 45964 6556
rect 45964 6500 45968 6556
rect 45904 6496 45968 6500
rect 6541 6012 6605 6016
rect 6541 5956 6545 6012
rect 6545 5956 6601 6012
rect 6601 5956 6605 6012
rect 6541 5952 6605 5956
rect 6621 6012 6685 6016
rect 6621 5956 6625 6012
rect 6625 5956 6681 6012
rect 6681 5956 6685 6012
rect 6621 5952 6685 5956
rect 6701 6012 6765 6016
rect 6701 5956 6705 6012
rect 6705 5956 6761 6012
rect 6761 5956 6765 6012
rect 6701 5952 6765 5956
rect 6781 6012 6845 6016
rect 6781 5956 6785 6012
rect 6785 5956 6841 6012
rect 6841 5956 6845 6012
rect 6781 5952 6845 5956
rect 17719 6012 17783 6016
rect 17719 5956 17723 6012
rect 17723 5956 17779 6012
rect 17779 5956 17783 6012
rect 17719 5952 17783 5956
rect 17799 6012 17863 6016
rect 17799 5956 17803 6012
rect 17803 5956 17859 6012
rect 17859 5956 17863 6012
rect 17799 5952 17863 5956
rect 17879 6012 17943 6016
rect 17879 5956 17883 6012
rect 17883 5956 17939 6012
rect 17939 5956 17943 6012
rect 17879 5952 17943 5956
rect 17959 6012 18023 6016
rect 17959 5956 17963 6012
rect 17963 5956 18019 6012
rect 18019 5956 18023 6012
rect 17959 5952 18023 5956
rect 28897 6012 28961 6016
rect 28897 5956 28901 6012
rect 28901 5956 28957 6012
rect 28957 5956 28961 6012
rect 28897 5952 28961 5956
rect 28977 6012 29041 6016
rect 28977 5956 28981 6012
rect 28981 5956 29037 6012
rect 29037 5956 29041 6012
rect 28977 5952 29041 5956
rect 29057 6012 29121 6016
rect 29057 5956 29061 6012
rect 29061 5956 29117 6012
rect 29117 5956 29121 6012
rect 29057 5952 29121 5956
rect 29137 6012 29201 6016
rect 29137 5956 29141 6012
rect 29141 5956 29197 6012
rect 29197 5956 29201 6012
rect 29137 5952 29201 5956
rect 40075 6012 40139 6016
rect 40075 5956 40079 6012
rect 40079 5956 40135 6012
rect 40135 5956 40139 6012
rect 40075 5952 40139 5956
rect 40155 6012 40219 6016
rect 40155 5956 40159 6012
rect 40159 5956 40215 6012
rect 40215 5956 40219 6012
rect 40155 5952 40219 5956
rect 40235 6012 40299 6016
rect 40235 5956 40239 6012
rect 40239 5956 40295 6012
rect 40295 5956 40299 6012
rect 40235 5952 40299 5956
rect 40315 6012 40379 6016
rect 40315 5956 40319 6012
rect 40319 5956 40375 6012
rect 40375 5956 40379 6012
rect 40315 5952 40379 5956
rect 12130 5468 12194 5472
rect 12130 5412 12134 5468
rect 12134 5412 12190 5468
rect 12190 5412 12194 5468
rect 12130 5408 12194 5412
rect 12210 5468 12274 5472
rect 12210 5412 12214 5468
rect 12214 5412 12270 5468
rect 12270 5412 12274 5468
rect 12210 5408 12274 5412
rect 12290 5468 12354 5472
rect 12290 5412 12294 5468
rect 12294 5412 12350 5468
rect 12350 5412 12354 5468
rect 12290 5408 12354 5412
rect 12370 5468 12434 5472
rect 12370 5412 12374 5468
rect 12374 5412 12430 5468
rect 12430 5412 12434 5468
rect 12370 5408 12434 5412
rect 23308 5468 23372 5472
rect 23308 5412 23312 5468
rect 23312 5412 23368 5468
rect 23368 5412 23372 5468
rect 23308 5408 23372 5412
rect 23388 5468 23452 5472
rect 23388 5412 23392 5468
rect 23392 5412 23448 5468
rect 23448 5412 23452 5468
rect 23388 5408 23452 5412
rect 23468 5468 23532 5472
rect 23468 5412 23472 5468
rect 23472 5412 23528 5468
rect 23528 5412 23532 5468
rect 23468 5408 23532 5412
rect 23548 5468 23612 5472
rect 23548 5412 23552 5468
rect 23552 5412 23608 5468
rect 23608 5412 23612 5468
rect 23548 5408 23612 5412
rect 34486 5468 34550 5472
rect 34486 5412 34490 5468
rect 34490 5412 34546 5468
rect 34546 5412 34550 5468
rect 34486 5408 34550 5412
rect 34566 5468 34630 5472
rect 34566 5412 34570 5468
rect 34570 5412 34626 5468
rect 34626 5412 34630 5468
rect 34566 5408 34630 5412
rect 34646 5468 34710 5472
rect 34646 5412 34650 5468
rect 34650 5412 34706 5468
rect 34706 5412 34710 5468
rect 34646 5408 34710 5412
rect 34726 5468 34790 5472
rect 34726 5412 34730 5468
rect 34730 5412 34786 5468
rect 34786 5412 34790 5468
rect 34726 5408 34790 5412
rect 45664 5468 45728 5472
rect 45664 5412 45668 5468
rect 45668 5412 45724 5468
rect 45724 5412 45728 5468
rect 45664 5408 45728 5412
rect 45744 5468 45808 5472
rect 45744 5412 45748 5468
rect 45748 5412 45804 5468
rect 45804 5412 45808 5468
rect 45744 5408 45808 5412
rect 45824 5468 45888 5472
rect 45824 5412 45828 5468
rect 45828 5412 45884 5468
rect 45884 5412 45888 5468
rect 45824 5408 45888 5412
rect 45904 5468 45968 5472
rect 45904 5412 45908 5468
rect 45908 5412 45964 5468
rect 45964 5412 45968 5468
rect 45904 5408 45968 5412
rect 6541 4924 6605 4928
rect 6541 4868 6545 4924
rect 6545 4868 6601 4924
rect 6601 4868 6605 4924
rect 6541 4864 6605 4868
rect 6621 4924 6685 4928
rect 6621 4868 6625 4924
rect 6625 4868 6681 4924
rect 6681 4868 6685 4924
rect 6621 4864 6685 4868
rect 6701 4924 6765 4928
rect 6701 4868 6705 4924
rect 6705 4868 6761 4924
rect 6761 4868 6765 4924
rect 6701 4864 6765 4868
rect 6781 4924 6845 4928
rect 6781 4868 6785 4924
rect 6785 4868 6841 4924
rect 6841 4868 6845 4924
rect 6781 4864 6845 4868
rect 17719 4924 17783 4928
rect 17719 4868 17723 4924
rect 17723 4868 17779 4924
rect 17779 4868 17783 4924
rect 17719 4864 17783 4868
rect 17799 4924 17863 4928
rect 17799 4868 17803 4924
rect 17803 4868 17859 4924
rect 17859 4868 17863 4924
rect 17799 4864 17863 4868
rect 17879 4924 17943 4928
rect 17879 4868 17883 4924
rect 17883 4868 17939 4924
rect 17939 4868 17943 4924
rect 17879 4864 17943 4868
rect 17959 4924 18023 4928
rect 17959 4868 17963 4924
rect 17963 4868 18019 4924
rect 18019 4868 18023 4924
rect 17959 4864 18023 4868
rect 28897 4924 28961 4928
rect 28897 4868 28901 4924
rect 28901 4868 28957 4924
rect 28957 4868 28961 4924
rect 28897 4864 28961 4868
rect 28977 4924 29041 4928
rect 28977 4868 28981 4924
rect 28981 4868 29037 4924
rect 29037 4868 29041 4924
rect 28977 4864 29041 4868
rect 29057 4924 29121 4928
rect 29057 4868 29061 4924
rect 29061 4868 29117 4924
rect 29117 4868 29121 4924
rect 29057 4864 29121 4868
rect 29137 4924 29201 4928
rect 29137 4868 29141 4924
rect 29141 4868 29197 4924
rect 29197 4868 29201 4924
rect 29137 4864 29201 4868
rect 40075 4924 40139 4928
rect 40075 4868 40079 4924
rect 40079 4868 40135 4924
rect 40135 4868 40139 4924
rect 40075 4864 40139 4868
rect 40155 4924 40219 4928
rect 40155 4868 40159 4924
rect 40159 4868 40215 4924
rect 40215 4868 40219 4924
rect 40155 4864 40219 4868
rect 40235 4924 40299 4928
rect 40235 4868 40239 4924
rect 40239 4868 40295 4924
rect 40295 4868 40299 4924
rect 40235 4864 40299 4868
rect 40315 4924 40379 4928
rect 40315 4868 40319 4924
rect 40319 4868 40375 4924
rect 40375 4868 40379 4924
rect 40315 4864 40379 4868
rect 12130 4380 12194 4384
rect 12130 4324 12134 4380
rect 12134 4324 12190 4380
rect 12190 4324 12194 4380
rect 12130 4320 12194 4324
rect 12210 4380 12274 4384
rect 12210 4324 12214 4380
rect 12214 4324 12270 4380
rect 12270 4324 12274 4380
rect 12210 4320 12274 4324
rect 12290 4380 12354 4384
rect 12290 4324 12294 4380
rect 12294 4324 12350 4380
rect 12350 4324 12354 4380
rect 12290 4320 12354 4324
rect 12370 4380 12434 4384
rect 12370 4324 12374 4380
rect 12374 4324 12430 4380
rect 12430 4324 12434 4380
rect 12370 4320 12434 4324
rect 23308 4380 23372 4384
rect 23308 4324 23312 4380
rect 23312 4324 23368 4380
rect 23368 4324 23372 4380
rect 23308 4320 23372 4324
rect 23388 4380 23452 4384
rect 23388 4324 23392 4380
rect 23392 4324 23448 4380
rect 23448 4324 23452 4380
rect 23388 4320 23452 4324
rect 23468 4380 23532 4384
rect 23468 4324 23472 4380
rect 23472 4324 23528 4380
rect 23528 4324 23532 4380
rect 23468 4320 23532 4324
rect 23548 4380 23612 4384
rect 23548 4324 23552 4380
rect 23552 4324 23608 4380
rect 23608 4324 23612 4380
rect 23548 4320 23612 4324
rect 34486 4380 34550 4384
rect 34486 4324 34490 4380
rect 34490 4324 34546 4380
rect 34546 4324 34550 4380
rect 34486 4320 34550 4324
rect 34566 4380 34630 4384
rect 34566 4324 34570 4380
rect 34570 4324 34626 4380
rect 34626 4324 34630 4380
rect 34566 4320 34630 4324
rect 34646 4380 34710 4384
rect 34646 4324 34650 4380
rect 34650 4324 34706 4380
rect 34706 4324 34710 4380
rect 34646 4320 34710 4324
rect 34726 4380 34790 4384
rect 34726 4324 34730 4380
rect 34730 4324 34786 4380
rect 34786 4324 34790 4380
rect 34726 4320 34790 4324
rect 45664 4380 45728 4384
rect 45664 4324 45668 4380
rect 45668 4324 45724 4380
rect 45724 4324 45728 4380
rect 45664 4320 45728 4324
rect 45744 4380 45808 4384
rect 45744 4324 45748 4380
rect 45748 4324 45804 4380
rect 45804 4324 45808 4380
rect 45744 4320 45808 4324
rect 45824 4380 45888 4384
rect 45824 4324 45828 4380
rect 45828 4324 45884 4380
rect 45884 4324 45888 4380
rect 45824 4320 45888 4324
rect 45904 4380 45968 4384
rect 45904 4324 45908 4380
rect 45908 4324 45964 4380
rect 45964 4324 45968 4380
rect 45904 4320 45968 4324
rect 6541 3836 6605 3840
rect 6541 3780 6545 3836
rect 6545 3780 6601 3836
rect 6601 3780 6605 3836
rect 6541 3776 6605 3780
rect 6621 3836 6685 3840
rect 6621 3780 6625 3836
rect 6625 3780 6681 3836
rect 6681 3780 6685 3836
rect 6621 3776 6685 3780
rect 6701 3836 6765 3840
rect 6701 3780 6705 3836
rect 6705 3780 6761 3836
rect 6761 3780 6765 3836
rect 6701 3776 6765 3780
rect 6781 3836 6845 3840
rect 6781 3780 6785 3836
rect 6785 3780 6841 3836
rect 6841 3780 6845 3836
rect 6781 3776 6845 3780
rect 17719 3836 17783 3840
rect 17719 3780 17723 3836
rect 17723 3780 17779 3836
rect 17779 3780 17783 3836
rect 17719 3776 17783 3780
rect 17799 3836 17863 3840
rect 17799 3780 17803 3836
rect 17803 3780 17859 3836
rect 17859 3780 17863 3836
rect 17799 3776 17863 3780
rect 17879 3836 17943 3840
rect 17879 3780 17883 3836
rect 17883 3780 17939 3836
rect 17939 3780 17943 3836
rect 17879 3776 17943 3780
rect 17959 3836 18023 3840
rect 17959 3780 17963 3836
rect 17963 3780 18019 3836
rect 18019 3780 18023 3836
rect 17959 3776 18023 3780
rect 28897 3836 28961 3840
rect 28897 3780 28901 3836
rect 28901 3780 28957 3836
rect 28957 3780 28961 3836
rect 28897 3776 28961 3780
rect 28977 3836 29041 3840
rect 28977 3780 28981 3836
rect 28981 3780 29037 3836
rect 29037 3780 29041 3836
rect 28977 3776 29041 3780
rect 29057 3836 29121 3840
rect 29057 3780 29061 3836
rect 29061 3780 29117 3836
rect 29117 3780 29121 3836
rect 29057 3776 29121 3780
rect 29137 3836 29201 3840
rect 29137 3780 29141 3836
rect 29141 3780 29197 3836
rect 29197 3780 29201 3836
rect 29137 3776 29201 3780
rect 40075 3836 40139 3840
rect 40075 3780 40079 3836
rect 40079 3780 40135 3836
rect 40135 3780 40139 3836
rect 40075 3776 40139 3780
rect 40155 3836 40219 3840
rect 40155 3780 40159 3836
rect 40159 3780 40215 3836
rect 40215 3780 40219 3836
rect 40155 3776 40219 3780
rect 40235 3836 40299 3840
rect 40235 3780 40239 3836
rect 40239 3780 40295 3836
rect 40295 3780 40299 3836
rect 40235 3776 40299 3780
rect 40315 3836 40379 3840
rect 40315 3780 40319 3836
rect 40319 3780 40375 3836
rect 40375 3780 40379 3836
rect 40315 3776 40379 3780
rect 12130 3292 12194 3296
rect 12130 3236 12134 3292
rect 12134 3236 12190 3292
rect 12190 3236 12194 3292
rect 12130 3232 12194 3236
rect 12210 3292 12274 3296
rect 12210 3236 12214 3292
rect 12214 3236 12270 3292
rect 12270 3236 12274 3292
rect 12210 3232 12274 3236
rect 12290 3292 12354 3296
rect 12290 3236 12294 3292
rect 12294 3236 12350 3292
rect 12350 3236 12354 3292
rect 12290 3232 12354 3236
rect 12370 3292 12434 3296
rect 12370 3236 12374 3292
rect 12374 3236 12430 3292
rect 12430 3236 12434 3292
rect 12370 3232 12434 3236
rect 23308 3292 23372 3296
rect 23308 3236 23312 3292
rect 23312 3236 23368 3292
rect 23368 3236 23372 3292
rect 23308 3232 23372 3236
rect 23388 3292 23452 3296
rect 23388 3236 23392 3292
rect 23392 3236 23448 3292
rect 23448 3236 23452 3292
rect 23388 3232 23452 3236
rect 23468 3292 23532 3296
rect 23468 3236 23472 3292
rect 23472 3236 23528 3292
rect 23528 3236 23532 3292
rect 23468 3232 23532 3236
rect 23548 3292 23612 3296
rect 23548 3236 23552 3292
rect 23552 3236 23608 3292
rect 23608 3236 23612 3292
rect 23548 3232 23612 3236
rect 34486 3292 34550 3296
rect 34486 3236 34490 3292
rect 34490 3236 34546 3292
rect 34546 3236 34550 3292
rect 34486 3232 34550 3236
rect 34566 3292 34630 3296
rect 34566 3236 34570 3292
rect 34570 3236 34626 3292
rect 34626 3236 34630 3292
rect 34566 3232 34630 3236
rect 34646 3292 34710 3296
rect 34646 3236 34650 3292
rect 34650 3236 34706 3292
rect 34706 3236 34710 3292
rect 34646 3232 34710 3236
rect 34726 3292 34790 3296
rect 34726 3236 34730 3292
rect 34730 3236 34786 3292
rect 34786 3236 34790 3292
rect 34726 3232 34790 3236
rect 45664 3292 45728 3296
rect 45664 3236 45668 3292
rect 45668 3236 45724 3292
rect 45724 3236 45728 3292
rect 45664 3232 45728 3236
rect 45744 3292 45808 3296
rect 45744 3236 45748 3292
rect 45748 3236 45804 3292
rect 45804 3236 45808 3292
rect 45744 3232 45808 3236
rect 45824 3292 45888 3296
rect 45824 3236 45828 3292
rect 45828 3236 45884 3292
rect 45884 3236 45888 3292
rect 45824 3232 45888 3236
rect 45904 3292 45968 3296
rect 45904 3236 45908 3292
rect 45908 3236 45964 3292
rect 45964 3236 45968 3292
rect 45904 3232 45968 3236
rect 6541 2748 6605 2752
rect 6541 2692 6545 2748
rect 6545 2692 6601 2748
rect 6601 2692 6605 2748
rect 6541 2688 6605 2692
rect 6621 2748 6685 2752
rect 6621 2692 6625 2748
rect 6625 2692 6681 2748
rect 6681 2692 6685 2748
rect 6621 2688 6685 2692
rect 6701 2748 6765 2752
rect 6701 2692 6705 2748
rect 6705 2692 6761 2748
rect 6761 2692 6765 2748
rect 6701 2688 6765 2692
rect 6781 2748 6845 2752
rect 6781 2692 6785 2748
rect 6785 2692 6841 2748
rect 6841 2692 6845 2748
rect 6781 2688 6845 2692
rect 17719 2748 17783 2752
rect 17719 2692 17723 2748
rect 17723 2692 17779 2748
rect 17779 2692 17783 2748
rect 17719 2688 17783 2692
rect 17799 2748 17863 2752
rect 17799 2692 17803 2748
rect 17803 2692 17859 2748
rect 17859 2692 17863 2748
rect 17799 2688 17863 2692
rect 17879 2748 17943 2752
rect 17879 2692 17883 2748
rect 17883 2692 17939 2748
rect 17939 2692 17943 2748
rect 17879 2688 17943 2692
rect 17959 2748 18023 2752
rect 17959 2692 17963 2748
rect 17963 2692 18019 2748
rect 18019 2692 18023 2748
rect 17959 2688 18023 2692
rect 28897 2748 28961 2752
rect 28897 2692 28901 2748
rect 28901 2692 28957 2748
rect 28957 2692 28961 2748
rect 28897 2688 28961 2692
rect 28977 2748 29041 2752
rect 28977 2692 28981 2748
rect 28981 2692 29037 2748
rect 29037 2692 29041 2748
rect 28977 2688 29041 2692
rect 29057 2748 29121 2752
rect 29057 2692 29061 2748
rect 29061 2692 29117 2748
rect 29117 2692 29121 2748
rect 29057 2688 29121 2692
rect 29137 2748 29201 2752
rect 29137 2692 29141 2748
rect 29141 2692 29197 2748
rect 29197 2692 29201 2748
rect 29137 2688 29201 2692
rect 40075 2748 40139 2752
rect 40075 2692 40079 2748
rect 40079 2692 40135 2748
rect 40135 2692 40139 2748
rect 40075 2688 40139 2692
rect 40155 2748 40219 2752
rect 40155 2692 40159 2748
rect 40159 2692 40215 2748
rect 40215 2692 40219 2748
rect 40155 2688 40219 2692
rect 40235 2748 40299 2752
rect 40235 2692 40239 2748
rect 40239 2692 40295 2748
rect 40295 2692 40299 2748
rect 40235 2688 40299 2692
rect 40315 2748 40379 2752
rect 40315 2692 40319 2748
rect 40319 2692 40375 2748
rect 40375 2692 40379 2748
rect 40315 2688 40379 2692
rect 12130 2204 12194 2208
rect 12130 2148 12134 2204
rect 12134 2148 12190 2204
rect 12190 2148 12194 2204
rect 12130 2144 12194 2148
rect 12210 2204 12274 2208
rect 12210 2148 12214 2204
rect 12214 2148 12270 2204
rect 12270 2148 12274 2204
rect 12210 2144 12274 2148
rect 12290 2204 12354 2208
rect 12290 2148 12294 2204
rect 12294 2148 12350 2204
rect 12350 2148 12354 2204
rect 12290 2144 12354 2148
rect 12370 2204 12434 2208
rect 12370 2148 12374 2204
rect 12374 2148 12430 2204
rect 12430 2148 12434 2204
rect 12370 2144 12434 2148
rect 23308 2204 23372 2208
rect 23308 2148 23312 2204
rect 23312 2148 23368 2204
rect 23368 2148 23372 2204
rect 23308 2144 23372 2148
rect 23388 2204 23452 2208
rect 23388 2148 23392 2204
rect 23392 2148 23448 2204
rect 23448 2148 23452 2204
rect 23388 2144 23452 2148
rect 23468 2204 23532 2208
rect 23468 2148 23472 2204
rect 23472 2148 23528 2204
rect 23528 2148 23532 2204
rect 23468 2144 23532 2148
rect 23548 2204 23612 2208
rect 23548 2148 23552 2204
rect 23552 2148 23608 2204
rect 23608 2148 23612 2204
rect 23548 2144 23612 2148
rect 34486 2204 34550 2208
rect 34486 2148 34490 2204
rect 34490 2148 34546 2204
rect 34546 2148 34550 2204
rect 34486 2144 34550 2148
rect 34566 2204 34630 2208
rect 34566 2148 34570 2204
rect 34570 2148 34626 2204
rect 34626 2148 34630 2204
rect 34566 2144 34630 2148
rect 34646 2204 34710 2208
rect 34646 2148 34650 2204
rect 34650 2148 34706 2204
rect 34706 2148 34710 2204
rect 34646 2144 34710 2148
rect 34726 2204 34790 2208
rect 34726 2148 34730 2204
rect 34730 2148 34786 2204
rect 34786 2148 34790 2204
rect 34726 2144 34790 2148
rect 45664 2204 45728 2208
rect 45664 2148 45668 2204
rect 45668 2148 45724 2204
rect 45724 2148 45728 2204
rect 45664 2144 45728 2148
rect 45744 2204 45808 2208
rect 45744 2148 45748 2204
rect 45748 2148 45804 2204
rect 45804 2148 45808 2204
rect 45744 2144 45808 2148
rect 45824 2204 45888 2208
rect 45824 2148 45828 2204
rect 45828 2148 45884 2204
rect 45884 2148 45888 2204
rect 45824 2144 45888 2148
rect 45904 2204 45968 2208
rect 45904 2148 45908 2204
rect 45908 2148 45964 2204
rect 45964 2148 45968 2204
rect 45904 2144 45968 2148
rect 6541 1660 6605 1664
rect 6541 1604 6545 1660
rect 6545 1604 6601 1660
rect 6601 1604 6605 1660
rect 6541 1600 6605 1604
rect 6621 1660 6685 1664
rect 6621 1604 6625 1660
rect 6625 1604 6681 1660
rect 6681 1604 6685 1660
rect 6621 1600 6685 1604
rect 6701 1660 6765 1664
rect 6701 1604 6705 1660
rect 6705 1604 6761 1660
rect 6761 1604 6765 1660
rect 6701 1600 6765 1604
rect 6781 1660 6845 1664
rect 6781 1604 6785 1660
rect 6785 1604 6841 1660
rect 6841 1604 6845 1660
rect 6781 1600 6845 1604
rect 17719 1660 17783 1664
rect 17719 1604 17723 1660
rect 17723 1604 17779 1660
rect 17779 1604 17783 1660
rect 17719 1600 17783 1604
rect 17799 1660 17863 1664
rect 17799 1604 17803 1660
rect 17803 1604 17859 1660
rect 17859 1604 17863 1660
rect 17799 1600 17863 1604
rect 17879 1660 17943 1664
rect 17879 1604 17883 1660
rect 17883 1604 17939 1660
rect 17939 1604 17943 1660
rect 17879 1600 17943 1604
rect 17959 1660 18023 1664
rect 17959 1604 17963 1660
rect 17963 1604 18019 1660
rect 18019 1604 18023 1660
rect 17959 1600 18023 1604
rect 28897 1660 28961 1664
rect 28897 1604 28901 1660
rect 28901 1604 28957 1660
rect 28957 1604 28961 1660
rect 28897 1600 28961 1604
rect 28977 1660 29041 1664
rect 28977 1604 28981 1660
rect 28981 1604 29037 1660
rect 29037 1604 29041 1660
rect 28977 1600 29041 1604
rect 29057 1660 29121 1664
rect 29057 1604 29061 1660
rect 29061 1604 29117 1660
rect 29117 1604 29121 1660
rect 29057 1600 29121 1604
rect 29137 1660 29201 1664
rect 29137 1604 29141 1660
rect 29141 1604 29197 1660
rect 29197 1604 29201 1660
rect 29137 1600 29201 1604
rect 40075 1660 40139 1664
rect 40075 1604 40079 1660
rect 40079 1604 40135 1660
rect 40135 1604 40139 1660
rect 40075 1600 40139 1604
rect 40155 1660 40219 1664
rect 40155 1604 40159 1660
rect 40159 1604 40215 1660
rect 40215 1604 40219 1660
rect 40155 1600 40219 1604
rect 40235 1660 40299 1664
rect 40235 1604 40239 1660
rect 40239 1604 40295 1660
rect 40295 1604 40299 1660
rect 40235 1600 40299 1604
rect 40315 1660 40379 1664
rect 40315 1604 40319 1660
rect 40319 1604 40375 1660
rect 40375 1604 40379 1660
rect 40315 1600 40379 1604
rect 12130 1116 12194 1120
rect 12130 1060 12134 1116
rect 12134 1060 12190 1116
rect 12190 1060 12194 1116
rect 12130 1056 12194 1060
rect 12210 1116 12274 1120
rect 12210 1060 12214 1116
rect 12214 1060 12270 1116
rect 12270 1060 12274 1116
rect 12210 1056 12274 1060
rect 12290 1116 12354 1120
rect 12290 1060 12294 1116
rect 12294 1060 12350 1116
rect 12350 1060 12354 1116
rect 12290 1056 12354 1060
rect 12370 1116 12434 1120
rect 12370 1060 12374 1116
rect 12374 1060 12430 1116
rect 12430 1060 12434 1116
rect 12370 1056 12434 1060
rect 23308 1116 23372 1120
rect 23308 1060 23312 1116
rect 23312 1060 23368 1116
rect 23368 1060 23372 1116
rect 23308 1056 23372 1060
rect 23388 1116 23452 1120
rect 23388 1060 23392 1116
rect 23392 1060 23448 1116
rect 23448 1060 23452 1116
rect 23388 1056 23452 1060
rect 23468 1116 23532 1120
rect 23468 1060 23472 1116
rect 23472 1060 23528 1116
rect 23528 1060 23532 1116
rect 23468 1056 23532 1060
rect 23548 1116 23612 1120
rect 23548 1060 23552 1116
rect 23552 1060 23608 1116
rect 23608 1060 23612 1116
rect 23548 1056 23612 1060
rect 34486 1116 34550 1120
rect 34486 1060 34490 1116
rect 34490 1060 34546 1116
rect 34546 1060 34550 1116
rect 34486 1056 34550 1060
rect 34566 1116 34630 1120
rect 34566 1060 34570 1116
rect 34570 1060 34626 1116
rect 34626 1060 34630 1116
rect 34566 1056 34630 1060
rect 34646 1116 34710 1120
rect 34646 1060 34650 1116
rect 34650 1060 34706 1116
rect 34706 1060 34710 1116
rect 34646 1056 34710 1060
rect 34726 1116 34790 1120
rect 34726 1060 34730 1116
rect 34730 1060 34786 1116
rect 34786 1060 34790 1116
rect 34726 1056 34790 1060
rect 45664 1116 45728 1120
rect 45664 1060 45668 1116
rect 45668 1060 45724 1116
rect 45724 1060 45728 1116
rect 45664 1056 45728 1060
rect 45744 1116 45808 1120
rect 45744 1060 45748 1116
rect 45748 1060 45804 1116
rect 45804 1060 45808 1116
rect 45744 1056 45808 1060
rect 45824 1116 45888 1120
rect 45824 1060 45828 1116
rect 45828 1060 45884 1116
rect 45884 1060 45888 1116
rect 45824 1056 45888 1060
rect 45904 1116 45968 1120
rect 45904 1060 45908 1116
rect 45908 1060 45964 1116
rect 45964 1060 45968 1116
rect 45904 1056 45968 1060
<< metal4 >>
rect 20667 9212 20733 9213
rect 20667 9148 20668 9212
rect 20732 9148 20733 9212
rect 20667 9147 20733 9148
rect 6533 8192 6853 8752
rect 6533 8128 6541 8192
rect 6605 8128 6621 8192
rect 6685 8128 6701 8192
rect 6765 8128 6781 8192
rect 6845 8128 6853 8192
rect 6533 7104 6853 8128
rect 6533 7040 6541 7104
rect 6605 7040 6621 7104
rect 6685 7040 6701 7104
rect 6765 7040 6781 7104
rect 6845 7040 6853 7104
rect 6533 6016 6853 7040
rect 6533 5952 6541 6016
rect 6605 5952 6621 6016
rect 6685 5952 6701 6016
rect 6765 5952 6781 6016
rect 6845 5952 6853 6016
rect 6533 4928 6853 5952
rect 6533 4864 6541 4928
rect 6605 4864 6621 4928
rect 6685 4864 6701 4928
rect 6765 4864 6781 4928
rect 6845 4864 6853 4928
rect 6533 3840 6853 4864
rect 6533 3776 6541 3840
rect 6605 3776 6621 3840
rect 6685 3776 6701 3840
rect 6765 3776 6781 3840
rect 6845 3776 6853 3840
rect 6533 2752 6853 3776
rect 6533 2688 6541 2752
rect 6605 2688 6621 2752
rect 6685 2688 6701 2752
rect 6765 2688 6781 2752
rect 6845 2688 6853 2752
rect 6533 1664 6853 2688
rect 6533 1600 6541 1664
rect 6605 1600 6621 1664
rect 6685 1600 6701 1664
rect 6765 1600 6781 1664
rect 6845 1600 6853 1664
rect 6533 1040 6853 1600
rect 12122 8736 12442 8752
rect 12122 8672 12130 8736
rect 12194 8672 12210 8736
rect 12274 8672 12290 8736
rect 12354 8672 12370 8736
rect 12434 8672 12442 8736
rect 12122 7648 12442 8672
rect 12122 7584 12130 7648
rect 12194 7584 12210 7648
rect 12274 7584 12290 7648
rect 12354 7584 12370 7648
rect 12434 7584 12442 7648
rect 12122 6560 12442 7584
rect 12122 6496 12130 6560
rect 12194 6496 12210 6560
rect 12274 6496 12290 6560
rect 12354 6496 12370 6560
rect 12434 6496 12442 6560
rect 12122 5472 12442 6496
rect 12122 5408 12130 5472
rect 12194 5408 12210 5472
rect 12274 5408 12290 5472
rect 12354 5408 12370 5472
rect 12434 5408 12442 5472
rect 12122 4384 12442 5408
rect 12122 4320 12130 4384
rect 12194 4320 12210 4384
rect 12274 4320 12290 4384
rect 12354 4320 12370 4384
rect 12434 4320 12442 4384
rect 12122 3296 12442 4320
rect 12122 3232 12130 3296
rect 12194 3232 12210 3296
rect 12274 3232 12290 3296
rect 12354 3232 12370 3296
rect 12434 3232 12442 3296
rect 12122 2208 12442 3232
rect 12122 2144 12130 2208
rect 12194 2144 12210 2208
rect 12274 2144 12290 2208
rect 12354 2144 12370 2208
rect 12434 2144 12442 2208
rect 12122 1120 12442 2144
rect 12122 1056 12130 1120
rect 12194 1056 12210 1120
rect 12274 1056 12290 1120
rect 12354 1056 12370 1120
rect 12434 1056 12442 1120
rect 12122 1040 12442 1056
rect 17711 8192 18031 8752
rect 17711 8128 17719 8192
rect 17783 8128 17799 8192
rect 17863 8128 17879 8192
rect 17943 8128 17959 8192
rect 18023 8128 18031 8192
rect 17711 7104 18031 8128
rect 20670 7853 20730 9147
rect 23300 8736 23620 8752
rect 23300 8672 23308 8736
rect 23372 8672 23388 8736
rect 23452 8672 23468 8736
rect 23532 8672 23548 8736
rect 23612 8672 23620 8736
rect 20667 7852 20733 7853
rect 20667 7788 20668 7852
rect 20732 7788 20733 7852
rect 20667 7787 20733 7788
rect 17711 7040 17719 7104
rect 17783 7040 17799 7104
rect 17863 7040 17879 7104
rect 17943 7040 17959 7104
rect 18023 7040 18031 7104
rect 17711 6016 18031 7040
rect 17711 5952 17719 6016
rect 17783 5952 17799 6016
rect 17863 5952 17879 6016
rect 17943 5952 17959 6016
rect 18023 5952 18031 6016
rect 17711 4928 18031 5952
rect 17711 4864 17719 4928
rect 17783 4864 17799 4928
rect 17863 4864 17879 4928
rect 17943 4864 17959 4928
rect 18023 4864 18031 4928
rect 17711 3840 18031 4864
rect 17711 3776 17719 3840
rect 17783 3776 17799 3840
rect 17863 3776 17879 3840
rect 17943 3776 17959 3840
rect 18023 3776 18031 3840
rect 17711 2752 18031 3776
rect 17711 2688 17719 2752
rect 17783 2688 17799 2752
rect 17863 2688 17879 2752
rect 17943 2688 17959 2752
rect 18023 2688 18031 2752
rect 17711 1664 18031 2688
rect 17711 1600 17719 1664
rect 17783 1600 17799 1664
rect 17863 1600 17879 1664
rect 17943 1600 17959 1664
rect 18023 1600 18031 1664
rect 17711 1040 18031 1600
rect 23300 7648 23620 8672
rect 23300 7584 23308 7648
rect 23372 7584 23388 7648
rect 23452 7584 23468 7648
rect 23532 7584 23548 7648
rect 23612 7584 23620 7648
rect 23300 6560 23620 7584
rect 23300 6496 23308 6560
rect 23372 6496 23388 6560
rect 23452 6496 23468 6560
rect 23532 6496 23548 6560
rect 23612 6496 23620 6560
rect 23300 5472 23620 6496
rect 23300 5408 23308 5472
rect 23372 5408 23388 5472
rect 23452 5408 23468 5472
rect 23532 5408 23548 5472
rect 23612 5408 23620 5472
rect 23300 4384 23620 5408
rect 23300 4320 23308 4384
rect 23372 4320 23388 4384
rect 23452 4320 23468 4384
rect 23532 4320 23548 4384
rect 23612 4320 23620 4384
rect 23300 3296 23620 4320
rect 23300 3232 23308 3296
rect 23372 3232 23388 3296
rect 23452 3232 23468 3296
rect 23532 3232 23548 3296
rect 23612 3232 23620 3296
rect 23300 2208 23620 3232
rect 23300 2144 23308 2208
rect 23372 2144 23388 2208
rect 23452 2144 23468 2208
rect 23532 2144 23548 2208
rect 23612 2144 23620 2208
rect 23300 1120 23620 2144
rect 23300 1056 23308 1120
rect 23372 1056 23388 1120
rect 23452 1056 23468 1120
rect 23532 1056 23548 1120
rect 23612 1056 23620 1120
rect 23300 1040 23620 1056
rect 28889 8192 29209 8752
rect 28889 8128 28897 8192
rect 28961 8128 28977 8192
rect 29041 8128 29057 8192
rect 29121 8128 29137 8192
rect 29201 8128 29209 8192
rect 28889 7104 29209 8128
rect 28889 7040 28897 7104
rect 28961 7040 28977 7104
rect 29041 7040 29057 7104
rect 29121 7040 29137 7104
rect 29201 7040 29209 7104
rect 28889 6016 29209 7040
rect 28889 5952 28897 6016
rect 28961 5952 28977 6016
rect 29041 5952 29057 6016
rect 29121 5952 29137 6016
rect 29201 5952 29209 6016
rect 28889 4928 29209 5952
rect 28889 4864 28897 4928
rect 28961 4864 28977 4928
rect 29041 4864 29057 4928
rect 29121 4864 29137 4928
rect 29201 4864 29209 4928
rect 28889 3840 29209 4864
rect 28889 3776 28897 3840
rect 28961 3776 28977 3840
rect 29041 3776 29057 3840
rect 29121 3776 29137 3840
rect 29201 3776 29209 3840
rect 28889 2752 29209 3776
rect 28889 2688 28897 2752
rect 28961 2688 28977 2752
rect 29041 2688 29057 2752
rect 29121 2688 29137 2752
rect 29201 2688 29209 2752
rect 28889 1664 29209 2688
rect 28889 1600 28897 1664
rect 28961 1600 28977 1664
rect 29041 1600 29057 1664
rect 29121 1600 29137 1664
rect 29201 1600 29209 1664
rect 28889 1040 29209 1600
rect 34478 8736 34798 8752
rect 34478 8672 34486 8736
rect 34550 8672 34566 8736
rect 34630 8672 34646 8736
rect 34710 8672 34726 8736
rect 34790 8672 34798 8736
rect 34478 7648 34798 8672
rect 34478 7584 34486 7648
rect 34550 7584 34566 7648
rect 34630 7584 34646 7648
rect 34710 7584 34726 7648
rect 34790 7584 34798 7648
rect 34478 6560 34798 7584
rect 34478 6496 34486 6560
rect 34550 6496 34566 6560
rect 34630 6496 34646 6560
rect 34710 6496 34726 6560
rect 34790 6496 34798 6560
rect 34478 5472 34798 6496
rect 34478 5408 34486 5472
rect 34550 5408 34566 5472
rect 34630 5408 34646 5472
rect 34710 5408 34726 5472
rect 34790 5408 34798 5472
rect 34478 4384 34798 5408
rect 34478 4320 34486 4384
rect 34550 4320 34566 4384
rect 34630 4320 34646 4384
rect 34710 4320 34726 4384
rect 34790 4320 34798 4384
rect 34478 3296 34798 4320
rect 34478 3232 34486 3296
rect 34550 3232 34566 3296
rect 34630 3232 34646 3296
rect 34710 3232 34726 3296
rect 34790 3232 34798 3296
rect 34478 2208 34798 3232
rect 34478 2144 34486 2208
rect 34550 2144 34566 2208
rect 34630 2144 34646 2208
rect 34710 2144 34726 2208
rect 34790 2144 34798 2208
rect 34478 1120 34798 2144
rect 34478 1056 34486 1120
rect 34550 1056 34566 1120
rect 34630 1056 34646 1120
rect 34710 1056 34726 1120
rect 34790 1056 34798 1120
rect 34478 1040 34798 1056
rect 40067 8192 40387 8752
rect 40067 8128 40075 8192
rect 40139 8128 40155 8192
rect 40219 8128 40235 8192
rect 40299 8128 40315 8192
rect 40379 8128 40387 8192
rect 40067 7104 40387 8128
rect 40067 7040 40075 7104
rect 40139 7040 40155 7104
rect 40219 7040 40235 7104
rect 40299 7040 40315 7104
rect 40379 7040 40387 7104
rect 40067 6016 40387 7040
rect 40067 5952 40075 6016
rect 40139 5952 40155 6016
rect 40219 5952 40235 6016
rect 40299 5952 40315 6016
rect 40379 5952 40387 6016
rect 40067 4928 40387 5952
rect 40067 4864 40075 4928
rect 40139 4864 40155 4928
rect 40219 4864 40235 4928
rect 40299 4864 40315 4928
rect 40379 4864 40387 4928
rect 40067 3840 40387 4864
rect 40067 3776 40075 3840
rect 40139 3776 40155 3840
rect 40219 3776 40235 3840
rect 40299 3776 40315 3840
rect 40379 3776 40387 3840
rect 40067 2752 40387 3776
rect 40067 2688 40075 2752
rect 40139 2688 40155 2752
rect 40219 2688 40235 2752
rect 40299 2688 40315 2752
rect 40379 2688 40387 2752
rect 40067 1664 40387 2688
rect 40067 1600 40075 1664
rect 40139 1600 40155 1664
rect 40219 1600 40235 1664
rect 40299 1600 40315 1664
rect 40379 1600 40387 1664
rect 40067 1040 40387 1600
rect 45656 8736 45976 8752
rect 45656 8672 45664 8736
rect 45728 8672 45744 8736
rect 45808 8672 45824 8736
rect 45888 8672 45904 8736
rect 45968 8672 45976 8736
rect 45656 7648 45976 8672
rect 45656 7584 45664 7648
rect 45728 7584 45744 7648
rect 45808 7584 45824 7648
rect 45888 7584 45904 7648
rect 45968 7584 45976 7648
rect 45656 6560 45976 7584
rect 45656 6496 45664 6560
rect 45728 6496 45744 6560
rect 45808 6496 45824 6560
rect 45888 6496 45904 6560
rect 45968 6496 45976 6560
rect 45656 5472 45976 6496
rect 45656 5408 45664 5472
rect 45728 5408 45744 5472
rect 45808 5408 45824 5472
rect 45888 5408 45904 5472
rect 45968 5408 45976 5472
rect 45656 4384 45976 5408
rect 45656 4320 45664 4384
rect 45728 4320 45744 4384
rect 45808 4320 45824 4384
rect 45888 4320 45904 4384
rect 45968 4320 45976 4384
rect 45656 3296 45976 4320
rect 45656 3232 45664 3296
rect 45728 3232 45744 3296
rect 45808 3232 45824 3296
rect 45888 3232 45904 3296
rect 45968 3232 45976 3296
rect 45656 2208 45976 3232
rect 45656 2144 45664 2208
rect 45728 2144 45744 2208
rect 45808 2144 45824 2208
rect 45888 2144 45904 2208
rect 45968 2144 45976 2208
rect 45656 1120 45976 2144
rect 45656 1056 45664 1120
rect 45728 1056 45744 1120
rect 45808 1056 45824 1120
rect 45888 1056 45904 1120
rect 45968 1056 45976 1120
rect 45656 1040 45976 1056
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 2024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_7 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1748 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1688980957
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_32
timestamp 1688980957
transform 1 0 4048 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_44
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_69 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_75
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_79 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8372 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_97 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_103
timestamp 1688980957
transform 1 0 10580 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_121
timestamp 1688980957
transform 1 0 12236 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_127
timestamp 1688980957
transform 1 0 12788 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_147
timestamp 1688980957
transform 1 0 14628 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_151
timestamp 1688980957
transform 1 0 14996 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_163
timestamp 1688980957
transform 1 0 16100 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1688980957
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_175
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_187
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1688980957
transform 1 0 19044 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_200
timestamp 1688980957
transform 1 0 19504 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_212
timestamp 1688980957
transform 1 0 20608 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_243
timestamp 1688980957
transform 1 0 23460 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_247
timestamp 1688980957
transform 1 0 23828 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_271
timestamp 1688980957
transform 1 0 26036 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_289
timestamp 1688980957
transform 1 0 27692 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_295
timestamp 1688980957
transform 1 0 28244 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_315
timestamp 1688980957
transform 1 0 30084 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_319
timestamp 1688980957
transform 1 0 30452 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_331
timestamp 1688980957
transform 1 0 31556 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1688980957
transform 1 0 31924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_343
timestamp 1688980957
transform 1 0 32660 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_355
timestamp 1688980957
transform 1 0 33764 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_363
timestamp 1688980957
transform 1 0 34500 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_368
timestamp 1688980957
transform 1 0 34960 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_380
timestamp 1688980957
transform 1 0 36064 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_391
timestamp 1688980957
transform 1 0 37076 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_405
timestamp 1688980957
transform 1 0 38364 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_411
timestamp 1688980957
transform 1 0 38916 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_415
timestamp 1688980957
transform 1 0 39284 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_419
timestamp 1688980957
transform 1 0 39652 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_439
timestamp 1688980957
transform 1 0 41492 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_447
timestamp 1688980957
transform 1 0 42228 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_457
timestamp 1688980957
transform 1 0 43148 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_463
timestamp 1688980957
transform 1 0 43700 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_475
timestamp 1688980957
transform 1 0 44804 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_477
timestamp 1688980957
transform 1 0 44988 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_204
timestamp 1688980957
transform 1 0 19872 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_216
timestamp 1688980957
transform 1 0 20976 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_236 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22816 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_244
timestamp 1688980957
transform 1 0 23552 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_250
timestamp 1688980957
transform 1 0 24104 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_254
timestamp 1688980957
transform 1 0 24472 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_266
timestamp 1688980957
transform 1 0 25576 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_278
timestamp 1688980957
transform 1 0 26680 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_326
timestamp 1688980957
transform 1 0 31096 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_334
timestamp 1688980957
transform 1 0 31832 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_396
timestamp 1688980957
transform 1 0 37536 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_408
timestamp 1688980957
transform 1 0 38640 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_420
timestamp 1688980957
transform 1 0 39744 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_432
timestamp 1688980957
transform 1 0 40848 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_440
timestamp 1688980957
transform 1 0 41584 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_445
timestamp 1688980957
transform 1 0 42044 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_461
timestamp 1688980957
transform 1 0 43516 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_468
timestamp 1688980957
transform 1 0 44160 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_472
timestamp 1688980957
transform 1 0 44528 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_476
timestamp 1688980957
transform 1 0 44896 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_482
timestamp 1688980957
transform 1 0 45448 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_215
timestamp 1688980957
transform 1 0 20884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_227
timestamp 1688980957
transform 1 0 21988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_241
timestamp 1688980957
transform 1 0 23276 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 1688980957
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_257
timestamp 1688980957
transform 1 0 24748 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_261
timestamp 1688980957
transform 1 0 25116 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_273
timestamp 1688980957
transform 1 0 26220 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_285
timestamp 1688980957
transform 1 0 27324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_297
timestamp 1688980957
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_302
timestamp 1688980957
transform 1 0 28888 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_329
timestamp 1688980957
transform 1 0 31372 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_406
timestamp 1688980957
transform 1 0 38456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_418
timestamp 1688980957
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_469
timestamp 1688980957
transform 1 0 44252 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_247
timestamp 1688980957
transform 1 0 23828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_259
timestamp 1688980957
transform 1 0 24932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_271
timestamp 1688980957
transform 1 0 26036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_278
timestamp 1688980957
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_309
timestamp 1688980957
transform 1 0 29532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_321
timestamp 1688980957
transform 1 0 30636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_333
timestamp 1688980957
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_421
timestamp 1688980957
transform 1 0 39836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_433
timestamp 1688980957
transform 1 0 40940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_445
timestamp 1688980957
transform 1 0 42044 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_473
timestamp 1688980957
transform 1 0 44620 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_481
timestamp 1688980957
transform 1 0 45356 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_230
timestamp 1688980957
transform 1 0 22264 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_242
timestamp 1688980957
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_246
timestamp 1688980957
transform 1 0 23736 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1688980957
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_350
timestamp 1688980957
transform 1 0 33304 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_362
timestamp 1688980957
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1688980957
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_477
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_233
timestamp 1688980957
transform 1 0 22540 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_240
timestamp 1688980957
transform 1 0 23184 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_244
timestamp 1688980957
transform 1 0 23552 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_248
timestamp 1688980957
transform 1 0 23920 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_260
timestamp 1688980957
transform 1 0 25024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_272
timestamp 1688980957
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_285
timestamp 1688980957
transform 1 0 27324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_297
timestamp 1688980957
transform 1 0 28428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_309
timestamp 1688980957
transform 1 0 29532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_321
timestamp 1688980957
transform 1 0 30636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_333
timestamp 1688980957
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_353
timestamp 1688980957
transform 1 0 33580 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_357
timestamp 1688980957
transform 1 0 33948 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_369
timestamp 1688980957
transform 1 0 35052 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_374
timestamp 1688980957
transform 1 0 35512 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_386
timestamp 1688980957
transform 1 0 36616 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_469
timestamp 1688980957
transform 1 0 44252 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_473
timestamp 1688980957
transform 1 0 44620 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_481
timestamp 1688980957
transform 1 0 45356 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_241
timestamp 1688980957
transform 1 0 23276 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_247
timestamp 1688980957
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_381
timestamp 1688980957
transform 1 0 36156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_393
timestamp 1688980957
transform 1 0 37260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_405
timestamp 1688980957
transform 1 0 38364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_417
timestamp 1688980957
transform 1 0 39468 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_469
timestamp 1688980957
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 1688980957
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_473
timestamp 1688980957
transform 1 0 44620 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_481
timestamp 1688980957
transform 1 0 45356 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 1688980957
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_477
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_473
timestamp 1688980957
transform 1 0 44620 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_481
timestamp 1688980957
transform 1 0 45356 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_240
timestamp 1688980957
transform 1 0 23184 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_469
timestamp 1688980957
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 1688980957
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_13
timestamp 1688980957
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_25
timestamp 1688980957
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_37
timestamp 1688980957
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_49
timestamp 1688980957
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_199
timestamp 1688980957
transform 1 0 19412 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_203
timestamp 1688980957
transform 1 0 19780 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_207
timestamp 1688980957
transform 1 0 20148 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_215
timestamp 1688980957
transform 1 0 20884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_219
timestamp 1688980957
transform 1 0 21252 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_243
timestamp 1688980957
transform 1 0 23460 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_251
timestamp 1688980957
transform 1 0 24196 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_263
timestamp 1688980957
transform 1 0 25300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_275
timestamp 1688980957
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_461
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_481
timestamp 1688980957
transform 1 0 45356 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_22
timestamp 1688980957
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_40
timestamp 1688980957
transform 1 0 4784 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_52
timestamp 1688980957
transform 1 0 5888 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_68
timestamp 1688980957
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 1688980957
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_92
timestamp 1688980957
transform 1 0 9568 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_100
timestamp 1688980957
transform 1 0 10304 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_112
timestamp 1688980957
transform 1 0 11408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_120
timestamp 1688980957
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_128
timestamp 1688980957
transform 1 0 12880 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_148
timestamp 1688980957
transform 1 0 14720 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_160
timestamp 1688980957
transform 1 0 15824 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_172
timestamp 1688980957
transform 1 0 16928 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_178
timestamp 1688980957
transform 1 0 17480 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_192
timestamp 1688980957
transform 1 0 18768 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_279
timestamp 1688980957
transform 1 0 26772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_283
timestamp 1688980957
transform 1 0 27140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_287
timestamp 1688980957
transform 1 0 27508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_291
timestamp 1688980957
transform 1 0 27876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_295
timestamp 1688980957
transform 1 0 28244 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_299
timestamp 1688980957
transform 1 0 28612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_303
timestamp 1688980957
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_437
timestamp 1688980957
transform 1 0 41308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_449
timestamp 1688980957
transform 1 0 42412 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_461
timestamp 1688980957
transform 1 0 43516 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_474
timestamp 1688980957
transform 1 0 44712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_8
timestamp 1688980957
transform 1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_12
timestamp 1688980957
transform 1 0 2208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_46
timestamp 1688980957
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_50
timestamp 1688980957
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_64
timestamp 1688980957
transform 1 0 6992 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_124
timestamp 1688980957
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_156
timestamp 1688980957
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_190
timestamp 1688980957
transform 1 0 18584 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_197
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_210
timestamp 1688980957
transform 1 0 20424 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_250
timestamp 1688980957
transform 1 0 24104 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_259
timestamp 1688980957
transform 1 0 24932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_263
timestamp 1688980957
transform 1 0 25300 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_267
timestamp 1688980957
transform 1 0 25668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_271
timestamp 1688980957
transform 1 0 26036 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_275
timestamp 1688980957
transform 1 0 26404 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_287
timestamp 1688980957
transform 1 0 27508 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_291
timestamp 1688980957
transform 1 0 27876 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_295
timestamp 1688980957
transform 1 0 28244 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_299
timestamp 1688980957
transform 1 0 28612 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_303
timestamp 1688980957
transform 1 0 28980 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_307
timestamp 1688980957
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_315
timestamp 1688980957
transform 1 0 30084 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_319
timestamp 1688980957
transform 1 0 30452 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_323
timestamp 1688980957
transform 1 0 30820 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_327
timestamp 1688980957
transform 1 0 31188 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_331
timestamp 1688980957
transform 1 0 31556 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_343
timestamp 1688980957
transform 1 0 32660 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_347
timestamp 1688980957
transform 1 0 33028 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_351
timestamp 1688980957
transform 1 0 33396 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_355
timestamp 1688980957
transform 1 0 33764 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_359
timestamp 1688980957
transform 1 0 34132 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_363
timestamp 1688980957
transform 1 0 34500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_371
timestamp 1688980957
transform 1 0 35236 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_375
timestamp 1688980957
transform 1 0 35604 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_379
timestamp 1688980957
transform 1 0 35972 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_383
timestamp 1688980957
transform 1 0 36340 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_387
timestamp 1688980957
transform 1 0 36708 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_399
timestamp 1688980957
transform 1 0 37812 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_403
timestamp 1688980957
transform 1 0 38180 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_407
timestamp 1688980957
transform 1 0 38548 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_411
timestamp 1688980957
transform 1 0 38916 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1688980957
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_475
timestamp 1688980957
transform 1 0 44804 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25760 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 27968 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 30176 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 32384 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 34684 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 36800 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 39008 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 41216 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 43424 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 45264 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 5888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 8096 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 10304 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 12512 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 14720 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 16928 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 21344 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 23552 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 19872 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 20332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 22172 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 22724 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 23276 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 25024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 25392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 25760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 26128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 26496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 27232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 30912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 31280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 31648 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 32752 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 27600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform 1 0 27968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 28336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 28704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 29072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 29532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 29808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 30176 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 30544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform 1 0 33120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1688980957
transform 1 0 36800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1688980957
transform 1 0 37536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform 1 0 37904 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1688980957
transform 1 0 38272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1688980957
transform 1 0 38640 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1688980957
transform 1 0 33488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1688980957
transform 1 0 33856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1688980957
transform 1 0 34224 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1688980957
transform 1 0 34684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1688980957
transform 1 0 34960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1688980957
transform 1 0 35328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1688980957
transform 1 0 35696 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1688980957
transform 1 0 36064 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1688980957
transform 1 0 36432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1688980957
transform 1 0 1472 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22448 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__00_
timestamp 1688980957
transform 1 0 26220 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__01_
timestamp 1688980957
transform 1 0 25944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__02_
timestamp 1688980957
transform 1 0 25668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__03_
timestamp 1688980957
transform 1 0 25392 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__04_
timestamp 1688980957
transform 1 0 24840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__05_
timestamp 1688980957
transform 1 0 25116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__06_
timestamp 1688980957
transform 1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__07_
timestamp 1688980957
transform 1 0 23552 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__08_
timestamp 1688980957
transform 1 0 22356 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__09_
timestamp 1688980957
transform 1 0 22356 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__10_
timestamp 1688980957
transform 1 0 21528 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__11_
timestamp 1688980957
transform 1 0 22080 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__12_
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__13_
timestamp 1688980957
transform 1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__14_
timestamp 1688980957
transform 1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__15_
timestamp 1688980957
transform 1 0 20424 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__16_
timestamp 1688980957
transform 1 0 22632 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__17_
timestamp 1688980957
transform 1 0 22908 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__18_
timestamp 1688980957
transform 1 0 28336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__19_
timestamp 1688980957
transform 1 0 27968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__20_
timestamp 1688980957
transform 1 0 27600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__21_
timestamp 1688980957
transform 1 0 27232 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__22_
timestamp 1688980957
transform 1 0 26864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__23_
timestamp 1688980957
transform 1 0 26496 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__24_
timestamp 1688980957
transform 1 0 23644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__25_
timestamp 1688980957
transform 1 0 23184 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__26_
timestamp 1688980957
transform 1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__27_
timestamp 1688980957
transform 1 0 23828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__28_
timestamp 1688980957
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__29_
timestamp 1688980957
transform 1 0 23736 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__30_
timestamp 1688980957
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__31_
timestamp 1688980957
transform 1 0 28704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__32_
timestamp 1688980957
transform 1 0 23000 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__33_
timestamp 1688980957
transform 1 0 22080 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__34_
timestamp 1688980957
transform 1 0 17848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__35_
timestamp 1688980957
transform 1 0 17572 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__36_
timestamp 1688980957
transform 1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__37_
timestamp 1688980957
transform 1 0 19136 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__38_
timestamp 1688980957
transform 1 0 19504 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__39_
timestamp 1688980957
transform 1 0 19596 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__40_
timestamp 1688980957
transform 1 0 23184 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__41_
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__42_
timestamp 1688980957
transform 1 0 22448 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__43_
timestamp 1688980957
transform 1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__44_
timestamp 1688980957
transform 1 0 22908 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__45_
timestamp 1688980957
transform 1 0 21804 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__46_
timestamp 1688980957
transform 1 0 21252 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__47_
timestamp 1688980957
transform 1 0 20976 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__48_
timestamp 1688980957
transform 1 0 20148 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__49_
timestamp 1688980957
transform 1 0 19872 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__50_
timestamp 1688980957
transform 1 0 19320 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__51_
timestamp 1688980957
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39376 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1688980957
transform 1 0 43884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1688980957
transform 1 0 43884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output77 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44252 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 44988 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 44988 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 44252 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 44804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 44160 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 43608 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 39836 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 40388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1688980957
transform 1 0 40940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 41308 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1688980957
transform 1 0 41860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 42780 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 43332 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 1656 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output96
timestamp 1688980957
transform 1 0 2208 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1688980957
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1688980957
transform 1 0 1472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 2392 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform 1 0 2944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1688980957
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 3864 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 3864 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1688980957
transform 1 0 4416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1688980957
transform 1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 4784 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 5336 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1688980957
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 6440 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 6440 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1688980957
transform 1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1688980957
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1688980957
transform 1 0 7544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 11592 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1688980957
transform 1 0 11592 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 11960 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1688980957
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1688980957
transform 1 0 12696 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1688980957
transform 1 0 13064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 7912 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1688980957
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 9016 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1688980957
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1688980957
transform 1 0 9936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1688980957
transform 1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 10304 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1688980957
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 18032 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1688980957
transform 1 0 18400 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1688980957
transform 1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 19872 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 19320 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 14168 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1688980957
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1688980957
transform 1 0 14536 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1688980957
transform 1 0 15456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1688980957
transform 1 0 15640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1688980957
transform 1 0 16928 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1688980957
transform 1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1688980957
transform 1 0 39008 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 45816 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 45816 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 45816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 45816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 45816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 45816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 45816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 45816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 45816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 45816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 45816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 45816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 45816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 45816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 23000 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform 1 0 23276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform 1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform 1 0 22724 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 23276 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 22172 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform 1 0 19596 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 21988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 24196 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 26404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 30820 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 33028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 35236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 37260 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 39560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 41768 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 43884 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 44620 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 23552 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 23644 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 23368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 20516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 27048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 29256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 31464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 33672 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 35880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 44344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 44896 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 37168 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 44896 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 3606 0 3662 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 25686 0 25742 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 27894 0 27950 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 30102 0 30158 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 32310 0 32366 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 34518 0 34574 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 36726 0 36782 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 38934 0 38990 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 41142 0 41198 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 43350 0 43406 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 45558 0 45614 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 5814 0 5870 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 8022 0 8078 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 10230 0 10286 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 12438 0 12494 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 14646 0 14702 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 16854 0 16910 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 19062 0 19118 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 21270 0 21326 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 23478 0 23534 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 39302 9840 39358 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 42982 9840 43038 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 43350 9840 43406 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 43718 9840 43774 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 44086 9840 44142 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 44454 9840 44510 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 44822 9840 44878 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 45190 9840 45246 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 45558 9840 45614 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 45926 9840 45982 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 46294 9840 46350 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 39670 9840 39726 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 40038 9840 40094 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 40406 9840 40462 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 40774 9840 40830 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 41142 9840 41198 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 41510 9840 41566 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 41878 9840 41934 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 42246 9840 42302 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 42614 9840 42670 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 662 9840 718 10000 0 FreeSans 224 90 0 0 N1BEG[0]
port 40 nsew signal tristate
flabel metal2 s 1030 9840 1086 10000 0 FreeSans 224 90 0 0 N1BEG[1]
port 41 nsew signal tristate
flabel metal2 s 1398 9840 1454 10000 0 FreeSans 224 90 0 0 N1BEG[2]
port 42 nsew signal tristate
flabel metal2 s 1766 9840 1822 10000 0 FreeSans 224 90 0 0 N1BEG[3]
port 43 nsew signal tristate
flabel metal2 s 2134 9840 2190 10000 0 FreeSans 224 90 0 0 N2BEG[0]
port 44 nsew signal tristate
flabel metal2 s 2502 9840 2558 10000 0 FreeSans 224 90 0 0 N2BEG[1]
port 45 nsew signal tristate
flabel metal2 s 2870 9840 2926 10000 0 FreeSans 224 90 0 0 N2BEG[2]
port 46 nsew signal tristate
flabel metal2 s 3238 9840 3294 10000 0 FreeSans 224 90 0 0 N2BEG[3]
port 47 nsew signal tristate
flabel metal2 s 3606 9840 3662 10000 0 FreeSans 224 90 0 0 N2BEG[4]
port 48 nsew signal tristate
flabel metal2 s 3974 9840 4030 10000 0 FreeSans 224 90 0 0 N2BEG[5]
port 49 nsew signal tristate
flabel metal2 s 4342 9840 4398 10000 0 FreeSans 224 90 0 0 N2BEG[6]
port 50 nsew signal tristate
flabel metal2 s 4710 9840 4766 10000 0 FreeSans 224 90 0 0 N2BEG[7]
port 51 nsew signal tristate
flabel metal2 s 5078 9840 5134 10000 0 FreeSans 224 90 0 0 N2BEGb[0]
port 52 nsew signal tristate
flabel metal2 s 5446 9840 5502 10000 0 FreeSans 224 90 0 0 N2BEGb[1]
port 53 nsew signal tristate
flabel metal2 s 5814 9840 5870 10000 0 FreeSans 224 90 0 0 N2BEGb[2]
port 54 nsew signal tristate
flabel metal2 s 6182 9840 6238 10000 0 FreeSans 224 90 0 0 N2BEGb[3]
port 55 nsew signal tristate
flabel metal2 s 6550 9840 6606 10000 0 FreeSans 224 90 0 0 N2BEGb[4]
port 56 nsew signal tristate
flabel metal2 s 6918 9840 6974 10000 0 FreeSans 224 90 0 0 N2BEGb[5]
port 57 nsew signal tristate
flabel metal2 s 7286 9840 7342 10000 0 FreeSans 224 90 0 0 N2BEGb[6]
port 58 nsew signal tristate
flabel metal2 s 7654 9840 7710 10000 0 FreeSans 224 90 0 0 N2BEGb[7]
port 59 nsew signal tristate
flabel metal2 s 8022 9840 8078 10000 0 FreeSans 224 90 0 0 N4BEG[0]
port 60 nsew signal tristate
flabel metal2 s 11702 9840 11758 10000 0 FreeSans 224 90 0 0 N4BEG[10]
port 61 nsew signal tristate
flabel metal2 s 12070 9840 12126 10000 0 FreeSans 224 90 0 0 N4BEG[11]
port 62 nsew signal tristate
flabel metal2 s 12438 9840 12494 10000 0 FreeSans 224 90 0 0 N4BEG[12]
port 63 nsew signal tristate
flabel metal2 s 12806 9840 12862 10000 0 FreeSans 224 90 0 0 N4BEG[13]
port 64 nsew signal tristate
flabel metal2 s 13174 9840 13230 10000 0 FreeSans 224 90 0 0 N4BEG[14]
port 65 nsew signal tristate
flabel metal2 s 13542 9840 13598 10000 0 FreeSans 224 90 0 0 N4BEG[15]
port 66 nsew signal tristate
flabel metal2 s 8390 9840 8446 10000 0 FreeSans 224 90 0 0 N4BEG[1]
port 67 nsew signal tristate
flabel metal2 s 8758 9840 8814 10000 0 FreeSans 224 90 0 0 N4BEG[2]
port 68 nsew signal tristate
flabel metal2 s 9126 9840 9182 10000 0 FreeSans 224 90 0 0 N4BEG[3]
port 69 nsew signal tristate
flabel metal2 s 9494 9840 9550 10000 0 FreeSans 224 90 0 0 N4BEG[4]
port 70 nsew signal tristate
flabel metal2 s 9862 9840 9918 10000 0 FreeSans 224 90 0 0 N4BEG[5]
port 71 nsew signal tristate
flabel metal2 s 10230 9840 10286 10000 0 FreeSans 224 90 0 0 N4BEG[6]
port 72 nsew signal tristate
flabel metal2 s 10598 9840 10654 10000 0 FreeSans 224 90 0 0 N4BEG[7]
port 73 nsew signal tristate
flabel metal2 s 10966 9840 11022 10000 0 FreeSans 224 90 0 0 N4BEG[8]
port 74 nsew signal tristate
flabel metal2 s 11334 9840 11390 10000 0 FreeSans 224 90 0 0 N4BEG[9]
port 75 nsew signal tristate
flabel metal2 s 13910 9840 13966 10000 0 FreeSans 224 90 0 0 NN4BEG[0]
port 76 nsew signal tristate
flabel metal2 s 17590 9840 17646 10000 0 FreeSans 224 90 0 0 NN4BEG[10]
port 77 nsew signal tristate
flabel metal2 s 17958 9840 18014 10000 0 FreeSans 224 90 0 0 NN4BEG[11]
port 78 nsew signal tristate
flabel metal2 s 18326 9840 18382 10000 0 FreeSans 224 90 0 0 NN4BEG[12]
port 79 nsew signal tristate
flabel metal2 s 18694 9840 18750 10000 0 FreeSans 224 90 0 0 NN4BEG[13]
port 80 nsew signal tristate
flabel metal2 s 19062 9840 19118 10000 0 FreeSans 224 90 0 0 NN4BEG[14]
port 81 nsew signal tristate
flabel metal2 s 19430 9840 19486 10000 0 FreeSans 224 90 0 0 NN4BEG[15]
port 82 nsew signal tristate
flabel metal2 s 14278 9840 14334 10000 0 FreeSans 224 90 0 0 NN4BEG[1]
port 83 nsew signal tristate
flabel metal2 s 14646 9840 14702 10000 0 FreeSans 224 90 0 0 NN4BEG[2]
port 84 nsew signal tristate
flabel metal2 s 15014 9840 15070 10000 0 FreeSans 224 90 0 0 NN4BEG[3]
port 85 nsew signal tristate
flabel metal2 s 15382 9840 15438 10000 0 FreeSans 224 90 0 0 NN4BEG[4]
port 86 nsew signal tristate
flabel metal2 s 15750 9840 15806 10000 0 FreeSans 224 90 0 0 NN4BEG[5]
port 87 nsew signal tristate
flabel metal2 s 16118 9840 16174 10000 0 FreeSans 224 90 0 0 NN4BEG[6]
port 88 nsew signal tristate
flabel metal2 s 16486 9840 16542 10000 0 FreeSans 224 90 0 0 NN4BEG[7]
port 89 nsew signal tristate
flabel metal2 s 16854 9840 16910 10000 0 FreeSans 224 90 0 0 NN4BEG[8]
port 90 nsew signal tristate
flabel metal2 s 17222 9840 17278 10000 0 FreeSans 224 90 0 0 NN4BEG[9]
port 91 nsew signal tristate
flabel metal2 s 19798 9840 19854 10000 0 FreeSans 224 90 0 0 S1END[0]
port 92 nsew signal input
flabel metal2 s 20166 9840 20222 10000 0 FreeSans 224 90 0 0 S1END[1]
port 93 nsew signal input
flabel metal2 s 20534 9840 20590 10000 0 FreeSans 224 90 0 0 S1END[2]
port 94 nsew signal input
flabel metal2 s 20902 9840 20958 10000 0 FreeSans 224 90 0 0 S1END[3]
port 95 nsew signal input
flabel metal2 s 21270 9840 21326 10000 0 FreeSans 224 90 0 0 S2END[0]
port 96 nsew signal input
flabel metal2 s 21638 9840 21694 10000 0 FreeSans 224 90 0 0 S2END[1]
port 97 nsew signal input
flabel metal2 s 22006 9840 22062 10000 0 FreeSans 224 90 0 0 S2END[2]
port 98 nsew signal input
flabel metal2 s 22374 9840 22430 10000 0 FreeSans 224 90 0 0 S2END[3]
port 99 nsew signal input
flabel metal2 s 22742 9840 22798 10000 0 FreeSans 224 90 0 0 S2END[4]
port 100 nsew signal input
flabel metal2 s 23110 9840 23166 10000 0 FreeSans 224 90 0 0 S2END[5]
port 101 nsew signal input
flabel metal2 s 23478 9840 23534 10000 0 FreeSans 224 90 0 0 S2END[6]
port 102 nsew signal input
flabel metal2 s 23846 9840 23902 10000 0 FreeSans 224 90 0 0 S2END[7]
port 103 nsew signal input
flabel metal2 s 24214 9840 24270 10000 0 FreeSans 224 90 0 0 S2MID[0]
port 104 nsew signal input
flabel metal2 s 24582 9840 24638 10000 0 FreeSans 224 90 0 0 S2MID[1]
port 105 nsew signal input
flabel metal2 s 24950 9840 25006 10000 0 FreeSans 224 90 0 0 S2MID[2]
port 106 nsew signal input
flabel metal2 s 25318 9840 25374 10000 0 FreeSans 224 90 0 0 S2MID[3]
port 107 nsew signal input
flabel metal2 s 25686 9840 25742 10000 0 FreeSans 224 90 0 0 S2MID[4]
port 108 nsew signal input
flabel metal2 s 26054 9840 26110 10000 0 FreeSans 224 90 0 0 S2MID[5]
port 109 nsew signal input
flabel metal2 s 26422 9840 26478 10000 0 FreeSans 224 90 0 0 S2MID[6]
port 110 nsew signal input
flabel metal2 s 26790 9840 26846 10000 0 FreeSans 224 90 0 0 S2MID[7]
port 111 nsew signal input
flabel metal2 s 27158 9840 27214 10000 0 FreeSans 224 90 0 0 S4END[0]
port 112 nsew signal input
flabel metal2 s 30838 9840 30894 10000 0 FreeSans 224 90 0 0 S4END[10]
port 113 nsew signal input
flabel metal2 s 31206 9840 31262 10000 0 FreeSans 224 90 0 0 S4END[11]
port 114 nsew signal input
flabel metal2 s 31574 9840 31630 10000 0 FreeSans 224 90 0 0 S4END[12]
port 115 nsew signal input
flabel metal2 s 31942 9840 31998 10000 0 FreeSans 224 90 0 0 S4END[13]
port 116 nsew signal input
flabel metal2 s 32310 9840 32366 10000 0 FreeSans 224 90 0 0 S4END[14]
port 117 nsew signal input
flabel metal2 s 32678 9840 32734 10000 0 FreeSans 224 90 0 0 S4END[15]
port 118 nsew signal input
flabel metal2 s 27526 9840 27582 10000 0 FreeSans 224 90 0 0 S4END[1]
port 119 nsew signal input
flabel metal2 s 27894 9840 27950 10000 0 FreeSans 224 90 0 0 S4END[2]
port 120 nsew signal input
flabel metal2 s 28262 9840 28318 10000 0 FreeSans 224 90 0 0 S4END[3]
port 121 nsew signal input
flabel metal2 s 28630 9840 28686 10000 0 FreeSans 224 90 0 0 S4END[4]
port 122 nsew signal input
flabel metal2 s 28998 9840 29054 10000 0 FreeSans 224 90 0 0 S4END[5]
port 123 nsew signal input
flabel metal2 s 29366 9840 29422 10000 0 FreeSans 224 90 0 0 S4END[6]
port 124 nsew signal input
flabel metal2 s 29734 9840 29790 10000 0 FreeSans 224 90 0 0 S4END[7]
port 125 nsew signal input
flabel metal2 s 30102 9840 30158 10000 0 FreeSans 224 90 0 0 S4END[8]
port 126 nsew signal input
flabel metal2 s 30470 9840 30526 10000 0 FreeSans 224 90 0 0 S4END[9]
port 127 nsew signal input
flabel metal2 s 33046 9840 33102 10000 0 FreeSans 224 90 0 0 SS4END[0]
port 128 nsew signal input
flabel metal2 s 36726 9840 36782 10000 0 FreeSans 224 90 0 0 SS4END[10]
port 129 nsew signal input
flabel metal2 s 37094 9840 37150 10000 0 FreeSans 224 90 0 0 SS4END[11]
port 130 nsew signal input
flabel metal2 s 37462 9840 37518 10000 0 FreeSans 224 90 0 0 SS4END[12]
port 131 nsew signal input
flabel metal2 s 37830 9840 37886 10000 0 FreeSans 224 90 0 0 SS4END[13]
port 132 nsew signal input
flabel metal2 s 38198 9840 38254 10000 0 FreeSans 224 90 0 0 SS4END[14]
port 133 nsew signal input
flabel metal2 s 38566 9840 38622 10000 0 FreeSans 224 90 0 0 SS4END[15]
port 134 nsew signal input
flabel metal2 s 33414 9840 33470 10000 0 FreeSans 224 90 0 0 SS4END[1]
port 135 nsew signal input
flabel metal2 s 33782 9840 33838 10000 0 FreeSans 224 90 0 0 SS4END[2]
port 136 nsew signal input
flabel metal2 s 34150 9840 34206 10000 0 FreeSans 224 90 0 0 SS4END[3]
port 137 nsew signal input
flabel metal2 s 34518 9840 34574 10000 0 FreeSans 224 90 0 0 SS4END[4]
port 138 nsew signal input
flabel metal2 s 34886 9840 34942 10000 0 FreeSans 224 90 0 0 SS4END[5]
port 139 nsew signal input
flabel metal2 s 35254 9840 35310 10000 0 FreeSans 224 90 0 0 SS4END[6]
port 140 nsew signal input
flabel metal2 s 35622 9840 35678 10000 0 FreeSans 224 90 0 0 SS4END[7]
port 141 nsew signal input
flabel metal2 s 35990 9840 36046 10000 0 FreeSans 224 90 0 0 SS4END[8]
port 142 nsew signal input
flabel metal2 s 36358 9840 36414 10000 0 FreeSans 224 90 0 0 SS4END[9]
port 143 nsew signal input
flabel metal2 s 1398 0 1454 160 0 FreeSans 224 90 0 0 UserCLK
port 144 nsew signal input
flabel metal2 s 38934 9840 38990 10000 0 FreeSans 224 90 0 0 UserCLKo
port 145 nsew signal tristate
flabel metal4 s 6533 1040 6853 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 17711 1040 18031 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 28889 1040 29209 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 40067 1040 40387 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 12122 1040 12442 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 23300 1040 23620 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 34478 1040 34798 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 45656 1040 45976 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
rlabel metal1 23460 8160 23460 8160 0 vccd1
rlabel via1 23540 8704 23540 8704 0 vssd1
rlabel metal2 3733 68 3733 68 0 FrameStrobe[0]
rlabel metal2 25859 68 25859 68 0 FrameStrobe[10]
rlabel metal2 28067 68 28067 68 0 FrameStrobe[11]
rlabel metal2 30275 68 30275 68 0 FrameStrobe[12]
rlabel metal2 32483 68 32483 68 0 FrameStrobe[13]
rlabel metal2 34737 68 34737 68 0 FrameStrobe[14]
rlabel metal2 36899 68 36899 68 0 FrameStrobe[15]
rlabel metal2 39107 68 39107 68 0 FrameStrobe[16]
rlabel metal2 41315 68 41315 68 0 FrameStrobe[17]
rlabel metal2 43523 68 43523 68 0 FrameStrobe[18]
rlabel metal2 45586 704 45586 704 0 FrameStrobe[19]
rlabel metal2 5895 68 5895 68 0 FrameStrobe[1]
rlabel metal2 8103 68 8103 68 0 FrameStrobe[2]
rlabel metal2 10311 68 10311 68 0 FrameStrobe[3]
rlabel metal2 12519 68 12519 68 0 FrameStrobe[4]
rlabel metal2 14727 68 14727 68 0 FrameStrobe[5]
rlabel metal2 17027 68 17027 68 0 FrameStrobe[6]
rlabel metal2 19281 68 19281 68 0 FrameStrobe[7]
rlabel metal2 21443 68 21443 68 0 FrameStrobe[8]
rlabel metal2 23506 143 23506 143 0 FrameStrobe[9]
rlabel metal1 39468 8602 39468 8602 0 FrameStrobe_O[0]
rlabel metal1 44114 8432 44114 8432 0 FrameStrobe_O[10]
rlabel metal1 43746 7514 43746 7514 0 FrameStrobe_O[11]
rlabel metal2 43746 9224 43746 9224 0 FrameStrobe_O[12]
rlabel metal1 44758 6834 44758 6834 0 FrameStrobe_O[13]
rlabel metal2 44482 8952 44482 8952 0 FrameStrobe_O[14]
rlabel metal2 44850 9224 44850 9224 0 FrameStrobe_O[15]
rlabel metal1 44988 7446 44988 7446 0 FrameStrobe_O[16]
rlabel metal2 45586 8680 45586 8680 0 FrameStrobe_O[17]
rlabel metal2 45954 9377 45954 9377 0 FrameStrobe_O[18]
rlabel metal2 46322 8850 46322 8850 0 FrameStrobe_O[19]
rlabel metal2 39698 9224 39698 9224 0 FrameStrobe_O[1]
rlabel metal2 40066 9462 40066 9462 0 FrameStrobe_O[2]
rlabel metal1 40802 8330 40802 8330 0 FrameStrobe_O[3]
rlabel metal1 40986 8058 40986 8058 0 FrameStrobe_O[4]
rlabel metal2 41170 9224 41170 9224 0 FrameStrobe_O[5]
rlabel metal1 41814 8330 41814 8330 0 FrameStrobe_O[6]
rlabel metal1 42274 8602 42274 8602 0 FrameStrobe_O[7]
rlabel metal2 42274 9190 42274 9190 0 FrameStrobe_O[8]
rlabel metal2 42642 9088 42642 9088 0 FrameStrobe_O[9]
rlabel metal1 23460 1802 23460 1802 0 FrameStrobe_O_i\[0\]
rlabel metal1 26772 3162 26772 3162 0 FrameStrobe_O_i\[10\]
rlabel metal1 28980 2618 28980 2618 0 FrameStrobe_O_i\[11\]
rlabel metal1 31188 2074 31188 2074 0 FrameStrobe_O_i\[12\]
rlabel metal1 33396 3706 33396 3706 0 FrameStrobe_O_i\[13\]
rlabel metal2 35926 4284 35926 4284 0 FrameStrobe_O_i\[14\]
rlabel metal1 37766 2074 37766 2074 0 FrameStrobe_O_i\[15\]
rlabel metal1 42090 3162 42090 3162 0 FrameStrobe_O_i\[16\]
rlabel metal2 41814 2244 41814 2244 0 FrameStrobe_O_i\[17\]
rlabel metal2 43930 2210 43930 2210 0 FrameStrobe_O_i\[18\]
rlabel metal1 45080 2074 45080 2074 0 FrameStrobe_O_i\[19\]
rlabel metal1 23322 3978 23322 3978 0 FrameStrobe_O_i\[1\]
rlabel metal1 23276 3162 23276 3162 0 FrameStrobe_O_i\[2\]
rlabel metal2 23046 3332 23046 3332 0 FrameStrobe_O_i\[3\]
rlabel metal1 23184 2550 23184 2550 0 FrameStrobe_O_i\[4\]
rlabel metal1 23276 2074 23276 2074 0 FrameStrobe_O_i\[5\]
rlabel metal1 22632 2074 22632 2074 0 FrameStrobe_O_i\[6\]
rlabel metal1 20148 2074 20148 2074 0 FrameStrobe_O_i\[7\]
rlabel metal2 22678 3910 22678 3910 0 FrameStrobe_O_i\[8\]
rlabel metal1 24564 2074 24564 2074 0 FrameStrobe_O_i\[9\]
rlabel metal2 690 8952 690 8952 0 N1BEG[0]
rlabel metal2 1058 8680 1058 8680 0 N1BEG[1]
rlabel metal2 1426 8918 1426 8918 0 N1BEG[2]
rlabel metal1 1978 7514 1978 7514 0 N1BEG[3]
rlabel metal2 2162 8952 2162 8952 0 N2BEG[0]
rlabel metal1 2116 8602 2116 8602 0 N2BEG[1]
rlabel metal1 2852 8602 2852 8602 0 N2BEG[2]
rlabel metal1 3220 8602 3220 8602 0 N2BEG[3]
rlabel metal1 3588 8602 3588 8602 0 N2BEG[4]
rlabel metal2 4002 8918 4002 8918 0 N2BEG[5]
rlabel metal1 4324 8602 4324 8602 0 N2BEG[6]
rlabel metal1 4692 8058 4692 8058 0 N2BEG[7]
rlabel metal1 4876 8602 4876 8602 0 N2BEGb[0]
rlabel metal1 5336 8602 5336 8602 0 N2BEGb[1]
rlabel metal1 5796 8058 5796 8058 0 N2BEGb[2]
rlabel metal1 6164 8602 6164 8602 0 N2BEGb[3]
rlabel metal2 6578 9309 6578 9309 0 N2BEGb[4]
rlabel metal2 6854 8823 6854 8823 0 N2BEGb[5]
rlabel metal1 7268 8058 7268 8058 0 N2BEGb[6]
rlabel metal1 7544 8602 7544 8602 0 N2BEGb[7]
rlabel metal1 7912 8602 7912 8602 0 N4BEG[0]
rlabel metal2 11730 8952 11730 8952 0 N4BEG[10]
rlabel metal1 11914 8602 11914 8602 0 N4BEG[11]
rlabel metal2 12466 9513 12466 9513 0 N4BEG[12]
rlabel metal1 12788 8058 12788 8058 0 N4BEG[13]
rlabel metal1 13064 8602 13064 8602 0 N4BEG[14]
rlabel metal1 13432 8602 13432 8602 0 N4BEG[15]
rlabel metal1 8372 8602 8372 8602 0 N4BEG[1]
rlabel metal1 8740 8602 8740 8602 0 N4BEG[2]
rlabel metal2 9154 8952 9154 8952 0 N4BEG[3]
rlabel metal1 9384 8602 9384 8602 0 N4BEG[4]
rlabel metal1 9844 8602 9844 8602 0 N4BEG[5]
rlabel metal1 10212 8058 10212 8058 0 N4BEG[6]
rlabel metal1 10396 8602 10396 8602 0 N4BEG[7]
rlabel metal1 10856 8602 10856 8602 0 N4BEG[8]
rlabel metal1 11316 8602 11316 8602 0 N4BEG[9]
rlabel metal1 13892 8602 13892 8602 0 NN4BEG[0]
rlabel metal1 17756 8602 17756 8602 0 NN4BEG[10]
rlabel metal2 17986 9224 17986 9224 0 NN4BEG[11]
rlabel metal1 18492 8058 18492 8058 0 NN4BEG[12]
rlabel metal1 18860 8602 18860 8602 0 NN4BEG[13]
rlabel metal2 19090 9785 19090 9785 0 NN4BEG[14]
rlabel metal2 19458 9224 19458 9224 0 NN4BEG[15]
rlabel metal2 14306 9326 14306 9326 0 NN4BEG[1]
rlabel metal1 14536 8602 14536 8602 0 NN4BEG[2]
rlabel metal1 14904 8602 14904 8602 0 NN4BEG[3]
rlabel metal1 15364 8602 15364 8602 0 NN4BEG[4]
rlabel metal1 15732 8058 15732 8058 0 NN4BEG[5]
rlabel metal1 16008 8602 16008 8602 0 NN4BEG[6]
rlabel metal1 16468 8602 16468 8602 0 NN4BEG[7]
rlabel metal1 17020 8602 17020 8602 0 NN4BEG[8]
rlabel metal1 17388 8602 17388 8602 0 NN4BEG[9]
rlabel metal2 19826 8612 19826 8612 0 S1END[0]
rlabel metal2 20194 9785 20194 9785 0 S1END[1]
rlabel metal2 20562 8612 20562 8612 0 S1END[2]
rlabel metal2 20930 9241 20930 9241 0 S1END[3]
rlabel metal2 21298 9190 21298 9190 0 S2END[0]
rlabel metal2 21666 9122 21666 9122 0 S2END[1]
rlabel metal2 22034 9190 22034 9190 0 S2END[2]
rlabel metal1 21666 8432 21666 8432 0 S2END[3]
rlabel metal2 22770 9190 22770 9190 0 S2END[4]
rlabel metal2 23138 9122 23138 9122 0 S2END[5]
rlabel metal2 23506 9785 23506 9785 0 S2END[6]
rlabel metal2 23874 9173 23874 9173 0 S2END[7]
rlabel metal2 24242 9156 24242 9156 0 S2MID[0]
rlabel metal2 24610 9785 24610 9785 0 S2MID[1]
rlabel metal2 24978 9156 24978 9156 0 S2MID[2]
rlabel metal2 25346 9156 25346 9156 0 S2MID[3]
rlabel metal2 25714 9156 25714 9156 0 S2MID[4]
rlabel metal2 26082 9156 26082 9156 0 S2MID[5]
rlabel metal2 26450 9156 26450 9156 0 S2MID[6]
rlabel metal2 26818 9156 26818 9156 0 S2MID[7]
rlabel metal2 27186 9785 27186 9785 0 S4END[0]
rlabel metal2 30866 9156 30866 9156 0 S4END[10]
rlabel metal2 31234 9156 31234 9156 0 S4END[11]
rlabel metal2 31602 9156 31602 9156 0 S4END[12]
rlabel metal2 31970 9156 31970 9156 0 S4END[13]
rlabel metal2 32338 9156 32338 9156 0 S4END[14]
rlabel metal2 32706 9156 32706 9156 0 S4END[15]
rlabel metal2 27554 9156 27554 9156 0 S4END[1]
rlabel metal2 27922 9156 27922 9156 0 S4END[2]
rlabel metal2 28290 9156 28290 9156 0 S4END[3]
rlabel metal2 28658 9156 28658 9156 0 S4END[4]
rlabel metal2 29026 9156 29026 9156 0 S4END[5]
rlabel metal2 29394 9156 29394 9156 0 S4END[6]
rlabel metal2 29762 9785 29762 9785 0 S4END[7]
rlabel metal2 30130 9156 30130 9156 0 S4END[8]
rlabel metal2 30498 9156 30498 9156 0 S4END[9]
rlabel metal2 33074 9156 33074 9156 0 SS4END[0]
rlabel metal2 36754 9156 36754 9156 0 SS4END[10]
rlabel metal2 37122 9156 37122 9156 0 SS4END[11]
rlabel metal2 37490 9156 37490 9156 0 SS4END[12]
rlabel metal2 37858 9156 37858 9156 0 SS4END[13]
rlabel metal2 38226 9156 38226 9156 0 SS4END[14]
rlabel metal2 38594 9156 38594 9156 0 SS4END[15]
rlabel metal2 33442 9156 33442 9156 0 SS4END[1]
rlabel metal2 33810 9156 33810 9156 0 SS4END[2]
rlabel metal2 34178 9156 34178 9156 0 SS4END[3]
rlabel metal2 34546 9377 34546 9377 0 SS4END[4]
rlabel metal2 34914 9156 34914 9156 0 SS4END[5]
rlabel metal2 35282 9156 35282 9156 0 SS4END[6]
rlabel metal2 35650 9156 35650 9156 0 SS4END[7]
rlabel metal2 36018 9156 36018 9156 0 SS4END[8]
rlabel metal2 36386 9156 36386 9156 0 SS4END[9]
rlabel metal2 1479 68 1479 68 0 UserCLK
rlabel metal1 39100 8602 39100 8602 0 UserCLKo
rlabel metal1 4002 1224 4002 1224 0 net1
rlabel metal1 43792 1530 43792 1530 0 net10
rlabel metal1 2622 8466 2622 8466 0 net100
rlabel metal2 2990 7667 2990 7667 0 net101
rlabel metal2 7038 7497 7038 7497 0 net102
rlabel metal2 4002 7242 4002 7242 0 net103
rlabel metal1 4094 9554 4094 9554 0 net104
rlabel metal2 4462 8772 4462 8772 0 net105
rlabel metal1 17250 8364 17250 8364 0 net106
rlabel metal1 12558 8568 12558 8568 0 net107
rlabel metal2 21758 6749 21758 6749 0 net108
rlabel metal2 17066 8568 17066 8568 0 net109
rlabel metal1 45080 1530 45080 1530 0 net11
rlabel metal1 21850 7514 21850 7514 0 net110
rlabel metal2 21574 7667 21574 7667 0 net111
rlabel metal1 17894 7480 17894 7480 0 net112
rlabel metal1 20562 7718 20562 7718 0 net113
rlabel metal2 17158 8959 17158 8959 0 net114
rlabel metal2 28566 7225 28566 7225 0 net115
rlabel metal2 28198 8653 28198 8653 0 net116
rlabel metal1 12650 8500 12650 8500 0 net117
rlabel via2 25530 7973 25530 7973 0 net118
rlabel metal2 12742 9010 12742 9010 0 net119
rlabel metal2 6118 1088 6118 1088 0 net12
rlabel metal2 13110 9112 13110 9112 0 net120
rlabel metal1 16606 9384 16606 9384 0 net121
rlabel metal1 14030 8976 14030 8976 0 net122
rlabel metal1 15410 7344 15410 7344 0 net123
rlabel via2 21758 9469 21758 9469 0 net124
rlabel metal1 9798 8840 9798 8840 0 net125
rlabel metal1 17986 7990 17986 7990 0 net126
rlabel metal1 17434 9928 17434 9928 0 net127
rlabel metal2 17526 9554 17526 9554 0 net128
rlabel metal2 15134 8653 15134 8653 0 net129
rlabel metal1 8326 680 8326 680 0 net13
rlabel metal2 14122 8704 14122 8704 0 net130
rlabel metal1 17756 8058 17756 8058 0 net131
rlabel metal1 17572 7718 17572 7718 0 net132
rlabel metal1 18446 7888 18446 7888 0 net133
rlabel metal1 18998 7242 18998 7242 0 net134
rlabel metal1 19780 7514 19780 7514 0 net135
rlabel metal1 19550 8058 19550 8058 0 net136
rlabel metal1 18722 8024 18722 8024 0 net137
rlabel via2 19090 7157 19090 7157 0 net138
rlabel metal2 15226 7667 15226 7667 0 net139
rlabel metal1 16790 952 16790 952 0 net14
rlabel metal2 15594 8551 15594 8551 0 net140
rlabel metal1 21942 7378 21942 7378 0 net141
rlabel metal2 16606 7548 16606 7548 0 net142
rlabel metal1 21620 8058 21620 8058 0 net143
rlabel metal1 21206 8058 21206 8058 0 net144
rlabel metal1 18538 7956 18538 7956 0 net145
rlabel metal1 22954 2006 22954 2006 0 net146
rlabel metal1 17066 1292 17066 1292 0 net15
rlabel metal2 16882 1088 16882 1088 0 net16
rlabel metal1 18952 1190 18952 1190 0 net17
rlabel metal1 19550 1530 19550 1530 0 net18
rlabel metal2 21390 2346 21390 2346 0 net19
rlabel metal1 26220 3026 26220 3026 0 net2
rlabel metal1 24012 1530 24012 1530 0 net20
rlabel metal1 19596 7174 19596 7174 0 net21
rlabel metal1 19136 7514 19136 7514 0 net22
rlabel metal1 20286 7242 20286 7242 0 net23
rlabel metal1 20286 7514 20286 7514 0 net24
rlabel metal1 20562 7854 20562 7854 0 net25
rlabel metal1 20838 7854 20838 7854 0 net26
rlabel metal1 21298 7378 21298 7378 0 net27
rlabel metal1 21850 7412 21850 7412 0 net28
rlabel metal2 22310 7854 22310 7854 0 net29
rlabel metal1 28428 1530 28428 1530 0 net3
rlabel metal2 21850 8228 21850 8228 0 net30
rlabel metal1 22586 7378 22586 7378 0 net31
rlabel metal1 22402 7888 22402 7888 0 net32
rlabel metal1 23598 8432 23598 8432 0 net33
rlabel metal1 23506 7820 23506 7820 0 net34
rlabel metal1 25116 7854 25116 7854 0 net35
rlabel metal1 24886 7888 24886 7888 0 net36
rlabel metal1 25530 7854 25530 7854 0 net37
rlabel metal1 25806 7854 25806 7854 0 net38
rlabel metal1 26036 7854 26036 7854 0 net39
rlabel metal1 30636 1530 30636 1530 0 net4
rlabel metal1 26358 7854 26358 7854 0 net40
rlabel metal1 26680 7854 26680 7854 0 net41
rlabel metal1 24012 8466 24012 8466 0 net42
rlabel metal1 25760 7378 25760 7378 0 net43
rlabel metal2 30682 7820 30682 7820 0 net44
rlabel metal2 31050 8908 31050 8908 0 net45
rlabel metal1 32614 8568 32614 8568 0 net46
rlabel metal2 32982 9112 32982 9112 0 net47
rlabel metal1 27048 7854 27048 7854 0 net48
rlabel metal1 27324 7854 27324 7854 0 net49
rlabel metal2 32430 2346 32430 2346 0 net5
rlabel metal1 27784 7854 27784 7854 0 net50
rlabel metal1 28014 7922 28014 7922 0 net51
rlabel metal1 28382 7888 28382 7888 0 net52
rlabel metal1 29164 7854 29164 7854 0 net53
rlabel metal1 24610 7888 24610 7888 0 net54
rlabel metal1 23782 7922 23782 7922 0 net55
rlabel metal1 24288 7854 24288 7854 0 net56
rlabel metal2 33350 7752 33350 7752 0 net57
rlabel metal1 37030 8568 37030 8568 0 net58
rlabel metal1 37352 8602 37352 8602 0 net59
rlabel metal1 35098 1190 35098 1190 0 net6
rlabel metal2 37766 8704 37766 8704 0 net60
rlabel metal2 38134 8075 38134 8075 0 net61
rlabel metal2 38502 7803 38502 7803 0 net62
rlabel metal2 38870 9078 38870 9078 0 net63
rlabel metal2 33718 7582 33718 7582 0 net64
rlabel metal2 31970 7871 31970 7871 0 net65
rlabel metal1 33626 8602 33626 8602 0 net66
rlabel metal1 34914 8568 34914 8568 0 net67
rlabel metal2 35190 8976 35190 8976 0 net68
rlabel metal2 34178 7650 34178 7650 0 net69
rlabel metal1 37168 1190 37168 1190 0 net7
rlabel metal1 35926 8398 35926 8398 0 net70
rlabel via1 31786 8381 31786 8381 0 net71
rlabel metal2 36662 7548 36662 7548 0 net72
rlabel metal2 1702 1700 1702 1700 0 net73
rlabel metal1 24518 2550 24518 2550 0 net74
rlabel metal1 43516 8398 43516 8398 0 net75
rlabel metal1 42688 7378 42688 7378 0 net76
rlabel metal1 40066 2414 40066 2414 0 net77
rlabel metal2 42826 5202 42826 5202 0 net78
rlabel metal1 40020 4726 40020 4726 0 net79
rlabel metal2 39054 2108 39054 2108 0 net8
rlabel metal1 41768 2278 41768 2278 0 net80
rlabel metal2 44390 5644 44390 5644 0 net81
rlabel metal1 44804 2618 44804 2618 0 net82
rlabel metal1 44666 7786 44666 7786 0 net83
rlabel metal1 44758 2550 44758 2550 0 net84
rlabel metal2 39974 6494 39974 6494 0 net85
rlabel metal1 39330 8534 39330 8534 0 net86
rlabel metal2 40986 8840 40986 8840 0 net87
rlabel metal2 40986 5406 40986 5406 0 net88
rlabel metal1 23782 2278 23782 2278 0 net89
rlabel metal1 41630 1530 41630 1530 0 net9
rlabel metal2 41906 5508 41906 5508 0 net90
rlabel metal1 42458 8942 42458 8942 0 net91
rlabel metal1 36018 8330 36018 8330 0 net92
rlabel metal1 40434 9146 40434 9146 0 net93
rlabel metal1 1794 7888 1794 7888 0 net94
rlabel metal1 1518 7344 1518 7344 0 net95
rlabel metal2 2346 7514 2346 7514 0 net96
rlabel metal2 17710 7616 17710 7616 0 net97
rlabel metal2 8326 6885 8326 6885 0 net98
rlabel metal2 1518 8840 1518 8840 0 net99
<< properties >>
string FIXED_BBOX 0 0 47000 10000
<< end >>
