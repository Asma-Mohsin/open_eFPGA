magic
tech sky130A
magscale 1 2
timestamp 1733394399
<< obsli1 >>
rect 1104 1071 45816 8721
<< obsm1 >>
rect 658 8 45986 9036
<< metal2 >>
rect 1398 9840 1454 10000
rect 3606 9840 3662 10000
rect 5814 9840 5870 10000
rect 8022 9840 8078 10000
rect 10230 9840 10286 10000
rect 12438 9840 12494 10000
rect 14646 9840 14702 10000
rect 16854 9840 16910 10000
rect 19062 9840 19118 10000
rect 21270 9840 21326 10000
rect 23478 9840 23534 10000
rect 25686 9840 25742 10000
rect 27894 9840 27950 10000
rect 30102 9840 30158 10000
rect 32310 9840 32366 10000
rect 34518 9840 34574 10000
rect 36726 9840 36782 10000
rect 38934 9840 38990 10000
rect 41142 9840 41198 10000
rect 43350 9840 43406 10000
rect 45558 9840 45614 10000
rect 662 0 718 160
rect 1030 0 1086 160
rect 1398 0 1454 160
rect 1766 0 1822 160
rect 2134 0 2190 160
rect 2502 0 2558 160
rect 2870 0 2926 160
rect 3238 0 3294 160
rect 3606 0 3662 160
rect 3974 0 4030 160
rect 4342 0 4398 160
rect 4710 0 4766 160
rect 5078 0 5134 160
rect 5446 0 5502 160
rect 5814 0 5870 160
rect 6182 0 6238 160
rect 6550 0 6606 160
rect 6918 0 6974 160
rect 7286 0 7342 160
rect 7654 0 7710 160
rect 8022 0 8078 160
rect 8390 0 8446 160
rect 8758 0 8814 160
rect 9126 0 9182 160
rect 9494 0 9550 160
rect 9862 0 9918 160
rect 10230 0 10286 160
rect 10598 0 10654 160
rect 10966 0 11022 160
rect 11334 0 11390 160
rect 11702 0 11758 160
rect 12070 0 12126 160
rect 12438 0 12494 160
rect 12806 0 12862 160
rect 13174 0 13230 160
rect 13542 0 13598 160
rect 13910 0 13966 160
rect 14278 0 14334 160
rect 14646 0 14702 160
rect 15014 0 15070 160
rect 15382 0 15438 160
rect 15750 0 15806 160
rect 16118 0 16174 160
rect 16486 0 16542 160
rect 16854 0 16910 160
rect 17222 0 17278 160
rect 17590 0 17646 160
rect 17958 0 18014 160
rect 18326 0 18382 160
rect 18694 0 18750 160
rect 19062 0 19118 160
rect 19430 0 19486 160
rect 19798 0 19854 160
rect 20166 0 20222 160
rect 20534 0 20590 160
rect 20902 0 20958 160
rect 21270 0 21326 160
rect 21638 0 21694 160
rect 22006 0 22062 160
rect 22374 0 22430 160
rect 22742 0 22798 160
rect 23110 0 23166 160
rect 23478 0 23534 160
rect 23846 0 23902 160
rect 24214 0 24270 160
rect 24582 0 24638 160
rect 24950 0 25006 160
rect 25318 0 25374 160
rect 25686 0 25742 160
rect 26054 0 26110 160
rect 26422 0 26478 160
rect 26790 0 26846 160
rect 27158 0 27214 160
rect 27526 0 27582 160
rect 27894 0 27950 160
rect 28262 0 28318 160
rect 28630 0 28686 160
rect 28998 0 29054 160
rect 29366 0 29422 160
rect 29734 0 29790 160
rect 30102 0 30158 160
rect 30470 0 30526 160
rect 30838 0 30894 160
rect 31206 0 31262 160
rect 31574 0 31630 160
rect 31942 0 31998 160
rect 32310 0 32366 160
rect 32678 0 32734 160
rect 33046 0 33102 160
rect 33414 0 33470 160
rect 33782 0 33838 160
rect 34150 0 34206 160
rect 34518 0 34574 160
rect 34886 0 34942 160
rect 35254 0 35310 160
rect 35622 0 35678 160
rect 35990 0 36046 160
rect 36358 0 36414 160
rect 36726 0 36782 160
rect 37094 0 37150 160
rect 37462 0 37518 160
rect 37830 0 37886 160
rect 38198 0 38254 160
rect 38566 0 38622 160
rect 38934 0 38990 160
rect 39302 0 39358 160
rect 39670 0 39726 160
rect 40038 0 40094 160
rect 40406 0 40462 160
rect 40774 0 40830 160
rect 41142 0 41198 160
rect 41510 0 41566 160
rect 41878 0 41934 160
rect 42246 0 42302 160
rect 42614 0 42670 160
rect 42982 0 43038 160
rect 43350 0 43406 160
rect 43718 0 43774 160
rect 44086 0 44142 160
rect 44454 0 44510 160
rect 44822 0 44878 160
rect 45190 0 45246 160
rect 45558 0 45614 160
rect 45926 0 45982 160
rect 46294 0 46350 160
<< obsm2 >>
rect 664 9784 1342 9874
rect 1510 9784 3550 9874
rect 3718 9784 5758 9874
rect 5926 9784 7966 9874
rect 8134 9784 10174 9874
rect 10342 9784 12382 9874
rect 12550 9784 14590 9874
rect 14758 9784 16798 9874
rect 16966 9784 19006 9874
rect 19174 9784 21214 9874
rect 21382 9784 23422 9874
rect 23590 9784 25630 9874
rect 25798 9784 27838 9874
rect 28006 9784 30046 9874
rect 30214 9784 32254 9874
rect 32422 9784 34462 9874
rect 34630 9784 36670 9874
rect 36838 9784 38878 9874
rect 39046 9784 41086 9874
rect 41254 9784 43294 9874
rect 43462 9784 45502 9874
rect 45670 9784 46294 9874
rect 664 216 46294 9784
rect 774 2 974 216
rect 1142 2 1342 216
rect 1510 2 1710 216
rect 1878 2 2078 216
rect 2246 2 2446 216
rect 2614 2 2814 216
rect 2982 2 3182 216
rect 3350 2 3550 216
rect 3718 2 3918 216
rect 4086 2 4286 216
rect 4454 2 4654 216
rect 4822 2 5022 216
rect 5190 2 5390 216
rect 5558 2 5758 216
rect 5926 2 6126 216
rect 6294 2 6494 216
rect 6662 2 6862 216
rect 7030 2 7230 216
rect 7398 2 7598 216
rect 7766 2 7966 216
rect 8134 2 8334 216
rect 8502 2 8702 216
rect 8870 2 9070 216
rect 9238 2 9438 216
rect 9606 2 9806 216
rect 9974 2 10174 216
rect 10342 2 10542 216
rect 10710 2 10910 216
rect 11078 2 11278 216
rect 11446 2 11646 216
rect 11814 2 12014 216
rect 12182 2 12382 216
rect 12550 2 12750 216
rect 12918 2 13118 216
rect 13286 2 13486 216
rect 13654 2 13854 216
rect 14022 2 14222 216
rect 14390 2 14590 216
rect 14758 2 14958 216
rect 15126 2 15326 216
rect 15494 2 15694 216
rect 15862 2 16062 216
rect 16230 2 16430 216
rect 16598 2 16798 216
rect 16966 2 17166 216
rect 17334 2 17534 216
rect 17702 2 17902 216
rect 18070 2 18270 216
rect 18438 2 18638 216
rect 18806 2 19006 216
rect 19174 2 19374 216
rect 19542 2 19742 216
rect 19910 2 20110 216
rect 20278 2 20478 216
rect 20646 2 20846 216
rect 21014 2 21214 216
rect 21382 2 21582 216
rect 21750 2 21950 216
rect 22118 2 22318 216
rect 22486 2 22686 216
rect 22854 2 23054 216
rect 23222 2 23422 216
rect 23590 2 23790 216
rect 23958 2 24158 216
rect 24326 2 24526 216
rect 24694 2 24894 216
rect 25062 2 25262 216
rect 25430 2 25630 216
rect 25798 2 25998 216
rect 26166 2 26366 216
rect 26534 2 26734 216
rect 26902 2 27102 216
rect 27270 2 27470 216
rect 27638 2 27838 216
rect 28006 2 28206 216
rect 28374 2 28574 216
rect 28742 2 28942 216
rect 29110 2 29310 216
rect 29478 2 29678 216
rect 29846 2 30046 216
rect 30214 2 30414 216
rect 30582 2 30782 216
rect 30950 2 31150 216
rect 31318 2 31518 216
rect 31686 2 31886 216
rect 32054 2 32254 216
rect 32422 2 32622 216
rect 32790 2 32990 216
rect 33158 2 33358 216
rect 33526 2 33726 216
rect 33894 2 34094 216
rect 34262 2 34462 216
rect 34630 2 34830 216
rect 34998 2 35198 216
rect 35366 2 35566 216
rect 35734 2 35934 216
rect 36102 2 36302 216
rect 36470 2 36670 216
rect 36838 2 37038 216
rect 37206 2 37406 216
rect 37574 2 37774 216
rect 37942 2 38142 216
rect 38310 2 38510 216
rect 38678 2 38878 216
rect 39046 2 39246 216
rect 39414 2 39614 216
rect 39782 2 39982 216
rect 40150 2 40350 216
rect 40518 2 40718 216
rect 40886 2 41086 216
rect 41254 2 41454 216
rect 41622 2 41822 216
rect 41990 2 42190 216
rect 42358 2 42558 216
rect 42726 2 42926 216
rect 43094 2 43294 216
rect 43462 2 43662 216
rect 43830 2 44030 216
rect 44198 2 44398 216
rect 44566 2 44766 216
rect 44934 2 45134 216
rect 45302 2 45502 216
rect 45670 2 45870 216
rect 46038 2 46238 216
<< obsm3 >>
rect 2037 171 45974 8737
<< metal4 >>
rect 6533 1040 6853 8752
rect 12122 1040 12442 8752
rect 17711 1040 18031 8752
rect 23300 1040 23620 8752
rect 28889 1040 29209 8752
rect 34478 1040 34798 8752
rect 40067 1040 40387 8752
rect 45656 1040 45976 8752
<< labels >>
rlabel metal2 s 39302 0 39358 160 6 FrameStrobe[0]
port 1 nsew signal input
rlabel metal2 s 42982 0 43038 160 6 FrameStrobe[10]
port 2 nsew signal input
rlabel metal2 s 43350 0 43406 160 6 FrameStrobe[11]
port 3 nsew signal input
rlabel metal2 s 43718 0 43774 160 6 FrameStrobe[12]
port 4 nsew signal input
rlabel metal2 s 44086 0 44142 160 6 FrameStrobe[13]
port 5 nsew signal input
rlabel metal2 s 44454 0 44510 160 6 FrameStrobe[14]
port 6 nsew signal input
rlabel metal2 s 44822 0 44878 160 6 FrameStrobe[15]
port 7 nsew signal input
rlabel metal2 s 45190 0 45246 160 6 FrameStrobe[16]
port 8 nsew signal input
rlabel metal2 s 45558 0 45614 160 6 FrameStrobe[17]
port 9 nsew signal input
rlabel metal2 s 45926 0 45982 160 6 FrameStrobe[18]
port 10 nsew signal input
rlabel metal2 s 46294 0 46350 160 6 FrameStrobe[19]
port 11 nsew signal input
rlabel metal2 s 39670 0 39726 160 6 FrameStrobe[1]
port 12 nsew signal input
rlabel metal2 s 40038 0 40094 160 6 FrameStrobe[2]
port 13 nsew signal input
rlabel metal2 s 40406 0 40462 160 6 FrameStrobe[3]
port 14 nsew signal input
rlabel metal2 s 40774 0 40830 160 6 FrameStrobe[4]
port 15 nsew signal input
rlabel metal2 s 41142 0 41198 160 6 FrameStrobe[5]
port 16 nsew signal input
rlabel metal2 s 41510 0 41566 160 6 FrameStrobe[6]
port 17 nsew signal input
rlabel metal2 s 41878 0 41934 160 6 FrameStrobe[7]
port 18 nsew signal input
rlabel metal2 s 42246 0 42302 160 6 FrameStrobe[8]
port 19 nsew signal input
rlabel metal2 s 42614 0 42670 160 6 FrameStrobe[9]
port 20 nsew signal input
rlabel metal2 s 3606 9840 3662 10000 6 FrameStrobe_O[0]
port 21 nsew signal output
rlabel metal2 s 25686 9840 25742 10000 6 FrameStrobe_O[10]
port 22 nsew signal output
rlabel metal2 s 27894 9840 27950 10000 6 FrameStrobe_O[11]
port 23 nsew signal output
rlabel metal2 s 30102 9840 30158 10000 6 FrameStrobe_O[12]
port 24 nsew signal output
rlabel metal2 s 32310 9840 32366 10000 6 FrameStrobe_O[13]
port 25 nsew signal output
rlabel metal2 s 34518 9840 34574 10000 6 FrameStrobe_O[14]
port 26 nsew signal output
rlabel metal2 s 36726 9840 36782 10000 6 FrameStrobe_O[15]
port 27 nsew signal output
rlabel metal2 s 38934 9840 38990 10000 6 FrameStrobe_O[16]
port 28 nsew signal output
rlabel metal2 s 41142 9840 41198 10000 6 FrameStrobe_O[17]
port 29 nsew signal output
rlabel metal2 s 43350 9840 43406 10000 6 FrameStrobe_O[18]
port 30 nsew signal output
rlabel metal2 s 45558 9840 45614 10000 6 FrameStrobe_O[19]
port 31 nsew signal output
rlabel metal2 s 5814 9840 5870 10000 6 FrameStrobe_O[1]
port 32 nsew signal output
rlabel metal2 s 8022 9840 8078 10000 6 FrameStrobe_O[2]
port 33 nsew signal output
rlabel metal2 s 10230 9840 10286 10000 6 FrameStrobe_O[3]
port 34 nsew signal output
rlabel metal2 s 12438 9840 12494 10000 6 FrameStrobe_O[4]
port 35 nsew signal output
rlabel metal2 s 14646 9840 14702 10000 6 FrameStrobe_O[5]
port 36 nsew signal output
rlabel metal2 s 16854 9840 16910 10000 6 FrameStrobe_O[6]
port 37 nsew signal output
rlabel metal2 s 19062 9840 19118 10000 6 FrameStrobe_O[7]
port 38 nsew signal output
rlabel metal2 s 21270 9840 21326 10000 6 FrameStrobe_O[8]
port 39 nsew signal output
rlabel metal2 s 23478 9840 23534 10000 6 FrameStrobe_O[9]
port 40 nsew signal output
rlabel metal2 s 662 0 718 160 6 N1END[0]
port 41 nsew signal input
rlabel metal2 s 1030 0 1086 160 6 N1END[1]
port 42 nsew signal input
rlabel metal2 s 1398 0 1454 160 6 N1END[2]
port 43 nsew signal input
rlabel metal2 s 1766 0 1822 160 6 N1END[3]
port 44 nsew signal input
rlabel metal2 s 5078 0 5134 160 6 N2END[0]
port 45 nsew signal input
rlabel metal2 s 5446 0 5502 160 6 N2END[1]
port 46 nsew signal input
rlabel metal2 s 5814 0 5870 160 6 N2END[2]
port 47 nsew signal input
rlabel metal2 s 6182 0 6238 160 6 N2END[3]
port 48 nsew signal input
rlabel metal2 s 6550 0 6606 160 6 N2END[4]
port 49 nsew signal input
rlabel metal2 s 6918 0 6974 160 6 N2END[5]
port 50 nsew signal input
rlabel metal2 s 7286 0 7342 160 6 N2END[6]
port 51 nsew signal input
rlabel metal2 s 7654 0 7710 160 6 N2END[7]
port 52 nsew signal input
rlabel metal2 s 2134 0 2190 160 6 N2MID[0]
port 53 nsew signal input
rlabel metal2 s 2502 0 2558 160 6 N2MID[1]
port 54 nsew signal input
rlabel metal2 s 2870 0 2926 160 6 N2MID[2]
port 55 nsew signal input
rlabel metal2 s 3238 0 3294 160 6 N2MID[3]
port 56 nsew signal input
rlabel metal2 s 3606 0 3662 160 6 N2MID[4]
port 57 nsew signal input
rlabel metal2 s 3974 0 4030 160 6 N2MID[5]
port 58 nsew signal input
rlabel metal2 s 4342 0 4398 160 6 N2MID[6]
port 59 nsew signal input
rlabel metal2 s 4710 0 4766 160 6 N2MID[7]
port 60 nsew signal input
rlabel metal2 s 8022 0 8078 160 6 N4END[0]
port 61 nsew signal input
rlabel metal2 s 11702 0 11758 160 6 N4END[10]
port 62 nsew signal input
rlabel metal2 s 12070 0 12126 160 6 N4END[11]
port 63 nsew signal input
rlabel metal2 s 12438 0 12494 160 6 N4END[12]
port 64 nsew signal input
rlabel metal2 s 12806 0 12862 160 6 N4END[13]
port 65 nsew signal input
rlabel metal2 s 13174 0 13230 160 6 N4END[14]
port 66 nsew signal input
rlabel metal2 s 13542 0 13598 160 6 N4END[15]
port 67 nsew signal input
rlabel metal2 s 8390 0 8446 160 6 N4END[1]
port 68 nsew signal input
rlabel metal2 s 8758 0 8814 160 6 N4END[2]
port 69 nsew signal input
rlabel metal2 s 9126 0 9182 160 6 N4END[3]
port 70 nsew signal input
rlabel metal2 s 9494 0 9550 160 6 N4END[4]
port 71 nsew signal input
rlabel metal2 s 9862 0 9918 160 6 N4END[5]
port 72 nsew signal input
rlabel metal2 s 10230 0 10286 160 6 N4END[6]
port 73 nsew signal input
rlabel metal2 s 10598 0 10654 160 6 N4END[7]
port 74 nsew signal input
rlabel metal2 s 10966 0 11022 160 6 N4END[8]
port 75 nsew signal input
rlabel metal2 s 11334 0 11390 160 6 N4END[9]
port 76 nsew signal input
rlabel metal2 s 13910 0 13966 160 6 NN4END[0]
port 77 nsew signal input
rlabel metal2 s 17590 0 17646 160 6 NN4END[10]
port 78 nsew signal input
rlabel metal2 s 17958 0 18014 160 6 NN4END[11]
port 79 nsew signal input
rlabel metal2 s 18326 0 18382 160 6 NN4END[12]
port 80 nsew signal input
rlabel metal2 s 18694 0 18750 160 6 NN4END[13]
port 81 nsew signal input
rlabel metal2 s 19062 0 19118 160 6 NN4END[14]
port 82 nsew signal input
rlabel metal2 s 19430 0 19486 160 6 NN4END[15]
port 83 nsew signal input
rlabel metal2 s 14278 0 14334 160 6 NN4END[1]
port 84 nsew signal input
rlabel metal2 s 14646 0 14702 160 6 NN4END[2]
port 85 nsew signal input
rlabel metal2 s 15014 0 15070 160 6 NN4END[3]
port 86 nsew signal input
rlabel metal2 s 15382 0 15438 160 6 NN4END[4]
port 87 nsew signal input
rlabel metal2 s 15750 0 15806 160 6 NN4END[5]
port 88 nsew signal input
rlabel metal2 s 16118 0 16174 160 6 NN4END[6]
port 89 nsew signal input
rlabel metal2 s 16486 0 16542 160 6 NN4END[7]
port 90 nsew signal input
rlabel metal2 s 16854 0 16910 160 6 NN4END[8]
port 91 nsew signal input
rlabel metal2 s 17222 0 17278 160 6 NN4END[9]
port 92 nsew signal input
rlabel metal2 s 19798 0 19854 160 6 S1BEG[0]
port 93 nsew signal output
rlabel metal2 s 20166 0 20222 160 6 S1BEG[1]
port 94 nsew signal output
rlabel metal2 s 20534 0 20590 160 6 S1BEG[2]
port 95 nsew signal output
rlabel metal2 s 20902 0 20958 160 6 S1BEG[3]
port 96 nsew signal output
rlabel metal2 s 24214 0 24270 160 6 S2BEG[0]
port 97 nsew signal output
rlabel metal2 s 24582 0 24638 160 6 S2BEG[1]
port 98 nsew signal output
rlabel metal2 s 24950 0 25006 160 6 S2BEG[2]
port 99 nsew signal output
rlabel metal2 s 25318 0 25374 160 6 S2BEG[3]
port 100 nsew signal output
rlabel metal2 s 25686 0 25742 160 6 S2BEG[4]
port 101 nsew signal output
rlabel metal2 s 26054 0 26110 160 6 S2BEG[5]
port 102 nsew signal output
rlabel metal2 s 26422 0 26478 160 6 S2BEG[6]
port 103 nsew signal output
rlabel metal2 s 26790 0 26846 160 6 S2BEG[7]
port 104 nsew signal output
rlabel metal2 s 21270 0 21326 160 6 S2BEGb[0]
port 105 nsew signal output
rlabel metal2 s 21638 0 21694 160 6 S2BEGb[1]
port 106 nsew signal output
rlabel metal2 s 22006 0 22062 160 6 S2BEGb[2]
port 107 nsew signal output
rlabel metal2 s 22374 0 22430 160 6 S2BEGb[3]
port 108 nsew signal output
rlabel metal2 s 22742 0 22798 160 6 S2BEGb[4]
port 109 nsew signal output
rlabel metal2 s 23110 0 23166 160 6 S2BEGb[5]
port 110 nsew signal output
rlabel metal2 s 23478 0 23534 160 6 S2BEGb[6]
port 111 nsew signal output
rlabel metal2 s 23846 0 23902 160 6 S2BEGb[7]
port 112 nsew signal output
rlabel metal2 s 27158 0 27214 160 6 S4BEG[0]
port 113 nsew signal output
rlabel metal2 s 30838 0 30894 160 6 S4BEG[10]
port 114 nsew signal output
rlabel metal2 s 31206 0 31262 160 6 S4BEG[11]
port 115 nsew signal output
rlabel metal2 s 31574 0 31630 160 6 S4BEG[12]
port 116 nsew signal output
rlabel metal2 s 31942 0 31998 160 6 S4BEG[13]
port 117 nsew signal output
rlabel metal2 s 32310 0 32366 160 6 S4BEG[14]
port 118 nsew signal output
rlabel metal2 s 32678 0 32734 160 6 S4BEG[15]
port 119 nsew signal output
rlabel metal2 s 27526 0 27582 160 6 S4BEG[1]
port 120 nsew signal output
rlabel metal2 s 27894 0 27950 160 6 S4BEG[2]
port 121 nsew signal output
rlabel metal2 s 28262 0 28318 160 6 S4BEG[3]
port 122 nsew signal output
rlabel metal2 s 28630 0 28686 160 6 S4BEG[4]
port 123 nsew signal output
rlabel metal2 s 28998 0 29054 160 6 S4BEG[5]
port 124 nsew signal output
rlabel metal2 s 29366 0 29422 160 6 S4BEG[6]
port 125 nsew signal output
rlabel metal2 s 29734 0 29790 160 6 S4BEG[7]
port 126 nsew signal output
rlabel metal2 s 30102 0 30158 160 6 S4BEG[8]
port 127 nsew signal output
rlabel metal2 s 30470 0 30526 160 6 S4BEG[9]
port 128 nsew signal output
rlabel metal2 s 33046 0 33102 160 6 SS4BEG[0]
port 129 nsew signal output
rlabel metal2 s 36726 0 36782 160 6 SS4BEG[10]
port 130 nsew signal output
rlabel metal2 s 37094 0 37150 160 6 SS4BEG[11]
port 131 nsew signal output
rlabel metal2 s 37462 0 37518 160 6 SS4BEG[12]
port 132 nsew signal output
rlabel metal2 s 37830 0 37886 160 6 SS4BEG[13]
port 133 nsew signal output
rlabel metal2 s 38198 0 38254 160 6 SS4BEG[14]
port 134 nsew signal output
rlabel metal2 s 38566 0 38622 160 6 SS4BEG[15]
port 135 nsew signal output
rlabel metal2 s 33414 0 33470 160 6 SS4BEG[1]
port 136 nsew signal output
rlabel metal2 s 33782 0 33838 160 6 SS4BEG[2]
port 137 nsew signal output
rlabel metal2 s 34150 0 34206 160 6 SS4BEG[3]
port 138 nsew signal output
rlabel metal2 s 34518 0 34574 160 6 SS4BEG[4]
port 139 nsew signal output
rlabel metal2 s 34886 0 34942 160 6 SS4BEG[5]
port 140 nsew signal output
rlabel metal2 s 35254 0 35310 160 6 SS4BEG[6]
port 141 nsew signal output
rlabel metal2 s 35622 0 35678 160 6 SS4BEG[7]
port 142 nsew signal output
rlabel metal2 s 35990 0 36046 160 6 SS4BEG[8]
port 143 nsew signal output
rlabel metal2 s 36358 0 36414 160 6 SS4BEG[9]
port 144 nsew signal output
rlabel metal2 s 38934 0 38990 160 6 UserCLK
port 145 nsew signal input
rlabel metal2 s 1398 9840 1454 10000 6 UserCLKo
port 146 nsew signal output
rlabel metal4 s 6533 1040 6853 8752 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 17711 1040 18031 8752 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 28889 1040 29209 8752 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 40067 1040 40387 8752 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 12122 1040 12442 8752 6 vssd1
port 148 nsew ground bidirectional
rlabel metal4 s 23300 1040 23620 8752 6 vssd1
port 148 nsew ground bidirectional
rlabel metal4 s 34478 1040 34798 8752 6 vssd1
port 148 nsew ground bidirectional
rlabel metal4 s 45656 1040 45976 8752 6 vssd1
port 148 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 47000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 590188
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/N_term_single2/runs/24_12_05_10_25/results/signoff/N_term_single2.magic.gds
string GDS_START 50318
<< end >>

