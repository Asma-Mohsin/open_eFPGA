VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_1kbyte_1rw1r_32x256_8
   CLASS BLOCK ;
   SIZE 479.78 BY 397.5 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  106.76 0.0 107.14 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  112.88 0.0 113.26 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  118.32 0.0 118.7 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  125.12 0.0 125.5 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  130.56 0.0 130.94 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  136.0 0.0 136.38 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  141.44 0.0 141.82 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  148.24 0.0 148.62 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  153.68 0.0 154.06 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  159.12 0.0 159.5 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  165.24 0.0 165.62 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  170.68 0.0 171.06 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  177.48 0.0 177.86 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  182.92 0.0 183.3 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  188.36 0.0 188.74 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  194.48 0.0 194.86 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  201.28 0.0 201.66 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  206.72 0.0 207.1 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  212.16 0.0 212.54 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 0.0 217.98 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  224.4 0.0 224.78 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  229.84 0.0 230.22 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  235.28 0.0 235.66 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  241.4 0.0 241.78 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  246.84 0.0 247.22 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  253.64 0.0 254.02 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.08 0.0 259.46 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  264.52 0.0 264.9 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  269.96 0.0 270.34 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  276.08 0.0 276.46 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  282.88 0.0 283.26 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  288.32 0.0 288.7 1.06 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  77.52 0.0 77.9 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 128.52 1.06 128.9 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 137.36 1.06 137.74 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 142.12 1.06 142.5 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 150.28 1.06 150.66 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 155.72 1.06 156.1 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 164.56 1.06 164.94 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 170.68 1.06 171.06 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  397.12 396.44 397.5 397.5 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  478.72 82.96 479.78 83.34 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  478.72 74.8 479.78 75.18 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  478.72 68.0 479.78 68.38 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  415.48 0.0 415.86 1.06 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  413.44 0.0 413.82 1.06 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  414.12 0.0 414.5 1.06 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  414.8 0.0 415.18 1.06 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 27.88 1.06 28.26 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  478.72 382.16 479.78 382.54 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 36.04 1.06 36.42 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  29.24 0.0 29.62 1.06 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  450.16 396.44 450.54 397.5 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  83.64 0.0 84.02 1.06 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  89.08 0.0 89.46 1.06 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  95.88 0.0 96.26 1.06 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  100.64 0.0 101.02 1.06 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  139.4 0.0 139.78 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  146.2 0.0 146.58 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  151.64 0.0 152.02 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  159.8 0.0 160.18 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  165.92 0.0 166.3 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.04 0.0 172.42 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.16 0.0 178.54 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.28 0.0 184.66 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  189.04 0.0 189.42 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  196.52 0.0 196.9 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.32 0.0 203.7 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.44 0.0 209.82 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  215.56 0.0 215.94 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  221.68 0.0 222.06 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  227.8 0.0 228.18 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  233.24 0.0 233.62 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  239.36 0.0 239.74 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  245.48 0.0 245.86 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  252.96 0.0 253.34 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  257.04 0.0 257.42 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  265.88 0.0 266.26 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.0 0.0 272.38 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.12 0.0 278.5 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.24 0.0 284.62 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  289.0 0.0 289.38 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  296.48 0.0 296.86 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  302.6 0.0 302.98 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  309.4 0.0 309.78 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  315.52 0.0 315.9 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  321.64 0.0 322.02 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  327.76 0.0 328.14 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  333.88 0.0 334.26 1.06 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  140.76 396.44 141.14 397.5 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  147.56 396.44 147.94 397.5 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.0 396.44 153.38 397.5 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  159.8 396.44 160.18 397.5 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  165.92 396.44 166.3 397.5 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.72 396.44 173.1 397.5 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.84 396.44 179.22 397.5 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.28 396.44 184.66 397.5 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.08 396.44 191.46 397.5 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  196.52 396.44 196.9 397.5 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.32 396.44 203.7 397.5 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.44 396.44 209.82 397.5 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.24 396.44 216.62 397.5 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  221.68 396.44 222.06 397.5 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  227.8 396.44 228.18 397.5 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  234.6 396.44 234.98 397.5 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  240.72 396.44 241.1 397.5 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  247.52 396.44 247.9 397.5 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  252.96 396.44 253.34 397.5 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  259.76 396.44 260.14 397.5 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  265.2 396.44 265.58 397.5 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  271.32 396.44 271.7 397.5 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.12 396.44 278.5 397.5 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.24 396.44 284.62 397.5 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  291.04 396.44 291.42 397.5 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  296.48 396.44 296.86 397.5 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  303.28 396.44 303.66 397.5 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  309.4 396.44 309.78 397.5 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  316.2 396.44 316.58 397.5 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  321.64 396.44 322.02 397.5 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  327.76 396.44 328.14 397.5 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  334.56 396.44 334.94 397.5 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  473.28 4.76 475.02 392.74 ;
         LAYER met4 ;
         RECT  4.76 4.76 6.5 392.74 ;
         LAYER met3 ;
         RECT  4.76 4.76 475.02 6.5 ;
         LAYER met3 ;
         RECT  4.76 391.0 475.02 392.74 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  1.36 1.36 3.1 396.14 ;
         LAYER met3 ;
         RECT  1.36 394.4 478.42 396.14 ;
         LAYER met3 ;
         RECT  1.36 1.36 478.42 3.1 ;
         LAYER met4 ;
         RECT  476.68 1.36 478.42 396.14 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 479.16 396.88 ;
   LAYER  met2 ;
      RECT  0.62 0.62 479.16 396.88 ;
   LAYER  met3 ;
      RECT  1.66 127.92 479.16 129.5 ;
      RECT  0.62 129.5 1.66 136.76 ;
      RECT  0.62 138.34 1.66 141.52 ;
      RECT  0.62 143.1 1.66 149.68 ;
      RECT  0.62 151.26 1.66 155.12 ;
      RECT  0.62 156.7 1.66 163.96 ;
      RECT  0.62 165.54 1.66 170.08 ;
      RECT  1.66 82.36 478.12 83.94 ;
      RECT  1.66 83.94 478.12 127.92 ;
      RECT  478.12 83.94 479.16 127.92 ;
      RECT  478.12 75.78 479.16 82.36 ;
      RECT  478.12 68.98 479.16 74.2 ;
      RECT  1.66 129.5 478.12 381.56 ;
      RECT  1.66 381.56 478.12 383.14 ;
      RECT  478.12 129.5 479.16 381.56 ;
      RECT  0.62 28.86 1.66 35.44 ;
      RECT  0.62 37.02 1.66 127.92 ;
      RECT  1.66 4.16 4.16 7.1 ;
      RECT  1.66 7.1 4.16 82.36 ;
      RECT  4.16 7.1 475.62 82.36 ;
      RECT  475.62 4.16 478.12 7.1 ;
      RECT  475.62 7.1 478.12 82.36 ;
      RECT  1.66 383.14 4.16 390.4 ;
      RECT  1.66 390.4 4.16 393.34 ;
      RECT  4.16 383.14 475.62 390.4 ;
      RECT  475.62 383.14 478.12 390.4 ;
      RECT  475.62 390.4 478.12 393.34 ;
      RECT  0.62 171.66 0.76 393.8 ;
      RECT  0.62 393.8 0.76 396.74 ;
      RECT  0.62 396.74 0.76 396.88 ;
      RECT  0.76 171.66 1.66 393.8 ;
      RECT  0.76 396.74 1.66 396.88 ;
      RECT  478.12 383.14 479.02 393.8 ;
      RECT  478.12 396.74 479.02 396.88 ;
      RECT  479.02 383.14 479.16 393.8 ;
      RECT  479.02 393.8 479.16 396.74 ;
      RECT  479.02 396.74 479.16 396.88 ;
      RECT  1.66 393.34 4.16 393.8 ;
      RECT  1.66 396.74 4.16 396.88 ;
      RECT  4.16 393.34 475.62 393.8 ;
      RECT  4.16 396.74 475.62 396.88 ;
      RECT  475.62 393.34 478.12 393.8 ;
      RECT  475.62 396.74 478.12 396.88 ;
      RECT  478.12 0.62 479.02 0.76 ;
      RECT  478.12 3.7 479.02 67.4 ;
      RECT  479.02 0.62 479.16 0.76 ;
      RECT  479.02 0.76 479.16 3.7 ;
      RECT  479.02 3.7 479.16 67.4 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 27.28 ;
      RECT  0.76 0.62 1.66 0.76 ;
      RECT  0.76 3.7 1.66 27.28 ;
      RECT  1.66 0.62 4.16 0.76 ;
      RECT  1.66 3.7 4.16 4.16 ;
      RECT  4.16 0.62 475.62 0.76 ;
      RECT  4.16 3.7 475.62 4.16 ;
      RECT  475.62 0.62 478.12 0.76 ;
      RECT  475.62 3.7 478.12 4.16 ;
   LAYER  met4 ;
      RECT 10.880 389.150 11.260 391.380 ;
      RECT 19.720 389.150 20.100 391.380 ;
      RECT 27.200 389.150 27.580 391.380 ;
      RECT 36.040 389.150 36.420 391.380 ;
      RECT 44.880 389.150 45.260 391.380 ;
      RECT 52.360 389.150 52.740 391.380 ;
      RECT 61.200 389.150 61.580 391.380 ;
      RECT 70.040 389.150 70.420 391.380 ;
      RECT 78.200 389.150 78.580 391.380 ;
      RECT 87.040 389.150 87.420 391.380 ;
      RECT 94.520 389.150 94.900 391.380 ;
      RECT 103.360 389.150 103.740 391.380 ;
      RECT 110.840 389.150 111.220 391.380 ;
      RECT 119.680 389.150 120.060 391.380 ;
      RECT 128.520 389.150 128.900 391.380 ;
      RECT 137.360 389.150 137.740 391.380 ;
      RECT 10.905 388.985 11.235 389.150 ;
      RECT 19.745 388.985 20.075 389.150 ;
      RECT 27.225 388.985 27.555 389.150 ;
      RECT 36.065 388.985 36.395 389.150 ;
      RECT 44.905 388.985 45.235 389.150 ;
      RECT 52.385 388.985 52.715 389.150 ;
      RECT 61.225 388.985 61.555 389.150 ;
      RECT 70.065 388.985 70.395 389.150 ;
      RECT 78.225 388.985 78.555 389.150 ;
      RECT 87.065 388.985 87.395 389.150 ;
      RECT 94.545 388.985 94.875 389.150 ;
      RECT 103.385 388.985 103.715 389.150 ;
      RECT 110.865 388.985 111.195 389.150 ;
      RECT 119.705 388.985 120.035 389.150 ;
      RECT 128.545 388.985 128.875 389.150 ;
      RECT 137.385 388.985 137.715 389.150 ;
      RECT 140.760 370.790 141.140 396.440 ;
      RECT 144.840 389.150 145.220 391.380 ;
      RECT 144.865 388.985 145.195 389.150 ;
      RECT 147.560 370.790 147.940 396.440 ;
      RECT 148.945 388.470 149.275 388.635 ;
      RECT 140.785 370.625 141.115 370.790 ;
      RECT 147.585 370.625 147.915 370.790 ;
      RECT 148.920 369.240 149.300 388.470 ;
      RECT 153.000 370.790 153.380 396.440 ;
      RECT 154.360 389.150 154.740 391.380 ;
      RECT 154.385 388.985 154.715 389.150 ;
      RECT 159.800 370.790 160.180 396.440 ;
      RECT 162.520 389.150 162.900 391.380 ;
      RECT 162.545 388.985 162.875 389.150 ;
      RECT 165.920 370.790 166.300 396.440 ;
      RECT 170.680 389.150 171.060 391.380 ;
      RECT 170.705 388.985 171.035 389.150 ;
      RECT 172.720 370.790 173.100 396.440 ;
      RECT 177.480 389.150 177.860 391.380 ;
      RECT 177.505 388.985 177.835 389.150 ;
      RECT 178.840 370.790 179.220 396.440 ;
      RECT 184.280 370.790 184.660 396.440 ;
      RECT 187.000 389.150 187.380 391.380 ;
      RECT 187.025 388.985 187.355 389.150 ;
      RECT 191.080 370.790 191.460 396.440 ;
      RECT 195.840 389.150 196.220 391.380 ;
      RECT 195.865 388.985 196.195 389.150 ;
      RECT 196.520 370.790 196.900 396.440 ;
      RECT 202.640 389.150 203.020 391.380 ;
      RECT 202.665 388.985 202.995 389.150 ;
      RECT 203.320 370.790 203.700 396.440 ;
      RECT 209.440 370.790 209.820 396.440 ;
      RECT 212.160 389.150 212.540 391.380 ;
      RECT 212.185 388.985 212.515 389.150 ;
      RECT 216.240 370.790 216.620 396.440 ;
      RECT 221.000 389.150 221.380 391.380 ;
      RECT 221.025 388.985 221.355 389.150 ;
      RECT 221.680 370.790 222.060 396.440 ;
      RECT 227.800 370.790 228.180 396.440 ;
      RECT 229.160 389.150 229.540 391.380 ;
      RECT 229.185 388.985 229.515 389.150 ;
      RECT 234.600 370.790 234.980 396.440 ;
      RECT 237.320 389.150 237.700 391.380 ;
      RECT 237.345 388.985 237.675 389.150 ;
      RECT 240.720 370.790 241.100 396.440 ;
      RECT 246.160 389.150 246.540 391.380 ;
      RECT 246.185 388.985 246.515 389.150 ;
      RECT 247.520 370.790 247.900 396.440 ;
      RECT 252.960 370.790 253.340 396.440 ;
      RECT 253.640 389.150 254.020 391.380 ;
      RECT 253.665 388.985 253.995 389.150 ;
      RECT 259.760 370.790 260.140 396.440 ;
      RECT 263.160 389.150 263.540 391.380 ;
      RECT 263.185 388.985 263.515 389.150 ;
      RECT 265.200 370.790 265.580 396.440 ;
      RECT 270.640 389.150 271.020 391.380 ;
      RECT 270.665 388.985 270.995 389.150 ;
      RECT 271.320 370.790 271.700 396.440 ;
      RECT 278.120 370.790 278.500 396.440 ;
      RECT 279.480 389.150 279.860 391.380 ;
      RECT 279.505 388.985 279.835 389.150 ;
      RECT 284.240 370.790 284.620 396.440 ;
      RECT 288.320 389.150 288.700 391.380 ;
      RECT 288.345 388.985 288.675 389.150 ;
      RECT 291.040 370.790 291.420 396.440 ;
      RECT 295.800 389.150 296.180 391.380 ;
      RECT 295.825 388.985 296.155 389.150 ;
      RECT 296.480 370.790 296.860 396.440 ;
      RECT 303.280 370.790 303.660 396.440 ;
      RECT 304.640 389.150 305.020 391.380 ;
      RECT 304.665 388.985 304.995 389.150 ;
      RECT 309.400 370.790 309.780 396.440 ;
      RECT 313.480 389.150 313.860 391.380 ;
      RECT 313.505 388.985 313.835 389.150 ;
      RECT 316.200 370.790 316.580 396.440 ;
      RECT 320.280 389.150 320.660 391.380 ;
      RECT 320.305 388.985 320.635 389.150 ;
      RECT 321.640 370.790 322.020 396.440 ;
      RECT 327.760 370.790 328.140 396.440 ;
      RECT 329.800 389.150 330.180 391.380 ;
      RECT 329.825 388.985 330.155 389.150 ;
      RECT 334.560 370.790 334.940 396.440 ;
      RECT 338.640 389.150 339.020 391.380 ;
      RECT 346.120 389.150 346.500 391.380 ;
      RECT 355.640 389.150 356.020 391.380 ;
      RECT 363.800 389.150 364.180 391.380 ;
      RECT 371.960 389.150 372.340 391.380 ;
      RECT 380.800 389.150 381.180 391.380 ;
      RECT 388.280 389.150 388.660 391.380 ;
      RECT 338.665 388.985 338.995 389.150 ;
      RECT 346.145 388.985 346.475 389.150 ;
      RECT 355.665 388.985 355.995 389.150 ;
      RECT 363.825 388.985 364.155 389.150 ;
      RECT 371.985 388.985 372.315 389.150 ;
      RECT 380.825 388.985 381.155 389.150 ;
      RECT 388.305 388.985 388.635 389.150 ;
      RECT 394.400 382.350 394.780 394.780 ;
      RECT 396.440 389.150 396.820 391.380 ;
      RECT 396.465 388.985 396.795 389.150 ;
      RECT 394.425 382.185 394.755 382.350 ;
      RECT 396.440 375.550 396.820 388.660 ;
      RECT 397.120 379.630 397.500 396.440 ;
      RECT 405.960 389.150 406.340 391.380 ;
      RECT 405.985 388.985 406.315 389.150 ;
      RECT 409.385 388.470 409.715 388.635 ;
      RECT 397.145 379.465 397.475 379.630 ;
      RECT 409.360 378.760 409.740 388.470 ;
      RECT 410.720 385.750 411.100 394.780 ;
      RECT 413.440 389.150 413.820 391.380 ;
      RECT 422.280 389.150 422.660 391.380 ;
      RECT 431.120 389.150 431.500 391.380 ;
      RECT 438.600 389.150 438.980 391.380 ;
      RECT 448.120 389.150 448.500 391.380 ;
      RECT 413.465 388.985 413.795 389.150 ;
      RECT 422.305 388.985 422.635 389.150 ;
      RECT 431.145 388.985 431.475 389.150 ;
      RECT 438.625 388.985 438.955 389.150 ;
      RECT 448.145 388.985 448.475 389.150 ;
      RECT 410.745 385.585 411.075 385.750 ;
      RECT 410.065 385.070 410.395 385.235 ;
      RECT 396.465 375.385 396.795 375.550 ;
      RECT 153.025 370.625 153.355 370.790 ;
      RECT 159.825 370.625 160.155 370.790 ;
      RECT 165.945 370.625 166.275 370.790 ;
      RECT 172.745 370.625 173.075 370.790 ;
      RECT 178.865 370.625 179.195 370.790 ;
      RECT 184.305 370.625 184.635 370.790 ;
      RECT 191.105 370.625 191.435 370.790 ;
      RECT 196.545 370.625 196.875 370.790 ;
      RECT 203.345 370.625 203.675 370.790 ;
      RECT 209.465 370.625 209.795 370.790 ;
      RECT 216.265 370.625 216.595 370.790 ;
      RECT 221.705 370.625 222.035 370.790 ;
      RECT 227.825 370.625 228.155 370.790 ;
      RECT 234.625 370.625 234.955 370.790 ;
      RECT 240.745 370.625 241.075 370.790 ;
      RECT 247.545 370.625 247.875 370.790 ;
      RECT 252.985 370.625 253.315 370.790 ;
      RECT 259.785 370.625 260.115 370.790 ;
      RECT 265.225 370.625 265.555 370.790 ;
      RECT 271.345 370.625 271.675 370.790 ;
      RECT 278.145 370.625 278.475 370.790 ;
      RECT 284.265 370.625 284.595 370.790 ;
      RECT 291.065 370.625 291.395 370.790 ;
      RECT 296.505 370.625 296.835 370.790 ;
      RECT 303.305 370.625 303.635 370.790 ;
      RECT 309.425 370.625 309.755 370.790 ;
      RECT 316.225 370.625 316.555 370.790 ;
      RECT 321.665 370.625 321.995 370.790 ;
      RECT 327.785 370.625 328.115 370.790 ;
      RECT 334.585 370.625 334.915 370.790 ;
      RECT 155.745 370.110 156.075 370.275 ;
      RECT 142.800 365.350 143.180 368.940 ;
      RECT 148.920 365.350 149.300 368.940 ;
      RECT 155.040 365.350 155.420 368.940 ;
      RECT 142.825 365.185 143.155 365.350 ;
      RECT 148.945 365.185 149.275 365.350 ;
      RECT 155.065 365.185 155.395 365.350 ;
      RECT 142.825 361.270 143.155 361.435 ;
      RECT 142.800 352.240 143.180 361.270 ;
      RECT 138.040 340.870 138.420 351.940 ;
      RECT 154.360 344.950 154.740 364.180 ;
      RECT 155.720 361.080 156.100 370.110 ;
      RECT 160.480 365.350 160.860 368.940 ;
      RECT 167.280 365.350 167.660 368.940 ;
      RECT 173.400 365.350 173.780 368.940 ;
      RECT 180.200 365.350 180.580 368.940 ;
      RECT 186.320 365.350 186.700 368.940 ;
      RECT 192.440 365.350 192.820 368.940 ;
      RECT 198.560 365.350 198.940 368.940 ;
      RECT 204.000 365.350 204.380 368.940 ;
      RECT 210.145 368.750 210.475 368.915 ;
      RECT 160.505 365.185 160.835 365.350 ;
      RECT 167.305 365.185 167.635 365.350 ;
      RECT 173.425 365.185 173.755 365.350 ;
      RECT 180.225 365.185 180.555 365.350 ;
      RECT 186.345 365.185 186.675 365.350 ;
      RECT 192.465 365.185 192.795 365.350 ;
      RECT 198.585 365.185 198.915 365.350 ;
      RECT 204.025 365.185 204.355 365.350 ;
      RECT 210.120 365.160 210.500 368.750 ;
      RECT 211.480 365.350 211.860 368.940 ;
      RECT 216.920 365.350 217.300 368.940 ;
      RECT 223.720 365.350 224.100 368.940 ;
      RECT 229.840 365.350 230.220 368.940 ;
      RECT 235.960 365.350 236.340 368.940 ;
      RECT 242.760 365.350 243.140 368.940 ;
      RECT 248.880 365.350 249.260 368.940 ;
      RECT 255.000 365.350 255.380 368.940 ;
      RECT 260.440 365.350 260.820 368.940 ;
      RECT 267.240 365.350 267.620 368.940 ;
      RECT 273.360 365.350 273.740 368.940 ;
      RECT 280.160 365.350 280.540 368.940 ;
      RECT 286.280 365.350 286.660 368.940 ;
      RECT 292.400 365.350 292.780 368.940 ;
      RECT 298.520 365.350 298.900 368.940 ;
      RECT 303.960 365.350 304.340 368.940 ;
      RECT 310.760 365.350 311.140 368.940 ;
      RECT 317.560 365.350 317.940 368.940 ;
      RECT 323.680 365.350 324.060 368.940 ;
      RECT 329.800 365.350 330.180 368.940 ;
      RECT 335.920 365.350 336.300 368.940 ;
      RECT 211.505 365.185 211.835 365.350 ;
      RECT 216.945 365.185 217.275 365.350 ;
      RECT 223.745 365.185 224.075 365.350 ;
      RECT 229.865 365.185 230.195 365.350 ;
      RECT 235.985 365.185 236.315 365.350 ;
      RECT 242.785 365.185 243.115 365.350 ;
      RECT 248.905 365.185 249.235 365.350 ;
      RECT 255.025 365.185 255.355 365.350 ;
      RECT 260.465 365.185 260.795 365.350 ;
      RECT 267.265 365.185 267.595 365.350 ;
      RECT 273.385 365.185 273.715 365.350 ;
      RECT 280.185 365.185 280.515 365.350 ;
      RECT 286.305 365.185 286.635 365.350 ;
      RECT 292.425 365.185 292.755 365.350 ;
      RECT 298.545 365.185 298.875 365.350 ;
      RECT 303.985 365.185 304.315 365.350 ;
      RECT 310.785 365.185 311.115 365.350 ;
      RECT 317.585 365.185 317.915 365.350 ;
      RECT 323.705 365.185 324.035 365.350 ;
      RECT 329.825 365.185 330.155 365.350 ;
      RECT 335.945 365.185 336.275 365.350 ;
      RECT 374.025 364.670 374.355 364.835 ;
      RECT 409.360 364.670 409.740 378.460 ;
      RECT 410.040 371.280 410.420 385.070 ;
      RECT 450.160 382.350 450.540 396.440 ;
      RECT 456.280 389.150 456.660 391.380 ;
      RECT 464.440 389.150 464.820 391.380 ;
      RECT 456.305 388.985 456.635 389.150 ;
      RECT 464.465 388.985 464.795 389.150 ;
      RECT 450.185 382.185 450.515 382.350 ;
      RECT 344.785 351.750 345.115 351.915 ;
      RECT 154.385 344.785 154.715 344.950 ;
      RECT 141.465 343.590 141.795 343.755 ;
      RECT 146.225 343.590 146.555 343.755 ;
      RECT 141.440 341.360 141.820 343.590 ;
      RECT 138.065 340.705 138.395 340.870 ;
      RECT 146.200 340.680 146.580 343.590 ;
      RECT 151.640 341.550 152.020 343.780 ;
      RECT 153.025 343.590 153.355 343.755 ;
      RECT 151.665 341.385 151.995 341.550 ;
      RECT 153.000 341.360 153.380 343.590 ;
      RECT 157.760 341.550 158.140 343.780 ;
      RECT 158.465 343.590 158.795 343.755 ;
      RECT 157.785 341.385 158.115 341.550 ;
      RECT 158.440 341.360 158.820 343.590 ;
      RECT 163.880 341.550 164.260 343.780 ;
      RECT 166.625 343.590 166.955 343.755 ;
      RECT 163.905 341.385 164.235 341.550 ;
      RECT 166.600 341.360 166.980 343.590 ;
      RECT 170.680 341.550 171.060 343.780 ;
      RECT 176.120 341.550 176.500 343.780 ;
      RECT 178.865 343.590 179.195 343.755 ;
      RECT 170.705 341.385 171.035 341.550 ;
      RECT 176.145 341.385 176.475 341.550 ;
      RECT 178.840 341.360 179.220 343.590 ;
      RECT 182.920 341.550 183.300 343.780 ;
      RECT 189.040 341.550 189.420 343.780 ;
      RECT 191.785 343.590 192.115 343.755 ;
      RECT 182.945 341.385 183.275 341.550 ;
      RECT 189.065 341.385 189.395 341.550 ;
      RECT 191.760 341.360 192.140 343.590 ;
      RECT 195.160 341.550 195.540 343.780 ;
      RECT 196.545 343.590 196.875 343.755 ;
      RECT 195.185 341.385 195.515 341.550 ;
      RECT 196.520 341.360 196.900 343.590 ;
      RECT 201.280 341.550 201.660 343.780 ;
      RECT 209.440 341.550 209.820 343.780 ;
      RECT 214.200 341.550 214.580 343.780 ;
      RECT 216.945 343.590 217.275 343.755 ;
      RECT 201.305 341.385 201.635 341.550 ;
      RECT 209.465 341.385 209.795 341.550 ;
      RECT 214.225 341.385 214.555 341.550 ;
      RECT 216.920 341.360 217.300 343.590 ;
      RECT 220.320 341.550 220.700 343.780 ;
      RECT 229.185 343.590 229.515 343.755 ;
      RECT 220.345 341.385 220.675 341.550 ;
      RECT 229.160 341.360 229.540 343.590 ;
      RECT 232.560 341.550 232.940 343.780 ;
      RECT 235.305 343.590 235.635 343.755 ;
      RECT 232.585 341.385 232.915 341.550 ;
      RECT 235.280 341.360 235.660 343.590 ;
      RECT 238.680 341.550 239.060 343.780 ;
      RECT 244.800 341.550 245.180 343.780 ;
      RECT 252.960 341.550 253.340 343.780 ;
      RECT 257.720 341.550 258.100 343.780 ;
      RECT 260.465 343.590 260.795 343.755 ;
      RECT 238.705 341.385 239.035 341.550 ;
      RECT 244.825 341.385 245.155 341.550 ;
      RECT 252.985 341.385 253.315 341.550 ;
      RECT 257.745 341.385 258.075 341.550 ;
      RECT 260.440 341.360 260.820 343.590 ;
      RECT 263.840 341.550 264.220 343.780 ;
      RECT 265.225 343.590 265.555 343.755 ;
      RECT 263.865 341.385 264.195 341.550 ;
      RECT 265.200 341.360 265.580 343.590 ;
      RECT 269.960 341.550 270.340 343.780 ;
      RECT 276.080 341.550 276.460 343.780 ;
      RECT 278.825 343.590 279.155 343.755 ;
      RECT 269.985 341.385 270.315 341.550 ;
      RECT 276.105 341.385 276.435 341.550 ;
      RECT 278.800 341.360 279.180 343.590 ;
      RECT 284.240 341.550 284.620 343.780 ;
      RECT 289.000 341.550 289.380 343.780 ;
      RECT 289.705 343.590 290.035 343.755 ;
      RECT 284.265 341.385 284.595 341.550 ;
      RECT 289.025 341.385 289.355 341.550 ;
      RECT 289.680 341.360 290.060 343.590 ;
      RECT 295.120 341.550 295.500 343.780 ;
      RECT 297.865 343.590 298.195 343.755 ;
      RECT 295.145 341.385 295.475 341.550 ;
      RECT 297.840 341.360 298.220 343.590 ;
      RECT 301.240 341.550 301.620 343.780 ;
      RECT 303.985 343.590 304.315 343.755 ;
      RECT 301.265 341.385 301.595 341.550 ;
      RECT 303.960 341.360 304.340 343.590 ;
      RECT 307.360 341.550 307.740 343.780 ;
      RECT 313.480 341.550 313.860 343.780 ;
      RECT 320.280 341.550 320.660 343.780 ;
      RECT 326.400 341.550 326.780 343.780 ;
      RECT 332.520 341.550 332.900 343.780 ;
      RECT 335.265 343.590 335.595 343.755 ;
      RECT 307.385 341.385 307.715 341.550 ;
      RECT 313.505 341.385 313.835 341.550 ;
      RECT 320.305 341.385 320.635 341.550 ;
      RECT 326.425 341.385 326.755 341.550 ;
      RECT 332.545 341.385 332.875 341.550 ;
      RECT 335.240 341.360 335.620 343.590 ;
      RECT 338.640 341.550 339.020 343.780 ;
      RECT 341.385 343.590 341.715 343.755 ;
      RECT 338.665 341.385 338.995 341.550 ;
      RECT 341.360 341.360 341.740 343.590 ;
      RECT 134.665 340.190 134.995 340.355 ;
      RECT 134.640 338.640 135.020 340.190 ;
      RECT 344.760 338.640 345.140 351.750 ;
      RECT 351.585 341.550 351.915 341.715 ;
      RECT 346.800 338.830 347.180 340.380 ;
      RECT 351.560 340.000 351.940 341.550 ;
      RECT 369.265 338.830 369.595 338.995 ;
      RECT 346.825 338.665 347.155 338.830 ;
      RECT 369.240 336.600 369.620 338.830 ;
      RECT 372.640 336.790 373.020 351.260 ;
      RECT 373.320 340.190 373.700 358.060 ;
      RECT 374.000 351.560 374.380 364.670 ;
      RECT 409.385 364.505 409.715 364.670 ;
      RECT 410.040 357.870 410.420 370.980 ;
      RECT 410.745 363.990 411.075 364.155 ;
      RECT 410.065 357.705 410.395 357.870 ;
      RECT 410.065 357.190 410.395 357.355 ;
      RECT 410.040 343.400 410.420 357.190 ;
      RECT 410.720 350.200 411.100 363.990 ;
      RECT 470.585 357.190 470.915 357.355 ;
      RECT 470.560 354.960 470.940 357.190 ;
      RECT 462.425 349.710 462.755 349.875 ;
      RECT 373.345 340.025 373.675 340.190 ;
      RECT 372.665 336.625 372.995 336.790 ;
      RECT 102.000 333.390 102.380 334.940 ;
      RECT 104.720 334.750 105.100 336.300 ;
      RECT 105.400 334.750 105.780 336.300 ;
      RECT 106.785 336.110 107.115 336.275 ;
      RECT 108.825 336.110 109.155 336.275 ;
      RECT 110.185 336.110 110.515 336.275 ;
      RECT 369.945 336.110 370.275 336.275 ;
      RECT 104.745 334.585 105.075 334.750 ;
      RECT 105.425 334.585 105.755 334.750 ;
      RECT 106.760 334.560 107.140 336.110 ;
      RECT 108.800 334.560 109.180 336.110 ;
      RECT 110.160 334.560 110.540 336.110 ;
      RECT 102.025 333.225 102.355 333.390 ;
      RECT 108.120 332.710 108.500 334.260 ;
      RECT 110.160 332.710 110.540 334.260 ;
      RECT 136.000 334.070 136.380 335.620 ;
      RECT 345.440 334.070 345.820 335.620 ;
      RECT 369.920 334.560 370.300 336.110 ;
      RECT 371.960 334.750 372.340 336.300 ;
      RECT 373.345 336.110 373.675 336.275 ;
      RECT 371.985 334.585 372.315 334.750 ;
      RECT 373.320 334.560 373.700 336.110 ;
      RECT 462.400 335.920 462.780 349.710 ;
      RECT 467.120 347.985 467.450 348.315 ;
      RECT 462.400 335.240 463.460 335.620 ;
      RECT 369.945 334.070 370.275 334.235 ;
      RECT 136.025 333.905 136.355 334.070 ;
      RECT 345.465 333.905 345.795 334.070 ;
      RECT 108.145 332.545 108.475 332.710 ;
      RECT 110.185 332.545 110.515 332.710 ;
      RECT 102.680 329.310 103.060 330.860 ;
      RECT 344.760 329.990 345.140 331.540 ;
      RECT 345.440 331.350 345.820 332.900 ;
      RECT 369.920 332.520 370.300 334.070 ;
      RECT 371.280 332.710 371.660 334.260 ;
      RECT 378.080 333.390 378.460 334.940 ;
      RECT 378.105 333.225 378.435 333.390 ;
      RECT 371.305 332.545 371.635 332.710 ;
      RECT 345.465 331.185 345.795 331.350 ;
      RECT 375.360 330.670 375.740 332.220 ;
      RECT 375.385 330.505 375.715 330.670 ;
      RECT 344.785 329.825 345.115 329.990 ;
      RECT 134.665 329.310 134.995 329.475 ;
      RECT 344.785 329.310 345.115 329.475 ;
      RECT 377.400 329.310 377.780 330.860 ;
      RECT 102.705 329.145 103.035 329.310 ;
      RECT 102.000 327.270 102.380 328.820 ;
      RECT 104.040 327.270 104.420 328.820 ;
      RECT 134.640 327.760 135.020 329.310 ;
      RECT 344.760 327.760 345.140 329.310 ;
      RECT 377.425 329.145 377.755 329.310 ;
      RECT 373.345 328.630 373.675 328.795 ;
      RECT 102.025 327.105 102.355 327.270 ;
      RECT 104.065 327.105 104.395 327.270 ;
      RECT 102.000 325.230 102.380 326.780 ;
      RECT 108.800 325.230 109.180 326.780 ;
      RECT 110.160 325.230 110.540 326.780 ;
      RECT 136.000 325.910 136.380 327.460 ;
      RECT 373.320 327.080 373.700 328.630 ;
      RECT 374.680 327.270 375.060 328.820 ;
      RECT 377.425 328.630 377.755 328.795 ;
      RECT 374.705 327.105 375.035 327.270 ;
      RECT 377.400 327.080 377.780 328.630 ;
      RECT 369.265 326.590 369.595 326.755 ;
      RECT 136.025 325.745 136.355 325.910 ;
      RECT 102.025 325.065 102.355 325.230 ;
      RECT 108.825 325.065 109.155 325.230 ;
      RECT 110.185 325.065 110.515 325.230 ;
      RECT 369.240 325.040 369.620 326.590 ;
      RECT 371.280 325.230 371.660 326.780 ;
      RECT 378.105 326.590 378.435 326.755 ;
      RECT 371.305 325.065 371.635 325.230 ;
      RECT 378.080 325.040 378.460 326.590 ;
      RECT 102.025 324.550 102.355 324.715 ;
      RECT 102.000 323.000 102.380 324.550 ;
      RECT 107.440 323.190 107.820 324.740 ;
      RECT 108.825 324.550 109.155 324.715 ;
      RECT 110.185 324.550 110.515 324.715 ;
      RECT 107.465 323.025 107.795 323.190 ;
      RECT 108.800 323.000 109.180 324.550 ;
      RECT 110.160 323.000 110.540 324.550 ;
      RECT 369.920 323.190 370.300 324.740 ;
      RECT 371.305 324.550 371.635 324.715 ;
      RECT 375.385 324.550 375.715 324.715 ;
      RECT 377.425 324.550 377.755 324.715 ;
      RECT 369.945 323.025 370.275 323.190 ;
      RECT 371.280 323.000 371.660 324.550 ;
      RECT 375.360 323.000 375.740 324.550 ;
      RECT 377.400 323.000 377.780 324.550 ;
      RECT 102.680 321.150 103.060 322.700 ;
      RECT 104.065 322.510 104.395 322.675 ;
      RECT 102.705 320.985 103.035 321.150 ;
      RECT 104.040 320.960 104.420 322.510 ;
      RECT 107.440 321.150 107.820 322.700 ;
      RECT 108.120 321.150 108.500 322.700 ;
      RECT 110.185 322.510 110.515 322.675 ;
      RECT 369.265 322.510 369.595 322.675 ;
      RECT 107.465 320.985 107.795 321.150 ;
      RECT 108.145 320.985 108.475 321.150 ;
      RECT 110.160 320.960 110.540 322.510 ;
      RECT 369.240 320.960 369.620 322.510 ;
      RECT 371.960 321.150 372.340 322.700 ;
      RECT 374.000 321.150 374.380 322.700 ;
      RECT 378.080 321.150 378.460 322.700 ;
      RECT 462.400 322.510 462.780 335.240 ;
      RECT 462.425 322.345 462.755 322.510 ;
      RECT 371.985 320.985 372.315 321.150 ;
      RECT 374.025 320.985 374.355 321.150 ;
      RECT 378.105 320.985 378.435 321.150 ;
      RECT 102.680 319.110 103.060 320.660 ;
      RECT 104.720 319.110 105.100 320.660 ;
      RECT 105.400 319.110 105.780 320.660 ;
      RECT 106.105 320.470 106.435 320.635 ;
      RECT 102.705 318.945 103.035 319.110 ;
      RECT 104.745 318.945 105.075 319.110 ;
      RECT 105.425 318.945 105.755 319.110 ;
      RECT 106.080 318.920 106.460 320.470 ;
      RECT 108.800 319.110 109.180 320.660 ;
      RECT 110.160 319.110 110.540 320.660 ;
      RECT 369.920 319.110 370.300 320.660 ;
      RECT 371.985 320.470 372.315 320.635 ;
      RECT 378.105 320.470 378.435 320.635 ;
      RECT 108.825 318.945 109.155 319.110 ;
      RECT 110.185 318.945 110.515 319.110 ;
      RECT 369.945 318.945 370.275 319.110 ;
      RECT 371.960 318.920 372.340 320.470 ;
      RECT 378.080 318.920 378.460 320.470 ;
      RECT 102.705 318.430 103.035 318.595 ;
      RECT 102.680 316.880 103.060 318.430 ;
      RECT 104.040 317.070 104.420 318.620 ;
      RECT 108.825 318.430 109.155 318.595 ;
      RECT 110.185 318.430 110.515 318.595 ;
      RECT 369.945 318.430 370.275 318.595 ;
      RECT 371.305 318.430 371.635 318.595 ;
      RECT 104.065 316.905 104.395 317.070 ;
      RECT 108.800 316.880 109.180 318.430 ;
      RECT 110.160 316.880 110.540 318.430 ;
      RECT 369.920 316.880 370.300 318.430 ;
      RECT 371.280 316.880 371.660 318.430 ;
      RECT 374.680 317.070 375.060 318.620 ;
      RECT 378.080 317.070 378.460 318.620 ;
      RECT 374.705 316.905 375.035 317.070 ;
      RECT 378.105 316.905 378.435 317.070 ;
      RECT 104.065 316.390 104.395 316.555 ;
      RECT 107.465 316.390 107.795 316.555 ;
      RECT 104.040 314.840 104.420 316.390 ;
      RECT 107.440 314.840 107.820 316.390 ;
      RECT 108.120 315.030 108.500 316.580 ;
      RECT 110.840 315.030 111.220 316.580 ;
      RECT 369.265 316.390 369.595 316.555 ;
      RECT 136.025 315.710 136.355 315.875 ;
      RECT 108.145 314.865 108.475 315.030 ;
      RECT 110.865 314.865 111.195 315.030 ;
      RECT 108.825 314.350 109.155 314.515 ;
      RECT 108.800 312.800 109.180 314.350 ;
      RECT 110.840 312.990 111.220 314.540 ;
      RECT 110.865 312.825 111.195 312.990 ;
      RECT 102.680 309.590 103.060 311.140 ;
      RECT 104.040 310.950 104.420 312.500 ;
      RECT 104.065 310.785 104.395 310.950 ;
      RECT 134.640 310.270 135.020 311.820 ;
      RECT 135.320 311.630 135.700 314.540 ;
      RECT 136.000 314.160 136.380 315.710 ;
      RECT 369.240 314.840 369.620 316.390 ;
      RECT 371.960 315.030 372.340 316.580 ;
      RECT 374.000 315.030 374.380 316.580 ;
      RECT 376.040 315.030 376.420 316.580 ;
      RECT 371.985 314.865 372.315 315.030 ;
      RECT 374.025 314.865 374.355 315.030 ;
      RECT 376.065 314.865 376.395 315.030 ;
      RECT 369.920 312.990 370.300 314.540 ;
      RECT 371.960 312.990 372.340 314.540 ;
      RECT 369.945 312.825 370.275 312.990 ;
      RECT 371.985 312.825 372.315 312.990 ;
      RECT 135.345 311.465 135.675 311.630 ;
      RECT 374.680 310.950 375.060 312.500 ;
      RECT 378.105 310.950 378.435 311.115 ;
      RECT 374.705 310.785 375.035 310.950 ;
      RECT 134.665 310.105 134.995 310.270 ;
      RECT 134.665 309.590 134.995 309.755 ;
      RECT 102.705 309.425 103.035 309.590 ;
      RECT 102.025 308.910 102.355 309.075 ;
      RECT 104.745 308.910 105.075 309.075 ;
      RECT 105.425 308.910 105.755 309.075 ;
      RECT 102.000 307.360 102.380 308.910 ;
      RECT 104.720 307.360 105.100 308.910 ;
      RECT 105.400 307.360 105.780 308.910 ;
      RECT 134.640 308.040 135.020 309.590 ;
      RECT 344.760 308.230 345.140 309.780 ;
      RECT 378.080 309.400 378.460 310.950 ;
      RECT 373.345 308.910 373.675 309.075 ;
      RECT 344.785 308.065 345.115 308.230 ;
      RECT 102.705 306.870 103.035 307.035 ;
      RECT 102.680 305.320 103.060 306.870 ;
      RECT 108.120 305.510 108.500 307.060 ;
      RECT 110.160 305.510 110.540 307.060 ;
      RECT 136.000 306.190 136.380 307.740 ;
      RECT 373.320 307.360 373.700 308.910 ;
      RECT 375.360 307.550 375.740 309.100 ;
      RECT 377.400 307.550 377.780 309.100 ;
      RECT 375.385 307.385 375.715 307.550 ;
      RECT 377.425 307.385 377.755 307.550 ;
      RECT 369.945 306.870 370.275 307.035 ;
      RECT 136.025 306.025 136.355 306.190 ;
      RECT 108.145 305.345 108.475 305.510 ;
      RECT 110.185 305.345 110.515 305.510 ;
      RECT 369.920 305.320 370.300 306.870 ;
      RECT 371.280 305.510 371.660 307.060 ;
      RECT 378.080 305.510 378.460 307.060 ;
      RECT 371.305 305.345 371.635 305.510 ;
      RECT 378.105 305.345 378.435 305.510 ;
      RECT 102.025 304.830 102.355 304.995 ;
      RECT 102.000 303.280 102.380 304.830 ;
      RECT 105.400 303.470 105.780 305.020 ;
      RECT 106.760 303.470 107.140 305.020 ;
      RECT 108.145 304.830 108.475 304.995 ;
      RECT 105.425 303.305 105.755 303.470 ;
      RECT 106.785 303.305 107.115 303.470 ;
      RECT 108.120 303.280 108.500 304.830 ;
      RECT 110.160 303.470 110.540 305.020 ;
      RECT 369.920 303.470 370.300 305.020 ;
      RECT 371.305 304.830 371.635 304.995 ;
      RECT 110.185 303.305 110.515 303.470 ;
      RECT 369.945 303.305 370.275 303.470 ;
      RECT 371.280 303.280 371.660 304.830 ;
      RECT 375.360 303.470 375.740 305.020 ;
      RECT 378.105 304.830 378.435 304.995 ;
      RECT 375.385 303.305 375.715 303.470 ;
      RECT 378.080 303.280 378.460 304.830 ;
      RECT 102.680 301.430 103.060 302.980 ;
      RECT 104.745 302.790 105.075 302.955 ;
      RECT 105.425 302.790 105.755 302.955 ;
      RECT 102.705 301.265 103.035 301.430 ;
      RECT 104.720 301.240 105.100 302.790 ;
      RECT 105.400 301.240 105.780 302.790 ;
      RECT 108.800 301.430 109.180 302.980 ;
      RECT 110.185 302.790 110.515 302.955 ;
      RECT 369.945 302.790 370.275 302.955 ;
      RECT 108.825 301.265 109.155 301.430 ;
      RECT 110.160 301.240 110.540 302.790 ;
      RECT 369.920 301.240 370.300 302.790 ;
      RECT 371.960 301.430 372.340 302.980 ;
      RECT 373.345 302.790 373.675 302.955 ;
      RECT 371.985 301.265 372.315 301.430 ;
      RECT 373.320 301.240 373.700 302.790 ;
      RECT 374.680 301.430 375.060 302.980 ;
      RECT 377.400 301.430 377.780 302.980 ;
      RECT 374.705 301.265 375.035 301.430 ;
      RECT 377.425 301.265 377.755 301.430 ;
      RECT 102.680 299.390 103.060 300.940 ;
      RECT 106.785 300.750 107.115 300.915 ;
      RECT 102.705 299.225 103.035 299.390 ;
      RECT 106.760 299.200 107.140 300.750 ;
      RECT 108.120 299.390 108.500 300.940 ;
      RECT 110.840 299.390 111.220 300.940 ;
      RECT 369.240 299.390 369.620 300.940 ;
      RECT 371.305 300.750 371.635 300.915 ;
      RECT 374.025 300.750 374.355 300.915 ;
      RECT 108.145 299.225 108.475 299.390 ;
      RECT 110.865 299.225 111.195 299.390 ;
      RECT 369.265 299.225 369.595 299.390 ;
      RECT 371.280 299.200 371.660 300.750 ;
      RECT 374.000 299.200 374.380 300.750 ;
      RECT 378.080 299.390 378.460 300.940 ;
      RECT 378.105 299.225 378.435 299.390 ;
      RECT 102.680 297.350 103.060 298.900 ;
      RECT 104.065 298.710 104.395 298.875 ;
      RECT 102.705 297.185 103.035 297.350 ;
      RECT 104.040 297.160 104.420 298.710 ;
      RECT 105.400 297.350 105.780 298.900 ;
      RECT 107.440 297.350 107.820 298.900 ;
      RECT 108.145 298.710 108.475 298.875 ;
      RECT 105.425 297.185 105.755 297.350 ;
      RECT 107.465 297.185 107.795 297.350 ;
      RECT 108.120 297.160 108.500 298.710 ;
      RECT 110.160 297.350 110.540 298.900 ;
      RECT 369.265 298.710 369.595 298.875 ;
      RECT 110.185 297.185 110.515 297.350 ;
      RECT 369.240 297.160 369.620 298.710 ;
      RECT 371.960 297.350 372.340 298.900 ;
      RECT 373.320 297.350 373.700 298.900 ;
      RECT 378.105 298.710 378.435 298.875 ;
      RECT 371.985 297.185 372.315 297.350 ;
      RECT 373.345 297.185 373.675 297.350 ;
      RECT 378.080 297.160 378.460 298.710 ;
      RECT 104.745 296.670 105.075 296.835 ;
      RECT 105.425 296.670 105.755 296.835 ;
      RECT 104.720 295.120 105.100 296.670 ;
      RECT 105.400 295.120 105.780 296.670 ;
      RECT 108.120 295.310 108.500 296.860 ;
      RECT 110.185 296.670 110.515 296.835 ;
      RECT 108.145 295.145 108.475 295.310 ;
      RECT 110.160 295.120 110.540 296.670 ;
      RECT 369.240 295.310 369.620 296.860 ;
      RECT 371.985 296.670 372.315 296.835 ;
      RECT 375.385 296.670 375.715 296.835 ;
      RECT 369.265 295.145 369.595 295.310 ;
      RECT 371.960 295.120 372.340 296.670 ;
      RECT 375.360 295.120 375.740 296.670 ;
      RECT 108.120 293.270 108.500 294.820 ;
      RECT 110.840 293.270 111.220 294.820 ;
      RECT 369.265 294.630 369.595 294.795 ;
      RECT 371.305 294.630 371.635 294.795 ;
      RECT 108.145 293.105 108.475 293.270 ;
      RECT 110.865 293.105 111.195 293.270 ;
      RECT 369.240 293.080 369.620 294.630 ;
      RECT 371.280 293.080 371.660 294.630 ;
      RECT 459.680 293.950 460.060 307.740 ;
      RECT 467.135 297.140 467.435 347.985 ;
      RECT 470.560 343.590 470.940 345.820 ;
      RECT 470.585 343.425 470.915 343.590 ;
      RECT 470.585 314.350 470.915 314.515 ;
      RECT 470.560 312.800 470.940 314.350 ;
      RECT 470.560 301.430 470.940 304.340 ;
      RECT 470.585 301.265 470.915 301.430 ;
      RECT 467.120 296.810 467.450 297.140 ;
      RECT 459.705 293.785 460.035 293.950 ;
      RECT 104.065 292.590 104.395 292.755 ;
      RECT 105.425 292.590 105.755 292.755 ;
      RECT 102.025 291.230 102.355 291.395 ;
      RECT 102.000 289.680 102.380 291.230 ;
      RECT 104.040 291.040 104.420 292.590 ;
      RECT 105.400 291.040 105.780 292.590 ;
      RECT 108.800 291.230 109.180 292.780 ;
      RECT 110.840 291.230 111.220 292.780 ;
      RECT 108.825 291.065 109.155 291.230 ;
      RECT 110.865 291.065 111.195 291.230 ;
      RECT 134.640 290.550 135.020 292.100 ;
      RECT 344.785 291.910 345.115 292.075 ;
      RECT 136.025 290.550 136.355 290.715 ;
      RECT 134.665 290.385 134.995 290.550 ;
      RECT 102.680 287.830 103.060 289.380 ;
      RECT 104.065 289.190 104.395 289.355 ;
      RECT 102.705 287.665 103.035 287.830 ;
      RECT 104.040 287.640 104.420 289.190 ;
      RECT 136.000 288.320 136.380 290.550 ;
      RECT 344.760 290.360 345.140 291.910 ;
      RECT 369.920 291.230 370.300 292.780 ;
      RECT 371.960 291.230 372.340 292.780 ;
      RECT 373.320 291.230 373.700 292.780 ;
      RECT 369.945 291.065 370.275 291.230 ;
      RECT 371.985 291.065 372.315 291.230 ;
      RECT 373.345 291.065 373.675 291.230 ;
      RECT 345.440 288.510 345.820 290.060 ;
      RECT 374.680 289.190 375.060 290.740 ;
      RECT 378.080 289.870 378.460 291.420 ;
      RECT 378.105 289.705 378.435 289.870 ;
      RECT 376.065 289.190 376.395 289.355 ;
      RECT 378.105 289.190 378.435 289.355 ;
      RECT 374.705 289.025 375.035 289.190 ;
      RECT 345.465 288.345 345.795 288.510 ;
      RECT 376.040 287.640 376.420 289.190 ;
      RECT 378.080 287.640 378.460 289.190 ;
      RECT 102.680 285.790 103.060 287.340 ;
      RECT 377.400 285.790 377.780 287.340 ;
      RECT 102.705 285.625 103.035 285.790 ;
      RECT 377.425 285.625 377.755 285.790 ;
      RECT 102.705 285.110 103.035 285.275 ;
      RECT 107.465 285.110 107.795 285.275 ;
      RECT 102.680 283.560 103.060 285.110 ;
      RECT 107.440 283.560 107.820 285.110 ;
      RECT 108.120 283.750 108.500 285.300 ;
      RECT 110.865 285.110 111.195 285.275 ;
      RECT 108.145 283.585 108.475 283.750 ;
      RECT 110.840 283.560 111.220 285.110 ;
      RECT 102.000 281.710 102.380 283.260 ;
      RECT 104.720 281.710 105.100 283.260 ;
      RECT 108.145 283.070 108.475 283.235 ;
      RECT 102.025 281.545 102.355 281.710 ;
      RECT 104.745 281.545 105.075 281.710 ;
      RECT 108.120 281.520 108.500 283.070 ;
      RECT 110.160 281.710 110.540 283.260 ;
      RECT 136.000 282.390 136.380 283.940 ;
      RECT 369.240 283.750 369.620 285.300 ;
      RECT 371.280 283.750 371.660 285.300 ;
      RECT 374.000 283.750 374.380 285.300 ;
      RECT 374.680 283.750 375.060 285.300 ;
      RECT 377.425 285.110 377.755 285.275 ;
      RECT 369.265 283.585 369.595 283.750 ;
      RECT 371.305 283.585 371.635 283.750 ;
      RECT 374.025 283.585 374.355 283.750 ;
      RECT 374.705 283.585 375.035 283.750 ;
      RECT 377.400 283.560 377.780 285.110 ;
      RECT 369.265 283.070 369.595 283.235 ;
      RECT 371.985 283.070 372.315 283.235 ;
      RECT 376.065 283.070 376.395 283.235 ;
      RECT 378.105 283.070 378.435 283.235 ;
      RECT 136.025 282.225 136.355 282.390 ;
      RECT 110.185 281.545 110.515 281.710 ;
      RECT 369.240 281.520 369.620 283.070 ;
      RECT 371.960 281.520 372.340 283.070 ;
      RECT 376.040 281.520 376.420 283.070 ;
      RECT 378.080 281.520 378.460 283.070 ;
      RECT 102.025 281.030 102.355 281.195 ;
      RECT 104.745 281.030 105.075 281.195 ;
      RECT 105.425 281.030 105.755 281.195 ;
      RECT 108.825 281.030 109.155 281.195 ;
      RECT 110.185 281.030 110.515 281.195 ;
      RECT 102.000 279.480 102.380 281.030 ;
      RECT 104.720 279.480 105.100 281.030 ;
      RECT 105.400 279.480 105.780 281.030 ;
      RECT 108.800 279.480 109.180 281.030 ;
      RECT 110.160 279.480 110.540 281.030 ;
      RECT 369.920 279.670 370.300 281.220 ;
      RECT 371.960 279.670 372.340 281.220 ;
      RECT 373.345 281.030 373.675 281.195 ;
      RECT 369.945 279.505 370.275 279.670 ;
      RECT 371.985 279.505 372.315 279.670 ;
      RECT 373.320 279.480 373.700 281.030 ;
      RECT 375.360 279.670 375.740 281.220 ;
      RECT 377.400 279.670 377.780 281.220 ;
      RECT 375.385 279.505 375.715 279.670 ;
      RECT 377.425 279.505 377.755 279.670 ;
      RECT 102.025 278.990 102.355 279.155 ;
      RECT 102.000 277.440 102.380 278.990 ;
      RECT 104.040 277.630 104.420 279.180 ;
      RECT 108.120 277.630 108.500 279.180 ;
      RECT 110.185 278.990 110.515 279.155 ;
      RECT 369.265 278.990 369.595 279.155 ;
      RECT 371.305 278.990 371.635 279.155 ;
      RECT 104.065 277.465 104.395 277.630 ;
      RECT 108.145 277.465 108.475 277.630 ;
      RECT 110.160 277.440 110.540 278.990 ;
      RECT 369.240 277.440 369.620 278.990 ;
      RECT 371.280 277.440 371.660 278.990 ;
      RECT 378.080 277.630 378.460 279.180 ;
      RECT 378.105 277.465 378.435 277.630 ;
      RECT 104.065 276.950 104.395 277.115 ;
      RECT 104.040 275.400 104.420 276.950 ;
      RECT 105.400 275.590 105.780 277.140 ;
      RECT 107.440 275.590 107.820 277.140 ;
      RECT 108.145 276.950 108.475 277.115 ;
      RECT 110.865 276.950 111.195 277.115 ;
      RECT 105.425 275.425 105.755 275.590 ;
      RECT 107.465 275.425 107.795 275.590 ;
      RECT 108.120 275.400 108.500 276.950 ;
      RECT 110.840 275.400 111.220 276.950 ;
      RECT 369.920 275.590 370.300 277.140 ;
      RECT 371.985 276.950 372.315 277.115 ;
      RECT 376.065 276.950 376.395 277.115 ;
      RECT 369.945 275.425 370.275 275.590 ;
      RECT 371.960 275.400 372.340 276.950 ;
      RECT 376.040 275.400 376.420 276.950 ;
      RECT 102.000 273.550 102.380 275.100 ;
      RECT 104.745 274.910 105.075 275.075 ;
      RECT 105.425 274.910 105.755 275.075 ;
      RECT 102.025 273.385 102.355 273.550 ;
      RECT 104.720 273.360 105.100 274.910 ;
      RECT 105.400 273.360 105.780 274.910 ;
      RECT 108.120 273.550 108.500 275.100 ;
      RECT 110.160 273.550 110.540 275.100 ;
      RECT 369.240 273.550 369.620 275.100 ;
      RECT 371.280 273.550 371.660 275.100 ;
      RECT 373.345 274.910 373.675 275.075 ;
      RECT 108.145 273.385 108.475 273.550 ;
      RECT 110.185 273.385 110.515 273.550 ;
      RECT 369.265 273.385 369.595 273.550 ;
      RECT 371.305 273.385 371.635 273.550 ;
      RECT 373.320 273.360 373.700 274.910 ;
      RECT 378.080 273.550 378.460 275.100 ;
      RECT 378.105 273.385 378.435 273.550 ;
      RECT 107.465 272.870 107.795 273.035 ;
      RECT 108.145 272.870 108.475 273.035 ;
      RECT 110.185 272.870 110.515 273.035 ;
      RECT 369.265 272.870 369.595 273.035 ;
      RECT 371.305 272.870 371.635 273.035 ;
      RECT 376.065 272.870 376.395 273.035 ;
      RECT 102.000 270.150 102.380 271.700 ;
      RECT 107.440 271.320 107.820 272.870 ;
      RECT 108.120 271.320 108.500 272.870 ;
      RECT 110.160 271.320 110.540 272.870 ;
      RECT 369.240 271.320 369.620 272.870 ;
      RECT 371.280 271.320 371.660 272.870 ;
      RECT 376.040 271.320 376.420 272.870 ;
      RECT 102.025 269.985 102.355 270.150 ;
      RECT 102.705 269.470 103.035 269.635 ;
      RECT 102.680 267.920 103.060 269.470 ;
      RECT 107.440 268.110 107.820 269.660 ;
      RECT 107.465 267.945 107.795 268.110 ;
      RECT 102.680 266.070 103.060 267.620 ;
      RECT 134.640 266.750 135.020 268.300 ;
      RECT 135.320 268.110 135.700 270.340 ;
      RECT 136.025 270.150 136.355 270.315 ;
      RECT 136.000 268.600 136.380 270.150 ;
      RECT 344.760 268.790 345.140 270.340 ;
      RECT 377.400 270.150 377.780 271.700 ;
      RECT 377.425 269.985 377.755 270.150 ;
      RECT 344.785 268.625 345.115 268.790 ;
      RECT 135.345 267.945 135.675 268.110 ;
      RECT 345.440 266.750 345.820 268.300 ;
      RECT 373.320 268.110 373.700 269.660 ;
      RECT 375.385 269.470 375.715 269.635 ;
      RECT 377.425 269.470 377.755 269.635 ;
      RECT 373.345 267.945 373.675 268.110 ;
      RECT 375.360 267.920 375.740 269.470 ;
      RECT 377.400 267.920 377.780 269.470 ;
      RECT 374.705 267.430 375.035 267.595 ;
      RECT 134.665 266.585 134.995 266.750 ;
      RECT 345.465 266.585 345.795 266.750 ;
      RECT 102.705 265.905 103.035 266.070 ;
      RECT 374.680 265.880 375.060 267.430 ;
      RECT 378.080 266.070 378.460 267.620 ;
      RECT 378.105 265.905 378.435 266.070 ;
      RECT 102.025 265.390 102.355 265.555 ;
      RECT 102.000 263.840 102.380 265.390 ;
      RECT 104.720 264.030 105.100 265.580 ;
      RECT 105.400 264.030 105.780 265.580 ;
      RECT 108.800 264.030 109.180 265.580 ;
      RECT 110.185 265.390 110.515 265.555 ;
      RECT 104.745 263.865 105.075 264.030 ;
      RECT 105.425 263.865 105.755 264.030 ;
      RECT 108.825 263.865 109.155 264.030 ;
      RECT 110.160 263.840 110.540 265.390 ;
      RECT 102.680 261.990 103.060 263.540 ;
      RECT 108.120 261.990 108.500 263.540 ;
      RECT 110.160 261.990 110.540 263.540 ;
      RECT 136.000 262.670 136.380 264.220 ;
      RECT 345.440 262.670 345.820 264.220 ;
      RECT 369.920 264.030 370.300 265.580 ;
      RECT 371.305 265.390 371.635 265.555 ;
      RECT 373.345 265.390 373.675 265.555 ;
      RECT 377.425 265.390 377.755 265.555 ;
      RECT 369.945 263.865 370.275 264.030 ;
      RECT 371.280 263.840 371.660 265.390 ;
      RECT 373.320 263.840 373.700 265.390 ;
      RECT 377.400 263.840 377.780 265.390 ;
      RECT 136.025 262.505 136.355 262.670 ;
      RECT 345.465 262.505 345.795 262.670 ;
      RECT 369.240 261.990 369.620 263.540 ;
      RECT 371.985 263.350 372.315 263.515 ;
      RECT 102.705 261.825 103.035 261.990 ;
      RECT 108.145 261.825 108.475 261.990 ;
      RECT 110.185 261.825 110.515 261.990 ;
      RECT 369.265 261.825 369.595 261.990 ;
      RECT 371.960 261.800 372.340 263.350 ;
      RECT 374.000 261.990 374.380 263.540 ;
      RECT 377.425 263.350 377.755 263.515 ;
      RECT 374.025 261.825 374.355 261.990 ;
      RECT 377.400 261.800 377.780 263.350 ;
      RECT 102.705 261.310 103.035 261.475 ;
      RECT 102.680 259.760 103.060 261.310 ;
      RECT 104.720 259.950 105.100 261.500 ;
      RECT 105.400 259.950 105.780 261.500 ;
      RECT 106.105 261.310 106.435 261.475 ;
      RECT 108.145 261.310 108.475 261.475 ;
      RECT 110.185 261.310 110.515 261.475 ;
      RECT 104.745 259.785 105.075 259.950 ;
      RECT 105.425 259.785 105.755 259.950 ;
      RECT 106.080 259.760 106.460 261.310 ;
      RECT 108.120 259.760 108.500 261.310 ;
      RECT 110.160 259.760 110.540 261.310 ;
      RECT 369.920 259.950 370.300 261.500 ;
      RECT 371.280 259.950 371.660 261.500 ;
      RECT 373.320 259.950 373.700 261.500 ;
      RECT 377.400 259.950 377.780 261.500 ;
      RECT 369.945 259.785 370.275 259.950 ;
      RECT 371.305 259.785 371.635 259.950 ;
      RECT 373.345 259.785 373.675 259.950 ;
      RECT 377.425 259.785 377.755 259.950 ;
      RECT 102.680 257.910 103.060 259.460 ;
      RECT 107.440 257.910 107.820 259.460 ;
      RECT 108.825 259.270 109.155 259.435 ;
      RECT 102.705 257.745 103.035 257.910 ;
      RECT 107.465 257.745 107.795 257.910 ;
      RECT 108.800 257.720 109.180 259.270 ;
      RECT 110.840 257.910 111.220 259.460 ;
      RECT 369.945 259.270 370.275 259.435 ;
      RECT 110.865 257.745 111.195 257.910 ;
      RECT 369.920 257.720 370.300 259.270 ;
      RECT 371.960 257.910 372.340 259.460 ;
      RECT 374.705 259.270 375.035 259.435 ;
      RECT 371.985 257.745 372.315 257.910 ;
      RECT 374.680 257.720 375.060 259.270 ;
      RECT 377.400 257.910 377.780 259.460 ;
      RECT 377.425 257.745 377.755 257.910 ;
      RECT 104.065 257.230 104.395 257.395 ;
      RECT 106.785 257.230 107.115 257.395 ;
      RECT 104.040 255.680 104.420 257.230 ;
      RECT 106.760 255.680 107.140 257.230 ;
      RECT 108.120 255.870 108.500 257.420 ;
      RECT 110.185 257.230 110.515 257.395 ;
      RECT 369.265 257.230 369.595 257.395 ;
      RECT 108.145 255.705 108.475 255.870 ;
      RECT 110.160 255.680 110.540 257.230 ;
      RECT 369.240 255.680 369.620 257.230 ;
      RECT 371.960 255.870 372.340 257.420 ;
      RECT 374.000 255.870 374.380 257.420 ;
      RECT 371.985 255.705 372.315 255.870 ;
      RECT 374.025 255.705 374.355 255.870 ;
      RECT 102.000 253.830 102.380 255.380 ;
      RECT 104.065 255.190 104.395 255.355 ;
      RECT 102.025 253.665 102.355 253.830 ;
      RECT 104.040 253.640 104.420 255.190 ;
      RECT 105.400 253.830 105.780 255.380 ;
      RECT 108.145 255.190 108.475 255.355 ;
      RECT 105.425 253.665 105.755 253.830 ;
      RECT 108.120 253.640 108.500 255.190 ;
      RECT 110.160 253.830 110.540 255.380 ;
      RECT 369.265 255.190 369.595 255.355 ;
      RECT 371.985 255.190 372.315 255.355 ;
      RECT 376.065 255.190 376.395 255.355 ;
      RECT 378.105 255.190 378.435 255.355 ;
      RECT 110.185 253.665 110.515 253.830 ;
      RECT 369.240 253.640 369.620 255.190 ;
      RECT 371.960 253.640 372.340 255.190 ;
      RECT 376.040 253.640 376.420 255.190 ;
      RECT 378.080 253.640 378.460 255.190 ;
      RECT 106.105 253.150 106.435 253.315 ;
      RECT 108.825 253.150 109.155 253.315 ;
      RECT 110.865 253.150 111.195 253.315 ;
      RECT 102.025 251.790 102.355 251.955 ;
      RECT 102.000 250.240 102.380 251.790 ;
      RECT 106.080 251.600 106.460 253.150 ;
      RECT 108.800 251.600 109.180 253.150 ;
      RECT 110.840 251.600 111.220 253.150 ;
      RECT 369.240 251.790 369.620 253.340 ;
      RECT 371.305 253.150 371.635 253.315 ;
      RECT 369.265 251.625 369.595 251.790 ;
      RECT 371.280 251.600 371.660 253.150 ;
      RECT 374.000 251.790 374.380 253.340 ;
      RECT 375.385 253.150 375.715 253.315 ;
      RECT 374.025 251.625 374.355 251.790 ;
      RECT 375.360 251.600 375.740 253.150 ;
      RECT 378.105 251.790 378.435 251.955 ;
      RECT 108.120 249.750 108.500 251.300 ;
      RECT 110.840 249.750 111.220 251.300 ;
      RECT 369.265 251.110 369.595 251.275 ;
      RECT 371.305 251.110 371.635 251.275 ;
      RECT 108.145 249.585 108.475 249.750 ;
      RECT 110.865 249.585 111.195 249.750 ;
      RECT 102.025 247.710 102.355 247.875 ;
      RECT 106.760 247.710 107.140 249.260 ;
      RECT 102.000 246.160 102.380 247.710 ;
      RECT 106.785 247.545 107.115 247.710 ;
      RECT 136.000 247.030 136.380 248.580 ;
      RECT 344.785 248.390 345.115 248.555 ;
      RECT 345.440 248.390 345.820 249.940 ;
      RECT 369.240 249.560 369.620 251.110 ;
      RECT 371.280 249.560 371.660 251.110 ;
      RECT 378.080 250.240 378.460 251.790 ;
      RECT 136.025 246.865 136.355 247.030 ;
      RECT 344.760 246.840 345.140 248.390 ;
      RECT 345.465 248.225 345.795 248.390 ;
      RECT 375.360 247.710 375.740 249.260 ;
      RECT 375.385 247.545 375.715 247.710 ;
      RECT 378.080 246.350 378.460 247.900 ;
      RECT 378.105 246.185 378.435 246.350 ;
      RECT 102.680 244.310 103.060 245.860 ;
      RECT 106.105 245.670 106.435 245.835 ;
      RECT 376.065 245.670 376.395 245.835 ;
      RECT 102.705 244.145 103.035 244.310 ;
      RECT 106.080 244.120 106.460 245.670 ;
      RECT 345.465 244.310 345.795 244.475 ;
      RECT 102.680 242.270 103.060 243.820 ;
      RECT 108.825 243.630 109.155 243.795 ;
      RECT 110.185 243.630 110.515 243.795 ;
      RECT 102.705 242.105 103.035 242.270 ;
      RECT 108.800 242.080 109.180 243.630 ;
      RECT 110.160 242.080 110.540 243.630 ;
      RECT 345.440 242.760 345.820 244.310 ;
      RECT 376.040 244.120 376.420 245.670 ;
      RECT 378.080 244.310 378.460 245.860 ;
      RECT 378.105 244.145 378.435 244.310 ;
      RECT 369.920 242.270 370.300 243.820 ;
      RECT 371.960 242.270 372.340 243.820 ;
      RECT 377.400 242.270 377.780 243.820 ;
      RECT 369.945 242.105 370.275 242.270 ;
      RECT 371.985 242.105 372.315 242.270 ;
      RECT 377.425 242.105 377.755 242.270 ;
      RECT 102.705 241.590 103.035 241.755 ;
      RECT 102.680 240.040 103.060 241.590 ;
      RECT 104.040 240.230 104.420 241.780 ;
      RECT 107.465 241.590 107.795 241.755 ;
      RECT 108.825 241.590 109.155 241.755 ;
      RECT 104.065 240.065 104.395 240.230 ;
      RECT 107.440 240.040 107.820 241.590 ;
      RECT 108.800 240.040 109.180 241.590 ;
      RECT 110.160 240.230 110.540 241.780 ;
      RECT 369.240 240.230 369.620 241.780 ;
      RECT 371.985 241.590 372.315 241.755 ;
      RECT 110.185 240.065 110.515 240.230 ;
      RECT 369.265 240.065 369.595 240.230 ;
      RECT 371.960 240.040 372.340 241.590 ;
      RECT 374.000 240.230 374.380 241.780 ;
      RECT 378.080 240.230 378.460 241.780 ;
      RECT 374.025 240.065 374.355 240.230 ;
      RECT 378.105 240.065 378.435 240.230 ;
      RECT 102.000 238.190 102.380 239.740 ;
      RECT 105.400 238.190 105.780 239.740 ;
      RECT 106.760 238.190 107.140 239.740 ;
      RECT 108.800 238.190 109.180 239.740 ;
      RECT 110.160 238.190 110.540 239.740 ;
      RECT 369.920 238.190 370.300 239.740 ;
      RECT 371.985 239.550 372.315 239.715 ;
      RECT 102.025 238.025 102.355 238.190 ;
      RECT 105.425 238.025 105.755 238.190 ;
      RECT 106.785 238.025 107.115 238.190 ;
      RECT 108.825 238.025 109.155 238.190 ;
      RECT 110.185 238.025 110.515 238.190 ;
      RECT 369.945 238.025 370.275 238.190 ;
      RECT 371.960 238.000 372.340 239.550 ;
      RECT 375.360 238.190 375.740 239.740 ;
      RECT 378.105 239.550 378.435 239.715 ;
      RECT 375.385 238.025 375.715 238.190 ;
      RECT 378.080 238.000 378.460 239.550 ;
      RECT 102.680 236.150 103.060 237.700 ;
      RECT 105.425 237.510 105.755 237.675 ;
      RECT 108.825 237.510 109.155 237.675 ;
      RECT 102.705 235.985 103.035 236.150 ;
      RECT 105.400 235.960 105.780 237.510 ;
      RECT 108.800 235.960 109.180 237.510 ;
      RECT 110.840 236.150 111.220 237.700 ;
      RECT 369.945 237.510 370.275 237.675 ;
      RECT 110.865 235.985 111.195 236.150 ;
      RECT 369.920 235.960 370.300 237.510 ;
      RECT 371.960 236.150 372.340 237.700 ;
      RECT 373.345 237.510 373.675 237.675 ;
      RECT 371.985 235.985 372.315 236.150 ;
      RECT 373.320 235.960 373.700 237.510 ;
      RECT 377.400 236.150 377.780 237.700 ;
      RECT 377.425 235.985 377.755 236.150 ;
      RECT 102.025 235.470 102.355 235.635 ;
      RECT 104.065 235.470 104.395 235.635 ;
      RECT 102.000 233.920 102.380 235.470 ;
      RECT 104.040 233.920 104.420 235.470 ;
      RECT 107.440 234.110 107.820 235.660 ;
      RECT 108.120 234.110 108.500 235.660 ;
      RECT 110.185 235.470 110.515 235.635 ;
      RECT 107.465 233.945 107.795 234.110 ;
      RECT 108.145 233.945 108.475 234.110 ;
      RECT 110.160 233.920 110.540 235.470 ;
      RECT 369.240 234.110 369.620 235.660 ;
      RECT 371.305 235.470 371.635 235.635 ;
      RECT 369.265 233.945 369.595 234.110 ;
      RECT 371.280 233.920 371.660 235.470 ;
      RECT 374.000 234.110 374.380 235.660 ;
      RECT 374.680 234.110 375.060 235.660 ;
      RECT 378.105 235.470 378.435 235.635 ;
      RECT 374.025 233.945 374.355 234.110 ;
      RECT 374.705 233.945 375.035 234.110 ;
      RECT 378.080 233.920 378.460 235.470 ;
      RECT 104.065 233.430 104.395 233.595 ;
      RECT 104.040 231.880 104.420 233.430 ;
      RECT 108.800 232.070 109.180 233.620 ;
      RECT 110.865 233.430 111.195 233.595 ;
      RECT 108.825 231.905 109.155 232.070 ;
      RECT 110.840 231.880 111.220 233.430 ;
      RECT 344.785 232.750 345.115 232.915 ;
      RECT 108.825 231.390 109.155 231.555 ;
      RECT 108.800 229.840 109.180 231.390 ;
      RECT 110.160 230.030 110.540 231.580 ;
      RECT 344.760 231.200 345.140 232.750 ;
      RECT 369.920 232.070 370.300 233.620 ;
      RECT 371.280 232.070 371.660 233.620 ;
      RECT 373.320 232.070 373.700 233.620 ;
      RECT 369.945 231.905 370.275 232.070 ;
      RECT 371.305 231.905 371.635 232.070 ;
      RECT 373.345 231.905 373.675 232.070 ;
      RECT 369.945 231.390 370.275 231.555 ;
      RECT 371.305 231.390 371.635 231.555 ;
      RECT 110.185 229.865 110.515 230.030 ;
      RECT 102.705 227.990 103.035 228.155 ;
      RECT 107.440 227.990 107.820 229.540 ;
      RECT 344.760 228.670 345.140 230.220 ;
      RECT 369.920 229.840 370.300 231.390 ;
      RECT 371.280 229.840 371.660 231.390 ;
      RECT 374.025 229.350 374.355 229.515 ;
      RECT 374.705 229.350 375.035 229.515 ;
      RECT 345.465 228.670 345.795 228.835 ;
      RECT 344.785 228.505 345.115 228.670 ;
      RECT 102.680 226.440 103.060 227.990 ;
      RECT 107.465 227.825 107.795 227.990 ;
      RECT 102.705 225.950 103.035 226.115 ;
      RECT 105.400 225.950 105.780 227.500 ;
      RECT 345.440 227.120 345.820 228.670 ;
      RECT 374.000 227.800 374.380 229.350 ;
      RECT 374.680 227.800 375.060 229.350 ;
      RECT 372.665 227.310 372.995 227.475 ;
      RECT 106.785 225.950 107.115 226.115 ;
      RECT 102.680 224.400 103.060 225.950 ;
      RECT 105.425 225.785 105.755 225.950 ;
      RECT 106.760 224.400 107.140 225.950 ;
      RECT 136.000 225.270 136.380 226.820 ;
      RECT 344.785 226.630 345.115 226.795 ;
      RECT 136.025 225.105 136.355 225.270 ;
      RECT 344.760 225.080 345.140 226.630 ;
      RECT 372.640 225.080 373.020 227.310 ;
      RECT 377.400 226.630 377.780 228.180 ;
      RECT 377.425 226.465 377.755 226.630 ;
      RECT 375.385 225.950 375.715 226.115 ;
      RECT 377.425 225.950 377.755 226.115 ;
      RECT 102.025 223.910 102.355 224.075 ;
      RECT 102.000 222.360 102.380 223.910 ;
      RECT 108.120 222.550 108.500 224.100 ;
      RECT 110.840 222.550 111.220 224.100 ;
      RECT 345.440 223.230 345.820 224.780 ;
      RECT 375.360 224.400 375.740 225.950 ;
      RECT 377.400 224.400 377.780 225.950 ;
      RECT 345.465 223.065 345.795 223.230 ;
      RECT 369.240 222.550 369.620 224.100 ;
      RECT 371.305 223.910 371.635 224.075 ;
      RECT 374.705 223.910 375.035 224.075 ;
      RECT 108.145 222.385 108.475 222.550 ;
      RECT 110.865 222.385 111.195 222.550 ;
      RECT 369.265 222.385 369.595 222.550 ;
      RECT 371.280 222.360 371.660 223.910 ;
      RECT 374.680 222.360 375.060 223.910 ;
      RECT 378.080 222.550 378.460 224.100 ;
      RECT 378.105 222.385 378.435 222.550 ;
      RECT 102.680 220.510 103.060 222.060 ;
      RECT 108.800 220.510 109.180 222.060 ;
      RECT 110.185 221.870 110.515 222.035 ;
      RECT 369.945 221.870 370.275 222.035 ;
      RECT 102.705 220.345 103.035 220.510 ;
      RECT 108.825 220.345 109.155 220.510 ;
      RECT 110.160 220.320 110.540 221.870 ;
      RECT 102.000 218.470 102.380 220.020 ;
      RECT 105.425 219.830 105.755 219.995 ;
      RECT 108.825 219.830 109.155 219.995 ;
      RECT 102.025 218.305 102.355 218.470 ;
      RECT 105.400 218.280 105.780 219.830 ;
      RECT 108.800 218.280 109.180 219.830 ;
      RECT 110.160 218.470 110.540 220.020 ;
      RECT 345.440 219.150 345.820 220.700 ;
      RECT 369.920 220.320 370.300 221.870 ;
      RECT 371.960 220.510 372.340 222.060 ;
      RECT 373.345 221.870 373.675 222.035 ;
      RECT 377.425 221.870 377.755 222.035 ;
      RECT 371.985 220.345 372.315 220.510 ;
      RECT 373.320 220.320 373.700 221.870 ;
      RECT 377.400 220.320 377.780 221.870 ;
      RECT 369.945 219.830 370.275 219.995 ;
      RECT 371.985 219.830 372.315 219.995 ;
      RECT 345.465 218.985 345.795 219.150 ;
      RECT 110.185 218.305 110.515 218.470 ;
      RECT 369.920 218.280 370.300 219.830 ;
      RECT 371.960 218.280 372.340 219.830 ;
      RECT 374.000 218.470 374.380 220.020 ;
      RECT 378.080 218.470 378.460 220.020 ;
      RECT 374.025 218.305 374.355 218.470 ;
      RECT 378.105 218.305 378.435 218.470 ;
      RECT 102.000 216.430 102.380 217.980 ;
      RECT 104.720 216.430 105.100 217.980 ;
      RECT 105.400 216.430 105.780 217.980 ;
      RECT 108.800 216.430 109.180 217.980 ;
      RECT 110.185 217.790 110.515 217.955 ;
      RECT 102.025 216.265 102.355 216.430 ;
      RECT 104.745 216.265 105.075 216.430 ;
      RECT 105.425 216.265 105.755 216.430 ;
      RECT 108.825 216.265 109.155 216.430 ;
      RECT 110.160 216.240 110.540 217.790 ;
      RECT 369.920 216.430 370.300 217.980 ;
      RECT 371.280 216.430 371.660 217.980 ;
      RECT 373.320 216.430 373.700 217.980 ;
      RECT 378.105 217.790 378.435 217.955 ;
      RECT 369.945 216.265 370.275 216.430 ;
      RECT 371.305 216.265 371.635 216.430 ;
      RECT 373.345 216.265 373.675 216.430 ;
      RECT 378.080 216.240 378.460 217.790 ;
      RECT 102.680 214.390 103.060 215.940 ;
      RECT 106.105 215.750 106.435 215.915 ;
      RECT 108.825 215.750 109.155 215.915 ;
      RECT 102.705 214.225 103.035 214.390 ;
      RECT 106.080 214.200 106.460 215.750 ;
      RECT 108.800 214.200 109.180 215.750 ;
      RECT 110.840 214.390 111.220 215.940 ;
      RECT 369.945 215.750 370.275 215.915 ;
      RECT 371.305 215.750 371.635 215.915 ;
      RECT 373.345 215.750 373.675 215.915 ;
      RECT 110.865 214.225 111.195 214.390 ;
      RECT 104.040 212.350 104.420 213.900 ;
      RECT 106.785 213.710 107.115 213.875 ;
      RECT 104.065 212.185 104.395 212.350 ;
      RECT 106.760 212.160 107.140 213.710 ;
      RECT 108.120 212.350 108.500 213.900 ;
      RECT 110.185 213.710 110.515 213.875 ;
      RECT 108.145 212.185 108.475 212.350 ;
      RECT 110.160 212.160 110.540 213.710 ;
      RECT 127.160 212.350 127.540 214.580 ;
      RECT 369.920 214.200 370.300 215.750 ;
      RECT 371.280 214.200 371.660 215.750 ;
      RECT 373.320 214.200 373.700 215.750 ;
      RECT 375.360 214.390 375.740 215.940 ;
      RECT 377.425 215.750 377.755 215.915 ;
      RECT 375.385 214.225 375.715 214.390 ;
      RECT 377.400 214.200 377.780 215.750 ;
      RECT 127.185 212.185 127.515 212.350 ;
      RECT 108.800 210.310 109.180 211.860 ;
      RECT 110.865 211.670 111.195 211.835 ;
      RECT 345.440 211.670 345.820 213.220 ;
      RECT 366.520 212.350 366.900 213.900 ;
      RECT 369.240 212.350 369.620 213.900 ;
      RECT 371.305 213.710 371.635 213.875 ;
      RECT 374.705 213.710 375.035 213.875 ;
      RECT 366.545 212.185 366.875 212.350 ;
      RECT 369.265 212.185 369.595 212.350 ;
      RECT 371.280 212.160 371.660 213.710 ;
      RECT 374.680 212.160 375.060 213.710 ;
      RECT 369.265 211.670 369.595 211.835 ;
      RECT 108.825 210.145 109.155 210.310 ;
      RECT 110.840 210.120 111.220 211.670 ;
      RECT 345.465 211.505 345.795 211.670 ;
      RECT 369.240 210.120 369.620 211.670 ;
      RECT 371.280 210.310 371.660 211.860 ;
      RECT 374.190 211.835 375.740 211.860 ;
      RECT 374.025 211.505 375.740 211.835 ;
      RECT 374.190 211.480 375.740 211.505 ;
      RECT 371.305 210.145 371.635 210.310 ;
      RECT 105.425 209.630 105.755 209.795 ;
      RECT 108.825 209.630 109.155 209.795 ;
      RECT 102.680 206.910 103.060 208.460 ;
      RECT 105.400 208.080 105.780 209.630 ;
      RECT 108.800 208.080 109.180 209.630 ;
      RECT 110.160 208.270 110.540 209.820 ;
      RECT 369.240 208.270 369.620 209.820 ;
      RECT 371.280 208.270 371.660 209.820 ;
      RECT 374.680 208.270 375.060 209.820 ;
      RECT 110.185 208.105 110.515 208.270 ;
      RECT 369.265 208.105 369.595 208.270 ;
      RECT 371.305 208.105 371.635 208.270 ;
      RECT 374.705 208.105 375.035 208.270 ;
      RECT 102.705 206.745 103.035 206.910 ;
      RECT 102.705 206.230 103.035 206.395 ;
      RECT 102.680 204.680 103.060 206.230 ;
      RECT 107.440 204.870 107.820 206.420 ;
      RECT 135.320 205.550 135.700 207.100 ;
      RECT 345.465 206.910 345.795 207.075 ;
      RECT 378.080 206.910 378.460 208.460 ;
      RECT 135.345 205.385 135.675 205.550 ;
      RECT 345.440 205.360 345.820 206.910 ;
      RECT 378.105 206.745 378.435 206.910 ;
      RECT 376.065 206.230 376.395 206.395 ;
      RECT 378.105 206.230 378.435 206.395 ;
      RECT 107.465 204.705 107.795 204.870 ;
      RECT 102.000 202.830 102.380 204.380 ;
      RECT 108.825 204.190 109.155 204.355 ;
      RECT 110.865 204.190 111.195 204.355 ;
      RECT 102.025 202.665 102.355 202.830 ;
      RECT 108.800 202.640 109.180 204.190 ;
      RECT 110.840 202.640 111.220 204.190 ;
      RECT 136.000 203.510 136.380 205.060 ;
      RECT 344.785 204.870 345.115 205.035 ;
      RECT 136.025 203.345 136.355 203.510 ;
      RECT 344.760 203.320 345.140 204.870 ;
      RECT 376.040 204.680 376.420 206.230 ;
      RECT 378.080 204.680 378.460 206.230 ;
      RECT 369.240 202.830 369.620 204.380 ;
      RECT 371.280 202.830 371.660 204.380 ;
      RECT 378.080 202.830 378.460 204.380 ;
      RECT 369.265 202.665 369.595 202.830 ;
      RECT 371.305 202.665 371.635 202.830 ;
      RECT 378.105 202.665 378.435 202.830 ;
      RECT 102.680 200.790 103.060 202.340 ;
      RECT 106.080 200.790 106.460 202.340 ;
      RECT 108.120 200.790 108.500 202.340 ;
      RECT 110.840 200.790 111.220 202.340 ;
      RECT 345.465 200.790 345.795 200.955 ;
      RECT 369.240 200.790 369.620 202.340 ;
      RECT 371.305 202.150 371.635 202.315 ;
      RECT 376.065 202.150 376.395 202.315 ;
      RECT 378.105 202.150 378.435 202.315 ;
      RECT 102.705 200.625 103.035 200.790 ;
      RECT 106.105 200.625 106.435 200.790 ;
      RECT 108.145 200.625 108.475 200.790 ;
      RECT 110.865 200.625 111.195 200.790 ;
      RECT 102.680 198.750 103.060 200.300 ;
      RECT 104.745 200.110 105.075 200.275 ;
      RECT 108.825 200.110 109.155 200.275 ;
      RECT 110.185 200.110 110.515 200.275 ;
      RECT 102.705 198.585 103.035 198.750 ;
      RECT 104.720 198.560 105.100 200.110 ;
      RECT 108.800 198.560 109.180 200.110 ;
      RECT 110.160 198.560 110.540 200.110 ;
      RECT 345.440 199.240 345.820 200.790 ;
      RECT 369.265 200.625 369.595 200.790 ;
      RECT 371.280 200.600 371.660 202.150 ;
      RECT 376.040 200.600 376.420 202.150 ;
      RECT 378.080 200.600 378.460 202.150 ;
      RECT 369.945 200.110 370.275 200.275 ;
      RECT 371.305 200.110 371.635 200.275 ;
      RECT 373.345 200.110 373.675 200.275 ;
      RECT 376.065 200.110 376.395 200.275 ;
      RECT 377.425 200.110 377.755 200.275 ;
      RECT 369.920 198.560 370.300 200.110 ;
      RECT 371.280 198.560 371.660 200.110 ;
      RECT 373.320 198.560 373.700 200.110 ;
      RECT 376.040 198.560 376.420 200.110 ;
      RECT 377.400 198.560 377.780 200.110 ;
      RECT 102.705 198.070 103.035 198.235 ;
      RECT 102.680 196.520 103.060 198.070 ;
      RECT 104.040 196.710 104.420 198.260 ;
      RECT 108.825 198.070 109.155 198.235 ;
      RECT 110.865 198.070 111.195 198.235 ;
      RECT 369.945 198.070 370.275 198.235 ;
      RECT 104.065 196.545 104.395 196.710 ;
      RECT 108.800 196.520 109.180 198.070 ;
      RECT 110.840 196.520 111.220 198.070 ;
      RECT 369.920 196.520 370.300 198.070 ;
      RECT 371.280 196.710 371.660 198.260 ;
      RECT 373.345 198.070 373.675 198.235 ;
      RECT 371.305 196.545 371.635 196.710 ;
      RECT 373.320 196.520 373.700 198.070 ;
      RECT 374.680 196.710 375.060 198.260 ;
      RECT 376.040 196.710 376.420 198.260 ;
      RECT 378.080 196.710 378.460 198.260 ;
      RECT 374.705 196.545 375.035 196.710 ;
      RECT 376.065 196.545 376.395 196.710 ;
      RECT 378.105 196.545 378.435 196.710 ;
      RECT 102.000 194.670 102.380 196.220 ;
      RECT 104.065 196.030 104.395 196.195 ;
      RECT 102.025 194.505 102.355 194.670 ;
      RECT 104.040 194.480 104.420 196.030 ;
      RECT 105.400 194.670 105.780 196.220 ;
      RECT 108.145 196.030 108.475 196.195 ;
      RECT 105.425 194.505 105.755 194.670 ;
      RECT 108.120 194.480 108.500 196.030 ;
      RECT 110.160 194.670 110.540 196.220 ;
      RECT 369.920 194.670 370.300 196.220 ;
      RECT 371.280 194.670 371.660 196.220 ;
      RECT 375.360 194.670 375.740 196.220 ;
      RECT 378.105 196.030 378.435 196.195 ;
      RECT 110.185 194.505 110.515 194.670 ;
      RECT 369.945 194.505 370.275 194.670 ;
      RECT 371.305 194.505 371.635 194.670 ;
      RECT 375.385 194.505 375.715 194.670 ;
      RECT 378.080 194.480 378.460 196.030 ;
      RECT 107.440 192.630 107.820 194.180 ;
      RECT 108.800 192.630 109.180 194.180 ;
      RECT 110.840 192.630 111.220 194.180 ;
      RECT 369.920 192.630 370.300 194.180 ;
      RECT 371.960 192.630 372.340 194.180 ;
      RECT 373.345 193.990 373.675 194.155 ;
      RECT 107.465 192.465 107.795 192.630 ;
      RECT 108.825 192.465 109.155 192.630 ;
      RECT 110.865 192.465 111.195 192.630 ;
      RECT 369.945 192.465 370.275 192.630 ;
      RECT 371.985 192.465 372.315 192.630 ;
      RECT 373.320 192.440 373.700 193.990 ;
      RECT 375.360 192.630 375.740 194.180 ;
      RECT 375.385 192.465 375.715 192.630 ;
      RECT 108.120 190.590 108.500 192.140 ;
      RECT 110.840 190.590 111.220 192.140 ;
      RECT 369.240 190.590 369.620 192.140 ;
      RECT 371.305 191.950 371.635 192.115 ;
      RECT 108.145 190.425 108.475 190.590 ;
      RECT 110.865 190.425 111.195 190.590 ;
      RECT 369.265 190.425 369.595 190.590 ;
      RECT 371.280 190.400 371.660 191.950 ;
      RECT 102.680 187.190 103.060 188.740 ;
      RECT 105.400 188.550 105.780 190.100 ;
      RECT 108.145 189.910 108.475 190.075 ;
      RECT 110.865 189.910 111.195 190.075 ;
      RECT 105.425 188.385 105.755 188.550 ;
      RECT 108.120 188.360 108.500 189.910 ;
      RECT 110.840 188.360 111.220 189.910 ;
      RECT 134.665 189.230 134.995 189.395 ;
      RECT 134.640 187.680 135.020 189.230 ;
      RECT 369.920 188.550 370.300 190.100 ;
      RECT 371.985 189.910 372.315 190.075 ;
      RECT 369.945 188.385 370.275 188.550 ;
      RECT 371.960 188.360 372.340 189.910 ;
      RECT 373.320 188.550 373.700 190.100 ;
      RECT 373.345 188.385 373.675 188.550 ;
      RECT 135.345 187.190 135.675 187.355 ;
      RECT 344.785 187.190 345.115 187.355 ;
      RECT 377.400 187.190 377.780 188.740 ;
      RECT 102.705 187.025 103.035 187.190 ;
      RECT 102.025 186.510 102.355 186.675 ;
      RECT 104.065 186.510 104.395 186.675 ;
      RECT 102.000 184.960 102.380 186.510 ;
      RECT 104.040 184.960 104.420 186.510 ;
      RECT 135.320 185.640 135.700 187.190 ;
      RECT 344.760 185.640 345.140 187.190 ;
      RECT 377.425 187.025 377.755 187.190 ;
      RECT 102.705 184.470 103.035 184.635 ;
      RECT 102.680 182.920 103.060 184.470 ;
      RECT 344.760 183.790 345.140 185.340 ;
      RECT 373.320 185.150 373.700 186.700 ;
      RECT 374.680 185.150 375.060 186.700 ;
      RECT 378.105 186.510 378.435 186.675 ;
      RECT 373.345 184.985 373.675 185.150 ;
      RECT 374.705 184.985 375.035 185.150 ;
      RECT 378.080 184.960 378.460 186.510 ;
      RECT 378.105 184.470 378.435 184.635 ;
      RECT 344.785 183.625 345.115 183.790 ;
      RECT 378.080 182.920 378.460 184.470 ;
      RECT 102.000 181.070 102.380 182.620 ;
      RECT 106.785 182.430 107.115 182.595 ;
      RECT 102.025 180.905 102.355 181.070 ;
      RECT 106.760 180.880 107.140 182.430 ;
      RECT 108.120 181.070 108.500 182.620 ;
      RECT 110.185 182.430 110.515 182.595 ;
      RECT 108.145 180.905 108.475 181.070 ;
      RECT 110.160 180.880 110.540 182.430 ;
      RECT 102.025 180.390 102.355 180.555 ;
      RECT 104.065 180.390 104.395 180.555 ;
      RECT 106.105 180.390 106.435 180.555 ;
      RECT 108.145 180.390 108.475 180.555 ;
      RECT 102.000 178.840 102.380 180.390 ;
      RECT 104.040 178.840 104.420 180.390 ;
      RECT 106.080 178.840 106.460 180.390 ;
      RECT 108.120 178.840 108.500 180.390 ;
      RECT 110.840 179.030 111.220 180.580 ;
      RECT 345.440 179.710 345.820 181.260 ;
      RECT 369.240 181.070 369.620 182.620 ;
      RECT 371.280 181.070 371.660 182.620 ;
      RECT 374.680 181.070 375.060 182.620 ;
      RECT 375.385 182.430 375.715 182.595 ;
      RECT 369.265 180.905 369.595 181.070 ;
      RECT 371.305 180.905 371.635 181.070 ;
      RECT 374.705 180.905 375.035 181.070 ;
      RECT 375.360 180.880 375.740 182.430 ;
      RECT 378.080 181.070 378.460 182.620 ;
      RECT 378.105 180.905 378.435 181.070 ;
      RECT 345.465 179.545 345.795 179.710 ;
      RECT 369.240 179.030 369.620 180.580 ;
      RECT 371.960 179.030 372.340 180.580 ;
      RECT 375.360 179.030 375.740 180.580 ;
      RECT 378.105 180.390 378.435 180.555 ;
      RECT 110.865 178.865 111.195 179.030 ;
      RECT 369.265 178.865 369.595 179.030 ;
      RECT 371.985 178.865 372.315 179.030 ;
      RECT 375.385 178.865 375.715 179.030 ;
      RECT 378.080 178.840 378.460 180.390 ;
      RECT 102.680 176.990 103.060 178.540 ;
      RECT 104.745 178.350 105.075 178.515 ;
      RECT 102.705 176.825 103.035 176.990 ;
      RECT 104.720 176.800 105.100 178.350 ;
      RECT 108.800 176.990 109.180 178.540 ;
      RECT 110.185 178.350 110.515 178.515 ;
      RECT 108.825 176.825 109.155 176.990 ;
      RECT 110.160 176.800 110.540 178.350 ;
      RECT 369.920 176.990 370.300 178.540 ;
      RECT 371.305 178.350 371.635 178.515 ;
      RECT 373.345 178.350 373.675 178.515 ;
      RECT 369.945 176.825 370.275 176.990 ;
      RECT 371.280 176.800 371.660 178.350 ;
      RECT 373.320 176.800 373.700 178.350 ;
      RECT 375.360 176.990 375.740 178.540 ;
      RECT 377.425 178.350 377.755 178.515 ;
      RECT 375.385 176.825 375.715 176.990 ;
      RECT 377.400 176.800 377.780 178.350 ;
      RECT 102.000 174.950 102.380 176.500 ;
      RECT 104.040 174.950 104.420 176.500 ;
      RECT 108.825 176.310 109.155 176.475 ;
      RECT 102.025 174.785 102.355 174.950 ;
      RECT 104.065 174.785 104.395 174.950 ;
      RECT 108.800 174.760 109.180 176.310 ;
      RECT 110.160 174.950 110.540 176.500 ;
      RECT 369.945 176.310 370.275 176.475 ;
      RECT 110.185 174.785 110.515 174.950 ;
      RECT 369.920 174.760 370.300 176.310 ;
      RECT 371.280 174.950 371.660 176.500 ;
      RECT 374.000 174.950 374.380 176.500 ;
      RECT 374.680 174.950 375.060 176.500 ;
      RECT 378.080 174.950 378.460 176.500 ;
      RECT 371.305 174.785 371.635 174.950 ;
      RECT 374.025 174.785 374.355 174.950 ;
      RECT 374.705 174.785 375.035 174.950 ;
      RECT 378.105 174.785 378.435 174.950 ;
      RECT 68.025 167.470 68.355 167.635 ;
      RECT 68.000 153.680 68.380 167.470 ;
      RECT 68.680 160.670 69.060 174.460 ;
      RECT 104.720 172.910 105.100 174.460 ;
      RECT 105.400 172.910 105.780 174.460 ;
      RECT 108.800 172.910 109.180 174.460 ;
      RECT 110.160 172.910 110.540 174.460 ;
      RECT 369.920 172.910 370.300 174.460 ;
      RECT 371.280 172.910 371.660 174.460 ;
      RECT 375.360 172.910 375.740 174.460 ;
      RECT 104.745 172.745 105.075 172.910 ;
      RECT 105.425 172.745 105.755 172.910 ;
      RECT 108.825 172.745 109.155 172.910 ;
      RECT 110.185 172.745 110.515 172.910 ;
      RECT 369.945 172.745 370.275 172.910 ;
      RECT 371.305 172.745 371.635 172.910 ;
      RECT 375.385 172.745 375.715 172.910 ;
      RECT 102.680 170.870 103.060 172.420 ;
      RECT 107.440 170.870 107.820 172.420 ;
      RECT 108.800 170.870 109.180 172.420 ;
      RECT 110.185 172.230 110.515 172.395 ;
      RECT 102.705 170.705 103.035 170.870 ;
      RECT 107.465 170.705 107.795 170.870 ;
      RECT 108.825 170.705 109.155 170.870 ;
      RECT 110.160 170.680 110.540 172.230 ;
      RECT 369.920 170.870 370.300 172.420 ;
      RECT 371.960 170.870 372.340 172.420 ;
      RECT 373.345 172.230 373.675 172.395 ;
      RECT 369.945 170.705 370.275 170.870 ;
      RECT 371.985 170.705 372.315 170.870 ;
      RECT 373.320 170.680 373.700 172.230 ;
      RECT 376.040 170.870 376.420 172.420 ;
      RECT 377.425 172.230 377.755 172.395 ;
      RECT 376.065 170.705 376.395 170.870 ;
      RECT 377.400 170.680 377.780 172.230 ;
      RECT 106.785 170.190 107.115 170.355 ;
      RECT 108.145 170.190 108.475 170.355 ;
      RECT 102.000 167.470 102.380 169.020 ;
      RECT 106.760 168.640 107.140 170.190 ;
      RECT 108.120 168.640 108.500 170.190 ;
      RECT 110.840 168.830 111.220 170.380 ;
      RECT 369.240 168.830 369.620 170.380 ;
      RECT 371.305 170.190 371.635 170.355 ;
      RECT 110.865 168.665 111.195 168.830 ;
      RECT 369.265 168.665 369.595 168.830 ;
      RECT 371.280 168.640 371.660 170.190 ;
      RECT 374.000 168.830 374.380 170.380 ;
      RECT 374.680 168.830 375.060 170.380 ;
      RECT 374.025 168.665 374.355 168.830 ;
      RECT 374.705 168.665 375.035 168.830 ;
      RECT 102.025 167.305 102.355 167.470 ;
      RECT 108.800 166.790 109.180 168.340 ;
      RECT 110.865 168.150 111.195 168.315 ;
      RECT 369.265 168.150 369.595 168.315 ;
      RECT 108.825 166.625 109.155 166.790 ;
      RECT 110.840 166.600 111.220 168.150 ;
      RECT 369.240 166.600 369.620 168.150 ;
      RECT 371.280 166.790 371.660 168.340 ;
      RECT 377.400 167.470 377.780 169.020 ;
      RECT 377.425 167.305 377.755 167.470 ;
      RECT 371.305 166.625 371.635 166.790 ;
      RECT 102.680 163.390 103.060 164.940 ;
      RECT 136.000 164.070 136.380 165.620 ;
      RECT 344.785 165.430 345.115 165.595 ;
      RECT 136.025 163.905 136.355 164.070 ;
      RECT 344.760 163.880 345.140 165.430 ;
      RECT 374.000 164.750 374.380 166.300 ;
      RECT 374.680 164.750 375.060 166.300 ;
      RECT 374.025 164.585 374.355 164.750 ;
      RECT 374.705 164.585 375.035 164.750 ;
      RECT 378.080 163.390 378.460 164.940 ;
      RECT 102.705 163.225 103.035 163.390 ;
      RECT 378.105 163.225 378.435 163.390 ;
      RECT 102.705 162.710 103.035 162.875 ;
      RECT 104.065 162.710 104.395 162.875 ;
      RECT 108.145 162.710 108.475 162.875 ;
      RECT 110.865 162.710 111.195 162.875 ;
      RECT 102.680 161.160 103.060 162.710 ;
      RECT 104.040 161.160 104.420 162.710 ;
      RECT 108.120 161.160 108.500 162.710 ;
      RECT 110.840 161.160 111.220 162.710 ;
      RECT 102.025 160.670 102.355 160.835 ;
      RECT 104.745 160.670 105.075 160.835 ;
      RECT 68.705 160.505 69.035 160.670 ;
      RECT 68.705 159.990 69.035 160.155 ;
      RECT 67.345 153.190 67.675 153.355 ;
      RECT 67.320 139.400 67.700 153.190 ;
      RECT 68.680 146.880 69.060 159.990 ;
      RECT 102.000 159.120 102.380 160.670 ;
      RECT 104.720 159.120 105.100 160.670 ;
      RECT 107.440 159.310 107.820 160.860 ;
      RECT 108.120 159.310 108.500 160.860 ;
      RECT 110.160 159.310 110.540 160.860 ;
      RECT 136.000 159.990 136.380 161.540 ;
      RECT 369.920 161.350 370.300 162.900 ;
      RECT 371.985 162.710 372.315 162.875 ;
      RECT 369.945 161.185 370.275 161.350 ;
      RECT 371.960 161.160 372.340 162.710 ;
      RECT 373.320 161.350 373.700 162.900 ;
      RECT 377.400 161.350 377.780 162.900 ;
      RECT 373.345 161.185 373.675 161.350 ;
      RECT 377.425 161.185 377.755 161.350 ;
      RECT 369.945 160.670 370.275 160.835 ;
      RECT 136.025 159.825 136.355 159.990 ;
      RECT 107.465 159.145 107.795 159.310 ;
      RECT 108.145 159.145 108.475 159.310 ;
      RECT 110.185 159.145 110.515 159.310 ;
      RECT 369.920 159.120 370.300 160.670 ;
      RECT 371.280 159.310 371.660 160.860 ;
      RECT 374.000 159.310 374.380 160.860 ;
      RECT 377.425 160.670 377.755 160.835 ;
      RECT 371.305 159.145 371.635 159.310 ;
      RECT 374.025 159.145 374.355 159.310 ;
      RECT 377.400 159.120 377.780 160.670 ;
      RECT 102.680 157.270 103.060 158.820 ;
      RECT 106.105 158.630 106.435 158.795 ;
      RECT 102.705 157.105 103.035 157.270 ;
      RECT 106.080 157.080 106.460 158.630 ;
      RECT 108.120 157.270 108.500 158.820 ;
      RECT 110.840 157.270 111.220 158.820 ;
      RECT 369.240 157.270 369.620 158.820 ;
      RECT 371.960 157.270 372.340 158.820 ;
      RECT 374.025 158.630 374.355 158.795 ;
      RECT 376.065 158.630 376.395 158.795 ;
      RECT 108.145 157.105 108.475 157.270 ;
      RECT 110.865 157.105 111.195 157.270 ;
      RECT 369.265 157.105 369.595 157.270 ;
      RECT 371.985 157.105 372.315 157.270 ;
      RECT 374.000 157.080 374.380 158.630 ;
      RECT 376.040 157.080 376.420 158.630 ;
      RECT 378.080 157.270 378.460 158.820 ;
      RECT 378.105 157.105 378.435 157.270 ;
      RECT 102.025 156.590 102.355 156.755 ;
      RECT 104.745 156.590 105.075 156.755 ;
      RECT 105.425 156.590 105.755 156.755 ;
      RECT 108.825 156.590 109.155 156.755 ;
      RECT 110.185 156.590 110.515 156.755 ;
      RECT 102.000 155.040 102.380 156.590 ;
      RECT 104.720 155.040 105.100 156.590 ;
      RECT 105.400 155.040 105.780 156.590 ;
      RECT 108.800 155.040 109.180 156.590 ;
      RECT 110.160 155.040 110.540 156.590 ;
      RECT 369.920 155.230 370.300 156.780 ;
      RECT 371.960 155.230 372.340 156.780 ;
      RECT 375.360 155.230 375.740 156.780 ;
      RECT 377.425 156.590 377.755 156.755 ;
      RECT 369.945 155.065 370.275 155.230 ;
      RECT 371.985 155.065 372.315 155.230 ;
      RECT 375.385 155.065 375.715 155.230 ;
      RECT 377.400 155.040 377.780 156.590 ;
      RECT 102.000 153.190 102.380 154.740 ;
      RECT 104.040 153.190 104.420 154.740 ;
      RECT 107.465 154.550 107.795 154.715 ;
      RECT 108.825 154.550 109.155 154.715 ;
      RECT 102.025 153.025 102.355 153.190 ;
      RECT 104.065 153.025 104.395 153.190 ;
      RECT 107.440 153.000 107.820 154.550 ;
      RECT 108.800 153.000 109.180 154.550 ;
      RECT 110.840 153.190 111.220 154.740 ;
      RECT 369.240 153.190 369.620 154.740 ;
      RECT 371.985 154.550 372.315 154.715 ;
      RECT 373.345 154.550 373.675 154.715 ;
      RECT 110.865 153.025 111.195 153.190 ;
      RECT 369.265 153.025 369.595 153.190 ;
      RECT 371.960 153.000 372.340 154.550 ;
      RECT 373.320 153.000 373.700 154.550 ;
      RECT 378.080 153.190 378.460 154.740 ;
      RECT 378.105 153.025 378.435 153.190 ;
      RECT 102.000 151.150 102.380 152.700 ;
      RECT 108.800 151.150 109.180 152.700 ;
      RECT 110.185 152.510 110.515 152.675 ;
      RECT 369.265 152.510 369.595 152.675 ;
      RECT 102.025 150.985 102.355 151.150 ;
      RECT 108.825 150.985 109.155 151.150 ;
      RECT 110.160 150.960 110.540 152.510 ;
      RECT 369.240 150.960 369.620 152.510 ;
      RECT 371.280 151.150 371.660 152.700 ;
      RECT 374.025 152.510 374.355 152.675 ;
      RECT 371.305 150.985 371.635 151.150 ;
      RECT 374.000 150.960 374.380 152.510 ;
      RECT 377.400 151.150 377.780 152.700 ;
      RECT 377.425 150.985 377.755 151.150 ;
      RECT 106.105 150.470 106.435 150.635 ;
      RECT 108.825 150.470 109.155 150.635 ;
      RECT 110.185 150.470 110.515 150.635 ;
      RECT 369.945 150.470 370.275 150.635 ;
      RECT 371.305 150.470 371.635 150.635 ;
      RECT 102.680 147.750 103.060 149.300 ;
      RECT 106.080 148.920 106.460 150.470 ;
      RECT 108.800 148.920 109.180 150.470 ;
      RECT 110.160 148.920 110.540 150.470 ;
      RECT 369.920 148.920 370.300 150.470 ;
      RECT 371.280 148.920 371.660 150.470 ;
      RECT 373.320 149.110 373.700 150.660 ;
      RECT 374.680 149.110 375.060 150.660 ;
      RECT 373.345 148.945 373.675 149.110 ;
      RECT 374.705 148.945 375.035 149.110 ;
      RECT 108.145 148.430 108.475 148.595 ;
      RECT 102.705 147.585 103.035 147.750 ;
      RECT 108.120 146.880 108.500 148.430 ;
      RECT 110.840 147.070 111.220 148.620 ;
      RECT 369.240 147.070 369.620 148.620 ;
      RECT 371.960 147.070 372.340 148.620 ;
      RECT 378.080 147.750 378.460 149.300 ;
      RECT 378.105 147.585 378.435 147.750 ;
      RECT 110.865 146.905 111.195 147.070 ;
      RECT 369.265 146.905 369.595 147.070 ;
      RECT 371.985 146.905 372.315 147.070 ;
      RECT 68.000 132.790 68.380 146.580 ;
      RECT 102.025 145.030 102.355 145.195 ;
      RECT 105.400 145.030 105.780 146.580 ;
      RECT 102.000 143.480 102.380 145.030 ;
      RECT 105.425 144.865 105.755 145.030 ;
      RECT 104.745 144.350 105.075 144.515 ;
      RECT 136.000 144.350 136.380 145.900 ;
      RECT 344.785 145.710 345.115 145.875 ;
      RECT 104.720 143.860 105.100 144.350 ;
      RECT 136.025 144.185 136.355 144.350 ;
      RECT 344.760 144.160 345.140 145.710 ;
      RECT 373.320 145.030 373.700 146.580 ;
      RECT 377.425 145.030 377.755 145.195 ;
      RECT 373.345 144.865 373.675 145.030 ;
      RECT 104.720 143.480 105.780 143.860 ;
      RECT 135.345 143.670 135.675 143.835 ;
      RECT 102.680 141.630 103.060 143.180 ;
      RECT 104.065 142.990 104.395 143.155 ;
      RECT 102.705 141.465 103.035 141.630 ;
      RECT 104.040 141.440 104.420 142.990 ;
      RECT 135.320 142.120 135.700 143.670 ;
      RECT 344.760 142.310 345.140 143.860 ;
      RECT 344.785 142.145 345.115 142.310 ;
      RECT 345.440 141.630 345.820 143.860 ;
      RECT 377.400 143.480 377.780 145.030 ;
      RECT 374.705 142.990 375.035 143.155 ;
      RECT 378.105 142.990 378.435 143.155 ;
      RECT 345.465 141.465 345.795 141.630 ;
      RECT 374.680 141.440 375.060 142.990 ;
      RECT 378.080 141.440 378.460 142.990 ;
      RECT 102.705 140.950 103.035 141.115 ;
      RECT 102.680 139.400 103.060 140.950 ;
      RECT 108.800 139.590 109.180 141.140 ;
      RECT 110.160 139.590 110.540 141.140 ;
      RECT 369.920 139.590 370.300 141.140 ;
      RECT 371.280 139.590 371.660 141.140 ;
      RECT 378.105 140.950 378.435 141.115 ;
      RECT 108.825 139.425 109.155 139.590 ;
      RECT 110.185 139.425 110.515 139.590 ;
      RECT 369.945 139.425 370.275 139.590 ;
      RECT 371.305 139.425 371.635 139.590 ;
      RECT 378.080 139.400 378.460 140.950 ;
      RECT 68.025 132.625 68.355 132.790 ;
      RECT 68.680 125.310 69.060 139.100 ;
      RECT 102.000 137.550 102.380 139.100 ;
      RECT 107.440 137.550 107.820 139.100 ;
      RECT 108.120 137.550 108.500 139.100 ;
      RECT 110.185 138.910 110.515 139.075 ;
      RECT 369.945 138.910 370.275 139.075 ;
      RECT 102.025 137.385 102.355 137.550 ;
      RECT 107.465 137.385 107.795 137.550 ;
      RECT 108.145 137.385 108.475 137.550 ;
      RECT 110.160 137.360 110.540 138.910 ;
      RECT 135.345 137.550 135.675 137.715 ;
      RECT 102.680 135.510 103.060 137.060 ;
      RECT 104.065 136.870 104.395 137.035 ;
      RECT 102.705 135.345 103.035 135.510 ;
      RECT 104.040 135.320 104.420 136.870 ;
      RECT 105.400 135.510 105.780 137.060 ;
      RECT 108.145 136.870 108.475 137.035 ;
      RECT 110.185 136.870 110.515 137.035 ;
      RECT 105.425 135.345 105.755 135.510 ;
      RECT 108.120 135.320 108.500 136.870 ;
      RECT 110.160 135.320 110.540 136.870 ;
      RECT 135.320 136.000 135.700 137.550 ;
      RECT 345.440 136.190 345.820 137.740 ;
      RECT 369.920 137.360 370.300 138.910 ;
      RECT 371.280 137.550 371.660 139.100 ;
      RECT 373.345 138.910 373.675 139.075 ;
      RECT 377.425 138.910 377.755 139.075 ;
      RECT 371.305 137.385 371.635 137.550 ;
      RECT 373.320 137.360 373.700 138.910 ;
      RECT 377.400 137.360 377.780 138.910 ;
      RECT 369.265 136.870 369.595 137.035 ;
      RECT 371.305 136.870 371.635 137.035 ;
      RECT 376.065 136.870 376.395 137.035 ;
      RECT 345.465 136.025 345.795 136.190 ;
      RECT 369.240 135.320 369.620 136.870 ;
      RECT 371.280 135.320 371.660 136.870 ;
      RECT 376.040 135.320 376.420 136.870 ;
      RECT 378.080 135.510 378.460 137.060 ;
      RECT 378.105 135.345 378.435 135.510 ;
      RECT 102.025 134.830 102.355 134.995 ;
      RECT 102.000 133.280 102.380 134.830 ;
      RECT 104.720 133.470 105.100 135.020 ;
      RECT 105.425 134.830 105.755 134.995 ;
      RECT 104.745 133.305 105.075 133.470 ;
      RECT 105.400 133.280 105.780 134.830 ;
      RECT 108.800 133.470 109.180 135.020 ;
      RECT 110.185 134.830 110.515 134.995 ;
      RECT 369.945 134.830 370.275 134.995 ;
      RECT 371.305 134.830 371.635 134.995 ;
      RECT 373.345 134.830 373.675 134.995 ;
      RECT 108.825 133.305 109.155 133.470 ;
      RECT 110.160 133.280 110.540 134.830 ;
      RECT 369.920 133.280 370.300 134.830 ;
      RECT 371.280 133.280 371.660 134.830 ;
      RECT 373.320 133.280 373.700 134.830 ;
      RECT 375.360 133.470 375.740 135.020 ;
      RECT 377.425 134.830 377.755 134.995 ;
      RECT 375.385 133.305 375.715 133.470 ;
      RECT 377.400 133.280 377.780 134.830 ;
      RECT 102.705 132.790 103.035 132.955 ;
      RECT 87.065 132.110 87.395 132.275 ;
      RECT 68.705 125.145 69.035 125.310 ;
      RECT 77.545 124.630 77.875 124.795 ;
      RECT 12.800 113.020 13.130 113.350 ;
      RECT 11.560 77.710 11.940 81.300 ;
      RECT 11.585 77.545 11.915 77.710 ;
      RECT 12.815 76.315 13.115 113.020 ;
      RECT 77.520 111.520 77.900 124.630 ;
      RECT 87.040 123.760 87.420 132.110 ;
      RECT 102.680 131.240 103.060 132.790 ;
      RECT 104.040 131.430 104.420 132.980 ;
      RECT 107.465 132.790 107.795 132.955 ;
      RECT 108.825 132.790 109.155 132.955 ;
      RECT 104.065 131.265 104.395 131.430 ;
      RECT 107.440 131.240 107.820 132.790 ;
      RECT 108.800 131.240 109.180 132.790 ;
      RECT 110.160 131.430 110.540 132.980 ;
      RECT 369.240 131.430 369.620 132.980 ;
      RECT 371.280 131.430 371.660 132.980 ;
      RECT 373.345 132.790 373.675 132.955 ;
      RECT 110.185 131.265 110.515 131.430 ;
      RECT 369.265 131.265 369.595 131.430 ;
      RECT 371.305 131.265 371.635 131.430 ;
      RECT 373.320 131.240 373.700 132.790 ;
      RECT 374.680 131.430 375.060 132.980 ;
      RECT 378.080 131.430 378.460 132.980 ;
      RECT 374.705 131.265 375.035 131.430 ;
      RECT 378.105 131.265 378.435 131.430 ;
      RECT 108.800 129.390 109.180 130.940 ;
      RECT 110.865 130.750 111.195 130.915 ;
      RECT 369.265 130.750 369.595 130.915 ;
      RECT 108.825 129.225 109.155 129.390 ;
      RECT 110.840 129.200 111.220 130.750 ;
      RECT 108.825 128.710 109.155 128.875 ;
      RECT 108.800 127.160 109.180 128.710 ;
      RECT 110.840 127.350 111.220 128.900 ;
      RECT 136.000 128.710 136.380 130.260 ;
      RECT 369.240 129.200 369.620 130.750 ;
      RECT 371.280 129.390 371.660 130.940 ;
      RECT 375.360 129.390 375.740 130.940 ;
      RECT 371.305 129.225 371.635 129.390 ;
      RECT 375.385 129.225 375.715 129.390 ;
      RECT 369.945 128.710 370.275 128.875 ;
      RECT 371.305 128.710 371.635 128.875 ;
      RECT 136.025 128.545 136.355 128.710 ;
      RECT 110.865 127.185 111.195 127.350 ;
      RECT 369.920 127.160 370.300 128.710 ;
      RECT 371.280 127.160 371.660 128.710 ;
      RECT 102.000 123.950 102.380 125.500 ;
      RECT 102.025 123.785 102.355 123.950 ;
      RECT 85.680 119.870 86.060 123.460 ;
      RECT 86.360 119.870 86.740 121.420 ;
      RECT 89.760 119.870 90.140 123.460 ;
      RECT 91.825 122.590 92.155 122.755 ;
      RECT 93.185 122.590 93.515 122.755 ;
      RECT 91.145 121.230 91.475 121.395 ;
      RECT 85.705 119.705 86.035 119.870 ;
      RECT 86.385 119.705 86.715 119.870 ;
      RECT 89.785 119.705 90.115 119.870 ;
      RECT 91.120 119.680 91.500 121.230 ;
      RECT 91.800 119.680 92.180 122.590 ;
      RECT 93.160 119.680 93.540 122.590 ;
      RECT 102.680 121.910 103.060 123.460 ;
      RECT 104.040 122.590 104.420 126.860 ;
      RECT 106.785 126.670 107.115 126.835 ;
      RECT 108.145 126.670 108.475 126.835 ;
      RECT 110.185 126.670 110.515 126.835 ;
      RECT 369.265 126.670 369.595 126.835 ;
      RECT 106.760 125.120 107.140 126.670 ;
      RECT 108.120 125.120 108.500 126.670 ;
      RECT 110.160 125.120 110.540 126.670 ;
      RECT 369.240 125.120 369.620 126.670 ;
      RECT 371.960 125.310 372.340 126.860 ;
      RECT 374.000 125.310 374.380 126.860 ;
      RECT 374.680 125.310 375.060 126.860 ;
      RECT 378.105 125.310 378.435 125.475 ;
      RECT 371.985 125.145 372.315 125.310 ;
      RECT 374.025 125.145 374.355 125.310 ;
      RECT 374.705 125.145 375.035 125.310 ;
      RECT 134.665 123.950 134.995 124.115 ;
      RECT 344.785 123.950 345.115 124.115 ;
      RECT 107.465 123.270 107.795 123.435 ;
      RECT 104.065 122.425 104.395 122.590 ;
      RECT 102.705 121.745 103.035 121.910 ;
      RECT 107.440 121.720 107.820 123.270 ;
      RECT 134.640 122.400 135.020 123.950 ;
      RECT 344.760 122.400 345.140 123.950 ;
      RECT 378.080 123.760 378.460 125.310 ;
      RECT 373.345 123.270 373.675 123.435 ;
      RECT 344.785 121.910 345.115 122.075 ;
      RECT 102.025 121.230 102.355 121.395 ;
      RECT 108.145 121.230 108.475 121.395 ;
      RECT 102.000 119.680 102.380 121.230 ;
      RECT 108.120 119.680 108.500 121.230 ;
      RECT 110.840 119.870 111.220 121.420 ;
      RECT 344.760 120.360 345.140 121.910 ;
      RECT 373.320 121.720 373.700 123.270 ;
      RECT 377.400 121.910 377.780 123.460 ;
      RECT 390.345 123.270 390.675 123.435 ;
      RECT 386.265 122.590 386.595 122.755 ;
      RECT 377.425 121.745 377.755 121.910 ;
      RECT 369.265 121.230 369.595 121.395 ;
      RECT 110.865 119.705 111.195 119.870 ;
      RECT 85.705 119.190 86.035 119.355 ;
      RECT 91.825 119.190 92.155 119.355 ;
      RECT 102.705 119.190 103.035 119.355 ;
      RECT 104.065 119.190 104.395 119.355 ;
      RECT 85.680 115.600 86.060 119.190 ;
      RECT 89.105 118.510 89.435 118.675 ;
      RECT 89.080 115.600 89.460 118.510 ;
      RECT 91.800 115.600 92.180 119.190 ;
      RECT 102.680 117.640 103.060 119.190 ;
      RECT 104.040 117.640 104.420 119.190 ;
      RECT 108.800 117.830 109.180 119.380 ;
      RECT 110.160 117.830 110.540 119.380 ;
      RECT 135.320 117.830 135.700 120.060 ;
      RECT 369.240 119.680 369.620 121.230 ;
      RECT 371.960 119.870 372.340 121.420 ;
      RECT 371.985 119.705 372.315 119.870 ;
      RECT 344.785 117.830 345.115 117.995 ;
      RECT 369.920 117.830 370.300 119.380 ;
      RECT 371.985 119.190 372.315 119.355 ;
      RECT 374.680 119.190 375.060 120.740 ;
      RECT 378.080 119.870 378.460 121.420 ;
      RECT 378.105 119.705 378.435 119.870 ;
      RECT 386.240 119.680 386.620 122.590 ;
      RECT 388.960 119.870 389.340 122.780 ;
      RECT 388.985 119.705 389.315 119.870 ;
      RECT 390.320 119.680 390.700 123.270 ;
      RECT 395.080 119.870 395.460 123.460 ;
      RECT 395.105 119.705 395.435 119.870 ;
      RECT 376.065 119.190 376.395 119.355 ;
      RECT 108.825 117.665 109.155 117.830 ;
      RECT 110.185 117.665 110.515 117.830 ;
      RECT 135.345 117.665 135.675 117.830 ;
      RECT 102.025 117.150 102.355 117.315 ;
      RECT 104.745 117.150 105.075 117.315 ;
      RECT 102.000 115.600 102.380 117.150 ;
      RECT 104.720 115.600 105.100 117.150 ;
      RECT 107.440 115.790 107.820 117.340 ;
      RECT 108.825 117.150 109.155 117.315 ;
      RECT 107.465 115.625 107.795 115.790 ;
      RECT 108.800 115.600 109.180 117.150 ;
      RECT 110.160 115.790 110.540 117.340 ;
      RECT 344.760 116.280 345.140 117.830 ;
      RECT 369.945 117.665 370.275 117.830 ;
      RECT 371.960 117.640 372.340 119.190 ;
      RECT 374.705 119.025 375.035 119.190 ;
      RECT 376.040 117.640 376.420 119.190 ;
      RECT 377.400 117.830 377.780 119.380 ;
      RECT 377.425 117.665 377.755 117.830 ;
      RECT 369.945 117.150 370.275 117.315 ;
      RECT 371.305 117.150 371.635 117.315 ;
      RECT 110.185 115.625 110.515 115.790 ;
      RECT 369.920 115.600 370.300 117.150 ;
      RECT 371.280 115.600 371.660 117.150 ;
      RECT 374.000 115.790 374.380 117.340 ;
      RECT 377.425 117.150 377.755 117.315 ;
      RECT 374.025 115.625 374.355 115.790 ;
      RECT 377.400 115.600 377.780 117.150 ;
      RECT 388.280 116.470 388.660 119.380 ;
      RECT 388.985 119.190 389.315 119.355 ;
      RECT 391.705 119.190 392.035 119.355 ;
      RECT 388.305 116.305 388.635 116.470 ;
      RECT 388.960 115.600 389.340 119.190 ;
      RECT 391.680 115.600 392.060 119.190 ;
      RECT 395.080 115.790 395.460 119.380 ;
      RECT 395.105 115.625 395.435 115.790 ;
      RECT 85.000 111.710 85.380 115.300 ;
      RECT 88.400 111.710 88.780 115.300 ;
      RECT 91.800 111.710 92.180 115.300 ;
      RECT 93.840 111.710 94.220 115.300 ;
      RECT 102.680 113.750 103.060 115.300 ;
      RECT 104.040 113.750 104.420 115.300 ;
      RECT 108.120 113.750 108.500 115.300 ;
      RECT 110.185 115.110 110.515 115.275 ;
      RECT 102.705 113.585 103.035 113.750 ;
      RECT 104.065 113.585 104.395 113.750 ;
      RECT 108.145 113.585 108.475 113.750 ;
      RECT 110.160 113.560 110.540 115.110 ;
      RECT 369.240 113.750 369.620 115.300 ;
      RECT 371.960 113.750 372.340 115.300 ;
      RECT 376.065 115.110 376.395 115.275 ;
      RECT 378.105 115.110 378.435 115.275 ;
      RECT 369.265 113.585 369.595 113.750 ;
      RECT 371.985 113.585 372.315 113.750 ;
      RECT 376.040 113.560 376.420 115.110 ;
      RECT 378.080 113.560 378.460 115.110 ;
      RECT 102.025 113.070 102.355 113.235 ;
      RECT 85.025 111.545 85.355 111.710 ;
      RECT 88.425 111.545 88.755 111.710 ;
      RECT 91.825 111.545 92.155 111.710 ;
      RECT 93.865 111.545 94.195 111.710 ;
      RECT 102.000 111.520 102.380 113.070 ;
      RECT 108.800 111.710 109.180 113.260 ;
      RECT 110.185 113.070 110.515 113.235 ;
      RECT 108.825 111.545 109.155 111.710 ;
      RECT 110.160 111.520 110.540 113.070 ;
      RECT 369.920 111.710 370.300 113.260 ;
      RECT 371.305 113.070 371.635 113.235 ;
      RECT 373.345 113.070 373.675 113.235 ;
      RECT 369.945 111.545 370.275 111.710 ;
      RECT 371.280 111.520 371.660 113.070 ;
      RECT 373.320 111.520 373.700 113.070 ;
      RECT 375.360 111.710 375.740 113.260 ;
      RECT 377.400 111.710 377.780 113.260 ;
      RECT 386.240 111.710 386.620 115.300 ;
      RECT 388.985 115.110 389.315 115.275 ;
      RECT 375.385 111.545 375.715 111.710 ;
      RECT 377.425 111.545 377.755 111.710 ;
      RECT 386.265 111.545 386.595 111.710 ;
      RECT 388.960 111.520 389.340 115.110 ;
      RECT 393.040 111.710 393.420 115.300 ;
      RECT 394.425 115.110 394.755 115.275 ;
      RECT 393.065 111.545 393.395 111.710 ;
      RECT 394.400 111.520 394.780 115.110 ;
      RECT 86.385 111.030 86.715 111.195 ;
      RECT 92.505 111.030 92.835 111.195 ;
      RECT 86.360 104.040 86.740 111.030 ;
      RECT 92.480 108.120 92.860 111.030 ;
      RECT 93.160 104.230 93.540 111.220 ;
      RECT 104.040 109.670 104.420 111.220 ;
      RECT 107.465 111.030 107.795 111.195 ;
      RECT 108.825 111.030 109.155 111.195 ;
      RECT 110.865 111.030 111.195 111.195 ;
      RECT 104.065 109.505 104.395 109.670 ;
      RECT 107.440 109.480 107.820 111.030 ;
      RECT 108.800 109.480 109.180 111.030 ;
      RECT 110.840 109.480 111.220 111.030 ;
      RECT 108.800 107.630 109.180 109.180 ;
      RECT 110.160 107.630 110.540 109.180 ;
      RECT 134.640 108.990 135.020 110.540 ;
      RECT 369.240 109.670 369.620 111.220 ;
      RECT 371.280 109.670 371.660 111.220 ;
      RECT 374.000 109.670 374.380 111.220 ;
      RECT 374.680 109.670 375.060 111.220 ;
      RECT 376.040 109.670 376.420 111.220 ;
      RECT 369.265 109.505 369.595 109.670 ;
      RECT 371.305 109.505 371.635 109.670 ;
      RECT 374.025 109.505 374.355 109.670 ;
      RECT 374.705 109.505 375.035 109.670 ;
      RECT 376.065 109.505 376.395 109.670 ;
      RECT 345.465 108.990 345.795 109.155 ;
      RECT 369.265 108.990 369.595 109.155 ;
      RECT 371.985 108.990 372.315 109.155 ;
      RECT 134.665 108.825 134.995 108.990 ;
      RECT 108.825 107.465 109.155 107.630 ;
      RECT 110.185 107.465 110.515 107.630 ;
      RECT 105.425 106.950 105.755 107.115 ;
      RECT 102.705 105.590 103.035 105.755 ;
      RECT 93.185 104.065 93.515 104.230 ;
      RECT 102.680 104.040 103.060 105.590 ;
      RECT 105.400 105.400 105.780 106.950 ;
      RECT 108.800 105.590 109.180 107.140 ;
      RECT 110.185 106.950 110.515 107.115 ;
      RECT 108.825 105.425 109.155 105.590 ;
      RECT 110.160 105.400 110.540 106.950 ;
      RECT 344.760 105.590 345.140 107.820 ;
      RECT 345.440 106.760 345.820 108.990 ;
      RECT 369.240 107.440 369.620 108.990 ;
      RECT 371.960 107.440 372.340 108.990 ;
      RECT 369.945 106.950 370.275 107.115 ;
      RECT 344.785 105.425 345.115 105.590 ;
      RECT 369.920 105.400 370.300 106.950 ;
      RECT 371.960 105.590 372.340 107.140 ;
      RECT 375.360 105.590 375.740 107.140 ;
      RECT 377.425 105.590 377.755 105.755 ;
      RECT 371.985 105.425 372.315 105.590 ;
      RECT 375.385 105.425 375.715 105.590 ;
      RECT 136.025 104.230 136.355 104.395 ;
      RECT 345.465 104.230 345.795 104.395 ;
      RECT 19.040 88.590 19.420 102.380 ;
      RECT 82.280 100.150 82.660 103.060 ;
      RECT 87.040 100.150 87.420 103.060 ;
      RECT 89.080 100.150 89.460 103.060 ;
      RECT 91.800 100.150 92.180 103.060 ;
      RECT 93.840 100.150 94.220 103.060 ;
      RECT 102.000 102.190 102.380 103.740 ;
      RECT 107.465 103.550 107.795 103.715 ;
      RECT 102.025 102.025 102.355 102.190 ;
      RECT 107.440 102.000 107.820 103.550 ;
      RECT 134.665 102.190 134.995 102.355 ;
      RECT 102.025 101.510 102.355 101.675 ;
      RECT 82.305 99.985 82.635 100.150 ;
      RECT 87.065 99.985 87.395 100.150 ;
      RECT 89.105 99.985 89.435 100.150 ;
      RECT 91.825 99.985 92.155 100.150 ;
      RECT 93.865 99.985 94.195 100.150 ;
      RECT 102.000 99.960 102.380 101.510 ;
      RECT 134.640 100.640 135.020 102.190 ;
      RECT 136.000 102.000 136.380 104.230 ;
      RECT 345.440 102.680 345.820 104.230 ;
      RECT 377.400 104.040 377.780 105.590 ;
      RECT 386.920 104.230 387.300 111.220 ;
      RECT 392.385 110.350 392.715 110.515 ;
      RECT 386.945 104.065 387.275 104.230 ;
      RECT 392.360 104.040 392.740 110.350 ;
      RECT 373.320 102.190 373.700 103.740 ;
      RECT 377.400 102.190 377.780 103.740 ;
      RECT 373.345 102.025 373.675 102.190 ;
      RECT 377.425 102.025 377.755 102.190 ;
      RECT 377.425 101.510 377.755 101.675 ;
      RECT 91.145 99.470 91.475 99.635 ;
      RECT 93.185 99.470 93.515 99.635 ;
      RECT 102.025 99.470 102.355 99.635 ;
      RECT 104.065 99.470 104.395 99.635 ;
      RECT 91.120 91.800 91.500 99.470 ;
      RECT 93.160 91.800 93.540 99.470 ;
      RECT 102.000 97.920 102.380 99.470 ;
      RECT 104.040 97.920 104.420 99.470 ;
      RECT 107.440 98.110 107.820 99.660 ;
      RECT 108.120 98.110 108.500 99.660 ;
      RECT 110.185 99.470 110.515 99.635 ;
      RECT 135.320 99.470 135.700 101.020 ;
      RECT 107.465 97.945 107.795 98.110 ;
      RECT 108.145 97.945 108.475 98.110 ;
      RECT 110.160 97.920 110.540 99.470 ;
      RECT 135.345 99.305 135.675 99.470 ;
      RECT 345.440 98.110 345.820 100.340 ;
      RECT 377.400 99.960 377.780 101.510 ;
      RECT 388.280 100.150 388.660 103.060 ;
      RECT 391.000 100.150 391.380 103.060 ;
      RECT 393.040 100.150 393.420 103.060 ;
      RECT 397.145 102.190 397.475 102.355 ;
      RECT 388.305 99.985 388.635 100.150 ;
      RECT 391.025 99.985 391.355 100.150 ;
      RECT 393.065 99.985 393.395 100.150 ;
      RECT 397.120 99.960 397.500 102.190 ;
      RECT 369.240 98.110 369.620 99.660 ;
      RECT 371.305 99.470 371.635 99.635 ;
      RECT 378.105 99.470 378.435 99.635 ;
      RECT 345.465 97.945 345.795 98.110 ;
      RECT 369.265 97.945 369.595 98.110 ;
      RECT 371.280 97.920 371.660 99.470 ;
      RECT 378.080 97.920 378.460 99.470 ;
      RECT 102.000 96.070 102.380 97.620 ;
      RECT 104.720 96.070 105.100 97.620 ;
      RECT 108.145 97.430 108.475 97.595 ;
      RECT 110.865 97.430 111.195 97.595 ;
      RECT 369.265 97.430 369.595 97.595 ;
      RECT 102.025 95.905 102.355 96.070 ;
      RECT 104.745 95.905 105.075 96.070 ;
      RECT 108.120 95.880 108.500 97.430 ;
      RECT 110.840 95.880 111.220 97.430 ;
      RECT 369.240 95.880 369.620 97.430 ;
      RECT 371.280 96.070 371.660 97.620 ;
      RECT 376.065 97.430 376.395 97.595 ;
      RECT 371.305 95.905 371.635 96.070 ;
      RECT 376.040 95.880 376.420 97.430 ;
      RECT 377.400 96.070 377.780 97.620 ;
      RECT 377.425 95.905 377.755 96.070 ;
      RECT 102.025 95.390 102.355 95.555 ;
      RECT 106.785 95.390 107.115 95.555 ;
      RECT 102.000 93.840 102.380 95.390 ;
      RECT 106.760 93.840 107.140 95.390 ;
      RECT 108.120 94.030 108.500 95.580 ;
      RECT 110.160 94.030 110.540 95.580 ;
      RECT 369.240 94.030 369.620 95.580 ;
      RECT 371.280 94.030 371.660 95.580 ;
      RECT 374.000 94.030 374.380 95.580 ;
      RECT 377.425 95.390 377.755 95.555 ;
      RECT 108.145 93.865 108.475 94.030 ;
      RECT 110.185 93.865 110.515 94.030 ;
      RECT 369.265 93.865 369.595 94.030 ;
      RECT 371.305 93.865 371.635 94.030 ;
      RECT 374.025 93.865 374.355 94.030 ;
      RECT 377.400 93.840 377.780 95.390 ;
      RECT 102.025 93.350 102.355 93.515 ;
      RECT 104.065 93.350 104.395 93.515 ;
      RECT 106.105 93.350 106.435 93.515 ;
      RECT 102.000 91.800 102.380 93.350 ;
      RECT 104.040 91.800 104.420 93.350 ;
      RECT 106.080 91.800 106.460 93.350 ;
      RECT 108.120 91.990 108.500 93.540 ;
      RECT 110.185 93.350 110.515 93.515 ;
      RECT 369.265 93.350 369.595 93.515 ;
      RECT 371.305 93.350 371.635 93.515 ;
      RECT 108.145 91.825 108.475 91.990 ;
      RECT 110.160 91.800 110.540 93.350 ;
      RECT 369.240 91.800 369.620 93.350 ;
      RECT 371.280 91.800 371.660 93.350 ;
      RECT 375.360 91.990 375.740 93.540 ;
      RECT 378.080 91.990 378.460 93.540 ;
      RECT 389.640 91.990 390.020 93.540 ;
      RECT 391.000 91.990 391.380 99.660 ;
      RECT 393.065 99.470 393.395 99.635 ;
      RECT 392.385 93.350 392.715 93.515 ;
      RECT 375.385 91.825 375.715 91.990 ;
      RECT 378.105 91.825 378.435 91.990 ;
      RECT 389.665 91.825 389.995 91.990 ;
      RECT 391.025 91.825 391.355 91.990 ;
      RECT 392.360 91.800 392.740 93.350 ;
      RECT 393.040 91.800 393.420 99.470 ;
      RECT 19.065 88.425 19.395 88.590 ;
      RECT 12.800 75.985 13.130 76.315 ;
      RECT 19.040 73.630 19.420 88.100 ;
      RECT 87.720 87.910 88.100 91.500 ;
      RECT 91.120 87.910 91.500 91.500 ;
      RECT 93.865 91.310 94.195 91.475 ;
      RECT 87.745 87.745 88.075 87.910 ;
      RECT 91.145 87.745 91.475 87.910 ;
      RECT 93.840 87.720 94.220 91.310 ;
      RECT 104.720 89.950 105.100 91.500 ;
      RECT 108.825 91.310 109.155 91.475 ;
      RECT 104.745 89.785 105.075 89.950 ;
      RECT 108.800 89.760 109.180 91.310 ;
      RECT 110.840 89.950 111.220 91.500 ;
      RECT 369.920 89.950 370.300 91.500 ;
      RECT 371.960 89.950 372.340 91.500 ;
      RECT 373.345 91.310 373.675 91.475 ;
      RECT 375.385 91.310 375.715 91.475 ;
      RECT 110.865 89.785 111.195 89.950 ;
      RECT 369.945 89.785 370.275 89.950 ;
      RECT 371.985 89.785 372.315 89.950 ;
      RECT 373.320 89.760 373.700 91.310 ;
      RECT 375.360 89.760 375.740 91.310 ;
      RECT 102.680 87.910 103.060 89.460 ;
      RECT 108.120 87.910 108.500 89.460 ;
      RECT 110.865 89.270 111.195 89.435 ;
      RECT 102.705 87.745 103.035 87.910 ;
      RECT 108.145 87.745 108.475 87.910 ;
      RECT 110.840 87.720 111.220 89.270 ;
      RECT 369.240 87.910 369.620 89.460 ;
      RECT 371.280 87.910 371.660 89.460 ;
      RECT 374.000 87.910 374.380 89.460 ;
      RECT 374.680 87.910 375.060 89.460 ;
      RECT 378.080 87.910 378.460 89.460 ;
      RECT 386.920 87.910 387.300 91.500 ;
      RECT 393.065 91.310 393.395 91.475 ;
      RECT 369.265 87.745 369.595 87.910 ;
      RECT 371.305 87.745 371.635 87.910 ;
      RECT 374.025 87.745 374.355 87.910 ;
      RECT 374.705 87.745 375.035 87.910 ;
      RECT 378.105 87.745 378.435 87.910 ;
      RECT 386.945 87.745 387.275 87.910 ;
      RECT 393.040 87.720 393.420 91.310 ;
      RECT 397.145 90.630 397.475 90.795 ;
      RECT 397.120 87.720 397.500 90.630 ;
      RECT 80.920 81.790 81.300 87.420 ;
      RECT 80.945 81.625 81.275 81.790 ;
      RECT 19.065 73.465 19.395 73.630 ;
      RECT 19.720 73.140 20.100 73.820 ;
      RECT 19.040 72.760 20.100 73.140 ;
      RECT 15.665 68.870 15.995 69.035 ;
      RECT 15.640 67.320 16.020 68.870 ;
      RECT 19.040 60.030 19.420 72.760 ;
      RECT 19.065 59.865 19.395 60.030 ;
      RECT 70.040 53.230 70.420 67.020 ;
      RECT 70.720 60.030 71.100 73.820 ;
      RECT 71.400 67.510 71.780 81.300 ;
      RECT 82.960 74.310 83.340 87.420 ;
      RECT 103.385 87.230 103.715 87.395 ;
      RECT 110.185 87.230 110.515 87.395 ;
      RECT 114.265 87.230 114.595 87.395 ;
      RECT 398.505 87.230 398.835 87.395 ;
      RECT 412.105 87.230 412.435 87.395 ;
      RECT 82.985 74.145 83.315 74.310 ;
      RECT 103.360 73.440 103.740 87.230 ;
      RECT 110.160 85.000 110.540 87.230 ;
      RECT 114.240 85.000 114.620 87.230 ;
      RECT 142.825 85.190 143.155 85.355 ;
      RECT 105.425 72.950 105.755 73.115 ;
      RECT 71.425 67.345 71.755 67.510 ;
      RECT 70.745 59.865 71.075 60.030 ;
      RECT 71.425 59.350 71.755 59.515 ;
      RECT 70.065 53.065 70.395 53.230 ;
      RECT 70.065 52.550 70.395 52.715 ;
      RECT 70.040 38.760 70.420 52.550 ;
      RECT 71.400 46.240 71.780 59.350 ;
      RECT 105.400 59.160 105.780 72.950 ;
      RECT 110.160 66.150 110.540 84.700 ;
      RECT 132.625 84.510 132.955 84.675 ;
      RECT 132.600 82.960 132.980 84.510 ;
      RECT 141.440 80.430 141.820 82.660 ;
      RECT 141.465 80.265 141.795 80.430 ;
      RECT 142.800 72.760 143.180 85.190 ;
      RECT 146.200 80.430 146.580 82.660 ;
      RECT 152.320 80.430 152.700 83.340 ;
      RECT 157.785 82.470 158.115 82.635 ;
      RECT 146.225 80.265 146.555 80.430 ;
      RECT 152.345 80.265 152.675 80.430 ;
      RECT 157.760 80.240 158.140 82.470 ;
      RECT 160.480 80.430 160.860 82.660 ;
      RECT 163.905 82.470 164.235 82.635 ;
      RECT 160.505 80.265 160.835 80.430 ;
      RECT 163.880 80.240 164.260 82.470 ;
      RECT 166.600 80.430 166.980 82.660 ;
      RECT 170.705 82.470 171.035 82.635 ;
      RECT 166.625 80.265 166.955 80.430 ;
      RECT 170.680 80.240 171.060 82.470 ;
      RECT 172.720 80.430 173.100 82.660 ;
      RECT 178.840 80.430 179.220 82.660 ;
      RECT 182.945 82.470 183.275 82.635 ;
      RECT 172.745 80.265 173.075 80.430 ;
      RECT 178.865 80.265 179.195 80.430 ;
      RECT 182.920 80.240 183.300 82.470 ;
      RECT 191.760 80.430 192.140 82.660 ;
      RECT 195.185 82.470 195.515 82.635 ;
      RECT 191.785 80.265 192.115 80.430 ;
      RECT 195.160 80.240 195.540 82.470 ;
      RECT 197.880 80.430 198.260 82.660 ;
      RECT 201.305 82.470 201.635 82.635 ;
      RECT 197.905 80.265 198.235 80.430 ;
      RECT 201.280 80.240 201.660 82.470 ;
      RECT 204.000 80.430 204.380 82.660 ;
      RECT 210.120 80.430 210.500 82.660 ;
      RECT 214.225 82.470 214.555 82.635 ;
      RECT 204.025 80.265 204.355 80.430 ;
      RECT 210.145 80.265 210.475 80.430 ;
      RECT 214.200 80.240 214.580 82.470 ;
      RECT 223.040 80.430 223.420 82.660 ;
      RECT 226.465 82.470 226.795 82.635 ;
      RECT 223.065 80.265 223.395 80.430 ;
      RECT 226.440 80.240 226.820 82.470 ;
      RECT 229.160 80.430 229.540 82.660 ;
      RECT 232.585 82.470 232.915 82.635 ;
      RECT 229.185 80.265 229.515 80.430 ;
      RECT 232.560 80.240 232.940 82.470 ;
      RECT 235.280 80.430 235.660 82.660 ;
      RECT 238.705 82.470 239.035 82.635 ;
      RECT 235.305 80.265 235.635 80.430 ;
      RECT 238.680 80.240 239.060 82.470 ;
      RECT 241.400 80.430 241.780 82.660 ;
      RECT 246.865 82.470 247.195 82.635 ;
      RECT 251.625 82.470 251.955 82.635 ;
      RECT 241.425 80.265 241.755 80.430 ;
      RECT 246.840 80.240 247.220 82.470 ;
      RECT 251.600 80.240 251.980 82.470 ;
      RECT 253.640 80.430 254.020 82.660 ;
      RECT 257.745 82.470 258.075 82.635 ;
      RECT 253.665 80.265 253.995 80.430 ;
      RECT 257.720 80.240 258.100 82.470 ;
      RECT 259.760 80.430 260.140 82.660 ;
      RECT 266.560 80.430 266.940 82.660 ;
      RECT 269.985 82.470 270.315 82.635 ;
      RECT 259.785 80.265 260.115 80.430 ;
      RECT 266.585 80.265 266.915 80.430 ;
      RECT 269.960 80.240 270.340 82.470 ;
      RECT 272.680 80.430 273.060 82.660 ;
      RECT 276.785 82.470 277.115 82.635 ;
      RECT 272.705 80.265 273.035 80.430 ;
      RECT 276.760 80.240 277.140 82.470 ;
      RECT 278.800 80.430 279.180 82.660 ;
      RECT 282.225 82.470 282.555 82.635 ;
      RECT 278.825 80.265 279.155 80.430 ;
      RECT 282.200 80.240 282.580 82.470 ;
      RECT 284.920 80.430 285.300 82.660 ;
      RECT 289.025 82.470 289.355 82.635 ;
      RECT 284.945 80.265 285.275 80.430 ;
      RECT 289.000 80.240 289.380 82.470 ;
      RECT 289.680 80.430 290.060 82.660 ;
      RECT 295.145 82.470 295.475 82.635 ;
      RECT 289.705 80.265 290.035 80.430 ;
      RECT 295.120 80.240 295.500 82.470 ;
      RECT 297.840 80.430 298.220 82.660 ;
      RECT 301.265 82.470 301.595 82.635 ;
      RECT 297.865 80.265 298.195 80.430 ;
      RECT 301.240 80.240 301.620 82.470 ;
      RECT 303.960 80.430 304.340 82.660 ;
      RECT 310.080 80.430 310.460 82.660 ;
      RECT 316.200 80.430 316.580 82.660 ;
      RECT 320.960 80.430 321.340 83.340 ;
      RECT 326.425 82.470 326.755 82.635 ;
      RECT 303.985 80.265 304.315 80.430 ;
      RECT 310.105 80.265 310.435 80.430 ;
      RECT 316.225 80.265 316.555 80.430 ;
      RECT 320.985 80.265 321.315 80.430 ;
      RECT 326.400 80.240 326.780 82.470 ;
      RECT 328.440 80.430 328.820 82.660 ;
      RECT 332.545 82.470 332.875 82.635 ;
      RECT 328.465 80.265 328.795 80.430 ;
      RECT 332.520 80.240 332.900 82.470 ;
      RECT 335.240 80.430 335.620 82.660 ;
      RECT 338.665 82.470 338.995 82.635 ;
      RECT 335.265 80.265 335.595 80.430 ;
      RECT 338.640 80.240 339.020 82.470 ;
      RECT 341.360 80.430 341.740 82.660 ;
      RECT 341.385 80.265 341.715 80.430 ;
      RECT 110.185 65.985 110.515 66.150 ;
      RECT 155.720 63.430 156.100 71.780 ;
      RECT 155.745 63.265 156.075 63.430 ;
      RECT 290.360 60.030 290.740 79.940 ;
      RECT 398.480 78.880 398.860 87.230 ;
      RECT 412.080 85.680 412.460 87.230 ;
      RECT 412.080 72.270 412.460 85.380 ;
      RECT 412.785 78.390 413.115 78.555 ;
      RECT 412.105 72.105 412.435 72.270 ;
      RECT 411.425 70.910 411.755 71.075 ;
      RECT 290.385 59.865 290.715 60.030 ;
      RECT 142.145 59.350 142.475 59.515 ;
      RECT 148.945 59.350 149.275 59.515 ;
      RECT 155.065 59.350 155.395 59.515 ;
      RECT 160.505 59.350 160.835 59.515 ;
      RECT 167.305 59.350 167.635 59.515 ;
      RECT 173.425 59.350 173.755 59.515 ;
      RECT 180.225 59.350 180.555 59.515 ;
      RECT 185.665 59.350 185.995 59.515 ;
      RECT 192.465 59.350 192.795 59.515 ;
      RECT 198.585 59.350 198.915 59.515 ;
      RECT 204.025 59.350 204.355 59.515 ;
      RECT 210.825 59.350 211.155 59.515 ;
      RECT 216.945 59.350 217.275 59.515 ;
      RECT 223.745 59.350 224.075 59.515 ;
      RECT 229.185 59.350 229.515 59.515 ;
      RECT 235.985 59.350 236.315 59.515 ;
      RECT 242.105 59.350 242.435 59.515 ;
      RECT 248.905 59.350 249.235 59.515 ;
      RECT 255.025 59.350 255.355 59.515 ;
      RECT 260.465 59.350 260.795 59.515 ;
      RECT 267.265 59.350 267.595 59.515 ;
      RECT 272.705 59.350 273.035 59.515 ;
      RECT 280.185 59.350 280.515 59.515 ;
      RECT 285.625 59.350 285.955 59.515 ;
      RECT 292.425 59.350 292.755 59.515 ;
      RECT 298.545 59.350 298.875 59.515 ;
      RECT 303.985 59.350 304.315 59.515 ;
      RECT 310.785 59.350 311.115 59.515 ;
      RECT 316.905 59.350 317.235 59.515 ;
      RECT 142.120 55.760 142.500 59.350 ;
      RECT 148.920 55.760 149.300 59.350 ;
      RECT 155.040 55.760 155.420 59.350 ;
      RECT 160.480 55.760 160.860 59.350 ;
      RECT 167.280 55.760 167.660 59.350 ;
      RECT 173.400 55.760 173.780 59.350 ;
      RECT 180.200 55.760 180.580 59.350 ;
      RECT 185.640 55.760 186.020 59.350 ;
      RECT 192.440 55.760 192.820 59.350 ;
      RECT 198.560 55.760 198.940 59.350 ;
      RECT 204.000 55.760 204.380 59.350 ;
      RECT 210.800 55.760 211.180 59.350 ;
      RECT 216.920 55.760 217.300 59.350 ;
      RECT 223.720 55.760 224.100 59.350 ;
      RECT 229.160 55.760 229.540 59.350 ;
      RECT 235.960 55.760 236.340 59.350 ;
      RECT 242.080 55.760 242.460 59.350 ;
      RECT 248.880 55.760 249.260 59.350 ;
      RECT 255.000 55.760 255.380 59.350 ;
      RECT 260.440 55.760 260.820 59.350 ;
      RECT 267.240 55.760 267.620 59.350 ;
      RECT 272.680 55.760 273.060 59.350 ;
      RECT 280.160 55.760 280.540 59.350 ;
      RECT 285.600 55.760 285.980 59.350 ;
      RECT 292.400 55.760 292.780 59.350 ;
      RECT 298.520 55.760 298.900 59.350 ;
      RECT 303.960 55.760 304.340 59.350 ;
      RECT 310.760 55.760 311.140 59.350 ;
      RECT 316.880 55.760 317.260 59.350 ;
      RECT 323.000 55.460 323.380 63.620 ;
      RECT 323.705 59.350 324.035 59.515 ;
      RECT 329.145 59.350 329.475 59.515 ;
      RECT 335.945 59.350 336.275 59.515 ;
      RECT 323.680 55.760 324.060 59.350 ;
      RECT 329.120 55.760 329.500 59.350 ;
      RECT 335.920 55.760 336.300 59.350 ;
      RECT 411.400 57.800 411.780 70.910 ;
      RECT 412.760 64.600 413.140 78.390 ;
      RECT 412.105 64.110 412.435 64.275 ;
      RECT 139.425 53.230 139.755 53.395 ;
      RECT 12.945 34.870 13.275 35.035 ;
      RECT 12.920 31.960 13.300 34.870 ;
      RECT 70.720 32.150 71.100 45.940 ;
      RECT 71.425 38.270 71.755 38.435 ;
      RECT 70.745 31.985 71.075 32.150 ;
      RECT 29.265 27.390 29.595 27.555 ;
      RECT 10.905 8.350 11.235 8.515 ;
      RECT 19.745 8.350 20.075 8.515 ;
      RECT 27.225 8.350 27.555 8.515 ;
      RECT 10.880 6.120 11.260 8.350 ;
      RECT 19.720 6.120 20.100 8.350 ;
      RECT 27.200 6.120 27.580 8.350 ;
      RECT 29.240 1.060 29.620 27.390 ;
      RECT 71.400 25.160 71.780 38.270 ;
      RECT 138.720 35.550 139.100 44.580 ;
      RECT 138.745 35.385 139.075 35.550 ;
      RECT 79.585 31.470 79.915 31.635 ;
      RECT 79.560 19.040 79.940 31.470 ;
      RECT 117.720 31.065 118.050 31.395 ;
      RECT 100.200 29.845 100.530 30.175 ;
      RECT 88.520 27.405 88.850 27.735 ;
      RECT 80.265 23.990 80.595 24.155 ;
      RECT 77.545 14.470 77.875 14.635 ;
      RECT 36.065 8.350 36.395 8.515 ;
      RECT 44.905 8.350 45.235 8.515 ;
      RECT 52.385 8.350 52.715 8.515 ;
      RECT 61.225 8.350 61.555 8.515 ;
      RECT 70.065 8.350 70.395 8.515 ;
      RECT 36.040 6.120 36.420 8.350 ;
      RECT 44.880 6.120 45.260 8.350 ;
      RECT 52.360 6.120 52.740 8.350 ;
      RECT 61.200 6.120 61.580 8.350 ;
      RECT 70.040 6.120 70.420 8.350 ;
      RECT 77.520 1.060 77.900 14.470 ;
      RECT 80.240 12.240 80.620 23.990 ;
      RECT 86.385 18.550 86.715 18.715 ;
      RECT 83.665 14.470 83.995 14.635 ;
      RECT 78.905 8.350 79.235 8.515 ;
      RECT 78.880 6.120 79.260 8.350 ;
      RECT 83.640 1.060 84.020 14.470 ;
      RECT 86.360 8.840 86.740 18.550 ;
      RECT 88.535 15.410 88.835 27.405 ;
      RECT 94.360 20.085 94.690 20.415 ;
      RECT 94.375 15.410 94.675 20.085 ;
      RECT 100.215 15.410 100.515 29.845 ;
      RECT 111.880 28.625 112.210 28.955 ;
      RECT 106.040 21.305 106.370 21.635 ;
      RECT 106.055 15.410 106.355 21.305 ;
      RECT 111.895 15.410 112.195 28.625 ;
      RECT 117.735 15.410 118.035 31.065 ;
      RECT 135.240 24.965 135.570 25.295 ;
      RECT 129.400 23.745 129.730 24.075 ;
      RECT 123.560 22.525 123.890 22.855 ;
      RECT 123.575 15.410 123.875 22.525 ;
      RECT 129.415 15.410 129.715 23.745 ;
      RECT 135.255 15.410 135.555 24.965 ;
      RECT 88.520 15.080 88.850 15.410 ;
      RECT 94.360 15.080 94.690 15.410 ;
      RECT 100.200 15.080 100.530 15.410 ;
      RECT 106.040 15.080 106.370 15.410 ;
      RECT 111.880 15.080 112.210 15.410 ;
      RECT 117.720 15.080 118.050 15.410 ;
      RECT 123.560 15.080 123.890 15.410 ;
      RECT 129.400 15.080 129.730 15.410 ;
      RECT 135.240 15.080 135.570 15.410 ;
      RECT 89.105 14.470 89.435 14.635 ;
      RECT 95.905 14.470 96.235 14.635 ;
      RECT 100.665 14.470 100.995 14.635 ;
      RECT 106.785 14.470 107.115 14.635 ;
      RECT 112.905 14.470 113.235 14.635 ;
      RECT 118.345 14.470 118.675 14.635 ;
      RECT 125.145 14.470 125.475 14.635 ;
      RECT 130.585 14.470 130.915 14.635 ;
      RECT 136.025 14.470 136.355 14.635 ;
      RECT 87.065 8.350 87.395 8.515 ;
      RECT 87.040 6.120 87.420 8.350 ;
      RECT 89.080 1.060 89.460 14.470 ;
      RECT 94.545 8.350 94.875 8.515 ;
      RECT 94.520 6.120 94.900 8.350 ;
      RECT 95.880 1.060 96.260 14.470 ;
      RECT 100.640 1.060 101.020 14.470 ;
      RECT 103.385 8.350 103.715 8.515 ;
      RECT 103.360 6.120 103.740 8.350 ;
      RECT 106.760 1.060 107.140 14.470 ;
      RECT 112.225 8.350 112.555 8.515 ;
      RECT 112.200 6.120 112.580 8.350 ;
      RECT 112.880 1.060 113.260 14.470 ;
      RECT 118.320 1.060 118.700 14.470 ;
      RECT 119.705 8.350 120.035 8.515 ;
      RECT 119.680 6.120 120.060 8.350 ;
      RECT 125.120 1.060 125.500 14.470 ;
      RECT 128.545 8.350 128.875 8.515 ;
      RECT 128.520 6.120 128.900 8.350 ;
      RECT 130.560 1.060 130.940 14.470 ;
      RECT 133.305 11.750 133.635 11.915 ;
      RECT 133.280 2.720 133.660 11.750 ;
      RECT 136.000 1.060 136.380 14.470 ;
      RECT 137.385 8.350 137.715 8.515 ;
      RECT 137.360 6.120 137.740 8.350 ;
      RECT 139.400 1.060 139.780 53.230 ;
      RECT 142.800 50.510 143.180 53.420 ;
      RECT 146.225 53.230 146.555 53.395 ;
      RECT 142.825 50.345 143.155 50.510 ;
      RECT 142.145 49.150 142.475 49.315 ;
      RECT 141.465 47.110 141.795 47.275 ;
      RECT 140.760 40.990 141.140 43.220 ;
      RECT 141.440 42.840 141.820 47.110 ;
      RECT 142.120 46.240 142.500 49.150 ;
      RECT 141.815 41.830 142.145 42.160 ;
      RECT 140.785 40.825 141.115 40.990 ;
      RECT 140.390 36.230 140.720 36.560 ;
      RECT 140.405 27.735 140.705 36.230 ;
      RECT 141.830 28.955 142.130 41.830 ;
      RECT 141.815 28.625 142.145 28.955 ;
      RECT 140.390 27.405 140.720 27.735 ;
      RECT 141.080 26.185 141.410 26.515 ;
      RECT 141.095 15.410 141.395 26.185 ;
      RECT 141.080 15.080 141.410 15.410 ;
      RECT 141.465 14.470 141.795 14.635 ;
      RECT 141.440 1.060 141.820 14.470 ;
      RECT 144.865 8.350 145.195 8.515 ;
      RECT 144.840 6.120 145.220 8.350 ;
      RECT 146.200 1.060 146.580 53.230 ;
      RECT 148.920 50.510 149.300 53.420 ;
      RECT 151.665 53.230 151.995 53.395 ;
      RECT 148.945 50.345 149.275 50.510 ;
      RECT 148.945 49.150 149.275 49.315 ;
      RECT 148.265 47.110 148.595 47.275 ;
      RECT 148.240 42.840 148.620 47.110 ;
      RECT 148.920 46.240 149.300 49.150 ;
      RECT 148.055 41.830 148.385 42.160 ;
      RECT 148.070 31.395 148.370 41.830 ;
      RECT 148.055 31.065 148.385 31.395 ;
      RECT 146.920 27.405 147.250 27.735 ;
      RECT 146.935 15.410 147.235 27.405 ;
      RECT 146.920 15.080 147.250 15.410 ;
      RECT 148.265 14.470 148.595 14.635 ;
      RECT 148.240 1.060 148.620 14.470 ;
      RECT 151.640 1.060 152.020 53.230 ;
      RECT 154.360 50.510 154.740 53.420 ;
      RECT 159.825 53.230 160.155 53.395 ;
      RECT 154.385 50.345 154.715 50.510 ;
      RECT 154.385 49.150 154.715 49.315 ;
      RECT 153.705 47.110 154.035 47.275 ;
      RECT 153.680 42.840 154.060 47.110 ;
      RECT 154.360 46.240 154.740 49.150 ;
      RECT 154.295 41.830 154.625 42.160 ;
      RECT 152.760 28.625 153.090 28.955 ;
      RECT 152.775 15.410 153.075 28.625 ;
      RECT 154.310 22.855 154.610 41.830 ;
      RECT 154.295 22.525 154.625 22.855 ;
      RECT 158.600 22.525 158.930 22.855 ;
      RECT 158.615 15.410 158.915 22.525 ;
      RECT 152.760 15.080 153.090 15.410 ;
      RECT 158.600 15.080 158.930 15.410 ;
      RECT 153.705 14.470 154.035 14.635 ;
      RECT 159.145 14.470 159.475 14.635 ;
      RECT 153.025 8.350 153.355 8.515 ;
      RECT 153.000 6.120 153.380 8.350 ;
      RECT 153.680 1.060 154.060 14.470 ;
      RECT 159.120 1.060 159.500 14.470 ;
      RECT 159.800 1.060 160.180 53.230 ;
      RECT 161.160 50.510 161.540 53.420 ;
      RECT 165.945 53.230 166.275 53.395 ;
      RECT 161.185 50.345 161.515 50.510 ;
      RECT 161.865 49.150 162.195 49.315 ;
      RECT 161.185 47.110 161.515 47.275 ;
      RECT 161.160 42.840 161.540 47.110 ;
      RECT 161.840 46.240 162.220 49.150 ;
      RECT 160.535 41.830 160.865 42.160 ;
      RECT 160.550 24.075 160.850 41.830 ;
      RECT 160.535 23.745 160.865 24.075 ;
      RECT 164.440 23.745 164.770 24.075 ;
      RECT 164.455 15.410 164.755 23.745 ;
      RECT 164.440 15.080 164.770 15.410 ;
      RECT 165.265 14.470 165.595 14.635 ;
      RECT 161.865 8.350 162.195 8.515 ;
      RECT 161.840 6.120 162.220 8.350 ;
      RECT 165.240 1.060 165.620 14.470 ;
      RECT 165.920 1.060 166.300 53.230 ;
      RECT 167.280 50.510 167.660 53.420 ;
      RECT 172.065 53.230 172.395 53.395 ;
      RECT 167.305 50.345 167.635 50.510 ;
      RECT 167.985 49.150 168.315 49.315 ;
      RECT 167.305 47.110 167.635 47.275 ;
      RECT 167.280 42.840 167.660 47.110 ;
      RECT 167.960 46.240 168.340 49.150 ;
      RECT 166.775 41.830 167.105 42.160 ;
      RECT 166.790 25.295 167.090 41.830 ;
      RECT 166.775 24.965 167.105 25.295 ;
      RECT 170.280 24.965 170.610 25.295 ;
      RECT 170.295 15.410 170.595 24.965 ;
      RECT 170.280 15.080 170.610 15.410 ;
      RECT 170.705 14.470 171.035 14.635 ;
      RECT 170.025 8.350 170.355 8.515 ;
      RECT 170.000 6.120 170.380 8.350 ;
      RECT 170.680 1.060 171.060 14.470 ;
      RECT 172.040 1.060 172.420 53.230 ;
      RECT 174.080 50.510 174.460 53.420 ;
      RECT 178.185 53.230 178.515 53.395 ;
      RECT 174.105 50.345 174.435 50.510 ;
      RECT 174.105 49.150 174.435 49.315 ;
      RECT 173.425 47.110 173.755 47.275 ;
      RECT 173.400 42.840 173.780 47.110 ;
      RECT 174.080 46.240 174.460 49.150 ;
      RECT 173.015 41.830 173.345 42.160 ;
      RECT 173.030 26.515 173.330 41.830 ;
      RECT 173.015 26.185 173.345 26.515 ;
      RECT 176.120 26.185 176.450 26.515 ;
      RECT 176.135 15.410 176.435 26.185 ;
      RECT 176.120 15.080 176.450 15.410 ;
      RECT 177.505 14.470 177.835 14.635 ;
      RECT 177.480 1.060 177.860 14.470 ;
      RECT 178.160 1.060 178.540 53.230 ;
      RECT 180.200 50.510 180.580 53.420 ;
      RECT 184.305 53.230 184.635 53.395 ;
      RECT 180.225 50.345 180.555 50.510 ;
      RECT 180.225 49.150 180.555 49.315 ;
      RECT 179.545 47.110 179.875 47.275 ;
      RECT 179.520 42.840 179.900 47.110 ;
      RECT 180.200 46.240 180.580 49.150 ;
      RECT 179.255 41.830 179.585 42.160 ;
      RECT 179.270 27.735 179.570 41.830 ;
      RECT 179.255 27.405 179.585 27.735 ;
      RECT 181.960 27.405 182.290 27.735 ;
      RECT 181.975 15.410 182.275 27.405 ;
      RECT 181.960 15.080 182.290 15.410 ;
      RECT 182.945 14.470 183.275 14.635 ;
      RECT 178.865 8.350 179.195 8.515 ;
      RECT 178.840 6.120 179.220 8.350 ;
      RECT 182.920 1.060 183.300 14.470 ;
      RECT 184.280 1.060 184.660 53.230 ;
      RECT 185.640 50.510 186.020 53.420 ;
      RECT 189.065 53.230 189.395 53.395 ;
      RECT 185.665 50.345 185.995 50.510 ;
      RECT 186.345 49.150 186.675 49.315 ;
      RECT 185.665 47.110 185.995 47.275 ;
      RECT 185.640 42.840 186.020 47.110 ;
      RECT 186.320 46.240 186.700 49.150 ;
      RECT 185.495 41.830 185.825 42.160 ;
      RECT 185.510 28.955 185.810 41.830 ;
      RECT 185.495 28.625 185.825 28.955 ;
      RECT 187.800 28.625 188.130 28.955 ;
      RECT 187.815 15.410 188.115 28.625 ;
      RECT 187.800 15.080 188.130 15.410 ;
      RECT 188.385 14.470 188.715 14.635 ;
      RECT 187.025 8.350 187.355 8.515 ;
      RECT 187.000 6.120 187.380 8.350 ;
      RECT 188.360 1.060 188.740 14.470 ;
      RECT 189.040 1.060 189.420 53.230 ;
      RECT 191.105 49.150 191.435 49.315 ;
      RECT 191.080 46.240 191.460 49.150 ;
      RECT 192.440 47.790 192.820 55.460 ;
      RECT 323.000 55.080 324.060 55.460 ;
      RECT 323.680 53.910 324.060 55.080 ;
      RECT 323.705 53.745 324.035 53.910 ;
      RECT 193.120 50.510 193.500 53.420 ;
      RECT 196.545 53.230 196.875 53.395 ;
      RECT 193.145 50.345 193.475 50.510 ;
      RECT 192.465 47.625 192.795 47.790 ;
      RECT 191.785 47.110 192.115 47.275 ;
      RECT 191.760 42.840 192.140 47.110 ;
      RECT 191.735 41.830 192.065 42.160 ;
      RECT 190.310 36.230 190.640 36.560 ;
      RECT 190.325 20.415 190.625 36.230 ;
      RECT 191.750 22.855 192.050 41.830 ;
      RECT 193.640 31.065 193.970 31.395 ;
      RECT 191.735 22.525 192.065 22.855 ;
      RECT 190.310 20.085 190.640 20.415 ;
      RECT 193.655 15.410 193.955 31.065 ;
      RECT 193.640 15.080 193.970 15.410 ;
      RECT 194.505 14.470 194.835 14.635 ;
      RECT 194.480 1.060 194.860 14.470 ;
      RECT 195.865 8.350 196.195 8.515 ;
      RECT 195.840 6.120 196.220 8.350 ;
      RECT 196.520 1.060 196.900 53.230 ;
      RECT 198.560 50.510 198.940 53.420 ;
      RECT 203.345 53.230 203.675 53.395 ;
      RECT 198.585 50.345 198.915 50.510 ;
      RECT 198.585 49.150 198.915 49.315 ;
      RECT 197.905 47.110 198.235 47.275 ;
      RECT 197.880 42.840 198.260 47.110 ;
      RECT 198.560 46.240 198.940 49.150 ;
      RECT 197.975 41.830 198.305 42.160 ;
      RECT 197.990 24.075 198.290 41.830 ;
      RECT 199.480 32.285 199.810 32.615 ;
      RECT 197.975 23.745 198.305 24.075 ;
      RECT 199.495 15.410 199.795 32.285 ;
      RECT 199.480 15.080 199.810 15.410 ;
      RECT 201.305 14.470 201.635 14.635 ;
      RECT 201.280 1.060 201.660 14.470 ;
      RECT 202.665 8.350 202.995 8.515 ;
      RECT 202.640 6.120 203.020 8.350 ;
      RECT 203.320 1.060 203.700 53.230 ;
      RECT 204.680 50.510 205.060 53.420 ;
      RECT 208.785 53.230 209.115 53.395 ;
      RECT 209.465 53.230 209.795 53.395 ;
      RECT 204.705 50.345 205.035 50.510 ;
      RECT 208.760 50.320 209.140 53.230 ;
      RECT 205.385 49.150 205.715 49.315 ;
      RECT 204.705 47.110 205.035 47.275 ;
      RECT 204.680 42.840 205.060 47.110 ;
      RECT 205.360 46.240 205.740 49.150 ;
      RECT 204.215 41.830 204.545 42.160 ;
      RECT 204.230 25.295 204.530 41.830 ;
      RECT 204.215 24.965 204.545 25.295 ;
      RECT 205.320 20.085 205.650 20.415 ;
      RECT 205.335 15.410 205.635 20.085 ;
      RECT 205.320 15.080 205.650 15.410 ;
      RECT 206.745 14.470 207.075 14.635 ;
      RECT 206.720 1.060 207.100 14.470 ;
      RECT 209.440 1.060 209.820 53.230 ;
      RECT 211.480 50.510 211.860 53.420 ;
      RECT 215.585 53.230 215.915 53.395 ;
      RECT 211.505 50.345 211.835 50.510 ;
      RECT 211.505 49.150 211.835 49.315 ;
      RECT 210.825 47.110 211.155 47.275 ;
      RECT 210.800 42.840 211.180 47.110 ;
      RECT 211.480 46.240 211.860 49.150 ;
      RECT 210.455 41.830 210.785 42.160 ;
      RECT 210.470 26.515 210.770 41.830 ;
      RECT 210.455 26.185 210.785 26.515 ;
      RECT 211.160 22.525 211.490 22.855 ;
      RECT 211.175 15.410 211.475 22.525 ;
      RECT 211.160 15.080 211.490 15.410 ;
      RECT 212.185 14.470 212.515 14.635 ;
      RECT 211.505 8.350 211.835 8.515 ;
      RECT 211.480 6.120 211.860 8.350 ;
      RECT 212.160 1.060 212.540 14.470 ;
      RECT 215.560 1.060 215.940 53.230 ;
      RECT 217.600 50.510 217.980 53.420 ;
      RECT 221.705 53.230 222.035 53.395 ;
      RECT 217.625 50.345 217.955 50.510 ;
      RECT 216.945 47.110 217.275 47.275 ;
      RECT 216.920 42.840 217.300 47.110 ;
      RECT 217.600 45.070 217.980 49.340 ;
      RECT 217.625 44.905 217.955 45.070 ;
      RECT 216.695 41.830 217.025 42.160 ;
      RECT 216.710 27.735 217.010 41.830 ;
      RECT 216.695 27.405 217.025 27.735 ;
      RECT 217.000 23.745 217.330 24.075 ;
      RECT 217.015 15.410 217.315 23.745 ;
      RECT 217.000 15.080 217.330 15.410 ;
      RECT 217.625 14.470 217.955 14.635 ;
      RECT 217.600 1.060 217.980 14.470 ;
      RECT 221.025 8.350 221.355 8.515 ;
      RECT 221.000 6.120 221.380 8.350 ;
      RECT 221.680 1.060 222.060 53.230 ;
      RECT 223.720 50.510 224.100 53.420 ;
      RECT 226.465 53.230 226.795 53.395 ;
      RECT 227.825 53.230 228.155 53.395 ;
      RECT 223.745 50.345 224.075 50.510 ;
      RECT 226.440 50.320 226.820 53.230 ;
      RECT 223.745 49.150 224.075 49.315 ;
      RECT 223.065 47.110 223.395 47.275 ;
      RECT 223.040 42.840 223.420 47.110 ;
      RECT 223.720 46.240 224.100 49.150 ;
      RECT 222.935 41.830 223.265 42.160 ;
      RECT 222.950 28.955 223.250 41.830 ;
      RECT 222.935 28.625 223.265 28.955 ;
      RECT 222.840 24.965 223.170 25.295 ;
      RECT 222.855 15.410 223.155 24.965 ;
      RECT 222.840 15.080 223.170 15.410 ;
      RECT 224.425 14.470 224.755 14.635 ;
      RECT 224.400 1.060 224.780 14.470 ;
      RECT 227.800 1.060 228.180 53.230 ;
      RECT 229.840 50.510 230.220 53.420 ;
      RECT 233.265 53.230 233.595 53.395 ;
      RECT 229.865 50.345 230.195 50.510 ;
      RECT 229.865 49.150 230.195 49.315 ;
      RECT 229.185 47.110 229.515 47.275 ;
      RECT 229.160 42.840 229.540 47.110 ;
      RECT 229.840 46.240 230.220 49.150 ;
      RECT 229.175 41.830 229.505 42.160 ;
      RECT 229.190 31.395 229.490 41.830 ;
      RECT 229.175 31.065 229.505 31.395 ;
      RECT 228.680 26.185 229.010 26.515 ;
      RECT 228.695 15.410 228.995 26.185 ;
      RECT 228.680 15.080 229.010 15.410 ;
      RECT 229.865 14.470 230.195 14.635 ;
      RECT 229.185 8.350 229.515 8.515 ;
      RECT 229.160 6.120 229.540 8.350 ;
      RECT 229.840 1.060 230.220 14.470 ;
      RECT 233.240 1.060 233.620 53.230 ;
      RECT 235.960 50.510 236.340 53.420 ;
      RECT 238.705 53.230 239.035 53.395 ;
      RECT 239.385 53.230 239.715 53.395 ;
      RECT 235.985 50.345 236.315 50.510 ;
      RECT 238.680 50.320 239.060 53.230 ;
      RECT 235.985 49.150 236.315 49.315 ;
      RECT 235.305 47.110 235.635 47.275 ;
      RECT 235.280 42.840 235.660 47.110 ;
      RECT 235.960 46.240 236.340 49.150 ;
      RECT 235.415 41.830 235.745 42.160 ;
      RECT 235.430 32.615 235.730 41.830 ;
      RECT 235.415 32.285 235.745 32.615 ;
      RECT 234.520 27.405 234.850 27.735 ;
      RECT 234.535 15.410 234.835 27.405 ;
      RECT 234.520 15.080 234.850 15.410 ;
      RECT 235.305 14.470 235.635 14.635 ;
      RECT 235.280 1.060 235.660 14.470 ;
      RECT 237.345 8.350 237.675 8.515 ;
      RECT 237.320 6.120 237.700 8.350 ;
      RECT 239.360 1.060 239.740 53.230 ;
      RECT 242.080 50.510 242.460 53.420 ;
      RECT 244.825 53.230 245.155 53.395 ;
      RECT 245.505 53.230 245.835 53.395 ;
      RECT 244.800 51.680 245.180 53.230 ;
      RECT 242.105 50.345 242.435 50.510 ;
      RECT 242.105 49.150 242.435 49.315 ;
      RECT 241.425 47.110 241.755 47.275 ;
      RECT 241.400 42.840 241.780 47.110 ;
      RECT 242.080 46.240 242.460 49.150 ;
      RECT 241.655 41.830 241.985 42.160 ;
      RECT 240.230 36.230 240.560 36.560 ;
      RECT 240.245 30.175 240.545 36.230 ;
      RECT 240.230 29.845 240.560 30.175 ;
      RECT 240.360 28.625 240.690 28.955 ;
      RECT 240.375 15.410 240.675 28.625 ;
      RECT 241.670 20.415 241.970 41.830 ;
      RECT 241.655 20.085 241.985 20.415 ;
      RECT 240.360 15.080 240.690 15.410 ;
      RECT 241.425 14.470 241.755 14.635 ;
      RECT 241.400 1.060 241.780 14.470 ;
      RECT 244.825 8.350 245.155 8.515 ;
      RECT 244.800 6.120 245.180 8.350 ;
      RECT 245.480 1.060 245.860 53.230 ;
      RECT 248.200 51.870 248.580 53.420 ;
      RECT 248.225 51.705 248.555 51.870 ;
      RECT 248.880 50.510 249.260 53.420 ;
      RECT 252.985 53.230 253.315 53.395 ;
      RECT 248.905 50.345 249.235 50.510 ;
      RECT 248.905 49.150 249.235 49.315 ;
      RECT 248.225 47.110 248.555 47.275 ;
      RECT 248.200 42.840 248.580 47.110 ;
      RECT 248.880 46.240 249.260 49.150 ;
      RECT 247.895 41.830 248.225 42.160 ;
      RECT 247.910 22.855 248.210 41.830 ;
      RECT 247.895 22.525 248.225 22.855 ;
      RECT 252.040 22.525 252.370 22.855 ;
      RECT 246.200 20.085 246.530 20.415 ;
      RECT 246.215 15.410 246.515 20.085 ;
      RECT 252.055 15.410 252.355 22.525 ;
      RECT 246.200 15.080 246.530 15.410 ;
      RECT 252.040 15.080 252.370 15.410 ;
      RECT 246.865 14.470 247.195 14.635 ;
      RECT 246.840 1.060 247.220 14.470 ;
      RECT 252.960 1.060 253.340 53.230 ;
      RECT 255.000 50.510 255.380 53.420 ;
      RECT 257.065 53.230 257.395 53.395 ;
      RECT 255.025 50.345 255.355 50.510 ;
      RECT 254.345 49.150 254.675 49.315 ;
      RECT 253.665 47.110 253.995 47.275 ;
      RECT 253.640 42.840 254.020 47.110 ;
      RECT 254.320 46.240 254.700 49.150 ;
      RECT 254.135 41.830 254.465 42.160 ;
      RECT 254.150 24.075 254.450 41.830 ;
      RECT 254.135 23.745 254.465 24.075 ;
      RECT 253.665 14.470 253.995 14.635 ;
      RECT 253.640 1.060 254.020 14.470 ;
      RECT 255.025 8.350 255.355 8.515 ;
      RECT 255.000 6.120 255.380 8.350 ;
      RECT 257.040 1.060 257.420 53.230 ;
      RECT 261.120 50.510 261.500 53.420 ;
      RECT 265.905 53.230 266.235 53.395 ;
      RECT 261.145 50.345 261.475 50.510 ;
      RECT 259.785 47.110 260.115 47.275 ;
      RECT 259.760 42.840 260.140 47.110 ;
      RECT 260.440 45.070 260.820 49.340 ;
      RECT 260.465 44.905 260.795 45.070 ;
      RECT 260.375 41.830 260.705 42.160 ;
      RECT 260.390 25.295 260.690 41.830 ;
      RECT 260.375 24.965 260.705 25.295 ;
      RECT 263.720 24.965 264.050 25.295 ;
      RECT 257.880 23.745 258.210 24.075 ;
      RECT 257.895 15.410 258.195 23.745 ;
      RECT 263.735 15.410 264.035 24.965 ;
      RECT 257.880 15.080 258.210 15.410 ;
      RECT 263.720 15.080 264.050 15.410 ;
      RECT 259.105 14.470 259.435 14.635 ;
      RECT 264.545 14.470 264.875 14.635 ;
      RECT 259.080 1.060 259.460 14.470 ;
      RECT 263.185 8.350 263.515 8.515 ;
      RECT 263.160 6.120 263.540 8.350 ;
      RECT 264.520 1.060 264.900 14.470 ;
      RECT 265.880 1.060 266.260 53.230 ;
      RECT 267.240 50.510 267.620 53.420 ;
      RECT 272.025 53.230 272.355 53.395 ;
      RECT 267.265 50.345 267.595 50.510 ;
      RECT 267.945 49.150 268.275 49.315 ;
      RECT 267.265 47.110 267.595 47.275 ;
      RECT 267.240 42.840 267.620 47.110 ;
      RECT 267.920 46.240 268.300 49.150 ;
      RECT 266.615 41.830 266.945 42.160 ;
      RECT 266.630 26.515 266.930 41.830 ;
      RECT 266.615 26.185 266.945 26.515 ;
      RECT 269.560 26.185 269.890 26.515 ;
      RECT 269.575 15.410 269.875 26.185 ;
      RECT 269.560 15.080 269.890 15.410 ;
      RECT 269.985 14.470 270.315 14.635 ;
      RECT 269.960 1.060 270.340 14.470 ;
      RECT 271.345 8.350 271.675 8.515 ;
      RECT 271.320 6.120 271.700 8.350 ;
      RECT 272.000 1.060 272.380 53.230 ;
      RECT 273.360 50.510 273.740 53.420 ;
      RECT 278.145 53.230 278.475 53.395 ;
      RECT 273.385 50.345 273.715 50.510 ;
      RECT 273.385 49.150 273.715 49.315 ;
      RECT 272.705 47.110 273.035 47.275 ;
      RECT 272.680 42.840 273.060 47.110 ;
      RECT 273.360 46.240 273.740 49.150 ;
      RECT 272.855 41.830 273.185 42.160 ;
      RECT 272.870 27.735 273.170 41.830 ;
      RECT 272.855 27.405 273.185 27.735 ;
      RECT 275.400 27.405 275.730 27.735 ;
      RECT 275.415 15.410 275.715 27.405 ;
      RECT 275.400 15.080 275.730 15.410 ;
      RECT 276.105 14.470 276.435 14.635 ;
      RECT 276.080 1.060 276.460 14.470 ;
      RECT 278.120 1.060 278.500 53.230 ;
      RECT 279.480 50.510 279.860 53.420 ;
      RECT 284.265 53.230 284.595 53.395 ;
      RECT 279.505 50.345 279.835 50.510 ;
      RECT 280.185 49.150 280.515 49.315 ;
      RECT 279.505 47.110 279.835 47.275 ;
      RECT 279.480 42.840 279.860 47.110 ;
      RECT 280.160 46.240 280.540 49.150 ;
      RECT 283.560 46.430 283.940 49.340 ;
      RECT 283.585 46.265 283.915 46.430 ;
      RECT 279.095 41.830 279.425 42.160 ;
      RECT 279.110 28.955 279.410 41.830 ;
      RECT 279.095 28.625 279.425 28.955 ;
      RECT 281.240 28.625 281.570 28.955 ;
      RECT 281.255 15.410 281.555 28.625 ;
      RECT 281.240 15.080 281.570 15.410 ;
      RECT 282.905 14.470 283.235 14.635 ;
      RECT 279.505 8.350 279.835 8.515 ;
      RECT 279.480 6.120 279.860 8.350 ;
      RECT 282.880 1.060 283.260 14.470 ;
      RECT 284.240 1.060 284.620 53.230 ;
      RECT 286.280 50.510 286.660 53.420 ;
      RECT 289.025 53.230 289.355 53.395 ;
      RECT 286.305 50.345 286.635 50.510 ;
      RECT 285.625 49.150 285.955 49.315 ;
      RECT 284.945 47.110 285.275 47.275 ;
      RECT 284.920 42.840 285.300 47.110 ;
      RECT 285.600 46.240 285.980 49.150 ;
      RECT 285.335 41.830 285.665 42.160 ;
      RECT 285.350 20.415 285.650 41.830 ;
      RECT 285.335 20.085 285.665 20.415 ;
      RECT 287.080 20.085 287.410 20.415 ;
      RECT 287.095 15.410 287.395 20.085 ;
      RECT 287.080 15.080 287.410 15.410 ;
      RECT 288.345 14.470 288.675 14.635 ;
      RECT 287.665 8.350 287.995 8.515 ;
      RECT 287.640 6.120 288.020 8.350 ;
      RECT 288.320 1.060 288.700 14.470 ;
      RECT 289.000 1.060 289.380 53.230 ;
      RECT 292.400 50.510 292.780 53.420 ;
      RECT 295.825 53.230 296.155 53.395 ;
      RECT 296.505 53.230 296.835 53.395 ;
      RECT 292.425 50.345 292.755 50.510 ;
      RECT 295.800 50.320 296.180 53.230 ;
      RECT 292.425 49.150 292.755 49.315 ;
      RECT 291.745 47.110 292.075 47.275 ;
      RECT 291.720 42.840 292.100 47.110 ;
      RECT 292.400 46.240 292.780 49.150 ;
      RECT 291.575 41.830 291.905 42.160 ;
      RECT 290.150 36.230 290.480 36.560 ;
      RECT 290.165 21.635 290.465 36.230 ;
      RECT 291.590 22.855 291.890 41.830 ;
      RECT 291.575 22.525 291.905 22.855 ;
      RECT 290.150 21.305 290.480 21.635 ;
      RECT 292.920 21.305 293.250 21.635 ;
      RECT 292.935 15.410 293.235 21.305 ;
      RECT 292.920 15.080 293.250 15.410 ;
      RECT 295.825 8.350 296.155 8.515 ;
      RECT 295.800 6.120 296.180 8.350 ;
      RECT 296.480 1.060 296.860 53.230 ;
      RECT 298.520 50.510 298.900 53.420 ;
      RECT 302.625 53.230 302.955 53.395 ;
      RECT 298.545 50.345 298.875 50.510 ;
      RECT 298.545 49.150 298.875 49.315 ;
      RECT 297.865 47.110 298.195 47.275 ;
      RECT 297.840 42.840 298.220 47.110 ;
      RECT 298.520 46.240 298.900 49.150 ;
      RECT 297.815 41.830 298.145 42.160 ;
      RECT 297.830 24.075 298.130 41.830 ;
      RECT 297.815 23.745 298.145 24.075 ;
      RECT 302.600 1.060 302.980 53.230 ;
      RECT 304.640 50.510 305.020 53.420 ;
      RECT 308.745 53.230 309.075 53.395 ;
      RECT 309.425 53.230 309.755 53.395 ;
      RECT 304.665 50.345 304.995 50.510 ;
      RECT 308.720 50.320 309.100 53.230 ;
      RECT 304.665 49.150 304.995 49.315 ;
      RECT 303.985 47.110 304.315 47.275 ;
      RECT 303.960 42.840 304.340 47.110 ;
      RECT 304.640 46.240 305.020 49.150 ;
      RECT 304.055 41.830 304.385 42.160 ;
      RECT 304.070 25.295 304.370 41.830 ;
      RECT 304.055 24.965 304.385 25.295 ;
      RECT 304.665 8.350 304.995 8.515 ;
      RECT 304.640 6.120 305.020 8.350 ;
      RECT 309.400 1.060 309.780 53.230 ;
      RECT 310.760 50.510 311.140 53.420 ;
      RECT 314.865 53.230 315.195 53.395 ;
      RECT 315.545 53.230 315.875 53.395 ;
      RECT 310.785 50.345 311.115 50.510 ;
      RECT 314.840 50.320 315.220 53.230 ;
      RECT 311.465 49.150 311.795 49.315 ;
      RECT 310.785 47.110 311.115 47.275 ;
      RECT 310.760 42.840 311.140 47.110 ;
      RECT 311.440 46.240 311.820 49.150 ;
      RECT 310.295 41.830 310.625 42.160 ;
      RECT 310.310 26.515 310.610 41.830 ;
      RECT 310.295 26.185 310.625 26.515 ;
      RECT 313.505 8.350 313.835 8.515 ;
      RECT 313.480 6.120 313.860 8.350 ;
      RECT 315.520 1.060 315.900 53.230 ;
      RECT 317.560 50.510 317.940 53.420 ;
      RECT 321.665 53.230 321.995 53.395 ;
      RECT 317.585 50.345 317.915 50.510 ;
      RECT 317.585 49.150 317.915 49.315 ;
      RECT 316.905 47.110 317.235 47.275 ;
      RECT 316.880 42.840 317.260 47.110 ;
      RECT 317.560 46.240 317.940 49.150 ;
      RECT 316.535 41.830 316.865 42.160 ;
      RECT 316.550 27.735 316.850 41.830 ;
      RECT 316.535 27.405 316.865 27.735 ;
      RECT 320.305 8.350 320.635 8.515 ;
      RECT 320.280 6.120 320.660 8.350 ;
      RECT 321.640 1.060 322.020 53.230 ;
      RECT 323.680 50.510 324.060 53.420 ;
      RECT 327.105 53.230 327.435 53.395 ;
      RECT 327.785 53.230 328.115 53.395 ;
      RECT 323.705 50.345 324.035 50.510 ;
      RECT 327.080 50.320 327.460 53.230 ;
      RECT 323.025 47.110 323.355 47.275 ;
      RECT 323.000 42.840 323.380 47.110 ;
      RECT 323.680 45.070 324.060 49.340 ;
      RECT 323.705 44.905 324.035 45.070 ;
      RECT 322.775 41.830 323.105 42.160 ;
      RECT 322.790 28.955 323.090 41.830 ;
      RECT 322.775 28.625 323.105 28.955 ;
      RECT 327.760 1.060 328.140 53.230 ;
      RECT 329.800 50.510 330.180 53.420 ;
      RECT 333.905 53.230 334.235 53.395 ;
      RECT 329.825 50.345 330.155 50.510 ;
      RECT 329.145 49.150 329.475 49.315 ;
      RECT 328.465 47.110 328.795 47.275 ;
      RECT 328.440 42.840 328.820 47.110 ;
      RECT 329.120 46.240 329.500 49.150 ;
      RECT 329.015 41.830 329.345 42.160 ;
      RECT 329.030 20.415 329.330 41.830 ;
      RECT 329.015 20.085 329.345 20.415 ;
      RECT 329.825 8.350 330.155 8.515 ;
      RECT 329.800 6.120 330.180 8.350 ;
      RECT 333.880 1.060 334.260 53.230 ;
      RECT 335.240 50.510 335.620 53.420 ;
      RECT 335.265 50.345 335.595 50.510 ;
      RECT 412.080 50.320 412.460 64.110 ;
      RECT 415.505 60.030 415.835 60.195 ;
      RECT 335.945 49.150 336.275 49.315 ;
      RECT 335.265 47.110 335.595 47.275 ;
      RECT 335.240 42.840 335.620 47.110 ;
      RECT 335.920 46.240 336.300 49.150 ;
      RECT 340.025 44.390 340.355 44.555 ;
      RECT 339.345 43.030 339.675 43.195 ;
      RECT 335.255 41.830 335.585 42.160 ;
      RECT 335.270 21.635 335.570 41.830 ;
      RECT 339.320 40.800 339.700 43.030 ;
      RECT 340.000 35.360 340.380 44.390 ;
      RECT 412.080 36.910 412.460 50.020 ;
      RECT 412.760 43.710 413.140 57.500 ;
      RECT 413.465 54.590 413.795 54.755 ;
      RECT 412.785 43.545 413.115 43.710 ;
      RECT 412.105 36.745 412.435 36.910 ;
      RECT 335.255 21.305 335.585 21.635 ;
      RECT 338.665 8.350 338.995 8.515 ;
      RECT 346.145 8.350 346.475 8.515 ;
      RECT 354.985 8.350 355.315 8.515 ;
      RECT 363.145 8.350 363.475 8.515 ;
      RECT 371.305 8.350 371.635 8.515 ;
      RECT 380.825 8.350 381.155 8.515 ;
      RECT 388.305 8.350 388.635 8.515 ;
      RECT 397.145 8.350 397.475 8.515 ;
      RECT 405.985 8.350 406.315 8.515 ;
      RECT 412.785 8.350 413.115 8.515 ;
      RECT 338.640 6.120 339.020 8.350 ;
      RECT 346.120 6.120 346.500 8.350 ;
      RECT 354.960 6.120 355.340 8.350 ;
      RECT 363.120 6.120 363.500 8.350 ;
      RECT 371.280 6.120 371.660 8.350 ;
      RECT 380.800 6.120 381.180 8.350 ;
      RECT 388.280 6.120 388.660 8.350 ;
      RECT 397.120 6.120 397.500 8.350 ;
      RECT 405.960 6.120 406.340 8.350 ;
      RECT 412.760 6.120 413.140 8.350 ;
      RECT 413.440 1.060 413.820 54.590 ;
      RECT 414.145 45.750 414.475 45.915 ;
      RECT 414.120 1.060 414.500 45.750 ;
      RECT 414.825 40.310 415.155 40.475 ;
      RECT 414.800 1.060 415.180 40.310 ;
      RECT 415.480 1.060 415.860 60.030 ;
      RECT 422.305 8.350 422.635 8.515 ;
      RECT 431.145 8.350 431.475 8.515 ;
      RECT 438.625 8.350 438.955 8.515 ;
      RECT 447.465 8.350 447.795 8.515 ;
      RECT 455.625 8.350 455.955 8.515 ;
      RECT 463.785 8.350 464.115 8.515 ;
      RECT 422.280 6.120 422.660 8.350 ;
      RECT 431.120 6.120 431.500 8.350 ;
      RECT 438.600 6.120 438.980 8.350 ;
      RECT 447.440 6.120 447.820 8.350 ;
      RECT 455.600 6.120 455.980 8.350 ;
      RECT 463.760 6.120 464.140 8.350 ;
   END
END    sky130_sram_1kbyte_1rw1r_32x256_8
END    LIBRARY
