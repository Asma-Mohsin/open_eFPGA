magic
tech sky130A
magscale 1 2
timestamp 1733306364
<< viali >>
rect 2145 8585 2179 8619
rect 4169 8585 4203 8619
rect 6561 8585 6595 8619
rect 9137 8585 9171 8619
rect 10977 8585 11011 8619
rect 13185 8585 13219 8619
rect 15209 8585 15243 8619
rect 17601 8585 17635 8619
rect 19809 8585 19843 8619
rect 22017 8585 22051 8619
rect 24593 8585 24627 8619
rect 26249 8585 26283 8619
rect 28641 8585 28675 8619
rect 30849 8585 30883 8619
rect 33057 8585 33091 8619
rect 35265 8585 35299 8619
rect 37473 8585 37507 8619
rect 40049 8585 40083 8619
rect 41889 8585 41923 8619
rect 44097 8585 44131 8619
rect 46305 8585 46339 8619
rect 1961 8449 1995 8483
rect 4077 8449 4111 8483
rect 6377 8449 6411 8483
rect 8953 8449 8987 8483
rect 10793 8449 10827 8483
rect 13001 8449 13035 8483
rect 15117 8449 15151 8483
rect 17417 8449 17451 8483
rect 19625 8449 19659 8483
rect 21833 8449 21867 8483
rect 24409 8449 24443 8483
rect 26157 8449 26191 8483
rect 28457 8449 28491 8483
rect 30665 8449 30699 8483
rect 32873 8449 32907 8483
rect 35081 8449 35115 8483
rect 37381 8449 37415 8483
rect 39865 8449 39899 8483
rect 41705 8449 41739 8483
rect 43913 8449 43947 8483
rect 46121 8449 46155 8483
rect 17785 2601 17819 2635
rect 19441 2601 19475 2635
rect 19901 2601 19935 2635
rect 20637 2601 20671 2635
rect 21281 2601 21315 2635
rect 22109 2601 22143 2635
rect 24041 2601 24075 2635
rect 24777 2601 24811 2635
rect 24869 2601 24903 2635
rect 25329 2601 25363 2635
rect 26525 2601 26559 2635
rect 28733 2601 28767 2635
rect 31309 2601 31343 2635
rect 35357 2601 35391 2635
rect 37565 2601 37599 2635
rect 42073 2601 42107 2635
rect 44741 2601 44775 2635
rect 45017 2601 45051 2635
rect 45661 2601 45695 2635
rect 23765 2533 23799 2567
rect 25697 2533 25731 2567
rect 27813 2533 27847 2567
rect 30481 2533 30515 2567
rect 31033 2533 31067 2567
rect 17969 2397 18003 2431
rect 19625 2397 19659 2431
rect 20085 2397 20119 2431
rect 20361 2397 20395 2431
rect 20453 2397 20487 2431
rect 20913 2397 20947 2431
rect 21097 2397 21131 2431
rect 21649 2397 21683 2431
rect 22293 2397 22327 2431
rect 22845 2397 22879 2431
rect 22937 2397 22971 2431
rect 23397 2397 23431 2431
rect 23581 2397 23615 2431
rect 23857 2397 23891 2431
rect 24593 2397 24627 2431
rect 25053 2397 25087 2431
rect 25513 2397 25547 2431
rect 25973 2397 26007 2431
rect 26709 2397 26743 2431
rect 27353 2397 27387 2431
rect 27997 2397 28031 2431
rect 28273 2397 28307 2431
rect 28549 2397 28583 2431
rect 28917 2397 28951 2431
rect 30297 2397 30331 2431
rect 30665 2397 30699 2431
rect 30941 2397 30975 2431
rect 31217 2397 31251 2431
rect 31493 2397 31527 2431
rect 32321 2397 32355 2431
rect 32873 2397 32907 2431
rect 33333 2397 33367 2431
rect 35541 2397 35575 2431
rect 37749 2397 37783 2431
rect 38025 2397 38059 2431
rect 38393 2397 38427 2431
rect 42257 2397 42291 2431
rect 44557 2397 44591 2431
rect 45201 2397 45235 2431
rect 45845 2397 45879 2431
rect 25237 2329 25271 2363
rect 20177 2261 20211 2295
rect 20729 2261 20763 2295
rect 21465 2261 21499 2295
rect 22661 2261 22695 2295
rect 23121 2261 23155 2295
rect 23213 2261 23247 2295
rect 25789 2261 25823 2295
rect 27169 2261 27203 2295
rect 28089 2261 28123 2295
rect 28365 2261 28399 2295
rect 30113 2261 30147 2295
rect 30757 2261 30791 2295
rect 32137 2261 32171 2295
rect 32689 2261 32723 2295
rect 33149 2261 33183 2295
rect 37841 2261 37875 2295
rect 38577 2261 38611 2295
rect 4353 2057 4387 2091
rect 15945 2057 15979 2091
rect 16497 2057 16531 2091
rect 16957 2057 16991 2091
rect 17509 2057 17543 2091
rect 17601 2057 17635 2091
rect 18613 2057 18647 2091
rect 18889 2057 18923 2091
rect 19257 2057 19291 2091
rect 19809 2057 19843 2091
rect 20085 2057 20119 2091
rect 20545 2057 20579 2091
rect 21189 2057 21223 2091
rect 21925 2057 21959 2091
rect 23305 2057 23339 2091
rect 24317 2057 24351 2091
rect 24593 2057 24627 2091
rect 24961 2057 24995 2091
rect 25513 2057 25547 2091
rect 26525 2057 26559 2091
rect 26985 2057 27019 2091
rect 28089 2057 28123 2091
rect 29101 2057 29135 2091
rect 29285 2057 29319 2091
rect 30573 2057 30607 2091
rect 34529 2057 34563 2091
rect 35909 2057 35943 2091
rect 42441 2057 42475 2091
rect 45109 2057 45143 2091
rect 45385 2057 45419 2091
rect 45661 2057 45695 2091
rect 46305 2057 46339 2091
rect 31125 1989 31159 2023
rect 1409 1921 1443 1955
rect 4169 1921 4203 1955
rect 4537 1921 4571 1955
rect 15761 1921 15795 1955
rect 16037 1921 16071 1955
rect 16313 1921 16347 1955
rect 16773 1921 16807 1955
rect 17049 1921 17083 1955
rect 17325 1921 17359 1955
rect 17785 1921 17819 1955
rect 17877 1921 17911 1955
rect 18153 1921 18187 1955
rect 18429 1921 18463 1955
rect 18705 1921 18739 1955
rect 19165 1921 19199 1955
rect 19441 1921 19475 1955
rect 19533 1921 19567 1955
rect 19993 1921 20027 1955
rect 20269 1921 20303 1955
rect 20361 1921 20395 1955
rect 20637 1921 20671 1955
rect 21373 1921 21407 1955
rect 21649 1921 21683 1955
rect 22109 1921 22143 1955
rect 22385 1921 22419 1955
rect 22477 1921 22511 1955
rect 23213 1921 23247 1955
rect 23489 1921 23523 1955
rect 23581 1921 23615 1955
rect 24225 1921 24259 1955
rect 24501 1921 24535 1955
rect 24777 1921 24811 1955
rect 25145 1921 25179 1955
rect 25421 1921 25455 1955
rect 25697 1921 25731 1955
rect 25881 1921 25915 1955
rect 26433 1921 26467 1955
rect 26709 1921 26743 1955
rect 27169 1921 27203 1955
rect 27445 1921 27479 1955
rect 27721 1921 27755 1955
rect 27997 1921 28031 1955
rect 28273 1921 28307 1955
rect 28457 1921 28491 1955
rect 29009 1921 29043 1955
rect 29469 1921 29503 1955
rect 29745 1921 29779 1955
rect 29929 1921 29963 1955
rect 30481 1921 30515 1955
rect 30757 1921 30791 1955
rect 31585 1921 31619 1955
rect 32321 1921 32355 1955
rect 32597 1921 32631 1955
rect 32873 1921 32907 1955
rect 33425 1921 33459 1955
rect 33701 1921 33735 1955
rect 34161 1921 34195 1955
rect 34713 1921 34747 1955
rect 35449 1921 35483 1955
rect 36093 1921 36127 1955
rect 36277 1921 36311 1955
rect 37381 1921 37415 1955
rect 38117 1921 38151 1955
rect 38853 1921 38887 1955
rect 40509 1921 40543 1955
rect 40785 1921 40819 1955
rect 41061 1921 41095 1955
rect 41337 1921 41371 1955
rect 42625 1921 42659 1955
rect 45293 1921 45327 1955
rect 45569 1921 45603 1955
rect 45845 1921 45879 1955
rect 46213 1921 46247 1955
rect 46489 1921 46523 1955
rect 4721 1785 4755 1819
rect 18337 1785 18371 1819
rect 22201 1785 22235 1819
rect 25237 1785 25271 1819
rect 29561 1785 29595 1819
rect 31769 1785 31803 1819
rect 32413 1785 32447 1819
rect 40693 1785 40727 1819
rect 40969 1785 41003 1819
rect 41245 1785 41279 1819
rect 46029 1785 46063 1819
rect 1593 1717 1627 1751
rect 16221 1717 16255 1751
rect 17233 1717 17267 1751
rect 18061 1717 18095 1751
rect 18981 1717 19015 1751
rect 19717 1717 19751 1751
rect 20821 1717 20855 1751
rect 21465 1717 21499 1751
rect 22661 1717 22695 1751
rect 23029 1717 23063 1751
rect 23765 1717 23799 1751
rect 24041 1717 24075 1751
rect 26065 1717 26099 1751
rect 26249 1717 26283 1751
rect 27261 1717 27295 1751
rect 27537 1717 27571 1751
rect 27813 1717 27847 1751
rect 28641 1717 28675 1751
rect 30113 1717 30147 1751
rect 30297 1717 30331 1751
rect 31217 1717 31251 1751
rect 32137 1717 32171 1751
rect 33057 1717 33091 1751
rect 33241 1717 33275 1751
rect 33793 1717 33827 1751
rect 34345 1717 34379 1751
rect 35633 1717 35667 1751
rect 36369 1717 36403 1751
rect 37473 1717 37507 1751
rect 38393 1717 38427 1751
rect 38945 1717 38979 1751
rect 41521 1717 41555 1751
rect 6193 1513 6227 1547
rect 12449 1513 12483 1547
rect 15209 1513 15243 1547
rect 15485 1513 15519 1547
rect 16037 1513 16071 1547
rect 16681 1513 16715 1547
rect 17233 1513 17267 1547
rect 17509 1513 17543 1547
rect 18337 1513 18371 1547
rect 19257 1513 19291 1547
rect 24961 1513 24995 1547
rect 26433 1513 26467 1547
rect 27905 1513 27939 1547
rect 29009 1513 29043 1547
rect 29745 1513 29779 1547
rect 30481 1513 30515 1547
rect 32321 1513 32355 1547
rect 33425 1513 33459 1547
rect 33977 1513 34011 1547
rect 34897 1513 34931 1547
rect 36001 1513 36035 1547
rect 36553 1513 36587 1547
rect 38025 1513 38059 1547
rect 39129 1513 39163 1547
rect 40601 1513 40635 1547
rect 44833 1513 44867 1547
rect 45017 1513 45051 1547
rect 45753 1513 45787 1547
rect 16957 1445 16991 1479
rect 19717 1445 19751 1479
rect 32965 1445 32999 1479
rect 35541 1445 35575 1479
rect 38669 1445 38703 1479
rect 40141 1445 40175 1479
rect 44097 1445 44131 1479
rect 44465 1445 44499 1479
rect 20637 1377 20671 1411
rect 1593 1309 1627 1343
rect 1961 1309 1995 1343
rect 2329 1309 2363 1343
rect 2697 1309 2731 1343
rect 3157 1309 3191 1343
rect 3433 1309 3467 1343
rect 3801 1309 3835 1343
rect 4077 1309 4111 1343
rect 4905 1309 4939 1343
rect 5273 1309 5307 1343
rect 5641 1309 5675 1343
rect 6009 1309 6043 1343
rect 6377 1309 6411 1343
rect 6745 1309 6779 1343
rect 7113 1309 7147 1343
rect 7481 1309 7515 1343
rect 7849 1309 7883 1343
rect 8217 1309 8251 1343
rect 8585 1309 8619 1343
rect 8953 1309 8987 1343
rect 9321 1309 9355 1343
rect 9689 1309 9723 1343
rect 10057 1309 10091 1343
rect 10425 1309 10459 1343
rect 10793 1309 10827 1343
rect 11161 1309 11195 1343
rect 11529 1309 11563 1343
rect 11897 1309 11931 1343
rect 12265 1309 12299 1343
rect 12633 1309 12667 1343
rect 13001 1309 13035 1343
rect 13369 1309 13403 1343
rect 13737 1309 13771 1343
rect 14105 1309 14139 1343
rect 14657 1309 14691 1343
rect 15025 1309 15059 1343
rect 15393 1309 15427 1343
rect 15669 1309 15703 1343
rect 15945 1309 15979 1343
rect 16221 1309 16255 1343
rect 16497 1309 16531 1343
rect 16865 1309 16899 1343
rect 17141 1309 17175 1343
rect 17417 1309 17451 1343
rect 17693 1309 17727 1343
rect 17969 1309 18003 1343
rect 18245 1309 18279 1343
rect 18521 1309 18555 1343
rect 18797 1309 18831 1343
rect 18889 1309 18923 1343
rect 19441 1309 19475 1343
rect 19533 1309 19567 1343
rect 19901 1309 19935 1343
rect 21005 1309 21039 1343
rect 21373 1309 21407 1343
rect 22017 1309 22051 1343
rect 22201 1309 22235 1343
rect 22569 1309 22603 1343
rect 22845 1309 22879 1343
rect 23949 1309 23983 1343
rect 24409 1309 24443 1343
rect 25329 1309 25363 1343
rect 25697 1309 25731 1343
rect 26341 1309 26375 1343
rect 26985 1309 27019 1343
rect 27353 1309 27387 1343
rect 27813 1309 27847 1343
rect 28273 1309 28307 1343
rect 29653 1309 29687 1343
rect 30941 1309 30975 1343
rect 31309 1309 31343 1343
rect 31493 1309 31527 1343
rect 32781 1309 32815 1343
rect 33333 1309 33367 1343
rect 35357 1309 35391 1343
rect 38485 1309 38519 1343
rect 39037 1309 39071 1343
rect 39497 1309 39531 1343
rect 40969 1309 41003 1343
rect 41429 1309 41463 1343
rect 41705 1309 41739 1343
rect 42441 1309 42475 1343
rect 42717 1309 42751 1343
rect 42993 1309 43027 1343
rect 43269 1309 43303 1343
rect 43545 1309 43579 1343
rect 43913 1309 43947 1343
rect 44281 1309 44315 1343
rect 44649 1309 44683 1343
rect 45201 1309 45235 1343
rect 45569 1309 45603 1343
rect 45937 1309 45971 1343
rect 46305 1309 46339 1343
rect 20361 1241 20395 1275
rect 23305 1241 23339 1275
rect 24869 1241 24903 1275
rect 28917 1241 28951 1275
rect 30389 1241 30423 1275
rect 32229 1241 32263 1275
rect 33885 1241 33919 1275
rect 34805 1241 34839 1275
rect 35909 1241 35943 1275
rect 36461 1241 36495 1275
rect 37933 1241 37967 1275
rect 39957 1241 39991 1275
rect 40509 1241 40543 1275
rect 1777 1173 1811 1207
rect 2145 1173 2179 1207
rect 2513 1173 2547 1207
rect 2881 1173 2915 1207
rect 3341 1173 3375 1207
rect 3617 1173 3651 1207
rect 5089 1173 5123 1207
rect 5457 1173 5491 1207
rect 5825 1173 5859 1207
rect 6561 1173 6595 1207
rect 6929 1173 6963 1207
rect 7297 1173 7331 1207
rect 7665 1173 7699 1207
rect 8033 1173 8067 1207
rect 8401 1173 8435 1207
rect 8769 1173 8803 1207
rect 9137 1173 9171 1207
rect 9505 1173 9539 1207
rect 9873 1173 9907 1207
rect 10241 1173 10275 1207
rect 10609 1173 10643 1207
rect 10977 1173 11011 1207
rect 11345 1173 11379 1207
rect 11713 1173 11747 1207
rect 12081 1173 12115 1207
rect 12817 1173 12851 1207
rect 13185 1173 13219 1207
rect 13553 1173 13587 1207
rect 13921 1173 13955 1207
rect 14289 1173 14323 1207
rect 14473 1173 14507 1207
rect 14841 1173 14875 1207
rect 15761 1173 15795 1207
rect 16313 1173 16347 1207
rect 17785 1173 17819 1207
rect 18061 1173 18095 1207
rect 18613 1173 18647 1207
rect 19073 1173 19107 1207
rect 20085 1173 20119 1207
rect 21189 1173 21223 1207
rect 21557 1173 21591 1207
rect 21833 1173 21867 1207
rect 23029 1173 23063 1207
rect 23397 1173 23431 1207
rect 24133 1173 24167 1207
rect 24593 1173 24627 1207
rect 25513 1173 25547 1207
rect 25881 1173 25915 1207
rect 27169 1173 27203 1207
rect 27537 1173 27571 1207
rect 28457 1173 28491 1207
rect 31585 1173 31619 1207
rect 37473 1173 37507 1207
rect 39681 1173 39715 1207
rect 41153 1173 41187 1207
rect 42625 1173 42659 1207
rect 42901 1173 42935 1207
rect 43177 1173 43211 1207
rect 43453 1173 43487 1207
rect 43729 1173 43763 1207
rect 45385 1173 45419 1207
rect 46121 1173 46155 1207
<< metal1 >>
rect 23474 9024 23480 9036
rect 6380 8996 23480 9024
rect 6380 8832 6408 8996
rect 23474 8984 23480 8996
rect 23532 8984 23538 9036
rect 12986 8916 12992 8968
rect 13044 8956 13050 8968
rect 22186 8956 22192 8968
rect 13044 8928 22192 8956
rect 13044 8916 13050 8928
rect 22186 8916 22192 8928
rect 22244 8916 22250 8968
rect 25314 8888 25320 8900
rect 6472 8860 25320 8888
rect 6472 8832 6500 8860
rect 25314 8848 25320 8860
rect 25372 8848 25378 8900
rect 6362 8780 6368 8832
rect 6420 8780 6426 8832
rect 6454 8780 6460 8832
rect 6512 8780 6518 8832
rect 6546 8780 6552 8832
rect 6604 8820 6610 8832
rect 29178 8820 29184 8832
rect 6604 8792 29184 8820
rect 6604 8780 6610 8792
rect 29178 8780 29184 8792
rect 29236 8780 29242 8832
rect 1104 8730 46984 8752
rect 1104 8678 12380 8730
rect 12432 8678 12444 8730
rect 12496 8678 12508 8730
rect 12560 8678 12572 8730
rect 12624 8678 12636 8730
rect 12688 8678 23810 8730
rect 23862 8678 23874 8730
rect 23926 8678 23938 8730
rect 23990 8678 24002 8730
rect 24054 8678 24066 8730
rect 24118 8678 35240 8730
rect 35292 8678 35304 8730
rect 35356 8678 35368 8730
rect 35420 8678 35432 8730
rect 35484 8678 35496 8730
rect 35548 8678 46670 8730
rect 46722 8678 46734 8730
rect 46786 8678 46798 8730
rect 46850 8678 46862 8730
rect 46914 8678 46926 8730
rect 46978 8678 46984 8730
rect 1104 8656 46984 8678
rect 1854 8576 1860 8628
rect 1912 8616 1918 8628
rect 2133 8619 2191 8625
rect 2133 8616 2145 8619
rect 1912 8588 2145 8616
rect 1912 8576 1918 8588
rect 2133 8585 2145 8588
rect 2179 8585 2191 8619
rect 2133 8579 2191 8585
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 4157 8619 4215 8625
rect 4157 8616 4169 8619
rect 4120 8588 4169 8616
rect 4120 8576 4126 8588
rect 4157 8585 4169 8588
rect 4203 8585 4215 8619
rect 4157 8579 4215 8585
rect 6270 8576 6276 8628
rect 6328 8616 6334 8628
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 6328 8588 6561 8616
rect 6328 8576 6334 8588
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 6549 8579 6607 8585
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 9125 8619 9183 8625
rect 9125 8616 9137 8619
rect 8536 8588 9137 8616
rect 8536 8576 8542 8588
rect 9125 8585 9137 8588
rect 9171 8585 9183 8619
rect 9125 8579 9183 8585
rect 10686 8576 10692 8628
rect 10744 8616 10750 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10744 8588 10977 8616
rect 10744 8576 10750 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 10965 8579 11023 8585
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 13173 8619 13231 8625
rect 13173 8616 13185 8619
rect 12952 8588 13185 8616
rect 12952 8576 12958 8588
rect 13173 8585 13185 8588
rect 13219 8585 13231 8619
rect 13173 8579 13231 8585
rect 15102 8576 15108 8628
rect 15160 8616 15166 8628
rect 15197 8619 15255 8625
rect 15197 8616 15209 8619
rect 15160 8588 15209 8616
rect 15160 8576 15166 8588
rect 15197 8585 15209 8588
rect 15243 8585 15255 8619
rect 15197 8579 15255 8585
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 17589 8619 17647 8625
rect 17589 8616 17601 8619
rect 17368 8588 17601 8616
rect 17368 8576 17374 8588
rect 17589 8585 17601 8588
rect 17635 8585 17647 8619
rect 17589 8579 17647 8585
rect 19518 8576 19524 8628
rect 19576 8616 19582 8628
rect 19797 8619 19855 8625
rect 19797 8616 19809 8619
rect 19576 8588 19809 8616
rect 19576 8576 19582 8588
rect 19797 8585 19809 8588
rect 19843 8585 19855 8619
rect 19797 8579 19855 8585
rect 21726 8576 21732 8628
rect 21784 8616 21790 8628
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 21784 8588 22017 8616
rect 21784 8576 21790 8588
rect 22005 8585 22017 8588
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 24210 8576 24216 8628
rect 24268 8616 24274 8628
rect 24581 8619 24639 8625
rect 24581 8616 24593 8619
rect 24268 8588 24593 8616
rect 24268 8576 24274 8588
rect 24581 8585 24593 8588
rect 24627 8585 24639 8619
rect 24581 8579 24639 8585
rect 26142 8576 26148 8628
rect 26200 8616 26206 8628
rect 26237 8619 26295 8625
rect 26237 8616 26249 8619
rect 26200 8588 26249 8616
rect 26200 8576 26206 8588
rect 26237 8585 26249 8588
rect 26283 8585 26295 8619
rect 26237 8579 26295 8585
rect 28350 8576 28356 8628
rect 28408 8616 28414 8628
rect 28629 8619 28687 8625
rect 28629 8616 28641 8619
rect 28408 8588 28641 8616
rect 28408 8576 28414 8588
rect 28629 8585 28641 8588
rect 28675 8585 28687 8619
rect 28629 8579 28687 8585
rect 30558 8576 30564 8628
rect 30616 8616 30622 8628
rect 30837 8619 30895 8625
rect 30837 8616 30849 8619
rect 30616 8588 30849 8616
rect 30616 8576 30622 8588
rect 30837 8585 30849 8588
rect 30883 8585 30895 8619
rect 30837 8579 30895 8585
rect 32766 8576 32772 8628
rect 32824 8616 32830 8628
rect 33045 8619 33103 8625
rect 33045 8616 33057 8619
rect 32824 8588 33057 8616
rect 32824 8576 32830 8588
rect 33045 8585 33057 8588
rect 33091 8585 33103 8619
rect 33045 8579 33103 8585
rect 34974 8576 34980 8628
rect 35032 8616 35038 8628
rect 35253 8619 35311 8625
rect 35253 8616 35265 8619
rect 35032 8588 35265 8616
rect 35032 8576 35038 8588
rect 35253 8585 35265 8588
rect 35299 8585 35311 8619
rect 35253 8579 35311 8585
rect 37182 8576 37188 8628
rect 37240 8616 37246 8628
rect 37461 8619 37519 8625
rect 37461 8616 37473 8619
rect 37240 8588 37473 8616
rect 37240 8576 37246 8588
rect 37461 8585 37473 8588
rect 37507 8585 37519 8619
rect 37461 8579 37519 8585
rect 39390 8576 39396 8628
rect 39448 8616 39454 8628
rect 40037 8619 40095 8625
rect 40037 8616 40049 8619
rect 39448 8588 40049 8616
rect 39448 8576 39454 8588
rect 40037 8585 40049 8588
rect 40083 8585 40095 8619
rect 40037 8579 40095 8585
rect 41598 8576 41604 8628
rect 41656 8616 41662 8628
rect 41877 8619 41935 8625
rect 41877 8616 41889 8619
rect 41656 8588 41889 8616
rect 41656 8576 41662 8588
rect 41877 8585 41889 8588
rect 41923 8585 41935 8619
rect 41877 8579 41935 8585
rect 43806 8576 43812 8628
rect 43864 8616 43870 8628
rect 44085 8619 44143 8625
rect 44085 8616 44097 8619
rect 43864 8588 44097 8616
rect 43864 8576 43870 8588
rect 44085 8585 44097 8588
rect 44131 8585 44143 8619
rect 44085 8579 44143 8585
rect 46014 8576 46020 8628
rect 46072 8616 46078 8628
rect 46293 8619 46351 8625
rect 46293 8616 46305 8619
rect 46072 8588 46305 8616
rect 46072 8576 46078 8588
rect 46293 8585 46305 8588
rect 46339 8585 46351 8619
rect 46293 8579 46351 8585
rect 6454 8548 6460 8560
rect 4080 8520 6460 8548
rect 4080 8489 4108 8520
rect 6454 8508 6460 8520
rect 6512 8508 6518 8560
rect 24302 8548 24308 8560
rect 8956 8520 24308 8548
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 1964 8412 1992 8443
rect 6362 8440 6368 8492
rect 6420 8440 6426 8492
rect 8956 8489 8984 8520
rect 24302 8508 24308 8520
rect 24360 8508 24366 8560
rect 8941 8483 8999 8489
rect 8941 8449 8953 8483
rect 8987 8449 8999 8483
rect 8941 8443 8999 8449
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 6546 8412 6552 8424
rect 1964 8384 6552 8412
rect 6546 8372 6552 8384
rect 6604 8372 6610 8424
rect 10796 8344 10824 8443
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 15105 8483 15163 8489
rect 15105 8449 15117 8483
rect 15151 8480 15163 8483
rect 15151 8452 16574 8480
rect 15151 8449 15163 8452
rect 15105 8443 15163 8449
rect 16546 8412 16574 8452
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 19610 8440 19616 8492
rect 19668 8440 19674 8492
rect 21821 8483 21879 8489
rect 21821 8449 21833 8483
rect 21867 8480 21879 8483
rect 22094 8480 22100 8492
rect 21867 8452 22100 8480
rect 21867 8449 21879 8452
rect 21821 8443 21879 8449
rect 22094 8440 22100 8452
rect 22152 8440 22158 8492
rect 24397 8483 24455 8489
rect 24397 8449 24409 8483
rect 24443 8480 24455 8483
rect 24854 8480 24860 8492
rect 24443 8452 24860 8480
rect 24443 8449 24455 8452
rect 24397 8443 24455 8449
rect 24854 8440 24860 8452
rect 24912 8440 24918 8492
rect 26145 8483 26203 8489
rect 26145 8449 26157 8483
rect 26191 8480 26203 8483
rect 26510 8480 26516 8492
rect 26191 8452 26516 8480
rect 26191 8449 26203 8452
rect 26145 8443 26203 8449
rect 26510 8440 26516 8452
rect 26568 8440 26574 8492
rect 28442 8440 28448 8492
rect 28500 8440 28506 8492
rect 30650 8440 30656 8492
rect 30708 8440 30714 8492
rect 32861 8483 32919 8489
rect 32861 8449 32873 8483
rect 32907 8480 32919 8483
rect 33134 8480 33140 8492
rect 32907 8452 33140 8480
rect 32907 8449 32919 8452
rect 32861 8443 32919 8449
rect 33134 8440 33140 8452
rect 33192 8440 33198 8492
rect 35066 8440 35072 8492
rect 35124 8440 35130 8492
rect 37366 8440 37372 8492
rect 37424 8440 37430 8492
rect 39853 8483 39911 8489
rect 39853 8449 39865 8483
rect 39899 8449 39911 8483
rect 39853 8443 39911 8449
rect 21266 8412 21272 8424
rect 16546 8384 21272 8412
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 39868 8412 39896 8443
rect 41690 8440 41696 8492
rect 41748 8440 41754 8492
rect 43901 8483 43959 8489
rect 43901 8449 43913 8483
rect 43947 8480 43959 8483
rect 45002 8480 45008 8492
rect 43947 8452 45008 8480
rect 43947 8449 43959 8452
rect 43901 8443 43959 8449
rect 45002 8440 45008 8452
rect 45060 8440 45066 8492
rect 46106 8440 46112 8492
rect 46164 8440 46170 8492
rect 44726 8412 44732 8424
rect 39868 8384 44732 8412
rect 44726 8372 44732 8384
rect 44784 8372 44790 8424
rect 24670 8344 24676 8356
rect 10796 8316 24676 8344
rect 24670 8304 24676 8316
rect 24728 8304 24734 8356
rect 1104 8186 46828 8208
rect 1104 8134 6665 8186
rect 6717 8134 6729 8186
rect 6781 8134 6793 8186
rect 6845 8134 6857 8186
rect 6909 8134 6921 8186
rect 6973 8134 18095 8186
rect 18147 8134 18159 8186
rect 18211 8134 18223 8186
rect 18275 8134 18287 8186
rect 18339 8134 18351 8186
rect 18403 8134 29525 8186
rect 29577 8134 29589 8186
rect 29641 8134 29653 8186
rect 29705 8134 29717 8186
rect 29769 8134 29781 8186
rect 29833 8134 40955 8186
rect 41007 8134 41019 8186
rect 41071 8134 41083 8186
rect 41135 8134 41147 8186
rect 41199 8134 41211 8186
rect 41263 8134 46828 8186
rect 1104 8112 46828 8134
rect 1104 7642 46984 7664
rect 1104 7590 12380 7642
rect 12432 7590 12444 7642
rect 12496 7590 12508 7642
rect 12560 7590 12572 7642
rect 12624 7590 12636 7642
rect 12688 7590 23810 7642
rect 23862 7590 23874 7642
rect 23926 7590 23938 7642
rect 23990 7590 24002 7642
rect 24054 7590 24066 7642
rect 24118 7590 35240 7642
rect 35292 7590 35304 7642
rect 35356 7590 35368 7642
rect 35420 7590 35432 7642
rect 35484 7590 35496 7642
rect 35548 7590 46670 7642
rect 46722 7590 46734 7642
rect 46786 7590 46798 7642
rect 46850 7590 46862 7642
rect 46914 7590 46926 7642
rect 46978 7590 46984 7642
rect 1104 7568 46984 7590
rect 1104 7098 46828 7120
rect 1104 7046 6665 7098
rect 6717 7046 6729 7098
rect 6781 7046 6793 7098
rect 6845 7046 6857 7098
rect 6909 7046 6921 7098
rect 6973 7046 18095 7098
rect 18147 7046 18159 7098
rect 18211 7046 18223 7098
rect 18275 7046 18287 7098
rect 18339 7046 18351 7098
rect 18403 7046 29525 7098
rect 29577 7046 29589 7098
rect 29641 7046 29653 7098
rect 29705 7046 29717 7098
rect 29769 7046 29781 7098
rect 29833 7046 40955 7098
rect 41007 7046 41019 7098
rect 41071 7046 41083 7098
rect 41135 7046 41147 7098
rect 41199 7046 41211 7098
rect 41263 7046 46828 7098
rect 1104 7024 46828 7046
rect 1104 6554 46984 6576
rect 1104 6502 12380 6554
rect 12432 6502 12444 6554
rect 12496 6502 12508 6554
rect 12560 6502 12572 6554
rect 12624 6502 12636 6554
rect 12688 6502 23810 6554
rect 23862 6502 23874 6554
rect 23926 6502 23938 6554
rect 23990 6502 24002 6554
rect 24054 6502 24066 6554
rect 24118 6502 35240 6554
rect 35292 6502 35304 6554
rect 35356 6502 35368 6554
rect 35420 6502 35432 6554
rect 35484 6502 35496 6554
rect 35548 6502 46670 6554
rect 46722 6502 46734 6554
rect 46786 6502 46798 6554
rect 46850 6502 46862 6554
rect 46914 6502 46926 6554
rect 46978 6502 46984 6554
rect 1104 6480 46984 6502
rect 1104 6010 46828 6032
rect 1104 5958 6665 6010
rect 6717 5958 6729 6010
rect 6781 5958 6793 6010
rect 6845 5958 6857 6010
rect 6909 5958 6921 6010
rect 6973 5958 18095 6010
rect 18147 5958 18159 6010
rect 18211 5958 18223 6010
rect 18275 5958 18287 6010
rect 18339 5958 18351 6010
rect 18403 5958 29525 6010
rect 29577 5958 29589 6010
rect 29641 5958 29653 6010
rect 29705 5958 29717 6010
rect 29769 5958 29781 6010
rect 29833 5958 40955 6010
rect 41007 5958 41019 6010
rect 41071 5958 41083 6010
rect 41135 5958 41147 6010
rect 41199 5958 41211 6010
rect 41263 5958 46828 6010
rect 1104 5936 46828 5958
rect 1104 5466 46984 5488
rect 1104 5414 12380 5466
rect 12432 5414 12444 5466
rect 12496 5414 12508 5466
rect 12560 5414 12572 5466
rect 12624 5414 12636 5466
rect 12688 5414 23810 5466
rect 23862 5414 23874 5466
rect 23926 5414 23938 5466
rect 23990 5414 24002 5466
rect 24054 5414 24066 5466
rect 24118 5414 35240 5466
rect 35292 5414 35304 5466
rect 35356 5414 35368 5466
rect 35420 5414 35432 5466
rect 35484 5414 35496 5466
rect 35548 5414 46670 5466
rect 46722 5414 46734 5466
rect 46786 5414 46798 5466
rect 46850 5414 46862 5466
rect 46914 5414 46926 5466
rect 46978 5414 46984 5466
rect 1104 5392 46984 5414
rect 1104 4922 46828 4944
rect 1104 4870 6665 4922
rect 6717 4870 6729 4922
rect 6781 4870 6793 4922
rect 6845 4870 6857 4922
rect 6909 4870 6921 4922
rect 6973 4870 18095 4922
rect 18147 4870 18159 4922
rect 18211 4870 18223 4922
rect 18275 4870 18287 4922
rect 18339 4870 18351 4922
rect 18403 4870 29525 4922
rect 29577 4870 29589 4922
rect 29641 4870 29653 4922
rect 29705 4870 29717 4922
rect 29769 4870 29781 4922
rect 29833 4870 40955 4922
rect 41007 4870 41019 4922
rect 41071 4870 41083 4922
rect 41135 4870 41147 4922
rect 41199 4870 41211 4922
rect 41263 4870 46828 4922
rect 1104 4848 46828 4870
rect 7006 4496 7012 4548
rect 7064 4536 7070 4548
rect 26418 4536 26424 4548
rect 7064 4508 26424 4536
rect 7064 4496 7070 4508
rect 26418 4496 26424 4508
rect 26476 4496 26482 4548
rect 16942 4428 16948 4480
rect 17000 4468 17006 4480
rect 38102 4468 38108 4480
rect 17000 4440 38108 4468
rect 17000 4428 17006 4440
rect 38102 4428 38108 4440
rect 38160 4428 38166 4480
rect 1104 4378 46984 4400
rect 1104 4326 12380 4378
rect 12432 4326 12444 4378
rect 12496 4326 12508 4378
rect 12560 4326 12572 4378
rect 12624 4326 12636 4378
rect 12688 4326 23810 4378
rect 23862 4326 23874 4378
rect 23926 4326 23938 4378
rect 23990 4326 24002 4378
rect 24054 4326 24066 4378
rect 24118 4326 35240 4378
rect 35292 4326 35304 4378
rect 35356 4326 35368 4378
rect 35420 4326 35432 4378
rect 35484 4326 35496 4378
rect 35548 4326 46670 4378
rect 46722 4326 46734 4378
rect 46786 4326 46798 4378
rect 46850 4326 46862 4378
rect 46914 4326 46926 4378
rect 46978 4326 46984 4378
rect 1104 4304 46984 4326
rect 3970 4224 3976 4276
rect 4028 4264 4034 4276
rect 27430 4264 27436 4276
rect 4028 4236 27436 4264
rect 4028 4224 4034 4236
rect 27430 4224 27436 4236
rect 27488 4224 27494 4276
rect 2866 4156 2872 4208
rect 2924 4196 2930 4208
rect 27706 4196 27712 4208
rect 2924 4168 27712 4196
rect 2924 4156 2930 4168
rect 27706 4156 27712 4168
rect 27764 4156 27770 4208
rect 1104 3834 46828 3856
rect 1104 3782 6665 3834
rect 6717 3782 6729 3834
rect 6781 3782 6793 3834
rect 6845 3782 6857 3834
rect 6909 3782 6921 3834
rect 6973 3782 18095 3834
rect 18147 3782 18159 3834
rect 18211 3782 18223 3834
rect 18275 3782 18287 3834
rect 18339 3782 18351 3834
rect 18403 3782 29525 3834
rect 29577 3782 29589 3834
rect 29641 3782 29653 3834
rect 29705 3782 29717 3834
rect 29769 3782 29781 3834
rect 29833 3782 40955 3834
rect 41007 3782 41019 3834
rect 41071 3782 41083 3834
rect 41135 3782 41147 3834
rect 41199 3782 41211 3834
rect 41263 3782 46828 3834
rect 1104 3760 46828 3782
rect 13446 3476 13452 3528
rect 13504 3516 13510 3528
rect 21726 3516 21732 3528
rect 13504 3488 21732 3516
rect 13504 3476 13510 3488
rect 21726 3476 21732 3488
rect 21784 3476 21790 3528
rect 12710 3408 12716 3460
rect 12768 3448 12774 3460
rect 29362 3448 29368 3460
rect 12768 3420 29368 3448
rect 12768 3408 12774 3420
rect 29362 3408 29368 3420
rect 29420 3408 29426 3460
rect 15194 3340 15200 3392
rect 15252 3380 15258 3392
rect 25222 3380 25228 3392
rect 15252 3352 25228 3380
rect 15252 3340 15258 3352
rect 25222 3340 25228 3352
rect 25280 3340 25286 3392
rect 1104 3290 46984 3312
rect 1104 3238 12380 3290
rect 12432 3238 12444 3290
rect 12496 3238 12508 3290
rect 12560 3238 12572 3290
rect 12624 3238 12636 3290
rect 12688 3238 23810 3290
rect 23862 3238 23874 3290
rect 23926 3238 23938 3290
rect 23990 3238 24002 3290
rect 24054 3238 24066 3290
rect 24118 3238 35240 3290
rect 35292 3238 35304 3290
rect 35356 3238 35368 3290
rect 35420 3238 35432 3290
rect 35484 3238 35496 3290
rect 35548 3238 46670 3290
rect 46722 3238 46734 3290
rect 46786 3238 46798 3290
rect 46850 3238 46862 3290
rect 46914 3238 46926 3290
rect 46978 3238 46984 3290
rect 1104 3216 46984 3238
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 28166 3176 28172 3188
rect 8812 3148 28172 3176
rect 8812 3136 8818 3148
rect 28166 3136 28172 3148
rect 28224 3136 28230 3188
rect 5534 3068 5540 3120
rect 5592 3108 5598 3120
rect 19978 3108 19984 3120
rect 5592 3080 19984 3108
rect 5592 3068 5598 3080
rect 19978 3068 19984 3080
rect 20036 3068 20042 3120
rect 21634 3068 21640 3120
rect 21692 3108 21698 3120
rect 31110 3108 31116 3120
rect 21692 3080 31116 3108
rect 21692 3068 21698 3080
rect 31110 3068 31116 3080
rect 31168 3068 31174 3120
rect 17494 3000 17500 3052
rect 17552 3040 17558 3052
rect 33962 3040 33968 3052
rect 17552 3012 33968 3040
rect 17552 3000 17558 3012
rect 33962 3000 33968 3012
rect 34020 3000 34026 3052
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 20070 2972 20076 2984
rect 19392 2944 20076 2972
rect 19392 2932 19398 2944
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 5718 2864 5724 2916
rect 5776 2904 5782 2916
rect 20346 2904 20352 2916
rect 5776 2876 20352 2904
rect 5776 2864 5782 2876
rect 20346 2864 20352 2876
rect 20404 2864 20410 2916
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 37826 2904 37832 2916
rect 20680 2876 37832 2904
rect 20680 2864 20686 2876
rect 37826 2864 37832 2876
rect 37884 2864 37890 2916
rect 9582 2796 9588 2848
rect 9640 2836 9646 2848
rect 9674 2836 9680 2848
rect 9640 2808 9680 2836
rect 9640 2796 9646 2808
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 17126 2796 17132 2848
rect 17184 2836 17190 2848
rect 24762 2836 24768 2848
rect 17184 2808 24768 2836
rect 17184 2796 17190 2808
rect 24762 2796 24768 2808
rect 24820 2796 24826 2848
rect 32122 2796 32128 2848
rect 32180 2836 32186 2848
rect 38562 2836 38568 2848
rect 32180 2808 38568 2836
rect 32180 2796 32186 2808
rect 38562 2796 38568 2808
rect 38620 2796 38626 2848
rect 1104 2746 46828 2768
rect 1104 2694 6665 2746
rect 6717 2694 6729 2746
rect 6781 2694 6793 2746
rect 6845 2694 6857 2746
rect 6909 2694 6921 2746
rect 6973 2694 18095 2746
rect 18147 2694 18159 2746
rect 18211 2694 18223 2746
rect 18275 2694 18287 2746
rect 18339 2694 18351 2746
rect 18403 2694 29525 2746
rect 29577 2694 29589 2746
rect 29641 2694 29653 2746
rect 29705 2694 29717 2746
rect 29769 2694 29781 2746
rect 29833 2694 40955 2746
rect 41007 2694 41019 2746
rect 41071 2694 41083 2746
rect 41135 2694 41147 2746
rect 41199 2694 41211 2746
rect 41263 2694 46828 2746
rect 1104 2672 46828 2694
rect 17402 2592 17408 2644
rect 17460 2632 17466 2644
rect 17773 2635 17831 2641
rect 17773 2632 17785 2635
rect 17460 2604 17785 2632
rect 17460 2592 17466 2604
rect 17773 2601 17785 2604
rect 17819 2601 17831 2635
rect 17773 2595 17831 2601
rect 19429 2635 19487 2641
rect 19429 2601 19441 2635
rect 19475 2632 19487 2635
rect 19518 2632 19524 2644
rect 19475 2604 19524 2632
rect 19475 2601 19487 2604
rect 19429 2595 19487 2601
rect 19518 2592 19524 2604
rect 19576 2592 19582 2644
rect 19610 2592 19616 2644
rect 19668 2632 19674 2644
rect 19889 2635 19947 2641
rect 19889 2632 19901 2635
rect 19668 2604 19901 2632
rect 19668 2592 19674 2604
rect 19889 2601 19901 2604
rect 19935 2601 19947 2635
rect 19889 2595 19947 2601
rect 19996 2604 20576 2632
rect 8202 2524 8208 2576
rect 8260 2564 8266 2576
rect 19996 2564 20024 2604
rect 8260 2536 20024 2564
rect 20548 2564 20576 2604
rect 20622 2592 20628 2644
rect 20680 2592 20686 2644
rect 21266 2592 21272 2644
rect 21324 2592 21330 2644
rect 22094 2592 22100 2644
rect 22152 2592 22158 2644
rect 22186 2592 22192 2644
rect 22244 2592 22250 2644
rect 23474 2592 23480 2644
rect 23532 2632 23538 2644
rect 24029 2635 24087 2641
rect 24029 2632 24041 2635
rect 23532 2604 24041 2632
rect 23532 2592 23538 2604
rect 24029 2601 24041 2604
rect 24075 2601 24087 2635
rect 24029 2595 24087 2601
rect 24302 2592 24308 2644
rect 24360 2632 24366 2644
rect 24765 2635 24823 2641
rect 24765 2632 24777 2635
rect 24360 2604 24777 2632
rect 24360 2592 24366 2604
rect 24765 2601 24777 2604
rect 24811 2601 24823 2635
rect 24765 2595 24823 2601
rect 24854 2592 24860 2644
rect 24912 2592 24918 2644
rect 25314 2592 25320 2644
rect 25372 2592 25378 2644
rect 26510 2592 26516 2644
rect 26568 2592 26574 2644
rect 26620 2604 28120 2632
rect 21542 2564 21548 2576
rect 20548 2536 21548 2564
rect 8260 2524 8266 2536
rect 21542 2524 21548 2536
rect 21600 2524 21606 2576
rect 22204 2564 22232 2592
rect 23753 2567 23811 2573
rect 23753 2564 23765 2567
rect 22204 2536 23765 2564
rect 23753 2533 23765 2536
rect 23799 2533 23811 2567
rect 23753 2527 23811 2533
rect 24670 2524 24676 2576
rect 24728 2564 24734 2576
rect 25685 2567 25743 2573
rect 25685 2564 25697 2567
rect 24728 2536 25697 2564
rect 24728 2524 24734 2536
rect 25685 2533 25697 2536
rect 25731 2533 25743 2567
rect 25685 2527 25743 2533
rect 15378 2456 15384 2508
rect 15436 2496 15442 2508
rect 15436 2468 20484 2496
rect 15436 2456 15442 2468
rect 17954 2388 17960 2440
rect 18012 2388 18018 2440
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2424 19671 2431
rect 19978 2428 19984 2440
rect 19720 2424 19984 2428
rect 19659 2400 19984 2424
rect 19659 2397 19748 2400
rect 19613 2396 19748 2397
rect 19613 2391 19671 2396
rect 19978 2388 19984 2400
rect 20036 2388 20042 2440
rect 20070 2388 20076 2440
rect 20128 2388 20134 2440
rect 20346 2388 20352 2440
rect 20404 2388 20410 2440
rect 20456 2437 20484 2468
rect 20622 2456 20628 2508
rect 20680 2496 20686 2508
rect 26620 2496 26648 2604
rect 27801 2567 27859 2573
rect 27801 2533 27813 2567
rect 27847 2533 27859 2567
rect 27801 2527 27859 2533
rect 27816 2496 27844 2527
rect 20680 2468 22968 2496
rect 20680 2456 20686 2468
rect 20441 2431 20499 2437
rect 20441 2397 20453 2431
rect 20487 2397 20499 2431
rect 20441 2391 20499 2397
rect 20901 2431 20959 2437
rect 20901 2397 20913 2431
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 21085 2431 21143 2437
rect 21085 2397 21097 2431
rect 21131 2428 21143 2431
rect 21131 2400 21496 2428
rect 21131 2397 21143 2400
rect 21085 2391 21143 2397
rect 15102 2320 15108 2372
rect 15160 2360 15166 2372
rect 19886 2360 19892 2372
rect 15160 2332 19892 2360
rect 15160 2320 15166 2332
rect 19886 2320 19892 2332
rect 19944 2320 19950 2372
rect 20916 2360 20944 2391
rect 19996 2332 20944 2360
rect 13630 2252 13636 2304
rect 13688 2292 13694 2304
rect 19996 2292 20024 2332
rect 13688 2264 20024 2292
rect 20165 2295 20223 2301
rect 13688 2252 13694 2264
rect 20165 2261 20177 2295
rect 20211 2292 20223 2295
rect 20438 2292 20444 2304
rect 20211 2264 20444 2292
rect 20211 2261 20223 2264
rect 20165 2255 20223 2261
rect 20438 2252 20444 2264
rect 20496 2252 20502 2304
rect 20717 2295 20775 2301
rect 20717 2261 20729 2295
rect 20763 2292 20775 2295
rect 21082 2292 21088 2304
rect 20763 2264 21088 2292
rect 20763 2261 20775 2264
rect 20717 2255 20775 2261
rect 21082 2252 21088 2264
rect 21140 2252 21146 2304
rect 21468 2301 21496 2400
rect 21634 2388 21640 2440
rect 21692 2388 21698 2440
rect 22281 2431 22339 2437
rect 22281 2397 22293 2431
rect 22327 2428 22339 2431
rect 22327 2400 22692 2428
rect 22327 2397 22339 2400
rect 22281 2391 22339 2397
rect 21726 2320 21732 2372
rect 21784 2360 21790 2372
rect 21784 2332 22600 2360
rect 21784 2320 21790 2332
rect 22572 2304 22600 2332
rect 21453 2295 21511 2301
rect 21453 2261 21465 2295
rect 21499 2261 21511 2295
rect 21453 2255 21511 2261
rect 21542 2252 21548 2304
rect 21600 2292 21606 2304
rect 22370 2292 22376 2304
rect 21600 2264 22376 2292
rect 21600 2252 21606 2264
rect 22370 2252 22376 2264
rect 22428 2252 22434 2304
rect 22554 2252 22560 2304
rect 22612 2252 22618 2304
rect 22664 2301 22692 2400
rect 22830 2388 22836 2440
rect 22888 2388 22894 2440
rect 22940 2437 22968 2468
rect 25148 2468 26648 2496
rect 26712 2468 27844 2496
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 23382 2388 23388 2440
rect 23440 2388 23446 2440
rect 23566 2388 23572 2440
rect 23624 2388 23630 2440
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2428 23903 2431
rect 24302 2428 24308 2440
rect 23891 2400 24308 2428
rect 23891 2397 23903 2400
rect 23845 2391 23903 2397
rect 24302 2388 24308 2400
rect 24360 2388 24366 2440
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 25038 2388 25044 2440
rect 25096 2388 25102 2440
rect 24946 2360 24952 2372
rect 23124 2332 24952 2360
rect 23124 2301 23152 2332
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 22649 2295 22707 2301
rect 22649 2261 22661 2295
rect 22695 2261 22707 2295
rect 22649 2255 22707 2261
rect 23109 2295 23167 2301
rect 23109 2261 23121 2295
rect 23155 2261 23167 2295
rect 23109 2255 23167 2261
rect 23201 2295 23259 2301
rect 23201 2261 23213 2295
rect 23247 2292 23259 2295
rect 24210 2292 24216 2304
rect 23247 2264 24216 2292
rect 23247 2261 23259 2264
rect 23201 2255 23259 2261
rect 24210 2252 24216 2264
rect 24268 2252 24274 2304
rect 24486 2252 24492 2304
rect 24544 2292 24550 2304
rect 25148 2292 25176 2468
rect 25501 2431 25559 2437
rect 25501 2397 25513 2431
rect 25547 2428 25559 2431
rect 25866 2428 25872 2440
rect 25547 2400 25872 2428
rect 25547 2397 25559 2400
rect 25501 2391 25559 2397
rect 25866 2388 25872 2400
rect 25924 2388 25930 2440
rect 25958 2388 25964 2440
rect 26016 2388 26022 2440
rect 26712 2437 26740 2468
rect 26697 2431 26755 2437
rect 26697 2397 26709 2431
rect 26743 2397 26755 2431
rect 26697 2391 26755 2397
rect 27338 2388 27344 2440
rect 27396 2388 27402 2440
rect 27798 2388 27804 2440
rect 27856 2428 27862 2440
rect 27985 2431 28043 2437
rect 27985 2428 27997 2431
rect 27856 2400 27997 2428
rect 27856 2388 27862 2400
rect 27985 2397 27997 2400
rect 28031 2397 28043 2431
rect 27985 2391 28043 2397
rect 25225 2363 25283 2369
rect 25225 2329 25237 2363
rect 25271 2360 25283 2363
rect 26970 2360 26976 2372
rect 25271 2332 26976 2360
rect 25271 2329 25283 2332
rect 25225 2323 25283 2329
rect 26970 2320 26976 2332
rect 27028 2320 27034 2372
rect 28092 2360 28120 2604
rect 28442 2592 28448 2644
rect 28500 2632 28506 2644
rect 28721 2635 28779 2641
rect 28721 2632 28733 2635
rect 28500 2604 28733 2632
rect 28500 2592 28506 2604
rect 28721 2601 28733 2604
rect 28767 2601 28779 2635
rect 28721 2595 28779 2601
rect 28902 2592 28908 2644
rect 28960 2632 28966 2644
rect 30926 2632 30932 2644
rect 28960 2604 30932 2632
rect 28960 2592 28966 2604
rect 30926 2592 30932 2604
rect 30984 2592 30990 2644
rect 31297 2635 31355 2641
rect 31297 2632 31309 2635
rect 31220 2604 31309 2632
rect 31220 2576 31248 2604
rect 31297 2601 31309 2604
rect 31343 2601 31355 2635
rect 31297 2595 31355 2601
rect 35066 2592 35072 2644
rect 35124 2632 35130 2644
rect 35345 2635 35403 2641
rect 35345 2632 35357 2635
rect 35124 2604 35357 2632
rect 35124 2592 35130 2604
rect 35345 2601 35357 2604
rect 35391 2601 35403 2635
rect 35345 2595 35403 2601
rect 37366 2592 37372 2644
rect 37424 2632 37430 2644
rect 37553 2635 37611 2641
rect 37553 2632 37565 2635
rect 37424 2604 37565 2632
rect 37424 2592 37430 2604
rect 37553 2601 37565 2604
rect 37599 2601 37611 2635
rect 37553 2595 37611 2601
rect 37660 2604 41644 2632
rect 30469 2567 30527 2573
rect 30469 2533 30481 2567
rect 30515 2533 30527 2567
rect 30469 2527 30527 2533
rect 30484 2496 30512 2527
rect 31018 2524 31024 2576
rect 31076 2524 31082 2576
rect 31202 2524 31208 2576
rect 31260 2524 31266 2576
rect 37660 2564 37688 2604
rect 41506 2564 41512 2576
rect 32324 2536 34836 2564
rect 30834 2496 30840 2508
rect 30484 2468 30840 2496
rect 30834 2456 30840 2468
rect 30892 2456 30898 2508
rect 28258 2388 28264 2440
rect 28316 2388 28322 2440
rect 28534 2388 28540 2440
rect 28592 2388 28598 2440
rect 28905 2431 28963 2437
rect 28905 2397 28917 2431
rect 28951 2428 28963 2431
rect 30006 2428 30012 2440
rect 28951 2400 30012 2428
rect 28951 2397 28963 2400
rect 28905 2391 28963 2397
rect 30006 2388 30012 2400
rect 30064 2388 30070 2440
rect 30098 2388 30104 2440
rect 30156 2428 30162 2440
rect 30285 2431 30343 2437
rect 30285 2428 30297 2431
rect 30156 2400 30297 2428
rect 30156 2388 30162 2400
rect 30285 2397 30297 2400
rect 30331 2397 30343 2431
rect 30285 2391 30343 2397
rect 30374 2388 30380 2440
rect 30432 2428 30438 2440
rect 30653 2431 30711 2437
rect 30653 2428 30665 2431
rect 30432 2400 30665 2428
rect 30432 2388 30438 2400
rect 30653 2397 30665 2400
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 30929 2431 30987 2437
rect 30929 2428 30941 2431
rect 30800 2400 30941 2428
rect 30800 2388 30806 2400
rect 30929 2397 30941 2400
rect 30975 2397 30987 2431
rect 30929 2391 30987 2397
rect 31205 2431 31263 2437
rect 31205 2397 31217 2431
rect 31251 2397 31263 2431
rect 31205 2391 31263 2397
rect 31018 2360 31024 2372
rect 28092 2332 31024 2360
rect 31018 2320 31024 2332
rect 31076 2320 31082 2372
rect 31220 2360 31248 2391
rect 31478 2388 31484 2440
rect 31536 2388 31542 2440
rect 32324 2437 32352 2536
rect 34808 2496 34836 2536
rect 36004 2536 37688 2564
rect 38028 2536 41512 2564
rect 36004 2496 36032 2536
rect 34808 2468 36032 2496
rect 36078 2456 36084 2508
rect 36136 2496 36142 2508
rect 36136 2468 37964 2496
rect 36136 2456 36142 2468
rect 32309 2431 32367 2437
rect 32309 2397 32321 2431
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 32858 2388 32864 2440
rect 32916 2388 32922 2440
rect 33318 2388 33324 2440
rect 33376 2388 33382 2440
rect 35529 2431 35587 2437
rect 35529 2397 35541 2431
rect 35575 2428 35587 2431
rect 35894 2428 35900 2440
rect 35575 2400 35900 2428
rect 35575 2397 35587 2400
rect 35529 2391 35587 2397
rect 35894 2388 35900 2400
rect 35952 2388 35958 2440
rect 37737 2431 37795 2437
rect 37737 2397 37749 2431
rect 37783 2428 37795 2431
rect 37783 2400 37872 2428
rect 37783 2397 37795 2400
rect 37737 2391 37795 2397
rect 31220 2332 31754 2360
rect 24544 2264 25176 2292
rect 25777 2295 25835 2301
rect 24544 2252 24550 2264
rect 25777 2261 25789 2295
rect 25823 2292 25835 2295
rect 26510 2292 26516 2304
rect 25823 2264 26516 2292
rect 25823 2261 25835 2264
rect 25777 2255 25835 2261
rect 26510 2252 26516 2264
rect 26568 2252 26574 2304
rect 27154 2252 27160 2304
rect 27212 2252 27218 2304
rect 28074 2252 28080 2304
rect 28132 2252 28138 2304
rect 28353 2295 28411 2301
rect 28353 2261 28365 2295
rect 28399 2292 28411 2295
rect 28994 2292 29000 2304
rect 28399 2264 29000 2292
rect 28399 2261 28411 2264
rect 28353 2255 28411 2261
rect 28994 2252 29000 2264
rect 29052 2252 29058 2304
rect 30101 2295 30159 2301
rect 30101 2261 30113 2295
rect 30147 2292 30159 2295
rect 30650 2292 30656 2304
rect 30147 2264 30656 2292
rect 30147 2261 30159 2264
rect 30101 2255 30159 2261
rect 30650 2252 30656 2264
rect 30708 2252 30714 2304
rect 30745 2295 30803 2301
rect 30745 2261 30757 2295
rect 30791 2292 30803 2295
rect 31570 2292 31576 2304
rect 30791 2264 31576 2292
rect 30791 2261 30803 2264
rect 30745 2255 30803 2261
rect 31570 2252 31576 2264
rect 31628 2252 31634 2304
rect 31726 2292 31754 2332
rect 32125 2295 32183 2301
rect 32125 2292 32137 2295
rect 31726 2264 32137 2292
rect 32125 2261 32137 2264
rect 32171 2261 32183 2295
rect 32125 2255 32183 2261
rect 32677 2295 32735 2301
rect 32677 2261 32689 2295
rect 32723 2292 32735 2295
rect 32950 2292 32956 2304
rect 32723 2264 32956 2292
rect 32723 2261 32735 2264
rect 32677 2255 32735 2261
rect 32950 2252 32956 2264
rect 33008 2252 33014 2304
rect 33134 2252 33140 2304
rect 33192 2252 33198 2304
rect 37844 2301 37872 2400
rect 37936 2360 37964 2468
rect 38028 2437 38056 2536
rect 41506 2524 41512 2536
rect 41564 2524 41570 2576
rect 41616 2564 41644 2604
rect 41690 2592 41696 2644
rect 41748 2632 41754 2644
rect 42061 2635 42119 2641
rect 42061 2632 42073 2635
rect 41748 2604 42073 2632
rect 41748 2592 41754 2604
rect 42061 2601 42073 2604
rect 42107 2601 42119 2635
rect 42061 2595 42119 2601
rect 44726 2592 44732 2644
rect 44784 2592 44790 2644
rect 45002 2592 45008 2644
rect 45060 2592 45066 2644
rect 45649 2635 45707 2641
rect 45649 2601 45661 2635
rect 45695 2632 45707 2635
rect 46106 2632 46112 2644
rect 45695 2604 46112 2632
rect 45695 2601 45707 2604
rect 45649 2595 45707 2601
rect 46106 2592 46112 2604
rect 46164 2592 46170 2644
rect 44450 2564 44456 2576
rect 41616 2536 44456 2564
rect 44450 2524 44456 2536
rect 44508 2524 44514 2576
rect 38013 2431 38071 2437
rect 38013 2397 38025 2431
rect 38059 2397 38071 2431
rect 38013 2391 38071 2397
rect 38381 2431 38439 2437
rect 38381 2397 38393 2431
rect 38427 2397 38439 2431
rect 38381 2391 38439 2397
rect 38396 2360 38424 2391
rect 42242 2388 42248 2440
rect 42300 2388 42306 2440
rect 44542 2388 44548 2440
rect 44600 2388 44606 2440
rect 45186 2388 45192 2440
rect 45244 2388 45250 2440
rect 45830 2388 45836 2440
rect 45888 2388 45894 2440
rect 42794 2360 42800 2372
rect 37936 2332 38424 2360
rect 41386 2332 42800 2360
rect 37829 2295 37887 2301
rect 37829 2261 37841 2295
rect 37875 2261 37887 2295
rect 37829 2255 37887 2261
rect 38010 2252 38016 2304
rect 38068 2292 38074 2304
rect 38565 2295 38623 2301
rect 38565 2292 38577 2295
rect 38068 2264 38577 2292
rect 38068 2252 38074 2264
rect 38565 2261 38577 2264
rect 38611 2261 38623 2295
rect 38565 2255 38623 2261
rect 38654 2252 38660 2304
rect 38712 2292 38718 2304
rect 41386 2292 41414 2332
rect 42794 2320 42800 2332
rect 42852 2320 42858 2372
rect 38712 2264 41414 2292
rect 38712 2252 38718 2264
rect 1104 2202 46984 2224
rect 1104 2150 12380 2202
rect 12432 2150 12444 2202
rect 12496 2150 12508 2202
rect 12560 2150 12572 2202
rect 12624 2150 12636 2202
rect 12688 2150 23810 2202
rect 23862 2150 23874 2202
rect 23926 2150 23938 2202
rect 23990 2150 24002 2202
rect 24054 2150 24066 2202
rect 24118 2150 35240 2202
rect 35292 2150 35304 2202
rect 35356 2150 35368 2202
rect 35420 2150 35432 2202
rect 35484 2150 35496 2202
rect 35548 2150 46670 2202
rect 46722 2150 46734 2202
rect 46786 2150 46798 2202
rect 46850 2150 46862 2202
rect 46914 2150 46926 2202
rect 46978 2150 46984 2202
rect 1104 2128 46984 2150
rect 4341 2091 4399 2097
rect 4341 2057 4353 2091
rect 4387 2088 4399 2091
rect 15194 2088 15200 2100
rect 4387 2060 15200 2088
rect 4387 2057 4399 2060
rect 4341 2051 4399 2057
rect 15194 2048 15200 2060
rect 15252 2048 15258 2100
rect 15930 2048 15936 2100
rect 15988 2048 15994 2100
rect 16482 2048 16488 2100
rect 16540 2048 16546 2100
rect 16942 2048 16948 2100
rect 17000 2048 17006 2100
rect 17310 2048 17316 2100
rect 17368 2088 17374 2100
rect 17497 2091 17555 2097
rect 17497 2088 17509 2091
rect 17368 2060 17509 2088
rect 17368 2048 17374 2060
rect 17497 2057 17509 2060
rect 17543 2057 17555 2091
rect 17497 2051 17555 2057
rect 17589 2091 17647 2097
rect 17589 2057 17601 2091
rect 17635 2088 17647 2091
rect 17954 2088 17960 2100
rect 17635 2060 17960 2088
rect 17635 2057 17647 2060
rect 17589 2051 17647 2057
rect 17954 2048 17960 2060
rect 18012 2048 18018 2100
rect 18601 2091 18659 2097
rect 18601 2057 18613 2091
rect 18647 2057 18659 2091
rect 18601 2051 18659 2057
rect 17218 1980 17224 2032
rect 17276 2020 17282 2032
rect 18616 2020 18644 2051
rect 18874 2048 18880 2100
rect 18932 2048 18938 2100
rect 19245 2091 19303 2097
rect 19245 2057 19257 2091
rect 19291 2088 19303 2091
rect 19426 2088 19432 2100
rect 19291 2060 19432 2088
rect 19291 2057 19303 2060
rect 19245 2051 19303 2057
rect 19426 2048 19432 2060
rect 19484 2048 19490 2100
rect 19797 2091 19855 2097
rect 19797 2057 19809 2091
rect 19843 2088 19855 2091
rect 19978 2088 19984 2100
rect 19843 2060 19984 2088
rect 19843 2057 19855 2060
rect 19797 2051 19855 2057
rect 19978 2048 19984 2060
rect 20036 2048 20042 2100
rect 20073 2091 20131 2097
rect 20073 2057 20085 2091
rect 20119 2088 20131 2091
rect 20162 2088 20168 2100
rect 20119 2060 20168 2088
rect 20119 2057 20131 2060
rect 20073 2051 20131 2057
rect 20162 2048 20168 2060
rect 20220 2048 20226 2100
rect 20530 2048 20536 2100
rect 20588 2048 20594 2100
rect 21177 2091 21235 2097
rect 21177 2057 21189 2091
rect 21223 2057 21235 2091
rect 21177 2051 21235 2057
rect 21913 2091 21971 2097
rect 21913 2057 21925 2091
rect 21959 2088 21971 2091
rect 23293 2091 23351 2097
rect 21959 2060 22876 2088
rect 21959 2057 21971 2060
rect 21913 2051 21971 2057
rect 19610 2020 19616 2032
rect 17276 1992 17908 2020
rect 17276 1980 17282 1992
rect 1118 1912 1124 1964
rect 1176 1952 1182 1964
rect 1397 1955 1455 1961
rect 1397 1952 1409 1955
rect 1176 1924 1409 1952
rect 1176 1912 1182 1924
rect 1397 1921 1409 1924
rect 1443 1921 1455 1955
rect 1397 1915 1455 1921
rect 3970 1912 3976 1964
rect 4028 1952 4034 1964
rect 4157 1955 4215 1961
rect 4157 1952 4169 1955
rect 4028 1924 4169 1952
rect 4028 1912 4034 1924
rect 4157 1921 4169 1924
rect 4203 1921 4215 1955
rect 4157 1915 4215 1921
rect 4522 1912 4528 1964
rect 4580 1912 4586 1964
rect 15746 1912 15752 1964
rect 15804 1912 15810 1964
rect 16022 1912 16028 1964
rect 16080 1912 16086 1964
rect 16298 1912 16304 1964
rect 16356 1912 16362 1964
rect 16758 1912 16764 1964
rect 16816 1912 16822 1964
rect 17034 1912 17040 1964
rect 17092 1912 17098 1964
rect 17310 1912 17316 1964
rect 17368 1912 17374 1964
rect 17770 1912 17776 1964
rect 17828 1912 17834 1964
rect 17880 1961 17908 1992
rect 17972 1992 18460 2020
rect 18616 1992 19616 2020
rect 17972 1964 18000 1992
rect 17865 1955 17923 1961
rect 17865 1921 17877 1955
rect 17911 1921 17923 1955
rect 17865 1915 17923 1921
rect 17954 1912 17960 1964
rect 18012 1912 18018 1964
rect 18432 1961 18460 1992
rect 19610 1980 19616 1992
rect 19668 1980 19674 2032
rect 21192 2020 21220 2051
rect 22848 2020 22876 2060
rect 23293 2057 23305 2091
rect 23339 2088 23351 2091
rect 23566 2088 23572 2100
rect 23339 2060 23572 2088
rect 23339 2057 23351 2060
rect 23293 2051 23351 2057
rect 23566 2048 23572 2060
rect 23624 2048 23630 2100
rect 24302 2048 24308 2100
rect 24360 2048 24366 2100
rect 24581 2091 24639 2097
rect 24581 2057 24593 2091
rect 24627 2088 24639 2091
rect 24670 2088 24676 2100
rect 24627 2060 24676 2088
rect 24627 2057 24639 2060
rect 24581 2051 24639 2057
rect 24670 2048 24676 2060
rect 24728 2048 24734 2100
rect 24949 2091 25007 2097
rect 24949 2057 24961 2091
rect 24995 2057 25007 2091
rect 24949 2051 25007 2057
rect 24964 2020 24992 2051
rect 25038 2048 25044 2100
rect 25096 2088 25102 2100
rect 25501 2091 25559 2097
rect 25501 2088 25513 2091
rect 25096 2060 25513 2088
rect 25096 2048 25102 2060
rect 25501 2057 25513 2060
rect 25547 2057 25559 2091
rect 25501 2051 25559 2057
rect 25866 2048 25872 2100
rect 25924 2088 25930 2100
rect 26513 2091 26571 2097
rect 26513 2088 26525 2091
rect 25924 2060 26525 2088
rect 25924 2048 25930 2060
rect 26513 2057 26525 2060
rect 26559 2057 26571 2091
rect 26513 2051 26571 2057
rect 26970 2048 26976 2100
rect 27028 2048 27034 2100
rect 27154 2048 27160 2100
rect 27212 2088 27218 2100
rect 28077 2091 28135 2097
rect 27212 2060 28028 2088
rect 27212 2048 27218 2060
rect 28000 2020 28028 2060
rect 28077 2057 28089 2091
rect 28123 2088 28135 2091
rect 28902 2088 28908 2100
rect 28123 2060 28908 2088
rect 28123 2057 28135 2060
rect 28077 2051 28135 2057
rect 28902 2048 28908 2060
rect 28960 2048 28966 2100
rect 29089 2091 29147 2097
rect 29089 2057 29101 2091
rect 29135 2088 29147 2091
rect 29178 2088 29184 2100
rect 29135 2060 29184 2088
rect 29135 2057 29147 2060
rect 29089 2051 29147 2057
rect 29178 2048 29184 2060
rect 29236 2048 29242 2100
rect 29273 2091 29331 2097
rect 29273 2057 29285 2091
rect 29319 2088 29331 2091
rect 29319 2060 29960 2088
rect 29319 2057 29331 2060
rect 29273 2051 29331 2057
rect 21192 1992 22508 2020
rect 22848 1992 23612 2020
rect 24964 1992 25912 2020
rect 28000 1992 28488 2020
rect 18141 1955 18199 1961
rect 18141 1921 18153 1955
rect 18187 1921 18199 1955
rect 18141 1915 18199 1921
rect 18417 1955 18475 1961
rect 18417 1921 18429 1955
rect 18463 1921 18475 1955
rect 18417 1915 18475 1921
rect 14550 1844 14556 1896
rect 14608 1884 14614 1896
rect 14608 1856 17264 1884
rect 14608 1844 14614 1856
rect 4709 1819 4767 1825
rect 4709 1785 4721 1819
rect 4755 1816 4767 1819
rect 17126 1816 17132 1828
rect 4755 1788 17132 1816
rect 4755 1785 4767 1788
rect 4709 1779 4767 1785
rect 17126 1776 17132 1788
rect 17184 1776 17190 1828
rect 17236 1816 17264 1856
rect 17678 1844 17684 1896
rect 17736 1884 17742 1896
rect 18156 1884 18184 1915
rect 18690 1912 18696 1964
rect 18748 1912 18754 1964
rect 18874 1912 18880 1964
rect 18932 1952 18938 1964
rect 19153 1955 19211 1961
rect 19153 1952 19165 1955
rect 18932 1924 19165 1952
rect 18932 1912 18938 1924
rect 19153 1921 19165 1924
rect 19199 1921 19211 1955
rect 19153 1915 19211 1921
rect 19426 1912 19432 1964
rect 19484 1912 19490 1964
rect 19518 1912 19524 1964
rect 19576 1912 19582 1964
rect 19981 1955 20039 1961
rect 19981 1936 19993 1955
rect 19904 1921 19993 1936
rect 20027 1921 20039 1955
rect 19904 1915 20039 1921
rect 19904 1908 20024 1915
rect 20254 1912 20260 1964
rect 20312 1912 20318 1964
rect 20346 1912 20352 1964
rect 20404 1912 20410 1964
rect 20438 1912 20444 1964
rect 20496 1952 20502 1964
rect 20625 1955 20683 1961
rect 20625 1952 20637 1955
rect 20496 1924 20637 1952
rect 20496 1912 20502 1924
rect 20625 1921 20637 1924
rect 20671 1921 20683 1955
rect 20625 1915 20683 1921
rect 21358 1912 21364 1964
rect 21416 1912 21422 1964
rect 21634 1912 21640 1964
rect 21692 1912 21698 1964
rect 22094 1912 22100 1964
rect 22152 1912 22158 1964
rect 22370 1912 22376 1964
rect 22428 1912 22434 1964
rect 22480 1961 22508 1992
rect 22465 1955 22523 1961
rect 22465 1921 22477 1955
rect 22511 1921 22523 1955
rect 22465 1915 22523 1921
rect 22554 1912 22560 1964
rect 22612 1952 22618 1964
rect 23584 1961 23612 1992
rect 23201 1955 23259 1961
rect 23201 1952 23213 1955
rect 22612 1924 23213 1952
rect 22612 1912 22618 1924
rect 23201 1921 23213 1924
rect 23247 1921 23259 1955
rect 23201 1915 23259 1921
rect 23477 1955 23535 1961
rect 23477 1921 23489 1955
rect 23523 1921 23535 1955
rect 23477 1915 23535 1921
rect 23569 1955 23627 1961
rect 23569 1921 23581 1955
rect 23615 1921 23627 1955
rect 23569 1915 23627 1921
rect 19334 1884 19340 1896
rect 17736 1856 18184 1884
rect 18248 1856 19340 1884
rect 17736 1844 17742 1856
rect 18248 1816 18276 1856
rect 19334 1844 19340 1856
rect 19392 1844 19398 1896
rect 19702 1844 19708 1896
rect 19760 1884 19766 1896
rect 19904 1884 19932 1908
rect 19760 1856 19932 1884
rect 23492 1884 23520 1915
rect 23658 1912 23664 1964
rect 23716 1952 23722 1964
rect 24213 1955 24271 1961
rect 24213 1952 24225 1955
rect 23716 1924 24225 1952
rect 23716 1912 23722 1924
rect 24213 1921 24225 1924
rect 24259 1921 24271 1955
rect 24213 1915 24271 1921
rect 24486 1912 24492 1964
rect 24544 1912 24550 1964
rect 24762 1912 24768 1964
rect 24820 1912 24826 1964
rect 25130 1912 25136 1964
rect 25188 1912 25194 1964
rect 25406 1912 25412 1964
rect 25464 1912 25470 1964
rect 25682 1912 25688 1964
rect 25740 1912 25746 1964
rect 25884 1961 25912 1992
rect 25869 1955 25927 1961
rect 25869 1921 25881 1955
rect 25915 1921 25927 1955
rect 25869 1915 25927 1921
rect 26418 1912 26424 1964
rect 26476 1912 26482 1964
rect 26697 1955 26755 1961
rect 26697 1921 26709 1955
rect 26743 1952 26755 1955
rect 26878 1952 26884 1964
rect 26743 1924 26884 1952
rect 26743 1921 26755 1924
rect 26697 1915 26755 1921
rect 26878 1912 26884 1924
rect 26936 1912 26942 1964
rect 27157 1955 27215 1961
rect 27157 1936 27169 1955
rect 27080 1921 27169 1936
rect 27203 1921 27215 1955
rect 27080 1915 27215 1921
rect 27080 1908 27200 1915
rect 27246 1912 27252 1964
rect 27304 1952 27310 1964
rect 27304 1924 27384 1952
rect 27304 1912 27310 1924
rect 26602 1884 26608 1896
rect 23492 1856 26608 1884
rect 19760 1844 19766 1856
rect 26602 1844 26608 1856
rect 26660 1844 26666 1896
rect 17236 1788 18276 1816
rect 18325 1819 18383 1825
rect 18325 1785 18337 1819
rect 18371 1816 18383 1819
rect 21818 1816 21824 1828
rect 18371 1788 21824 1816
rect 18371 1785 18383 1788
rect 18325 1779 18383 1785
rect 21818 1776 21824 1788
rect 21876 1776 21882 1828
rect 22189 1819 22247 1825
rect 22189 1785 22201 1819
rect 22235 1816 22247 1819
rect 23474 1816 23480 1828
rect 22235 1788 23480 1816
rect 22235 1785 22247 1788
rect 22189 1779 22247 1785
rect 23474 1776 23480 1788
rect 23532 1776 23538 1828
rect 23676 1788 24532 1816
rect 1578 1708 1584 1760
rect 1636 1708 1642 1760
rect 16206 1708 16212 1760
rect 16264 1708 16270 1760
rect 17221 1751 17279 1757
rect 17221 1717 17233 1751
rect 17267 1748 17279 1751
rect 17494 1748 17500 1760
rect 17267 1720 17500 1748
rect 17267 1717 17279 1720
rect 17221 1711 17279 1717
rect 17494 1708 17500 1720
rect 17552 1708 17558 1760
rect 18049 1751 18107 1757
rect 18049 1717 18061 1751
rect 18095 1748 18107 1751
rect 18506 1748 18512 1760
rect 18095 1720 18512 1748
rect 18095 1717 18107 1720
rect 18049 1711 18107 1717
rect 18506 1708 18512 1720
rect 18564 1708 18570 1760
rect 18969 1751 19027 1757
rect 18969 1717 18981 1751
rect 19015 1748 19027 1751
rect 19150 1748 19156 1760
rect 19015 1720 19156 1748
rect 19015 1717 19027 1720
rect 18969 1711 19027 1717
rect 19150 1708 19156 1720
rect 19208 1708 19214 1760
rect 19705 1751 19763 1757
rect 19705 1717 19717 1751
rect 19751 1748 19763 1751
rect 20438 1748 20444 1760
rect 19751 1720 20444 1748
rect 19751 1717 19763 1720
rect 19705 1711 19763 1717
rect 20438 1708 20444 1720
rect 20496 1708 20502 1760
rect 20806 1708 20812 1760
rect 20864 1708 20870 1760
rect 21453 1751 21511 1757
rect 21453 1717 21465 1751
rect 21499 1748 21511 1751
rect 21910 1748 21916 1760
rect 21499 1720 21916 1748
rect 21499 1717 21511 1720
rect 21453 1711 21511 1717
rect 21910 1708 21916 1720
rect 21968 1708 21974 1760
rect 22646 1708 22652 1760
rect 22704 1708 22710 1760
rect 23017 1751 23075 1757
rect 23017 1717 23029 1751
rect 23063 1748 23075 1751
rect 23676 1748 23704 1788
rect 23063 1720 23704 1748
rect 23063 1717 23075 1720
rect 23017 1711 23075 1717
rect 23750 1708 23756 1760
rect 23808 1708 23814 1760
rect 24026 1708 24032 1760
rect 24084 1708 24090 1760
rect 24504 1748 24532 1788
rect 24578 1776 24584 1828
rect 24636 1816 24642 1828
rect 25225 1819 25283 1825
rect 25225 1816 25237 1819
rect 24636 1788 25237 1816
rect 24636 1776 24642 1788
rect 25225 1785 25237 1788
rect 25271 1785 25283 1819
rect 26786 1816 26792 1828
rect 25225 1779 25283 1785
rect 25976 1788 26792 1816
rect 24854 1748 24860 1760
rect 24504 1720 24860 1748
rect 24854 1708 24860 1720
rect 24912 1708 24918 1760
rect 24946 1708 24952 1760
rect 25004 1748 25010 1760
rect 25976 1748 26004 1788
rect 26786 1776 26792 1788
rect 26844 1776 26850 1828
rect 27080 1816 27108 1908
rect 27356 1884 27384 1924
rect 27430 1912 27436 1964
rect 27488 1912 27494 1964
rect 27706 1912 27712 1964
rect 27764 1912 27770 1964
rect 27985 1955 28043 1961
rect 27985 1921 27997 1955
rect 28031 1952 28043 1955
rect 28166 1952 28172 1964
rect 28031 1924 28172 1952
rect 28031 1921 28043 1924
rect 27985 1915 28043 1921
rect 28166 1912 28172 1924
rect 28224 1912 28230 1964
rect 28258 1912 28264 1964
rect 28316 1912 28322 1964
rect 28460 1961 28488 1992
rect 29362 1980 29368 2032
rect 29420 2020 29426 2032
rect 29420 1992 29776 2020
rect 29420 1980 29426 1992
rect 28445 1955 28503 1961
rect 28445 1921 28457 1955
rect 28491 1921 28503 1955
rect 28445 1915 28503 1921
rect 28997 1955 29055 1961
rect 28997 1921 29009 1955
rect 29043 1952 29055 1955
rect 29270 1952 29276 1964
rect 29043 1924 29276 1952
rect 29043 1921 29055 1924
rect 28997 1915 29055 1921
rect 29270 1912 29276 1924
rect 29328 1912 29334 1964
rect 29457 1955 29515 1961
rect 29457 1921 29469 1955
rect 29503 1952 29515 1955
rect 29638 1952 29644 1964
rect 29503 1924 29644 1952
rect 29503 1921 29515 1924
rect 29457 1915 29515 1921
rect 29638 1912 29644 1924
rect 29696 1912 29702 1964
rect 29748 1961 29776 1992
rect 29932 1961 29960 2060
rect 30006 2048 30012 2100
rect 30064 2088 30070 2100
rect 30561 2091 30619 2097
rect 30561 2088 30573 2091
rect 30064 2060 30573 2088
rect 30064 2048 30070 2060
rect 30561 2057 30573 2060
rect 30607 2057 30619 2091
rect 30561 2051 30619 2057
rect 30926 2048 30932 2100
rect 30984 2088 30990 2100
rect 30984 2060 32996 2088
rect 30984 2048 30990 2060
rect 31113 2023 31171 2029
rect 31113 1989 31125 2023
rect 31159 2020 31171 2023
rect 31202 2020 31208 2032
rect 31159 1992 31208 2020
rect 31159 1989 31171 1992
rect 31113 1983 31171 1989
rect 31202 1980 31208 1992
rect 31260 1980 31266 2032
rect 32968 2020 32996 2060
rect 33318 2048 33324 2100
rect 33376 2088 33382 2100
rect 34517 2091 34575 2097
rect 34517 2088 34529 2091
rect 33376 2060 34529 2088
rect 33376 2048 33382 2060
rect 34517 2057 34529 2060
rect 34563 2057 34575 2091
rect 34517 2051 34575 2057
rect 35894 2048 35900 2100
rect 35952 2048 35958 2100
rect 38654 2088 38660 2100
rect 36004 2060 38660 2088
rect 35526 2020 35532 2032
rect 32508 1992 32904 2020
rect 32968 1992 34192 2020
rect 29733 1955 29791 1961
rect 29733 1921 29745 1955
rect 29779 1921 29791 1955
rect 29733 1915 29791 1921
rect 29917 1955 29975 1961
rect 29917 1921 29929 1955
rect 29963 1921 29975 1955
rect 29917 1915 29975 1921
rect 30466 1912 30472 1964
rect 30524 1912 30530 1964
rect 30742 1912 30748 1964
rect 30800 1912 30806 1964
rect 31570 1912 31576 1964
rect 31628 1912 31634 1964
rect 32306 1912 32312 1964
rect 32364 1912 32370 1964
rect 32508 1952 32536 1992
rect 32416 1924 32536 1952
rect 32122 1884 32128 1896
rect 27356 1856 32128 1884
rect 32122 1844 32128 1856
rect 32180 1844 32186 1896
rect 29362 1816 29368 1828
rect 27080 1788 29368 1816
rect 29362 1776 29368 1788
rect 29420 1776 29426 1828
rect 29549 1819 29607 1825
rect 29549 1785 29561 1819
rect 29595 1816 29607 1819
rect 30374 1816 30380 1828
rect 29595 1788 30380 1816
rect 29595 1785 29607 1788
rect 29549 1779 29607 1785
rect 30374 1776 30380 1788
rect 30432 1776 30438 1828
rect 31662 1776 31668 1828
rect 31720 1816 31726 1828
rect 32416 1825 32444 1924
rect 32582 1912 32588 1964
rect 32640 1912 32646 1964
rect 32876 1961 32904 1992
rect 32861 1955 32919 1961
rect 32861 1921 32873 1955
rect 32907 1921 32919 1955
rect 32861 1915 32919 1921
rect 33410 1912 33416 1964
rect 33468 1912 33474 1964
rect 34164 1961 34192 1992
rect 34716 1992 35532 2020
rect 34716 1961 34744 1992
rect 35526 1980 35532 1992
rect 35584 1980 35590 2032
rect 35710 1980 35716 2032
rect 35768 2020 35774 2032
rect 36004 2020 36032 2060
rect 38654 2048 38660 2060
rect 38712 2048 38718 2100
rect 42242 2048 42248 2100
rect 42300 2088 42306 2100
rect 42429 2091 42487 2097
rect 42429 2088 42441 2091
rect 42300 2060 42441 2088
rect 42300 2048 42306 2060
rect 42429 2057 42441 2060
rect 42475 2057 42487 2091
rect 42429 2051 42487 2057
rect 44542 2048 44548 2100
rect 44600 2088 44606 2100
rect 45097 2091 45155 2097
rect 45097 2088 45109 2091
rect 44600 2060 45109 2088
rect 44600 2048 44606 2060
rect 45097 2057 45109 2060
rect 45143 2057 45155 2091
rect 45097 2051 45155 2057
rect 45186 2048 45192 2100
rect 45244 2088 45250 2100
rect 45373 2091 45431 2097
rect 45373 2088 45385 2091
rect 45244 2060 45385 2088
rect 45244 2048 45250 2060
rect 45373 2057 45385 2060
rect 45419 2057 45431 2091
rect 45373 2051 45431 2057
rect 45649 2091 45707 2097
rect 45649 2057 45661 2091
rect 45695 2088 45707 2091
rect 45830 2088 45836 2100
rect 45695 2060 45836 2088
rect 45695 2057 45707 2060
rect 45649 2051 45707 2057
rect 45830 2048 45836 2060
rect 45888 2048 45894 2100
rect 46293 2091 46351 2097
rect 46293 2057 46305 2091
rect 46339 2057 46351 2091
rect 46293 2051 46351 2057
rect 45002 2020 45008 2032
rect 35768 1992 36032 2020
rect 36188 1992 45008 2020
rect 35768 1980 35774 1992
rect 33689 1955 33747 1961
rect 33689 1921 33701 1955
rect 33735 1921 33747 1955
rect 33689 1915 33747 1921
rect 34149 1955 34207 1961
rect 34149 1921 34161 1955
rect 34195 1921 34207 1955
rect 34149 1915 34207 1921
rect 34701 1955 34759 1961
rect 34701 1921 34713 1955
rect 34747 1921 34759 1955
rect 35437 1955 35495 1961
rect 35437 1952 35449 1955
rect 34701 1915 34759 1921
rect 34808 1924 35449 1952
rect 32490 1844 32496 1896
rect 32548 1884 32554 1896
rect 33704 1884 33732 1915
rect 32548 1856 33732 1884
rect 32548 1844 32554 1856
rect 33778 1844 33784 1896
rect 33836 1884 33842 1896
rect 34808 1884 34836 1924
rect 35437 1921 35449 1924
rect 35483 1921 35495 1955
rect 35437 1915 35495 1921
rect 36081 1956 36139 1961
rect 36188 1956 36216 1992
rect 45002 1980 45008 1992
rect 45060 1980 45066 2032
rect 46308 2020 46336 2051
rect 45572 1992 46336 2020
rect 36081 1955 36216 1956
rect 36081 1921 36093 1955
rect 36127 1928 36216 1955
rect 36127 1921 36139 1928
rect 36081 1915 36139 1921
rect 36262 1912 36268 1964
rect 36320 1912 36326 1964
rect 37366 1912 37372 1964
rect 37424 1912 37430 1964
rect 38105 1955 38163 1961
rect 38105 1921 38117 1955
rect 38151 1952 38163 1955
rect 38194 1952 38200 1964
rect 38151 1924 38200 1952
rect 38151 1921 38163 1924
rect 38105 1915 38163 1921
rect 38194 1912 38200 1924
rect 38252 1912 38258 1964
rect 38746 1912 38752 1964
rect 38804 1952 38810 1964
rect 38841 1955 38899 1961
rect 38841 1952 38853 1955
rect 38804 1924 38853 1952
rect 38804 1912 38810 1924
rect 38841 1921 38853 1924
rect 38887 1921 38899 1955
rect 38841 1915 38899 1921
rect 40126 1912 40132 1964
rect 40184 1952 40190 1964
rect 40497 1955 40555 1961
rect 40497 1952 40509 1955
rect 40184 1924 40509 1952
rect 40184 1912 40190 1924
rect 40497 1921 40509 1924
rect 40543 1921 40555 1955
rect 40497 1915 40555 1921
rect 40586 1912 40592 1964
rect 40644 1952 40650 1964
rect 40773 1955 40831 1961
rect 40773 1952 40785 1955
rect 40644 1924 40785 1952
rect 40644 1912 40650 1924
rect 40773 1921 40785 1924
rect 40819 1921 40831 1955
rect 40773 1915 40831 1921
rect 41046 1912 41052 1964
rect 41104 1912 41110 1964
rect 41322 1912 41328 1964
rect 41380 1912 41386 1964
rect 42613 1955 42671 1961
rect 42613 1921 42625 1955
rect 42659 1952 42671 1955
rect 43990 1952 43996 1964
rect 42659 1924 43996 1952
rect 42659 1921 42671 1924
rect 42613 1915 42671 1921
rect 43990 1912 43996 1924
rect 44048 1912 44054 1964
rect 45572 1961 45600 1992
rect 45281 1955 45339 1961
rect 45281 1921 45293 1955
rect 45327 1921 45339 1955
rect 45281 1915 45339 1921
rect 45557 1955 45615 1961
rect 45557 1921 45569 1955
rect 45603 1921 45615 1955
rect 45557 1915 45615 1921
rect 45833 1955 45891 1961
rect 45833 1921 45845 1955
rect 45879 1952 45891 1955
rect 46201 1955 46259 1961
rect 45879 1924 46060 1952
rect 45879 1921 45891 1924
rect 45833 1915 45891 1921
rect 33836 1856 34836 1884
rect 33836 1844 33842 1856
rect 38562 1844 38568 1896
rect 38620 1884 38626 1896
rect 45296 1884 45324 1915
rect 45738 1884 45744 1896
rect 38620 1856 41276 1884
rect 45296 1856 45744 1884
rect 38620 1844 38626 1856
rect 31757 1819 31815 1825
rect 31757 1816 31769 1819
rect 31720 1788 31769 1816
rect 31720 1776 31726 1788
rect 31757 1785 31769 1788
rect 31803 1785 31815 1819
rect 31757 1779 31815 1785
rect 32401 1819 32459 1825
rect 32401 1785 32413 1819
rect 32447 1785 32459 1819
rect 32401 1779 32459 1785
rect 33410 1776 33416 1828
rect 33468 1816 33474 1828
rect 33468 1788 34376 1816
rect 33468 1776 33474 1788
rect 25004 1720 26004 1748
rect 25004 1708 25010 1720
rect 26050 1708 26056 1760
rect 26108 1708 26114 1760
rect 26234 1708 26240 1760
rect 26292 1708 26298 1760
rect 27246 1708 27252 1760
rect 27304 1708 27310 1760
rect 27522 1708 27528 1760
rect 27580 1708 27586 1760
rect 27801 1751 27859 1757
rect 27801 1717 27813 1751
rect 27847 1748 27859 1751
rect 27982 1748 27988 1760
rect 27847 1720 27988 1748
rect 27847 1717 27859 1720
rect 27801 1711 27859 1717
rect 27982 1708 27988 1720
rect 28040 1708 28046 1760
rect 28258 1708 28264 1760
rect 28316 1748 28322 1760
rect 28629 1751 28687 1757
rect 28629 1748 28641 1751
rect 28316 1720 28641 1748
rect 28316 1708 28322 1720
rect 28629 1717 28641 1720
rect 28675 1717 28687 1751
rect 28629 1711 28687 1717
rect 29086 1708 29092 1760
rect 29144 1748 29150 1760
rect 30101 1751 30159 1757
rect 30101 1748 30113 1751
rect 29144 1720 30113 1748
rect 29144 1708 29150 1720
rect 30101 1717 30113 1720
rect 30147 1717 30159 1751
rect 30101 1711 30159 1717
rect 30282 1708 30288 1760
rect 30340 1708 30346 1760
rect 30926 1708 30932 1760
rect 30984 1748 30990 1760
rect 31205 1751 31263 1757
rect 31205 1748 31217 1751
rect 30984 1720 31217 1748
rect 30984 1708 30990 1720
rect 31205 1717 31217 1720
rect 31251 1717 31263 1751
rect 31205 1711 31263 1717
rect 32122 1708 32128 1760
rect 32180 1708 32186 1760
rect 32490 1708 32496 1760
rect 32548 1748 32554 1760
rect 33045 1751 33103 1757
rect 33045 1748 33057 1751
rect 32548 1720 33057 1748
rect 32548 1708 32554 1720
rect 33045 1717 33057 1720
rect 33091 1717 33103 1751
rect 33045 1711 33103 1717
rect 33226 1708 33232 1760
rect 33284 1708 33290 1760
rect 33778 1708 33784 1760
rect 33836 1708 33842 1760
rect 34348 1757 34376 1788
rect 35986 1776 35992 1828
rect 36044 1816 36050 1828
rect 36044 1788 36584 1816
rect 36044 1776 36050 1788
rect 34333 1751 34391 1757
rect 34333 1717 34345 1751
rect 34379 1717 34391 1751
rect 34333 1711 34391 1717
rect 34606 1708 34612 1760
rect 34664 1748 34670 1760
rect 35621 1751 35679 1757
rect 35621 1748 35633 1751
rect 34664 1720 35633 1748
rect 34664 1708 34670 1720
rect 35621 1717 35633 1720
rect 35667 1717 35679 1751
rect 35621 1711 35679 1717
rect 36078 1708 36084 1760
rect 36136 1748 36142 1760
rect 36357 1751 36415 1757
rect 36357 1748 36369 1751
rect 36136 1720 36369 1748
rect 36136 1708 36142 1720
rect 36357 1717 36369 1720
rect 36403 1717 36415 1751
rect 36556 1748 36584 1788
rect 37274 1776 37280 1828
rect 37332 1816 37338 1828
rect 38194 1816 38200 1828
rect 37332 1788 38200 1816
rect 37332 1776 37338 1788
rect 38194 1776 38200 1788
rect 38252 1776 38258 1828
rect 38470 1776 38476 1828
rect 38528 1816 38534 1828
rect 40681 1819 40739 1825
rect 40681 1816 40693 1819
rect 38528 1788 40693 1816
rect 38528 1776 38534 1788
rect 40681 1785 40693 1788
rect 40727 1785 40739 1819
rect 40681 1779 40739 1785
rect 40770 1776 40776 1828
rect 40828 1816 40834 1828
rect 41248 1825 41276 1856
rect 45738 1844 45744 1856
rect 45796 1844 45802 1896
rect 46032 1825 46060 1924
rect 46201 1921 46213 1955
rect 46247 1921 46259 1955
rect 46201 1915 46259 1921
rect 46216 1884 46244 1915
rect 46474 1912 46480 1964
rect 46532 1912 46538 1964
rect 46566 1884 46572 1896
rect 46216 1856 46572 1884
rect 46566 1844 46572 1856
rect 46624 1844 46630 1896
rect 40957 1819 41015 1825
rect 40957 1816 40969 1819
rect 40828 1788 40969 1816
rect 40828 1776 40834 1788
rect 40957 1785 40969 1788
rect 41003 1785 41015 1819
rect 40957 1779 41015 1785
rect 41233 1819 41291 1825
rect 41233 1785 41245 1819
rect 41279 1785 41291 1819
rect 41233 1779 41291 1785
rect 46017 1819 46075 1825
rect 46017 1785 46029 1819
rect 46063 1785 46075 1819
rect 46017 1779 46075 1785
rect 37461 1751 37519 1757
rect 37461 1748 37473 1751
rect 36556 1720 37473 1748
rect 36357 1711 36415 1717
rect 37461 1717 37473 1720
rect 37507 1717 37519 1751
rect 37461 1711 37519 1717
rect 38378 1708 38384 1760
rect 38436 1708 38442 1760
rect 38930 1708 38936 1760
rect 38988 1708 38994 1760
rect 39114 1708 39120 1760
rect 39172 1748 39178 1760
rect 41509 1751 41567 1757
rect 41509 1748 41521 1751
rect 39172 1720 41521 1748
rect 39172 1708 39178 1720
rect 41509 1717 41521 1720
rect 41555 1717 41567 1751
rect 41509 1711 41567 1717
rect 1104 1658 46828 1680
rect 1104 1606 6665 1658
rect 6717 1606 6729 1658
rect 6781 1606 6793 1658
rect 6845 1606 6857 1658
rect 6909 1606 6921 1658
rect 6973 1606 18095 1658
rect 18147 1606 18159 1658
rect 18211 1606 18223 1658
rect 18275 1606 18287 1658
rect 18339 1606 18351 1658
rect 18403 1606 29525 1658
rect 29577 1606 29589 1658
rect 29641 1606 29653 1658
rect 29705 1606 29717 1658
rect 29769 1606 29781 1658
rect 29833 1606 40955 1658
rect 41007 1606 41019 1658
rect 41071 1606 41083 1658
rect 41135 1606 41147 1658
rect 41199 1606 41211 1658
rect 41263 1606 46828 1658
rect 1104 1584 46828 1606
rect 1578 1504 1584 1556
rect 1636 1544 1642 1556
rect 6181 1547 6239 1553
rect 1636 1516 2774 1544
rect 1636 1504 1642 1516
rect 2746 1476 2774 1516
rect 6181 1513 6193 1547
rect 6227 1544 6239 1547
rect 8202 1544 8208 1556
rect 6227 1516 8208 1544
rect 6227 1513 6239 1516
rect 6181 1507 6239 1513
rect 8202 1504 8208 1516
rect 8260 1504 8266 1556
rect 12437 1547 12495 1553
rect 12437 1513 12449 1547
rect 12483 1544 12495 1547
rect 12710 1544 12716 1556
rect 12483 1516 12716 1544
rect 12483 1513 12495 1516
rect 12437 1507 12495 1513
rect 12710 1504 12716 1516
rect 12768 1504 12774 1556
rect 15197 1547 15255 1553
rect 15197 1513 15209 1547
rect 15243 1544 15255 1547
rect 15378 1544 15384 1556
rect 15243 1516 15384 1544
rect 15243 1513 15255 1516
rect 15197 1507 15255 1513
rect 15378 1504 15384 1516
rect 15436 1504 15442 1556
rect 15473 1547 15531 1553
rect 15473 1513 15485 1547
rect 15519 1544 15531 1547
rect 15746 1544 15752 1556
rect 15519 1516 15752 1544
rect 15519 1513 15531 1516
rect 15473 1507 15531 1513
rect 15746 1504 15752 1516
rect 15804 1504 15810 1556
rect 16025 1547 16083 1553
rect 16025 1513 16037 1547
rect 16071 1544 16083 1547
rect 16298 1544 16304 1556
rect 16071 1516 16304 1544
rect 16071 1513 16083 1516
rect 16025 1507 16083 1513
rect 16298 1504 16304 1516
rect 16356 1504 16362 1556
rect 16669 1547 16727 1553
rect 16669 1513 16681 1547
rect 16715 1544 16727 1547
rect 17034 1544 17040 1556
rect 16715 1516 17040 1544
rect 16715 1513 16727 1516
rect 16669 1507 16727 1513
rect 17034 1504 17040 1516
rect 17092 1504 17098 1556
rect 17218 1504 17224 1556
rect 17276 1504 17282 1556
rect 17310 1504 17316 1556
rect 17368 1504 17374 1556
rect 17497 1547 17555 1553
rect 17497 1513 17509 1547
rect 17543 1544 17555 1547
rect 17678 1544 17684 1556
rect 17543 1516 17684 1544
rect 17543 1513 17555 1516
rect 17497 1507 17555 1513
rect 17678 1504 17684 1516
rect 17736 1504 17742 1556
rect 18325 1547 18383 1553
rect 18325 1513 18337 1547
rect 18371 1544 18383 1547
rect 18690 1544 18696 1556
rect 18371 1516 18696 1544
rect 18371 1513 18383 1516
rect 18325 1507 18383 1513
rect 18690 1504 18696 1516
rect 18748 1504 18754 1556
rect 19245 1547 19303 1553
rect 19245 1513 19257 1547
rect 19291 1544 19303 1547
rect 19518 1544 19524 1556
rect 19291 1516 19524 1544
rect 19291 1513 19303 1516
rect 19245 1507 19303 1513
rect 19518 1504 19524 1516
rect 19576 1504 19582 1556
rect 19628 1516 20024 1544
rect 16574 1476 16580 1488
rect 2746 1448 16580 1476
rect 16574 1436 16580 1448
rect 16632 1436 16638 1488
rect 16945 1479 17003 1485
rect 16945 1445 16957 1479
rect 16991 1476 17003 1479
rect 17328 1476 17356 1504
rect 19628 1476 19656 1516
rect 16991 1448 17356 1476
rect 18524 1448 19656 1476
rect 16991 1445 17003 1448
rect 16945 1439 17003 1445
rect 15102 1408 15108 1420
rect 6656 1380 6868 1408
rect 1578 1300 1584 1352
rect 1636 1300 1642 1352
rect 1946 1300 1952 1352
rect 2004 1300 2010 1352
rect 2314 1300 2320 1352
rect 2372 1300 2378 1352
rect 2682 1300 2688 1352
rect 2740 1300 2746 1352
rect 2866 1300 2872 1352
rect 2924 1300 2930 1352
rect 3142 1300 3148 1352
rect 3200 1300 3206 1352
rect 3418 1300 3424 1352
rect 3476 1300 3482 1352
rect 3789 1343 3847 1349
rect 3789 1309 3801 1343
rect 3835 1309 3847 1343
rect 3789 1303 3847 1309
rect 1762 1164 1768 1216
rect 1820 1164 1826 1216
rect 2130 1164 2136 1216
rect 2188 1164 2194 1216
rect 2498 1164 2504 1216
rect 2556 1164 2562 1216
rect 2884 1213 2912 1300
rect 2958 1232 2964 1284
rect 3016 1272 3022 1284
rect 3804 1272 3832 1303
rect 4062 1300 4068 1352
rect 4120 1300 4126 1352
rect 4890 1300 4896 1352
rect 4948 1300 4954 1352
rect 5258 1300 5264 1352
rect 5316 1300 5322 1352
rect 5626 1300 5632 1352
rect 5684 1300 5690 1352
rect 5994 1300 6000 1352
rect 6052 1300 6058 1352
rect 6362 1300 6368 1352
rect 6420 1300 6426 1352
rect 6656 1340 6684 1380
rect 6472 1312 6684 1340
rect 6472 1272 6500 1312
rect 6730 1300 6736 1352
rect 6788 1300 6794 1352
rect 6840 1340 6868 1380
rect 13648 1380 15108 1408
rect 7006 1340 7012 1352
rect 6840 1312 7012 1340
rect 7006 1300 7012 1312
rect 7064 1300 7070 1352
rect 7098 1300 7104 1352
rect 7156 1300 7162 1352
rect 7466 1300 7472 1352
rect 7524 1300 7530 1352
rect 7834 1300 7840 1352
rect 7892 1300 7898 1352
rect 8202 1300 8208 1352
rect 8260 1300 8266 1352
rect 8570 1300 8576 1352
rect 8628 1300 8634 1352
rect 8938 1300 8944 1352
rect 8996 1300 9002 1352
rect 9306 1300 9312 1352
rect 9364 1300 9370 1352
rect 9674 1300 9680 1352
rect 9732 1300 9738 1352
rect 10042 1300 10048 1352
rect 10100 1300 10106 1352
rect 10410 1300 10416 1352
rect 10468 1300 10474 1352
rect 10778 1300 10784 1352
rect 10836 1300 10842 1352
rect 11146 1300 11152 1352
rect 11204 1300 11210 1352
rect 11514 1300 11520 1352
rect 11572 1300 11578 1352
rect 11882 1300 11888 1352
rect 11940 1300 11946 1352
rect 12250 1300 12256 1352
rect 12308 1300 12314 1352
rect 12618 1300 12624 1352
rect 12676 1300 12682 1352
rect 12986 1300 12992 1352
rect 13044 1300 13050 1352
rect 13354 1300 13360 1352
rect 13412 1300 13418 1352
rect 7926 1272 7932 1284
rect 3016 1244 3832 1272
rect 5000 1244 6500 1272
rect 6564 1244 7932 1272
rect 3016 1232 3022 1244
rect 2869 1207 2927 1213
rect 2869 1173 2881 1207
rect 2915 1173 2927 1207
rect 2869 1167 2927 1173
rect 3326 1164 3332 1216
rect 3384 1164 3390 1216
rect 3605 1207 3663 1213
rect 3605 1173 3617 1207
rect 3651 1204 3663 1207
rect 5000 1204 5028 1244
rect 3651 1176 5028 1204
rect 3651 1173 3663 1176
rect 3605 1167 3663 1173
rect 5074 1164 5080 1216
rect 5132 1164 5138 1216
rect 5442 1164 5448 1216
rect 5500 1164 5506 1216
rect 5810 1164 5816 1216
rect 5868 1164 5874 1216
rect 6564 1213 6592 1244
rect 7926 1232 7932 1244
rect 7984 1232 7990 1284
rect 13648 1272 13676 1380
rect 15102 1368 15108 1380
rect 15160 1368 15166 1420
rect 18524 1408 18552 1448
rect 19702 1436 19708 1488
rect 19760 1436 19766 1488
rect 19794 1436 19800 1488
rect 19852 1436 19858 1488
rect 19242 1408 19248 1420
rect 15580 1380 18552 1408
rect 18800 1380 19248 1408
rect 13722 1300 13728 1352
rect 13780 1300 13786 1352
rect 13814 1300 13820 1352
rect 13872 1300 13878 1352
rect 14090 1300 14096 1352
rect 14148 1300 14154 1352
rect 14642 1300 14648 1352
rect 14700 1300 14706 1352
rect 15010 1300 15016 1352
rect 15068 1300 15074 1352
rect 15378 1300 15384 1352
rect 15436 1300 15442 1352
rect 8036 1244 13676 1272
rect 6549 1207 6607 1213
rect 6549 1173 6561 1207
rect 6595 1173 6607 1207
rect 6549 1167 6607 1173
rect 6914 1164 6920 1216
rect 6972 1164 6978 1216
rect 7282 1164 7288 1216
rect 7340 1164 7346 1216
rect 7650 1164 7656 1216
rect 7708 1164 7714 1216
rect 8036 1213 8064 1244
rect 8021 1207 8079 1213
rect 8021 1173 8033 1207
rect 8067 1173 8079 1207
rect 8021 1167 8079 1173
rect 8386 1164 8392 1216
rect 8444 1164 8450 1216
rect 8754 1164 8760 1216
rect 8812 1164 8818 1216
rect 9122 1164 9128 1216
rect 9180 1164 9186 1216
rect 9490 1164 9496 1216
rect 9548 1164 9554 1216
rect 9858 1164 9864 1216
rect 9916 1164 9922 1216
rect 10226 1164 10232 1216
rect 10284 1164 10290 1216
rect 10594 1164 10600 1216
rect 10652 1164 10658 1216
rect 10962 1164 10968 1216
rect 11020 1164 11026 1216
rect 11330 1164 11336 1216
rect 11388 1164 11394 1216
rect 11698 1164 11704 1216
rect 11756 1164 11762 1216
rect 12066 1164 12072 1216
rect 12124 1164 12130 1216
rect 12802 1164 12808 1216
rect 12860 1164 12866 1216
rect 13170 1164 13176 1216
rect 13228 1164 13234 1216
rect 13541 1207 13599 1213
rect 13541 1173 13553 1207
rect 13587 1204 13599 1207
rect 13832 1204 13860 1300
rect 15580 1272 15608 1380
rect 15654 1300 15660 1352
rect 15712 1300 15718 1352
rect 15930 1300 15936 1352
rect 15988 1300 15994 1352
rect 16022 1300 16028 1352
rect 16080 1300 16086 1352
rect 16206 1300 16212 1352
rect 16264 1300 16270 1352
rect 16485 1343 16543 1349
rect 16485 1309 16497 1343
rect 16531 1340 16543 1343
rect 16574 1340 16580 1352
rect 16531 1312 16580 1340
rect 16531 1309 16543 1312
rect 16485 1303 16543 1309
rect 16574 1300 16580 1312
rect 16632 1300 16638 1352
rect 16850 1300 16856 1352
rect 16908 1300 16914 1352
rect 17126 1300 17132 1352
rect 17184 1300 17190 1352
rect 17402 1300 17408 1352
rect 17460 1300 17466 1352
rect 17678 1300 17684 1352
rect 17736 1300 17742 1352
rect 17957 1343 18015 1349
rect 17957 1309 17969 1343
rect 18003 1309 18015 1343
rect 17957 1303 18015 1309
rect 16040 1272 16068 1300
rect 14476 1244 15608 1272
rect 15764 1244 16068 1272
rect 13587 1176 13860 1204
rect 13587 1173 13599 1176
rect 13541 1167 13599 1173
rect 13906 1164 13912 1216
rect 13964 1164 13970 1216
rect 14274 1164 14280 1216
rect 14332 1164 14338 1216
rect 14476 1213 14504 1244
rect 14461 1207 14519 1213
rect 14461 1173 14473 1207
rect 14507 1173 14519 1207
rect 14461 1167 14519 1173
rect 14826 1164 14832 1216
rect 14884 1164 14890 1216
rect 15764 1213 15792 1244
rect 16758 1232 16764 1284
rect 16816 1232 16822 1284
rect 17972 1272 18000 1303
rect 18230 1300 18236 1352
rect 18288 1300 18294 1352
rect 18506 1300 18512 1352
rect 18564 1300 18570 1352
rect 18800 1349 18828 1380
rect 19242 1368 19248 1380
rect 19300 1368 19306 1420
rect 19352 1380 19564 1408
rect 18785 1343 18843 1349
rect 18785 1309 18797 1343
rect 18831 1309 18843 1343
rect 18785 1303 18843 1309
rect 18877 1343 18935 1349
rect 18877 1309 18889 1343
rect 18923 1309 18935 1343
rect 19352 1340 19380 1380
rect 19536 1349 19564 1380
rect 18877 1303 18935 1309
rect 18984 1312 19380 1340
rect 19429 1343 19487 1349
rect 18414 1272 18420 1284
rect 17972 1244 18420 1272
rect 18414 1232 18420 1244
rect 18472 1232 18478 1284
rect 18892 1272 18920 1303
rect 18524 1244 18920 1272
rect 15749 1207 15807 1213
rect 15749 1173 15761 1207
rect 15795 1173 15807 1207
rect 15749 1167 15807 1173
rect 16301 1207 16359 1213
rect 16301 1173 16313 1207
rect 16347 1204 16359 1207
rect 16776 1204 16804 1232
rect 16347 1176 16804 1204
rect 17773 1207 17831 1213
rect 16347 1173 16359 1176
rect 16301 1167 16359 1173
rect 17773 1173 17785 1207
rect 17819 1204 17831 1207
rect 17954 1204 17960 1216
rect 17819 1176 17960 1204
rect 17819 1173 17831 1176
rect 17773 1167 17831 1173
rect 17954 1164 17960 1176
rect 18012 1164 18018 1216
rect 18049 1207 18107 1213
rect 18049 1173 18061 1207
rect 18095 1204 18107 1207
rect 18524 1204 18552 1244
rect 18095 1176 18552 1204
rect 18601 1207 18659 1213
rect 18095 1173 18107 1176
rect 18049 1167 18107 1173
rect 18601 1173 18613 1207
rect 18647 1204 18659 1207
rect 18984 1204 19012 1312
rect 19429 1309 19441 1343
rect 19475 1309 19487 1343
rect 19429 1303 19487 1309
rect 19521 1343 19579 1349
rect 19521 1309 19533 1343
rect 19567 1309 19579 1343
rect 19812 1340 19840 1436
rect 19996 1408 20024 1516
rect 20438 1504 20444 1556
rect 20496 1544 20502 1556
rect 24394 1544 24400 1556
rect 20496 1516 24400 1544
rect 20496 1504 20502 1516
rect 24394 1504 24400 1516
rect 24452 1504 24458 1556
rect 24670 1504 24676 1556
rect 24728 1544 24734 1556
rect 24949 1547 25007 1553
rect 24949 1544 24961 1547
rect 24728 1516 24961 1544
rect 24728 1504 24734 1516
rect 24949 1513 24961 1516
rect 24995 1513 25007 1547
rect 24949 1507 25007 1513
rect 26142 1504 26148 1556
rect 26200 1544 26206 1556
rect 26421 1547 26479 1553
rect 26421 1544 26433 1547
rect 26200 1516 26433 1544
rect 26200 1504 26206 1516
rect 26421 1513 26433 1516
rect 26467 1513 26479 1547
rect 26421 1507 26479 1513
rect 27614 1504 27620 1556
rect 27672 1544 27678 1556
rect 27893 1547 27951 1553
rect 27893 1544 27905 1547
rect 27672 1516 27905 1544
rect 27672 1504 27678 1516
rect 27893 1513 27905 1516
rect 27939 1513 27951 1547
rect 27893 1507 27951 1513
rect 28718 1504 28724 1556
rect 28776 1544 28782 1556
rect 28997 1547 29055 1553
rect 28997 1544 29009 1547
rect 28776 1516 29009 1544
rect 28776 1504 28782 1516
rect 28997 1513 29009 1516
rect 29043 1513 29055 1547
rect 28997 1507 29055 1513
rect 29733 1547 29791 1553
rect 29733 1513 29745 1547
rect 29779 1513 29791 1547
rect 29733 1507 29791 1513
rect 20162 1436 20168 1488
rect 20220 1476 20226 1488
rect 20220 1448 21404 1476
rect 20220 1436 20226 1448
rect 20530 1408 20536 1420
rect 19996 1380 20536 1408
rect 20530 1368 20536 1380
rect 20588 1368 20594 1420
rect 20622 1368 20628 1420
rect 20680 1368 20686 1420
rect 21376 1408 21404 1448
rect 21450 1436 21456 1488
rect 21508 1476 21514 1488
rect 23382 1476 23388 1488
rect 21508 1448 23388 1476
rect 21508 1436 21514 1448
rect 23382 1436 23388 1448
rect 23440 1436 23446 1488
rect 28902 1436 28908 1488
rect 28960 1476 28966 1488
rect 29748 1476 29776 1507
rect 29822 1504 29828 1556
rect 29880 1544 29886 1556
rect 30469 1547 30527 1553
rect 30469 1544 30481 1547
rect 29880 1516 30481 1544
rect 29880 1504 29886 1516
rect 30469 1513 30481 1516
rect 30515 1513 30527 1547
rect 30469 1507 30527 1513
rect 30834 1504 30840 1556
rect 30892 1544 30898 1556
rect 30892 1516 31248 1544
rect 30892 1504 30898 1516
rect 28960 1448 29776 1476
rect 31220 1476 31248 1516
rect 31294 1504 31300 1556
rect 31352 1544 31358 1556
rect 32309 1547 32367 1553
rect 32309 1544 32321 1547
rect 31352 1516 32321 1544
rect 31352 1504 31358 1516
rect 32309 1513 32321 1516
rect 32355 1513 32367 1547
rect 32309 1507 32367 1513
rect 32766 1504 32772 1556
rect 32824 1544 32830 1556
rect 33413 1547 33471 1553
rect 33413 1544 33425 1547
rect 32824 1516 33425 1544
rect 32824 1504 32830 1516
rect 33413 1513 33425 1516
rect 33459 1513 33471 1547
rect 33413 1507 33471 1513
rect 33965 1547 34023 1553
rect 33965 1513 33977 1547
rect 34011 1513 34023 1547
rect 33965 1507 34023 1513
rect 31220 1448 31616 1476
rect 28960 1436 28966 1448
rect 21376 1380 22232 1408
rect 19889 1343 19947 1349
rect 19889 1340 19901 1343
rect 19812 1312 19901 1340
rect 19521 1303 19579 1309
rect 19889 1309 19901 1312
rect 19935 1309 19947 1343
rect 19889 1303 19947 1309
rect 19150 1232 19156 1284
rect 19208 1232 19214 1284
rect 19444 1272 19472 1303
rect 19978 1300 19984 1352
rect 20036 1340 20042 1352
rect 20993 1343 21051 1349
rect 20993 1340 21005 1343
rect 20036 1312 21005 1340
rect 20036 1300 20042 1312
rect 20993 1309 21005 1312
rect 21039 1309 21051 1343
rect 20993 1303 21051 1309
rect 21082 1300 21088 1352
rect 21140 1340 21146 1352
rect 21361 1343 21419 1349
rect 21361 1340 21373 1343
rect 21140 1312 21373 1340
rect 21140 1300 21146 1312
rect 21361 1309 21373 1312
rect 21407 1309 21419 1343
rect 21361 1303 21419 1309
rect 22002 1300 22008 1352
rect 22060 1300 22066 1352
rect 22204 1349 22232 1380
rect 24044 1380 25360 1408
rect 24044 1352 24072 1380
rect 22189 1343 22247 1349
rect 22189 1309 22201 1343
rect 22235 1309 22247 1343
rect 22189 1303 22247 1309
rect 22278 1300 22284 1352
rect 22336 1340 22342 1352
rect 22557 1343 22615 1349
rect 22557 1340 22569 1343
rect 22336 1312 22569 1340
rect 22336 1300 22342 1312
rect 22557 1309 22569 1312
rect 22603 1309 22615 1343
rect 22557 1303 22615 1309
rect 22833 1343 22891 1349
rect 22833 1309 22845 1343
rect 22879 1309 22891 1343
rect 22833 1303 22891 1309
rect 19794 1272 19800 1284
rect 19444 1244 19800 1272
rect 19794 1232 19800 1244
rect 19852 1232 19858 1284
rect 20349 1275 20407 1281
rect 20349 1272 20361 1275
rect 19904 1244 20361 1272
rect 18647 1176 19012 1204
rect 18647 1173 18659 1176
rect 18601 1167 18659 1173
rect 19058 1164 19064 1216
rect 19116 1164 19122 1216
rect 19168 1204 19196 1232
rect 19904 1204 19932 1244
rect 20349 1241 20361 1244
rect 20395 1241 20407 1275
rect 22848 1272 22876 1303
rect 23474 1300 23480 1352
rect 23532 1340 23538 1352
rect 23937 1343 23995 1349
rect 23937 1340 23949 1343
rect 23532 1312 23949 1340
rect 23532 1300 23538 1312
rect 23937 1309 23949 1312
rect 23983 1309 23995 1343
rect 23937 1303 23995 1309
rect 24026 1300 24032 1352
rect 24084 1300 24090 1352
rect 24210 1300 24216 1352
rect 24268 1340 24274 1352
rect 24397 1343 24455 1349
rect 24397 1340 24409 1343
rect 24268 1312 24409 1340
rect 24268 1300 24274 1312
rect 24397 1309 24409 1312
rect 24443 1309 24455 1343
rect 24397 1303 24455 1309
rect 24762 1300 24768 1352
rect 24820 1340 24826 1352
rect 25332 1349 25360 1380
rect 25406 1368 25412 1420
rect 25464 1408 25470 1420
rect 30466 1408 30472 1420
rect 25464 1380 30472 1408
rect 25464 1368 25470 1380
rect 30466 1368 30472 1380
rect 30524 1368 30530 1420
rect 30650 1368 30656 1420
rect 30708 1408 30714 1420
rect 30708 1380 31524 1408
rect 30708 1368 30714 1380
rect 25317 1343 25375 1349
rect 24820 1312 25268 1340
rect 24820 1300 24826 1312
rect 23293 1275 23351 1281
rect 23293 1272 23305 1275
rect 20349 1235 20407 1241
rect 21836 1244 22876 1272
rect 22940 1244 23305 1272
rect 19168 1176 19932 1204
rect 20070 1164 20076 1216
rect 20128 1164 20134 1216
rect 21174 1164 21180 1216
rect 21232 1164 21238 1216
rect 21542 1164 21548 1216
rect 21600 1164 21606 1216
rect 21836 1213 21864 1244
rect 21821 1207 21879 1213
rect 21821 1173 21833 1207
rect 21867 1173 21879 1207
rect 21821 1167 21879 1173
rect 21910 1164 21916 1216
rect 21968 1204 21974 1216
rect 22940 1204 22968 1244
rect 23293 1241 23305 1244
rect 23339 1241 23351 1275
rect 23293 1235 23351 1241
rect 24854 1232 24860 1284
rect 24912 1232 24918 1284
rect 25240 1272 25268 1312
rect 25317 1309 25329 1343
rect 25363 1309 25375 1343
rect 25317 1303 25375 1309
rect 25685 1343 25743 1349
rect 25685 1309 25697 1343
rect 25731 1309 25743 1343
rect 25685 1303 25743 1309
rect 25700 1272 25728 1303
rect 26234 1300 26240 1352
rect 26292 1340 26298 1352
rect 26329 1343 26387 1349
rect 26329 1340 26341 1343
rect 26292 1312 26341 1340
rect 26292 1300 26298 1312
rect 26329 1309 26341 1312
rect 26375 1309 26387 1343
rect 26329 1303 26387 1309
rect 26510 1300 26516 1352
rect 26568 1340 26574 1352
rect 26973 1343 27031 1349
rect 26973 1340 26985 1343
rect 26568 1312 26985 1340
rect 26568 1300 26574 1312
rect 26973 1309 26985 1312
rect 27019 1309 27031 1343
rect 26973 1303 27031 1309
rect 27246 1300 27252 1352
rect 27304 1340 27310 1352
rect 27341 1343 27399 1349
rect 27341 1340 27353 1343
rect 27304 1312 27353 1340
rect 27304 1300 27310 1312
rect 27341 1309 27353 1312
rect 27387 1309 27399 1343
rect 27341 1303 27399 1309
rect 27522 1300 27528 1352
rect 27580 1340 27586 1352
rect 27801 1343 27859 1349
rect 27801 1340 27813 1343
rect 27580 1312 27813 1340
rect 27580 1300 27586 1312
rect 27801 1309 27813 1312
rect 27847 1309 27859 1343
rect 27801 1303 27859 1309
rect 27982 1300 27988 1352
rect 28040 1340 28046 1352
rect 28261 1343 28319 1349
rect 28261 1340 28273 1343
rect 28040 1312 28273 1340
rect 28040 1300 28046 1312
rect 28261 1309 28273 1312
rect 28307 1309 28319 1343
rect 28261 1303 28319 1309
rect 28994 1300 29000 1352
rect 29052 1340 29058 1352
rect 29641 1343 29699 1349
rect 29641 1340 29653 1343
rect 29052 1312 29653 1340
rect 29052 1300 29058 1312
rect 29641 1309 29653 1312
rect 29687 1309 29699 1343
rect 29641 1303 29699 1309
rect 30282 1300 30288 1352
rect 30340 1340 30346 1352
rect 30929 1343 30987 1349
rect 30929 1340 30941 1343
rect 30340 1312 30941 1340
rect 30340 1300 30346 1312
rect 30929 1309 30941 1312
rect 30975 1309 30987 1343
rect 30929 1303 30987 1309
rect 31018 1300 31024 1352
rect 31076 1340 31082 1352
rect 31496 1349 31524 1380
rect 31297 1343 31355 1349
rect 31297 1340 31309 1343
rect 31076 1312 31309 1340
rect 31076 1300 31082 1312
rect 31297 1309 31309 1312
rect 31343 1309 31355 1343
rect 31297 1303 31355 1309
rect 31481 1343 31539 1349
rect 31481 1309 31493 1343
rect 31527 1309 31539 1343
rect 31588 1340 31616 1448
rect 31662 1436 31668 1488
rect 31720 1476 31726 1488
rect 32953 1479 33011 1485
rect 32953 1476 32965 1479
rect 31720 1448 32965 1476
rect 31720 1436 31726 1448
rect 32953 1445 32965 1448
rect 32999 1445 33011 1479
rect 32953 1439 33011 1445
rect 33134 1436 33140 1488
rect 33192 1476 33198 1488
rect 33980 1476 34008 1507
rect 34146 1504 34152 1556
rect 34204 1544 34210 1556
rect 34885 1547 34943 1553
rect 34885 1544 34897 1547
rect 34204 1516 34897 1544
rect 34204 1504 34210 1516
rect 34885 1513 34897 1516
rect 34931 1513 34943 1547
rect 34885 1507 34943 1513
rect 34974 1504 34980 1556
rect 35032 1544 35038 1556
rect 35989 1547 36047 1553
rect 35989 1544 36001 1547
rect 35032 1516 36001 1544
rect 35032 1504 35038 1516
rect 35989 1513 36001 1516
rect 36035 1513 36047 1547
rect 35989 1507 36047 1513
rect 36541 1547 36599 1553
rect 36541 1513 36553 1547
rect 36587 1513 36599 1547
rect 36541 1507 36599 1513
rect 33192 1448 34008 1476
rect 33192 1436 33198 1448
rect 34330 1436 34336 1488
rect 34388 1476 34394 1488
rect 35529 1479 35587 1485
rect 35529 1476 35541 1479
rect 34388 1448 35541 1476
rect 34388 1436 34394 1448
rect 35529 1445 35541 1448
rect 35575 1445 35587 1479
rect 35529 1439 35587 1445
rect 35894 1436 35900 1488
rect 35952 1476 35958 1488
rect 36556 1476 36584 1507
rect 36814 1504 36820 1556
rect 36872 1544 36878 1556
rect 38013 1547 38071 1553
rect 38013 1544 38025 1547
rect 36872 1516 38025 1544
rect 36872 1504 36878 1516
rect 38013 1513 38025 1516
rect 38059 1513 38071 1547
rect 38013 1507 38071 1513
rect 38286 1504 38292 1556
rect 38344 1544 38350 1556
rect 39117 1547 39175 1553
rect 39117 1544 39129 1547
rect 38344 1516 39129 1544
rect 38344 1504 38350 1516
rect 39117 1513 39129 1516
rect 39163 1513 39175 1547
rect 39117 1507 39175 1513
rect 39298 1504 39304 1556
rect 39356 1544 39362 1556
rect 40589 1547 40647 1553
rect 40589 1544 40601 1547
rect 39356 1516 40601 1544
rect 39356 1504 39362 1516
rect 40589 1513 40601 1516
rect 40635 1513 40647 1547
rect 40589 1507 40647 1513
rect 40770 1504 40776 1556
rect 40828 1504 40834 1556
rect 41506 1504 41512 1556
rect 41564 1504 41570 1556
rect 42794 1504 42800 1556
rect 42852 1544 42858 1556
rect 44821 1547 44879 1553
rect 44821 1544 44833 1547
rect 42852 1516 44833 1544
rect 42852 1504 42858 1516
rect 44821 1513 44833 1516
rect 44867 1513 44879 1547
rect 44821 1507 44879 1513
rect 45002 1504 45008 1556
rect 45060 1504 45066 1556
rect 45738 1504 45744 1556
rect 45796 1504 45802 1556
rect 35952 1448 36584 1476
rect 35952 1436 35958 1448
rect 37090 1436 37096 1488
rect 37148 1476 37154 1488
rect 38657 1479 38715 1485
rect 38657 1476 38669 1479
rect 37148 1448 38669 1476
rect 37148 1436 37154 1448
rect 38657 1445 38669 1448
rect 38703 1445 38715 1479
rect 38657 1439 38715 1445
rect 38838 1436 38844 1488
rect 38896 1476 38902 1488
rect 40129 1479 40187 1485
rect 40129 1476 40141 1479
rect 38896 1448 40141 1476
rect 38896 1436 38902 1448
rect 40129 1445 40141 1448
rect 40175 1445 40187 1479
rect 40129 1439 40187 1445
rect 32490 1368 32496 1420
rect 32548 1408 32554 1420
rect 33594 1408 33600 1420
rect 32548 1380 33600 1408
rect 32548 1368 32554 1380
rect 33594 1368 33600 1380
rect 33652 1368 33658 1420
rect 33686 1368 33692 1420
rect 33744 1408 33750 1420
rect 40788 1408 40816 1504
rect 33744 1380 40816 1408
rect 41524 1408 41552 1504
rect 44082 1436 44088 1488
rect 44140 1436 44146 1488
rect 44450 1436 44456 1488
rect 44508 1436 44514 1488
rect 41524 1380 43116 1408
rect 33744 1368 33750 1380
rect 31588 1312 31892 1340
rect 31481 1303 31539 1309
rect 25240 1244 25728 1272
rect 28074 1232 28080 1284
rect 28132 1272 28138 1284
rect 28905 1275 28963 1281
rect 28905 1272 28917 1275
rect 28132 1244 28917 1272
rect 28132 1232 28138 1244
rect 28905 1241 28917 1244
rect 28951 1241 28963 1275
rect 28905 1235 28963 1241
rect 30374 1232 30380 1284
rect 30432 1232 30438 1284
rect 30466 1232 30472 1284
rect 30524 1272 30530 1284
rect 31864 1272 31892 1312
rect 32122 1300 32128 1352
rect 32180 1340 32186 1352
rect 32769 1343 32827 1349
rect 32769 1340 32781 1343
rect 32180 1312 32781 1340
rect 32180 1300 32186 1312
rect 32769 1309 32781 1312
rect 32815 1309 32827 1343
rect 32769 1303 32827 1309
rect 32950 1300 32956 1352
rect 33008 1300 33014 1352
rect 33226 1300 33232 1352
rect 33284 1340 33290 1352
rect 33321 1343 33379 1349
rect 33321 1340 33333 1343
rect 33284 1312 33333 1340
rect 33284 1300 33290 1312
rect 33321 1309 33333 1312
rect 33367 1309 33379 1343
rect 33321 1303 33379 1309
rect 34882 1300 34888 1352
rect 34940 1340 34946 1352
rect 35345 1343 35403 1349
rect 35345 1340 35357 1343
rect 34940 1312 35357 1340
rect 34940 1300 34946 1312
rect 35345 1309 35357 1312
rect 35391 1309 35403 1343
rect 35345 1303 35403 1309
rect 37734 1300 37740 1352
rect 37792 1340 37798 1352
rect 37792 1312 38056 1340
rect 37792 1300 37798 1312
rect 32217 1275 32275 1281
rect 32217 1272 32229 1275
rect 30524 1244 31754 1272
rect 31864 1244 32229 1272
rect 30524 1232 30530 1244
rect 21968 1176 22968 1204
rect 21968 1164 21974 1176
rect 23014 1164 23020 1216
rect 23072 1164 23078 1216
rect 23382 1164 23388 1216
rect 23440 1164 23446 1216
rect 24118 1164 24124 1216
rect 24176 1164 24182 1216
rect 24578 1164 24584 1216
rect 24636 1164 24642 1216
rect 25038 1164 25044 1216
rect 25096 1204 25102 1216
rect 25501 1207 25559 1213
rect 25501 1204 25513 1207
rect 25096 1176 25513 1204
rect 25096 1164 25102 1176
rect 25501 1173 25513 1176
rect 25547 1173 25559 1207
rect 25501 1167 25559 1173
rect 25590 1164 25596 1216
rect 25648 1204 25654 1216
rect 25869 1207 25927 1213
rect 25869 1204 25881 1207
rect 25648 1176 25881 1204
rect 25648 1164 25654 1176
rect 25869 1173 25881 1176
rect 25915 1173 25927 1207
rect 25869 1167 25927 1173
rect 26510 1164 26516 1216
rect 26568 1204 26574 1216
rect 27157 1207 27215 1213
rect 27157 1204 27169 1207
rect 26568 1176 27169 1204
rect 26568 1164 26574 1176
rect 27157 1173 27169 1176
rect 27203 1173 27215 1207
rect 27157 1167 27215 1173
rect 27246 1164 27252 1216
rect 27304 1204 27310 1216
rect 27525 1207 27583 1213
rect 27525 1204 27537 1207
rect 27304 1176 27537 1204
rect 27304 1164 27310 1176
rect 27525 1173 27537 1176
rect 27571 1173 27583 1207
rect 27525 1167 27583 1173
rect 27982 1164 27988 1216
rect 28040 1204 28046 1216
rect 28445 1207 28503 1213
rect 28445 1204 28457 1207
rect 28040 1176 28457 1204
rect 28040 1164 28046 1176
rect 28445 1173 28457 1176
rect 28491 1173 28503 1207
rect 28445 1167 28503 1173
rect 30282 1164 30288 1216
rect 30340 1204 30346 1216
rect 31573 1207 31631 1213
rect 31573 1204 31585 1207
rect 30340 1176 31585 1204
rect 30340 1164 30346 1176
rect 31573 1173 31585 1176
rect 31619 1173 31631 1207
rect 31726 1204 31754 1244
rect 32217 1241 32229 1244
rect 32263 1241 32275 1275
rect 32968 1272 32996 1300
rect 33873 1275 33931 1281
rect 33873 1272 33885 1275
rect 32968 1244 33885 1272
rect 32217 1235 32275 1241
rect 33873 1241 33885 1244
rect 33919 1241 33931 1275
rect 33873 1235 33931 1241
rect 34790 1232 34796 1284
rect 34848 1232 34854 1284
rect 35066 1232 35072 1284
rect 35124 1272 35130 1284
rect 35897 1275 35955 1281
rect 35897 1272 35909 1275
rect 35124 1244 35909 1272
rect 35124 1232 35130 1244
rect 35897 1241 35909 1244
rect 35943 1241 35955 1275
rect 35897 1235 35955 1241
rect 36449 1275 36507 1281
rect 36449 1241 36461 1275
rect 36495 1241 36507 1275
rect 36449 1235 36507 1241
rect 37921 1275 37979 1281
rect 37921 1241 37933 1275
rect 37967 1241 37979 1275
rect 38028 1272 38056 1312
rect 38102 1300 38108 1352
rect 38160 1340 38166 1352
rect 38473 1343 38531 1349
rect 38473 1340 38485 1343
rect 38160 1312 38485 1340
rect 38160 1300 38166 1312
rect 38473 1309 38485 1312
rect 38519 1309 38531 1343
rect 38473 1303 38531 1309
rect 39022 1300 39028 1352
rect 39080 1300 39086 1352
rect 39482 1300 39488 1352
rect 39540 1300 39546 1352
rect 40034 1300 40040 1352
rect 40092 1340 40098 1352
rect 40957 1343 41015 1349
rect 40957 1340 40969 1343
rect 40092 1312 40969 1340
rect 40092 1300 40098 1312
rect 40957 1309 40969 1312
rect 41003 1309 41015 1343
rect 40957 1303 41015 1309
rect 41417 1343 41475 1349
rect 41417 1309 41429 1343
rect 41463 1309 41475 1343
rect 41417 1303 41475 1309
rect 39945 1275 40003 1281
rect 39945 1272 39957 1275
rect 38028 1244 39957 1272
rect 37921 1235 37979 1241
rect 39945 1241 39957 1244
rect 39991 1241 40003 1275
rect 39945 1235 40003 1241
rect 36464 1204 36492 1235
rect 31726 1176 36492 1204
rect 31573 1167 31631 1173
rect 37458 1164 37464 1216
rect 37516 1204 37522 1216
rect 37936 1204 37964 1235
rect 40218 1232 40224 1284
rect 40276 1272 40282 1284
rect 40497 1275 40555 1281
rect 40497 1272 40509 1275
rect 40276 1244 40509 1272
rect 40276 1232 40282 1244
rect 40497 1241 40509 1244
rect 40543 1241 40555 1275
rect 41432 1272 41460 1303
rect 41690 1300 41696 1352
rect 41748 1300 41754 1352
rect 41874 1300 41880 1352
rect 41932 1340 41938 1352
rect 42429 1343 42487 1349
rect 42429 1340 42441 1343
rect 41932 1312 42441 1340
rect 41932 1300 41938 1312
rect 42429 1309 42441 1312
rect 42475 1309 42487 1343
rect 42705 1343 42763 1349
rect 42705 1340 42717 1343
rect 42429 1303 42487 1309
rect 42536 1312 42717 1340
rect 41966 1272 41972 1284
rect 41432 1244 41972 1272
rect 40497 1235 40555 1241
rect 41966 1232 41972 1244
rect 42024 1232 42030 1284
rect 42334 1232 42340 1284
rect 42392 1272 42398 1284
rect 42536 1272 42564 1312
rect 42705 1309 42717 1312
rect 42751 1309 42763 1343
rect 42705 1303 42763 1309
rect 42981 1343 43039 1349
rect 42981 1309 42993 1343
rect 43027 1309 43039 1343
rect 42981 1303 43039 1309
rect 42996 1272 43024 1303
rect 42392 1244 42564 1272
rect 42720 1244 43024 1272
rect 43088 1272 43116 1380
rect 43254 1300 43260 1352
rect 43312 1300 43318 1352
rect 43530 1300 43536 1352
rect 43588 1300 43594 1352
rect 43898 1300 43904 1352
rect 43956 1300 43962 1352
rect 44266 1300 44272 1352
rect 44324 1300 44330 1352
rect 44634 1300 44640 1352
rect 44692 1300 44698 1352
rect 45186 1300 45192 1352
rect 45244 1300 45250 1352
rect 45554 1300 45560 1352
rect 45612 1300 45618 1352
rect 45922 1300 45928 1352
rect 45980 1300 45986 1352
rect 46290 1300 46296 1352
rect 46348 1300 46354 1352
rect 43088 1244 43852 1272
rect 42392 1232 42398 1244
rect 42720 1216 42748 1244
rect 37516 1176 37964 1204
rect 37516 1164 37522 1176
rect 39666 1164 39672 1216
rect 39724 1164 39730 1216
rect 41138 1164 41144 1216
rect 41196 1164 41202 1216
rect 41230 1164 41236 1216
rect 41288 1204 41294 1216
rect 42613 1207 42671 1213
rect 42613 1204 42625 1207
rect 41288 1176 42625 1204
rect 41288 1164 41294 1176
rect 42613 1173 42625 1176
rect 42659 1173 42671 1207
rect 42613 1167 42671 1173
rect 42702 1164 42708 1216
rect 42760 1164 42766 1216
rect 42886 1164 42892 1216
rect 42944 1164 42950 1216
rect 43162 1164 43168 1216
rect 43220 1164 43226 1216
rect 43438 1164 43444 1216
rect 43496 1164 43502 1216
rect 43714 1164 43720 1216
rect 43772 1164 43778 1216
rect 43824 1204 43852 1244
rect 43990 1232 43996 1284
rect 44048 1272 44054 1284
rect 44048 1244 46152 1272
rect 44048 1232 44054 1244
rect 46124 1213 46152 1244
rect 45373 1207 45431 1213
rect 45373 1204 45385 1207
rect 43824 1176 45385 1204
rect 45373 1173 45385 1176
rect 45419 1173 45431 1207
rect 45373 1167 45431 1173
rect 46109 1207 46167 1213
rect 46109 1173 46121 1207
rect 46155 1173 46167 1207
rect 46109 1167 46167 1173
rect 1104 1114 46984 1136
rect 1104 1062 12380 1114
rect 12432 1062 12444 1114
rect 12496 1062 12508 1114
rect 12560 1062 12572 1114
rect 12624 1062 12636 1114
rect 12688 1062 23810 1114
rect 23862 1062 23874 1114
rect 23926 1062 23938 1114
rect 23990 1062 24002 1114
rect 24054 1062 24066 1114
rect 24118 1062 35240 1114
rect 35292 1062 35304 1114
rect 35356 1062 35368 1114
rect 35420 1062 35432 1114
rect 35484 1062 35496 1114
rect 35548 1062 46670 1114
rect 46722 1062 46734 1114
rect 46786 1062 46798 1114
rect 46850 1062 46862 1114
rect 46914 1062 46926 1114
rect 46978 1062 46984 1114
rect 1104 1040 46984 1062
rect 2130 960 2136 1012
rect 2188 1000 2194 1012
rect 2188 972 2774 1000
rect 2188 960 2194 972
rect 2746 728 2774 972
rect 7282 960 7288 1012
rect 7340 1000 7346 1012
rect 15102 1000 15108 1012
rect 7340 972 15108 1000
rect 7340 960 7346 972
rect 15102 960 15108 972
rect 15160 960 15166 1012
rect 15488 972 21496 1000
rect 7926 892 7932 944
rect 7984 932 7990 944
rect 7984 904 10180 932
rect 7984 892 7990 904
rect 3326 824 3332 876
rect 3384 864 3390 876
rect 9766 864 9772 876
rect 3384 836 9772 864
rect 3384 824 3390 836
rect 9766 824 9772 836
rect 9824 824 9830 876
rect 5074 756 5080 808
rect 5132 796 5138 808
rect 8662 796 8668 808
rect 5132 768 8668 796
rect 5132 756 5138 768
rect 8662 756 8668 768
rect 8720 756 8726 808
rect 2746 700 7052 728
rect 2498 552 2504 604
rect 2556 592 2562 604
rect 5534 592 5540 604
rect 2556 564 5540 592
rect 2556 552 2562 564
rect 5534 552 5540 564
rect 5592 552 5598 604
rect 1762 484 1768 536
rect 1820 524 1826 536
rect 5718 524 5724 536
rect 1820 496 5724 524
rect 1820 484 1826 496
rect 5718 484 5724 496
rect 5776 484 5782 536
rect 5810 484 5816 536
rect 5868 484 5874 536
rect 5442 416 5448 468
rect 5500 416 5506 468
rect 5460 116 5488 416
rect 5828 184 5856 484
rect 6914 416 6920 468
rect 6972 416 6978 468
rect 6932 252 6960 416
rect 7024 320 7052 700
rect 7650 688 7656 740
rect 7708 688 7714 740
rect 10152 728 10180 904
rect 11330 892 11336 944
rect 11388 892 11394 944
rect 11698 892 11704 944
rect 11756 932 11762 944
rect 15488 932 15516 972
rect 11756 904 15516 932
rect 11756 892 11762 904
rect 17494 892 17500 944
rect 17552 932 17558 944
rect 17552 904 19334 932
rect 17552 892 17558 904
rect 11348 796 11376 892
rect 17218 824 17224 876
rect 17276 864 17282 876
rect 18966 864 18972 876
rect 17276 836 18972 864
rect 17276 824 17282 836
rect 18966 824 18972 836
rect 19024 824 19030 876
rect 11348 768 17356 796
rect 17218 728 17224 740
rect 10152 700 17224 728
rect 17218 688 17224 700
rect 17276 688 17282 740
rect 17328 728 17356 768
rect 18506 756 18512 808
rect 18564 796 18570 808
rect 19150 796 19156 808
rect 18564 768 19156 796
rect 18564 756 18570 768
rect 19150 756 19156 768
rect 19208 756 19214 808
rect 19306 796 19334 904
rect 19426 892 19432 944
rect 19484 892 19490 944
rect 19444 864 19472 892
rect 20530 864 20536 876
rect 19444 836 20536 864
rect 20530 824 20536 836
rect 20588 824 20594 876
rect 21468 864 21496 972
rect 21818 960 21824 1012
rect 21876 1000 21882 1012
rect 30466 1000 30472 1012
rect 21876 972 30472 1000
rect 21876 960 21882 972
rect 30466 960 30472 972
rect 30524 960 30530 1012
rect 31110 960 31116 1012
rect 31168 1000 31174 1012
rect 41230 1000 41236 1012
rect 31168 972 41236 1000
rect 31168 960 31174 972
rect 41230 960 41236 972
rect 41288 960 41294 1012
rect 44082 960 44088 1012
rect 44140 960 44146 1012
rect 24302 892 24308 944
rect 24360 932 24366 944
rect 34790 932 34796 944
rect 24360 904 34796 932
rect 24360 892 24366 904
rect 34790 892 34796 904
rect 34848 892 34854 944
rect 35066 892 35072 944
rect 35124 892 35130 944
rect 39666 892 39672 944
rect 39724 892 39730 944
rect 21468 836 28672 864
rect 28534 796 28540 808
rect 19306 768 28540 796
rect 28534 756 28540 768
rect 28592 756 28598 808
rect 28350 728 28356 740
rect 17328 700 28356 728
rect 28350 688 28356 700
rect 28408 688 28414 740
rect 28644 728 28672 836
rect 28994 824 29000 876
rect 29052 864 29058 876
rect 35084 864 35112 892
rect 29052 836 35112 864
rect 29052 824 29058 836
rect 29270 756 29276 808
rect 29328 796 29334 808
rect 39684 796 39712 892
rect 29328 768 39712 796
rect 29328 756 29334 768
rect 30098 728 30104 740
rect 28644 700 30104 728
rect 30098 688 30104 700
rect 30156 688 30162 740
rect 30834 688 30840 740
rect 30892 728 30898 740
rect 31570 728 31576 740
rect 30892 700 31576 728
rect 30892 688 30898 700
rect 31570 688 31576 700
rect 31628 688 31634 740
rect 33962 688 33968 740
rect 34020 728 34026 740
rect 37458 728 37464 740
rect 34020 700 37464 728
rect 34020 688 34026 700
rect 37458 688 37464 700
rect 37516 688 37522 740
rect 7668 592 7696 688
rect 10226 620 10232 672
rect 10284 660 10290 672
rect 32214 660 32220 672
rect 10284 632 32220 660
rect 10284 620 10290 632
rect 32214 620 32220 632
rect 32272 620 32278 672
rect 44100 660 44128 960
rect 42996 632 44128 660
rect 14734 592 14740 604
rect 7668 564 14740 592
rect 14734 552 14740 564
rect 14792 552 14798 604
rect 32582 592 32588 604
rect 17236 564 32588 592
rect 8386 484 8392 536
rect 8444 484 8450 536
rect 9858 484 9864 536
rect 9916 524 9922 536
rect 17236 524 17264 564
rect 32582 552 32588 564
rect 32640 552 32646 604
rect 42886 592 42892 604
rect 41386 564 42892 592
rect 9916 496 17264 524
rect 9916 484 9922 496
rect 18230 484 18236 536
rect 18288 524 18294 536
rect 18782 524 18788 536
rect 18288 496 18788 524
rect 18288 484 18294 496
rect 18782 484 18788 496
rect 18840 484 18846 536
rect 20530 484 20536 536
rect 20588 524 20594 536
rect 41386 524 41414 564
rect 42886 552 42892 564
rect 42944 552 42950 604
rect 20588 496 41414 524
rect 20588 484 20594 496
rect 8404 388 8432 484
rect 13906 416 13912 468
rect 13964 456 13970 468
rect 27338 456 27344 468
rect 13964 428 27344 456
rect 13964 416 13970 428
rect 27338 416 27344 428
rect 27396 416 27402 468
rect 29362 416 29368 468
rect 29420 456 29426 468
rect 41138 456 41144 468
rect 29420 428 41144 456
rect 29420 416 29426 428
rect 41138 416 41144 428
rect 41196 416 41202 468
rect 13630 388 13636 400
rect 8404 360 13636 388
rect 13630 348 13636 360
rect 13688 348 13694 400
rect 14274 348 14280 400
rect 14332 388 14338 400
rect 28166 388 28172 400
rect 14332 360 28172 388
rect 14332 348 14338 360
rect 28166 348 28172 360
rect 28224 348 28230 400
rect 28350 348 28356 400
rect 28408 388 28414 400
rect 30558 388 30564 400
rect 28408 360 30564 388
rect 28408 348 28414 360
rect 30558 348 30564 360
rect 30616 348 30622 400
rect 30742 348 30748 400
rect 30800 388 30806 400
rect 42996 388 43024 632
rect 43438 552 43444 604
rect 43496 552 43502 604
rect 43714 552 43720 604
rect 43772 552 43778 604
rect 30800 360 43024 388
rect 30800 348 30806 360
rect 11238 320 11244 332
rect 7024 292 11244 320
rect 11238 280 11244 292
rect 11296 280 11302 332
rect 14550 320 14556 332
rect 11348 292 14556 320
rect 11348 252 11376 292
rect 14550 280 14556 292
rect 14608 280 14614 332
rect 14826 280 14832 332
rect 14884 320 14890 332
rect 20346 320 20352 332
rect 14884 292 20352 320
rect 14884 280 14890 292
rect 20346 280 20352 292
rect 20404 280 20410 332
rect 25682 280 25688 332
rect 25740 320 25746 332
rect 43456 320 43484 552
rect 25740 292 43484 320
rect 25740 280 25746 292
rect 12618 252 12624 264
rect 6932 224 11376 252
rect 12406 224 12624 252
rect 12406 184 12434 224
rect 12618 212 12624 224
rect 12676 212 12682 264
rect 12802 212 12808 264
rect 12860 252 12866 264
rect 12860 224 22094 252
rect 12860 212 12866 224
rect 5828 156 12434 184
rect 22066 184 22094 224
rect 27798 212 27804 264
rect 27856 252 27862 264
rect 43732 252 43760 552
rect 27856 224 43760 252
rect 27856 212 27862 224
rect 29914 184 29920 196
rect 22066 156 29920 184
rect 29914 144 29920 156
rect 29972 144 29978 196
rect 30098 144 30104 196
rect 30156 184 30162 196
rect 31018 184 31024 196
rect 30156 156 31024 184
rect 30156 144 30162 156
rect 31018 144 31024 156
rect 31076 144 31082 196
rect 40218 184 40224 196
rect 31726 156 40224 184
rect 13446 116 13452 128
rect 5460 88 13452 116
rect 13446 76 13452 88
rect 13504 76 13510 128
rect 26786 76 26792 128
rect 26844 116 26850 128
rect 31726 116 31754 156
rect 40218 144 40224 156
rect 40276 144 40282 196
rect 26844 88 31754 116
rect 26844 76 26850 88
<< via1 >>
rect 23480 8984 23532 9036
rect 12992 8916 13044 8968
rect 22192 8916 22244 8968
rect 25320 8848 25372 8900
rect 6368 8780 6420 8832
rect 6460 8780 6512 8832
rect 6552 8780 6604 8832
rect 29184 8780 29236 8832
rect 12380 8678 12432 8730
rect 12444 8678 12496 8730
rect 12508 8678 12560 8730
rect 12572 8678 12624 8730
rect 12636 8678 12688 8730
rect 23810 8678 23862 8730
rect 23874 8678 23926 8730
rect 23938 8678 23990 8730
rect 24002 8678 24054 8730
rect 24066 8678 24118 8730
rect 35240 8678 35292 8730
rect 35304 8678 35356 8730
rect 35368 8678 35420 8730
rect 35432 8678 35484 8730
rect 35496 8678 35548 8730
rect 46670 8678 46722 8730
rect 46734 8678 46786 8730
rect 46798 8678 46850 8730
rect 46862 8678 46914 8730
rect 46926 8678 46978 8730
rect 1860 8576 1912 8628
rect 4068 8576 4120 8628
rect 6276 8576 6328 8628
rect 8484 8576 8536 8628
rect 10692 8576 10744 8628
rect 12900 8576 12952 8628
rect 15108 8576 15160 8628
rect 17316 8576 17368 8628
rect 19524 8576 19576 8628
rect 21732 8576 21784 8628
rect 24216 8576 24268 8628
rect 26148 8576 26200 8628
rect 28356 8576 28408 8628
rect 30564 8576 30616 8628
rect 32772 8576 32824 8628
rect 34980 8576 35032 8628
rect 37188 8576 37240 8628
rect 39396 8576 39448 8628
rect 41604 8576 41656 8628
rect 43812 8576 43864 8628
rect 46020 8576 46072 8628
rect 6460 8508 6512 8560
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 24308 8508 24360 8560
rect 6552 8372 6604 8424
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 22100 8440 22152 8492
rect 24860 8440 24912 8492
rect 26516 8440 26568 8492
rect 28448 8483 28500 8492
rect 28448 8449 28457 8483
rect 28457 8449 28491 8483
rect 28491 8449 28500 8483
rect 28448 8440 28500 8449
rect 30656 8483 30708 8492
rect 30656 8449 30665 8483
rect 30665 8449 30699 8483
rect 30699 8449 30708 8483
rect 30656 8440 30708 8449
rect 33140 8440 33192 8492
rect 35072 8483 35124 8492
rect 35072 8449 35081 8483
rect 35081 8449 35115 8483
rect 35115 8449 35124 8483
rect 35072 8440 35124 8449
rect 37372 8483 37424 8492
rect 37372 8449 37381 8483
rect 37381 8449 37415 8483
rect 37415 8449 37424 8483
rect 37372 8440 37424 8449
rect 21272 8372 21324 8424
rect 41696 8483 41748 8492
rect 41696 8449 41705 8483
rect 41705 8449 41739 8483
rect 41739 8449 41748 8483
rect 41696 8440 41748 8449
rect 45008 8440 45060 8492
rect 46112 8483 46164 8492
rect 46112 8449 46121 8483
rect 46121 8449 46155 8483
rect 46155 8449 46164 8483
rect 46112 8440 46164 8449
rect 44732 8372 44784 8424
rect 24676 8304 24728 8356
rect 6665 8134 6717 8186
rect 6729 8134 6781 8186
rect 6793 8134 6845 8186
rect 6857 8134 6909 8186
rect 6921 8134 6973 8186
rect 18095 8134 18147 8186
rect 18159 8134 18211 8186
rect 18223 8134 18275 8186
rect 18287 8134 18339 8186
rect 18351 8134 18403 8186
rect 29525 8134 29577 8186
rect 29589 8134 29641 8186
rect 29653 8134 29705 8186
rect 29717 8134 29769 8186
rect 29781 8134 29833 8186
rect 40955 8134 41007 8186
rect 41019 8134 41071 8186
rect 41083 8134 41135 8186
rect 41147 8134 41199 8186
rect 41211 8134 41263 8186
rect 12380 7590 12432 7642
rect 12444 7590 12496 7642
rect 12508 7590 12560 7642
rect 12572 7590 12624 7642
rect 12636 7590 12688 7642
rect 23810 7590 23862 7642
rect 23874 7590 23926 7642
rect 23938 7590 23990 7642
rect 24002 7590 24054 7642
rect 24066 7590 24118 7642
rect 35240 7590 35292 7642
rect 35304 7590 35356 7642
rect 35368 7590 35420 7642
rect 35432 7590 35484 7642
rect 35496 7590 35548 7642
rect 46670 7590 46722 7642
rect 46734 7590 46786 7642
rect 46798 7590 46850 7642
rect 46862 7590 46914 7642
rect 46926 7590 46978 7642
rect 6665 7046 6717 7098
rect 6729 7046 6781 7098
rect 6793 7046 6845 7098
rect 6857 7046 6909 7098
rect 6921 7046 6973 7098
rect 18095 7046 18147 7098
rect 18159 7046 18211 7098
rect 18223 7046 18275 7098
rect 18287 7046 18339 7098
rect 18351 7046 18403 7098
rect 29525 7046 29577 7098
rect 29589 7046 29641 7098
rect 29653 7046 29705 7098
rect 29717 7046 29769 7098
rect 29781 7046 29833 7098
rect 40955 7046 41007 7098
rect 41019 7046 41071 7098
rect 41083 7046 41135 7098
rect 41147 7046 41199 7098
rect 41211 7046 41263 7098
rect 12380 6502 12432 6554
rect 12444 6502 12496 6554
rect 12508 6502 12560 6554
rect 12572 6502 12624 6554
rect 12636 6502 12688 6554
rect 23810 6502 23862 6554
rect 23874 6502 23926 6554
rect 23938 6502 23990 6554
rect 24002 6502 24054 6554
rect 24066 6502 24118 6554
rect 35240 6502 35292 6554
rect 35304 6502 35356 6554
rect 35368 6502 35420 6554
rect 35432 6502 35484 6554
rect 35496 6502 35548 6554
rect 46670 6502 46722 6554
rect 46734 6502 46786 6554
rect 46798 6502 46850 6554
rect 46862 6502 46914 6554
rect 46926 6502 46978 6554
rect 6665 5958 6717 6010
rect 6729 5958 6781 6010
rect 6793 5958 6845 6010
rect 6857 5958 6909 6010
rect 6921 5958 6973 6010
rect 18095 5958 18147 6010
rect 18159 5958 18211 6010
rect 18223 5958 18275 6010
rect 18287 5958 18339 6010
rect 18351 5958 18403 6010
rect 29525 5958 29577 6010
rect 29589 5958 29641 6010
rect 29653 5958 29705 6010
rect 29717 5958 29769 6010
rect 29781 5958 29833 6010
rect 40955 5958 41007 6010
rect 41019 5958 41071 6010
rect 41083 5958 41135 6010
rect 41147 5958 41199 6010
rect 41211 5958 41263 6010
rect 12380 5414 12432 5466
rect 12444 5414 12496 5466
rect 12508 5414 12560 5466
rect 12572 5414 12624 5466
rect 12636 5414 12688 5466
rect 23810 5414 23862 5466
rect 23874 5414 23926 5466
rect 23938 5414 23990 5466
rect 24002 5414 24054 5466
rect 24066 5414 24118 5466
rect 35240 5414 35292 5466
rect 35304 5414 35356 5466
rect 35368 5414 35420 5466
rect 35432 5414 35484 5466
rect 35496 5414 35548 5466
rect 46670 5414 46722 5466
rect 46734 5414 46786 5466
rect 46798 5414 46850 5466
rect 46862 5414 46914 5466
rect 46926 5414 46978 5466
rect 6665 4870 6717 4922
rect 6729 4870 6781 4922
rect 6793 4870 6845 4922
rect 6857 4870 6909 4922
rect 6921 4870 6973 4922
rect 18095 4870 18147 4922
rect 18159 4870 18211 4922
rect 18223 4870 18275 4922
rect 18287 4870 18339 4922
rect 18351 4870 18403 4922
rect 29525 4870 29577 4922
rect 29589 4870 29641 4922
rect 29653 4870 29705 4922
rect 29717 4870 29769 4922
rect 29781 4870 29833 4922
rect 40955 4870 41007 4922
rect 41019 4870 41071 4922
rect 41083 4870 41135 4922
rect 41147 4870 41199 4922
rect 41211 4870 41263 4922
rect 7012 4496 7064 4548
rect 26424 4496 26476 4548
rect 16948 4428 17000 4480
rect 38108 4428 38160 4480
rect 12380 4326 12432 4378
rect 12444 4326 12496 4378
rect 12508 4326 12560 4378
rect 12572 4326 12624 4378
rect 12636 4326 12688 4378
rect 23810 4326 23862 4378
rect 23874 4326 23926 4378
rect 23938 4326 23990 4378
rect 24002 4326 24054 4378
rect 24066 4326 24118 4378
rect 35240 4326 35292 4378
rect 35304 4326 35356 4378
rect 35368 4326 35420 4378
rect 35432 4326 35484 4378
rect 35496 4326 35548 4378
rect 46670 4326 46722 4378
rect 46734 4326 46786 4378
rect 46798 4326 46850 4378
rect 46862 4326 46914 4378
rect 46926 4326 46978 4378
rect 3976 4224 4028 4276
rect 27436 4224 27488 4276
rect 2872 4156 2924 4208
rect 27712 4156 27764 4208
rect 6665 3782 6717 3834
rect 6729 3782 6781 3834
rect 6793 3782 6845 3834
rect 6857 3782 6909 3834
rect 6921 3782 6973 3834
rect 18095 3782 18147 3834
rect 18159 3782 18211 3834
rect 18223 3782 18275 3834
rect 18287 3782 18339 3834
rect 18351 3782 18403 3834
rect 29525 3782 29577 3834
rect 29589 3782 29641 3834
rect 29653 3782 29705 3834
rect 29717 3782 29769 3834
rect 29781 3782 29833 3834
rect 40955 3782 41007 3834
rect 41019 3782 41071 3834
rect 41083 3782 41135 3834
rect 41147 3782 41199 3834
rect 41211 3782 41263 3834
rect 13452 3476 13504 3528
rect 21732 3476 21784 3528
rect 12716 3408 12768 3460
rect 29368 3408 29420 3460
rect 15200 3340 15252 3392
rect 25228 3340 25280 3392
rect 12380 3238 12432 3290
rect 12444 3238 12496 3290
rect 12508 3238 12560 3290
rect 12572 3238 12624 3290
rect 12636 3238 12688 3290
rect 23810 3238 23862 3290
rect 23874 3238 23926 3290
rect 23938 3238 23990 3290
rect 24002 3238 24054 3290
rect 24066 3238 24118 3290
rect 35240 3238 35292 3290
rect 35304 3238 35356 3290
rect 35368 3238 35420 3290
rect 35432 3238 35484 3290
rect 35496 3238 35548 3290
rect 46670 3238 46722 3290
rect 46734 3238 46786 3290
rect 46798 3238 46850 3290
rect 46862 3238 46914 3290
rect 46926 3238 46978 3290
rect 8760 3136 8812 3188
rect 28172 3136 28224 3188
rect 5540 3068 5592 3120
rect 19984 3068 20036 3120
rect 21640 3068 21692 3120
rect 31116 3068 31168 3120
rect 17500 3000 17552 3052
rect 33968 3000 34020 3052
rect 19340 2932 19392 2984
rect 20076 2932 20128 2984
rect 5724 2864 5776 2916
rect 20352 2864 20404 2916
rect 20628 2864 20680 2916
rect 37832 2864 37884 2916
rect 9588 2796 9640 2848
rect 9680 2796 9732 2848
rect 17132 2796 17184 2848
rect 24768 2796 24820 2848
rect 32128 2796 32180 2848
rect 38568 2796 38620 2848
rect 6665 2694 6717 2746
rect 6729 2694 6781 2746
rect 6793 2694 6845 2746
rect 6857 2694 6909 2746
rect 6921 2694 6973 2746
rect 18095 2694 18147 2746
rect 18159 2694 18211 2746
rect 18223 2694 18275 2746
rect 18287 2694 18339 2746
rect 18351 2694 18403 2746
rect 29525 2694 29577 2746
rect 29589 2694 29641 2746
rect 29653 2694 29705 2746
rect 29717 2694 29769 2746
rect 29781 2694 29833 2746
rect 40955 2694 41007 2746
rect 41019 2694 41071 2746
rect 41083 2694 41135 2746
rect 41147 2694 41199 2746
rect 41211 2694 41263 2746
rect 17408 2592 17460 2644
rect 19524 2592 19576 2644
rect 19616 2592 19668 2644
rect 8208 2524 8260 2576
rect 20628 2635 20680 2644
rect 20628 2601 20637 2635
rect 20637 2601 20671 2635
rect 20671 2601 20680 2635
rect 20628 2592 20680 2601
rect 21272 2635 21324 2644
rect 21272 2601 21281 2635
rect 21281 2601 21315 2635
rect 21315 2601 21324 2635
rect 21272 2592 21324 2601
rect 22100 2635 22152 2644
rect 22100 2601 22109 2635
rect 22109 2601 22143 2635
rect 22143 2601 22152 2635
rect 22100 2592 22152 2601
rect 22192 2592 22244 2644
rect 23480 2592 23532 2644
rect 24308 2592 24360 2644
rect 24860 2635 24912 2644
rect 24860 2601 24869 2635
rect 24869 2601 24903 2635
rect 24903 2601 24912 2635
rect 24860 2592 24912 2601
rect 25320 2635 25372 2644
rect 25320 2601 25329 2635
rect 25329 2601 25363 2635
rect 25363 2601 25372 2635
rect 25320 2592 25372 2601
rect 26516 2635 26568 2644
rect 26516 2601 26525 2635
rect 26525 2601 26559 2635
rect 26559 2601 26568 2635
rect 26516 2592 26568 2601
rect 21548 2524 21600 2576
rect 24676 2524 24728 2576
rect 15384 2456 15436 2508
rect 17960 2431 18012 2440
rect 17960 2397 17969 2431
rect 17969 2397 18003 2431
rect 18003 2397 18012 2431
rect 17960 2388 18012 2397
rect 19984 2388 20036 2440
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 20352 2431 20404 2440
rect 20352 2397 20361 2431
rect 20361 2397 20395 2431
rect 20395 2397 20404 2431
rect 20352 2388 20404 2397
rect 20628 2456 20680 2508
rect 15108 2320 15160 2372
rect 19892 2320 19944 2372
rect 13636 2252 13688 2304
rect 20444 2252 20496 2304
rect 21088 2252 21140 2304
rect 21640 2431 21692 2440
rect 21640 2397 21649 2431
rect 21649 2397 21683 2431
rect 21683 2397 21692 2431
rect 21640 2388 21692 2397
rect 21732 2320 21784 2372
rect 21548 2252 21600 2304
rect 22376 2252 22428 2304
rect 22560 2252 22612 2304
rect 22836 2431 22888 2440
rect 22836 2397 22845 2431
rect 22845 2397 22879 2431
rect 22879 2397 22888 2431
rect 22836 2388 22888 2397
rect 23388 2431 23440 2440
rect 23388 2397 23397 2431
rect 23397 2397 23431 2431
rect 23431 2397 23440 2431
rect 23388 2388 23440 2397
rect 23572 2431 23624 2440
rect 23572 2397 23581 2431
rect 23581 2397 23615 2431
rect 23615 2397 23624 2431
rect 23572 2388 23624 2397
rect 24308 2388 24360 2440
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 25044 2431 25096 2440
rect 25044 2397 25053 2431
rect 25053 2397 25087 2431
rect 25087 2397 25096 2431
rect 25044 2388 25096 2397
rect 24952 2320 25004 2372
rect 24216 2252 24268 2304
rect 24492 2252 24544 2304
rect 25872 2388 25924 2440
rect 25964 2431 26016 2440
rect 25964 2397 25973 2431
rect 25973 2397 26007 2431
rect 26007 2397 26016 2431
rect 25964 2388 26016 2397
rect 27344 2431 27396 2440
rect 27344 2397 27353 2431
rect 27353 2397 27387 2431
rect 27387 2397 27396 2431
rect 27344 2388 27396 2397
rect 27804 2388 27856 2440
rect 26976 2320 27028 2372
rect 28448 2592 28500 2644
rect 28908 2592 28960 2644
rect 30932 2592 30984 2644
rect 35072 2592 35124 2644
rect 37372 2592 37424 2644
rect 31024 2567 31076 2576
rect 31024 2533 31033 2567
rect 31033 2533 31067 2567
rect 31067 2533 31076 2567
rect 31024 2524 31076 2533
rect 31208 2524 31260 2576
rect 30840 2456 30892 2508
rect 28264 2431 28316 2440
rect 28264 2397 28273 2431
rect 28273 2397 28307 2431
rect 28307 2397 28316 2431
rect 28264 2388 28316 2397
rect 28540 2431 28592 2440
rect 28540 2397 28549 2431
rect 28549 2397 28583 2431
rect 28583 2397 28592 2431
rect 28540 2388 28592 2397
rect 30012 2388 30064 2440
rect 30104 2388 30156 2440
rect 30380 2388 30432 2440
rect 30748 2388 30800 2440
rect 31024 2320 31076 2372
rect 31484 2431 31536 2440
rect 31484 2397 31493 2431
rect 31493 2397 31527 2431
rect 31527 2397 31536 2431
rect 31484 2388 31536 2397
rect 36084 2456 36136 2508
rect 32864 2431 32916 2440
rect 32864 2397 32873 2431
rect 32873 2397 32907 2431
rect 32907 2397 32916 2431
rect 32864 2388 32916 2397
rect 33324 2431 33376 2440
rect 33324 2397 33333 2431
rect 33333 2397 33367 2431
rect 33367 2397 33376 2431
rect 33324 2388 33376 2397
rect 35900 2388 35952 2440
rect 26516 2252 26568 2304
rect 27160 2295 27212 2304
rect 27160 2261 27169 2295
rect 27169 2261 27203 2295
rect 27203 2261 27212 2295
rect 27160 2252 27212 2261
rect 28080 2295 28132 2304
rect 28080 2261 28089 2295
rect 28089 2261 28123 2295
rect 28123 2261 28132 2295
rect 28080 2252 28132 2261
rect 29000 2252 29052 2304
rect 30656 2252 30708 2304
rect 31576 2252 31628 2304
rect 32956 2252 33008 2304
rect 33140 2295 33192 2304
rect 33140 2261 33149 2295
rect 33149 2261 33183 2295
rect 33183 2261 33192 2295
rect 33140 2252 33192 2261
rect 41512 2524 41564 2576
rect 41696 2592 41748 2644
rect 44732 2635 44784 2644
rect 44732 2601 44741 2635
rect 44741 2601 44775 2635
rect 44775 2601 44784 2635
rect 44732 2592 44784 2601
rect 45008 2635 45060 2644
rect 45008 2601 45017 2635
rect 45017 2601 45051 2635
rect 45051 2601 45060 2635
rect 45008 2592 45060 2601
rect 46112 2592 46164 2644
rect 44456 2524 44508 2576
rect 42248 2431 42300 2440
rect 42248 2397 42257 2431
rect 42257 2397 42291 2431
rect 42291 2397 42300 2431
rect 42248 2388 42300 2397
rect 44548 2431 44600 2440
rect 44548 2397 44557 2431
rect 44557 2397 44591 2431
rect 44591 2397 44600 2431
rect 44548 2388 44600 2397
rect 45192 2431 45244 2440
rect 45192 2397 45201 2431
rect 45201 2397 45235 2431
rect 45235 2397 45244 2431
rect 45192 2388 45244 2397
rect 45836 2431 45888 2440
rect 45836 2397 45845 2431
rect 45845 2397 45879 2431
rect 45879 2397 45888 2431
rect 45836 2388 45888 2397
rect 38016 2252 38068 2304
rect 38660 2252 38712 2304
rect 42800 2320 42852 2372
rect 12380 2150 12432 2202
rect 12444 2150 12496 2202
rect 12508 2150 12560 2202
rect 12572 2150 12624 2202
rect 12636 2150 12688 2202
rect 23810 2150 23862 2202
rect 23874 2150 23926 2202
rect 23938 2150 23990 2202
rect 24002 2150 24054 2202
rect 24066 2150 24118 2202
rect 35240 2150 35292 2202
rect 35304 2150 35356 2202
rect 35368 2150 35420 2202
rect 35432 2150 35484 2202
rect 35496 2150 35548 2202
rect 46670 2150 46722 2202
rect 46734 2150 46786 2202
rect 46798 2150 46850 2202
rect 46862 2150 46914 2202
rect 46926 2150 46978 2202
rect 15200 2048 15252 2100
rect 15936 2091 15988 2100
rect 15936 2057 15945 2091
rect 15945 2057 15979 2091
rect 15979 2057 15988 2091
rect 15936 2048 15988 2057
rect 16488 2091 16540 2100
rect 16488 2057 16497 2091
rect 16497 2057 16531 2091
rect 16531 2057 16540 2091
rect 16488 2048 16540 2057
rect 16948 2091 17000 2100
rect 16948 2057 16957 2091
rect 16957 2057 16991 2091
rect 16991 2057 17000 2091
rect 16948 2048 17000 2057
rect 17316 2048 17368 2100
rect 17960 2048 18012 2100
rect 17224 1980 17276 2032
rect 18880 2091 18932 2100
rect 18880 2057 18889 2091
rect 18889 2057 18923 2091
rect 18923 2057 18932 2091
rect 18880 2048 18932 2057
rect 19432 2048 19484 2100
rect 19984 2048 20036 2100
rect 20168 2048 20220 2100
rect 20536 2091 20588 2100
rect 20536 2057 20545 2091
rect 20545 2057 20579 2091
rect 20579 2057 20588 2091
rect 20536 2048 20588 2057
rect 1124 1912 1176 1964
rect 3976 1912 4028 1964
rect 4528 1955 4580 1964
rect 4528 1921 4537 1955
rect 4537 1921 4571 1955
rect 4571 1921 4580 1955
rect 4528 1912 4580 1921
rect 15752 1955 15804 1964
rect 15752 1921 15761 1955
rect 15761 1921 15795 1955
rect 15795 1921 15804 1955
rect 15752 1912 15804 1921
rect 16028 1955 16080 1964
rect 16028 1921 16037 1955
rect 16037 1921 16071 1955
rect 16071 1921 16080 1955
rect 16028 1912 16080 1921
rect 16304 1955 16356 1964
rect 16304 1921 16313 1955
rect 16313 1921 16347 1955
rect 16347 1921 16356 1955
rect 16304 1912 16356 1921
rect 16764 1955 16816 1964
rect 16764 1921 16773 1955
rect 16773 1921 16807 1955
rect 16807 1921 16816 1955
rect 16764 1912 16816 1921
rect 17040 1955 17092 1964
rect 17040 1921 17049 1955
rect 17049 1921 17083 1955
rect 17083 1921 17092 1955
rect 17040 1912 17092 1921
rect 17316 1955 17368 1964
rect 17316 1921 17325 1955
rect 17325 1921 17359 1955
rect 17359 1921 17368 1955
rect 17316 1912 17368 1921
rect 17776 1955 17828 1964
rect 17776 1921 17785 1955
rect 17785 1921 17819 1955
rect 17819 1921 17828 1955
rect 17776 1912 17828 1921
rect 17960 1912 18012 1964
rect 19616 1980 19668 2032
rect 23572 2048 23624 2100
rect 24308 2091 24360 2100
rect 24308 2057 24317 2091
rect 24317 2057 24351 2091
rect 24351 2057 24360 2091
rect 24308 2048 24360 2057
rect 24676 2048 24728 2100
rect 25044 2048 25096 2100
rect 25872 2048 25924 2100
rect 26976 2091 27028 2100
rect 26976 2057 26985 2091
rect 26985 2057 27019 2091
rect 27019 2057 27028 2091
rect 26976 2048 27028 2057
rect 27160 2048 27212 2100
rect 28908 2048 28960 2100
rect 29184 2048 29236 2100
rect 14556 1844 14608 1896
rect 17132 1776 17184 1828
rect 17684 1844 17736 1896
rect 18696 1955 18748 1964
rect 18696 1921 18705 1955
rect 18705 1921 18739 1955
rect 18739 1921 18748 1955
rect 18696 1912 18748 1921
rect 18880 1912 18932 1964
rect 19432 1955 19484 1964
rect 19432 1921 19441 1955
rect 19441 1921 19475 1955
rect 19475 1921 19484 1955
rect 19432 1912 19484 1921
rect 19524 1955 19576 1964
rect 19524 1921 19533 1955
rect 19533 1921 19567 1955
rect 19567 1921 19576 1955
rect 19524 1912 19576 1921
rect 20260 1955 20312 1964
rect 20260 1921 20269 1955
rect 20269 1921 20303 1955
rect 20303 1921 20312 1955
rect 20260 1912 20312 1921
rect 20352 1955 20404 1964
rect 20352 1921 20361 1955
rect 20361 1921 20395 1955
rect 20395 1921 20404 1955
rect 20352 1912 20404 1921
rect 20444 1912 20496 1964
rect 21364 1955 21416 1964
rect 21364 1921 21373 1955
rect 21373 1921 21407 1955
rect 21407 1921 21416 1955
rect 21364 1912 21416 1921
rect 21640 1955 21692 1964
rect 21640 1921 21649 1955
rect 21649 1921 21683 1955
rect 21683 1921 21692 1955
rect 21640 1912 21692 1921
rect 22100 1955 22152 1964
rect 22100 1921 22109 1955
rect 22109 1921 22143 1955
rect 22143 1921 22152 1955
rect 22100 1912 22152 1921
rect 22376 1955 22428 1964
rect 22376 1921 22385 1955
rect 22385 1921 22419 1955
rect 22419 1921 22428 1955
rect 22376 1912 22428 1921
rect 22560 1912 22612 1964
rect 19340 1844 19392 1896
rect 19708 1844 19760 1896
rect 23664 1912 23716 1964
rect 24492 1955 24544 1964
rect 24492 1921 24501 1955
rect 24501 1921 24535 1955
rect 24535 1921 24544 1955
rect 24492 1912 24544 1921
rect 24768 1955 24820 1964
rect 24768 1921 24777 1955
rect 24777 1921 24811 1955
rect 24811 1921 24820 1955
rect 24768 1912 24820 1921
rect 25136 1955 25188 1964
rect 25136 1921 25145 1955
rect 25145 1921 25179 1955
rect 25179 1921 25188 1955
rect 25136 1912 25188 1921
rect 25412 1955 25464 1964
rect 25412 1921 25421 1955
rect 25421 1921 25455 1955
rect 25455 1921 25464 1955
rect 25412 1912 25464 1921
rect 25688 1955 25740 1964
rect 25688 1921 25697 1955
rect 25697 1921 25731 1955
rect 25731 1921 25740 1955
rect 25688 1912 25740 1921
rect 26424 1955 26476 1964
rect 26424 1921 26433 1955
rect 26433 1921 26467 1955
rect 26467 1921 26476 1955
rect 26424 1912 26476 1921
rect 26884 1912 26936 1964
rect 27252 1912 27304 1964
rect 26608 1844 26660 1896
rect 21824 1776 21876 1828
rect 23480 1776 23532 1828
rect 1584 1751 1636 1760
rect 1584 1717 1593 1751
rect 1593 1717 1627 1751
rect 1627 1717 1636 1751
rect 1584 1708 1636 1717
rect 16212 1751 16264 1760
rect 16212 1717 16221 1751
rect 16221 1717 16255 1751
rect 16255 1717 16264 1751
rect 16212 1708 16264 1717
rect 17500 1708 17552 1760
rect 18512 1708 18564 1760
rect 19156 1708 19208 1760
rect 20444 1708 20496 1760
rect 20812 1751 20864 1760
rect 20812 1717 20821 1751
rect 20821 1717 20855 1751
rect 20855 1717 20864 1751
rect 20812 1708 20864 1717
rect 21916 1708 21968 1760
rect 22652 1751 22704 1760
rect 22652 1717 22661 1751
rect 22661 1717 22695 1751
rect 22695 1717 22704 1751
rect 22652 1708 22704 1717
rect 23756 1751 23808 1760
rect 23756 1717 23765 1751
rect 23765 1717 23799 1751
rect 23799 1717 23808 1751
rect 23756 1708 23808 1717
rect 24032 1751 24084 1760
rect 24032 1717 24041 1751
rect 24041 1717 24075 1751
rect 24075 1717 24084 1751
rect 24032 1708 24084 1717
rect 24584 1776 24636 1828
rect 24860 1708 24912 1760
rect 24952 1708 25004 1760
rect 26792 1776 26844 1828
rect 27436 1955 27488 1964
rect 27436 1921 27445 1955
rect 27445 1921 27479 1955
rect 27479 1921 27488 1955
rect 27436 1912 27488 1921
rect 27712 1955 27764 1964
rect 27712 1921 27721 1955
rect 27721 1921 27755 1955
rect 27755 1921 27764 1955
rect 27712 1912 27764 1921
rect 28172 1912 28224 1964
rect 28264 1955 28316 1964
rect 28264 1921 28273 1955
rect 28273 1921 28307 1955
rect 28307 1921 28316 1955
rect 28264 1912 28316 1921
rect 29368 1980 29420 2032
rect 29276 1912 29328 1964
rect 29644 1912 29696 1964
rect 30012 2048 30064 2100
rect 30932 2048 30984 2100
rect 31208 1980 31260 2032
rect 33324 2048 33376 2100
rect 35900 2091 35952 2100
rect 35900 2057 35909 2091
rect 35909 2057 35943 2091
rect 35943 2057 35952 2091
rect 35900 2048 35952 2057
rect 30472 1955 30524 1964
rect 30472 1921 30481 1955
rect 30481 1921 30515 1955
rect 30515 1921 30524 1955
rect 30472 1912 30524 1921
rect 30748 1955 30800 1964
rect 30748 1921 30757 1955
rect 30757 1921 30791 1955
rect 30791 1921 30800 1955
rect 30748 1912 30800 1921
rect 31576 1955 31628 1964
rect 31576 1921 31585 1955
rect 31585 1921 31619 1955
rect 31619 1921 31628 1955
rect 31576 1912 31628 1921
rect 32312 1955 32364 1964
rect 32312 1921 32321 1955
rect 32321 1921 32355 1955
rect 32355 1921 32364 1955
rect 32312 1912 32364 1921
rect 32128 1844 32180 1896
rect 29368 1776 29420 1828
rect 30380 1776 30432 1828
rect 31668 1776 31720 1828
rect 32588 1955 32640 1964
rect 32588 1921 32597 1955
rect 32597 1921 32631 1955
rect 32631 1921 32640 1955
rect 32588 1912 32640 1921
rect 33416 1955 33468 1964
rect 33416 1921 33425 1955
rect 33425 1921 33459 1955
rect 33459 1921 33468 1955
rect 33416 1912 33468 1921
rect 35532 1980 35584 2032
rect 35716 1980 35768 2032
rect 38660 2048 38712 2100
rect 42248 2048 42300 2100
rect 44548 2048 44600 2100
rect 45192 2048 45244 2100
rect 45836 2048 45888 2100
rect 32496 1844 32548 1896
rect 33784 1844 33836 1896
rect 45008 1980 45060 2032
rect 36268 1955 36320 1964
rect 36268 1921 36277 1955
rect 36277 1921 36311 1955
rect 36311 1921 36320 1955
rect 36268 1912 36320 1921
rect 37372 1955 37424 1964
rect 37372 1921 37381 1955
rect 37381 1921 37415 1955
rect 37415 1921 37424 1955
rect 37372 1912 37424 1921
rect 38200 1912 38252 1964
rect 38752 1912 38804 1964
rect 40132 1912 40184 1964
rect 40592 1912 40644 1964
rect 41052 1955 41104 1964
rect 41052 1921 41061 1955
rect 41061 1921 41095 1955
rect 41095 1921 41104 1955
rect 41052 1912 41104 1921
rect 41328 1955 41380 1964
rect 41328 1921 41337 1955
rect 41337 1921 41371 1955
rect 41371 1921 41380 1955
rect 41328 1912 41380 1921
rect 43996 1912 44048 1964
rect 38568 1844 38620 1896
rect 33416 1776 33468 1828
rect 26056 1751 26108 1760
rect 26056 1717 26065 1751
rect 26065 1717 26099 1751
rect 26099 1717 26108 1751
rect 26056 1708 26108 1717
rect 26240 1751 26292 1760
rect 26240 1717 26249 1751
rect 26249 1717 26283 1751
rect 26283 1717 26292 1751
rect 26240 1708 26292 1717
rect 27252 1751 27304 1760
rect 27252 1717 27261 1751
rect 27261 1717 27295 1751
rect 27295 1717 27304 1751
rect 27252 1708 27304 1717
rect 27528 1751 27580 1760
rect 27528 1717 27537 1751
rect 27537 1717 27571 1751
rect 27571 1717 27580 1751
rect 27528 1708 27580 1717
rect 27988 1708 28040 1760
rect 28264 1708 28316 1760
rect 29092 1708 29144 1760
rect 30288 1751 30340 1760
rect 30288 1717 30297 1751
rect 30297 1717 30331 1751
rect 30331 1717 30340 1751
rect 30288 1708 30340 1717
rect 30932 1708 30984 1760
rect 32128 1751 32180 1760
rect 32128 1717 32137 1751
rect 32137 1717 32171 1751
rect 32171 1717 32180 1751
rect 32128 1708 32180 1717
rect 32496 1708 32548 1760
rect 33232 1751 33284 1760
rect 33232 1717 33241 1751
rect 33241 1717 33275 1751
rect 33275 1717 33284 1751
rect 33232 1708 33284 1717
rect 33784 1751 33836 1760
rect 33784 1717 33793 1751
rect 33793 1717 33827 1751
rect 33827 1717 33836 1751
rect 33784 1708 33836 1717
rect 35992 1776 36044 1828
rect 34612 1708 34664 1760
rect 36084 1708 36136 1760
rect 37280 1776 37332 1828
rect 38200 1776 38252 1828
rect 38476 1776 38528 1828
rect 40776 1776 40828 1828
rect 45744 1844 45796 1896
rect 46480 1955 46532 1964
rect 46480 1921 46489 1955
rect 46489 1921 46523 1955
rect 46523 1921 46532 1955
rect 46480 1912 46532 1921
rect 46572 1844 46624 1896
rect 38384 1751 38436 1760
rect 38384 1717 38393 1751
rect 38393 1717 38427 1751
rect 38427 1717 38436 1751
rect 38384 1708 38436 1717
rect 38936 1751 38988 1760
rect 38936 1717 38945 1751
rect 38945 1717 38979 1751
rect 38979 1717 38988 1751
rect 38936 1708 38988 1717
rect 39120 1708 39172 1760
rect 6665 1606 6717 1658
rect 6729 1606 6781 1658
rect 6793 1606 6845 1658
rect 6857 1606 6909 1658
rect 6921 1606 6973 1658
rect 18095 1606 18147 1658
rect 18159 1606 18211 1658
rect 18223 1606 18275 1658
rect 18287 1606 18339 1658
rect 18351 1606 18403 1658
rect 29525 1606 29577 1658
rect 29589 1606 29641 1658
rect 29653 1606 29705 1658
rect 29717 1606 29769 1658
rect 29781 1606 29833 1658
rect 40955 1606 41007 1658
rect 41019 1606 41071 1658
rect 41083 1606 41135 1658
rect 41147 1606 41199 1658
rect 41211 1606 41263 1658
rect 1584 1504 1636 1556
rect 8208 1504 8260 1556
rect 12716 1504 12768 1556
rect 15384 1504 15436 1556
rect 15752 1504 15804 1556
rect 16304 1504 16356 1556
rect 17040 1504 17092 1556
rect 17224 1547 17276 1556
rect 17224 1513 17233 1547
rect 17233 1513 17267 1547
rect 17267 1513 17276 1547
rect 17224 1504 17276 1513
rect 17316 1504 17368 1556
rect 17684 1504 17736 1556
rect 18696 1504 18748 1556
rect 19524 1504 19576 1556
rect 16580 1436 16632 1488
rect 1584 1343 1636 1352
rect 1584 1309 1593 1343
rect 1593 1309 1627 1343
rect 1627 1309 1636 1343
rect 1584 1300 1636 1309
rect 1952 1343 2004 1352
rect 1952 1309 1961 1343
rect 1961 1309 1995 1343
rect 1995 1309 2004 1343
rect 1952 1300 2004 1309
rect 2320 1343 2372 1352
rect 2320 1309 2329 1343
rect 2329 1309 2363 1343
rect 2363 1309 2372 1343
rect 2320 1300 2372 1309
rect 2688 1343 2740 1352
rect 2688 1309 2697 1343
rect 2697 1309 2731 1343
rect 2731 1309 2740 1343
rect 2688 1300 2740 1309
rect 2872 1300 2924 1352
rect 3148 1343 3200 1352
rect 3148 1309 3157 1343
rect 3157 1309 3191 1343
rect 3191 1309 3200 1343
rect 3148 1300 3200 1309
rect 3424 1343 3476 1352
rect 3424 1309 3433 1343
rect 3433 1309 3467 1343
rect 3467 1309 3476 1343
rect 3424 1300 3476 1309
rect 1768 1207 1820 1216
rect 1768 1173 1777 1207
rect 1777 1173 1811 1207
rect 1811 1173 1820 1207
rect 1768 1164 1820 1173
rect 2136 1207 2188 1216
rect 2136 1173 2145 1207
rect 2145 1173 2179 1207
rect 2179 1173 2188 1207
rect 2136 1164 2188 1173
rect 2504 1207 2556 1216
rect 2504 1173 2513 1207
rect 2513 1173 2547 1207
rect 2547 1173 2556 1207
rect 2504 1164 2556 1173
rect 2964 1232 3016 1284
rect 4068 1343 4120 1352
rect 4068 1309 4077 1343
rect 4077 1309 4111 1343
rect 4111 1309 4120 1343
rect 4068 1300 4120 1309
rect 4896 1343 4948 1352
rect 4896 1309 4905 1343
rect 4905 1309 4939 1343
rect 4939 1309 4948 1343
rect 4896 1300 4948 1309
rect 5264 1343 5316 1352
rect 5264 1309 5273 1343
rect 5273 1309 5307 1343
rect 5307 1309 5316 1343
rect 5264 1300 5316 1309
rect 5632 1343 5684 1352
rect 5632 1309 5641 1343
rect 5641 1309 5675 1343
rect 5675 1309 5684 1343
rect 5632 1300 5684 1309
rect 6000 1343 6052 1352
rect 6000 1309 6009 1343
rect 6009 1309 6043 1343
rect 6043 1309 6052 1343
rect 6000 1300 6052 1309
rect 6368 1343 6420 1352
rect 6368 1309 6377 1343
rect 6377 1309 6411 1343
rect 6411 1309 6420 1343
rect 6368 1300 6420 1309
rect 6736 1343 6788 1352
rect 6736 1309 6745 1343
rect 6745 1309 6779 1343
rect 6779 1309 6788 1343
rect 6736 1300 6788 1309
rect 7012 1300 7064 1352
rect 7104 1343 7156 1352
rect 7104 1309 7113 1343
rect 7113 1309 7147 1343
rect 7147 1309 7156 1343
rect 7104 1300 7156 1309
rect 7472 1343 7524 1352
rect 7472 1309 7481 1343
rect 7481 1309 7515 1343
rect 7515 1309 7524 1343
rect 7472 1300 7524 1309
rect 7840 1343 7892 1352
rect 7840 1309 7849 1343
rect 7849 1309 7883 1343
rect 7883 1309 7892 1343
rect 7840 1300 7892 1309
rect 8208 1343 8260 1352
rect 8208 1309 8217 1343
rect 8217 1309 8251 1343
rect 8251 1309 8260 1343
rect 8208 1300 8260 1309
rect 8576 1343 8628 1352
rect 8576 1309 8585 1343
rect 8585 1309 8619 1343
rect 8619 1309 8628 1343
rect 8576 1300 8628 1309
rect 8944 1343 8996 1352
rect 8944 1309 8953 1343
rect 8953 1309 8987 1343
rect 8987 1309 8996 1343
rect 8944 1300 8996 1309
rect 9312 1343 9364 1352
rect 9312 1309 9321 1343
rect 9321 1309 9355 1343
rect 9355 1309 9364 1343
rect 9312 1300 9364 1309
rect 9680 1343 9732 1352
rect 9680 1309 9689 1343
rect 9689 1309 9723 1343
rect 9723 1309 9732 1343
rect 9680 1300 9732 1309
rect 10048 1343 10100 1352
rect 10048 1309 10057 1343
rect 10057 1309 10091 1343
rect 10091 1309 10100 1343
rect 10048 1300 10100 1309
rect 10416 1343 10468 1352
rect 10416 1309 10425 1343
rect 10425 1309 10459 1343
rect 10459 1309 10468 1343
rect 10416 1300 10468 1309
rect 10784 1343 10836 1352
rect 10784 1309 10793 1343
rect 10793 1309 10827 1343
rect 10827 1309 10836 1343
rect 10784 1300 10836 1309
rect 11152 1343 11204 1352
rect 11152 1309 11161 1343
rect 11161 1309 11195 1343
rect 11195 1309 11204 1343
rect 11152 1300 11204 1309
rect 11520 1343 11572 1352
rect 11520 1309 11529 1343
rect 11529 1309 11563 1343
rect 11563 1309 11572 1343
rect 11520 1300 11572 1309
rect 11888 1343 11940 1352
rect 11888 1309 11897 1343
rect 11897 1309 11931 1343
rect 11931 1309 11940 1343
rect 11888 1300 11940 1309
rect 12256 1343 12308 1352
rect 12256 1309 12265 1343
rect 12265 1309 12299 1343
rect 12299 1309 12308 1343
rect 12256 1300 12308 1309
rect 12624 1343 12676 1352
rect 12624 1309 12633 1343
rect 12633 1309 12667 1343
rect 12667 1309 12676 1343
rect 12624 1300 12676 1309
rect 12992 1343 13044 1352
rect 12992 1309 13001 1343
rect 13001 1309 13035 1343
rect 13035 1309 13044 1343
rect 12992 1300 13044 1309
rect 13360 1343 13412 1352
rect 13360 1309 13369 1343
rect 13369 1309 13403 1343
rect 13403 1309 13412 1343
rect 13360 1300 13412 1309
rect 3332 1207 3384 1216
rect 3332 1173 3341 1207
rect 3341 1173 3375 1207
rect 3375 1173 3384 1207
rect 3332 1164 3384 1173
rect 5080 1207 5132 1216
rect 5080 1173 5089 1207
rect 5089 1173 5123 1207
rect 5123 1173 5132 1207
rect 5080 1164 5132 1173
rect 5448 1207 5500 1216
rect 5448 1173 5457 1207
rect 5457 1173 5491 1207
rect 5491 1173 5500 1207
rect 5448 1164 5500 1173
rect 5816 1207 5868 1216
rect 5816 1173 5825 1207
rect 5825 1173 5859 1207
rect 5859 1173 5868 1207
rect 5816 1164 5868 1173
rect 7932 1232 7984 1284
rect 15108 1368 15160 1420
rect 19708 1479 19760 1488
rect 19708 1445 19717 1479
rect 19717 1445 19751 1479
rect 19751 1445 19760 1479
rect 19708 1436 19760 1445
rect 19800 1436 19852 1488
rect 13728 1343 13780 1352
rect 13728 1309 13737 1343
rect 13737 1309 13771 1343
rect 13771 1309 13780 1343
rect 13728 1300 13780 1309
rect 13820 1300 13872 1352
rect 14096 1343 14148 1352
rect 14096 1309 14105 1343
rect 14105 1309 14139 1343
rect 14139 1309 14148 1343
rect 14096 1300 14148 1309
rect 14648 1343 14700 1352
rect 14648 1309 14657 1343
rect 14657 1309 14691 1343
rect 14691 1309 14700 1343
rect 14648 1300 14700 1309
rect 15016 1343 15068 1352
rect 15016 1309 15025 1343
rect 15025 1309 15059 1343
rect 15059 1309 15068 1343
rect 15016 1300 15068 1309
rect 15384 1343 15436 1352
rect 15384 1309 15393 1343
rect 15393 1309 15427 1343
rect 15427 1309 15436 1343
rect 15384 1300 15436 1309
rect 6920 1207 6972 1216
rect 6920 1173 6929 1207
rect 6929 1173 6963 1207
rect 6963 1173 6972 1207
rect 6920 1164 6972 1173
rect 7288 1207 7340 1216
rect 7288 1173 7297 1207
rect 7297 1173 7331 1207
rect 7331 1173 7340 1207
rect 7288 1164 7340 1173
rect 7656 1207 7708 1216
rect 7656 1173 7665 1207
rect 7665 1173 7699 1207
rect 7699 1173 7708 1207
rect 7656 1164 7708 1173
rect 8392 1207 8444 1216
rect 8392 1173 8401 1207
rect 8401 1173 8435 1207
rect 8435 1173 8444 1207
rect 8392 1164 8444 1173
rect 8760 1207 8812 1216
rect 8760 1173 8769 1207
rect 8769 1173 8803 1207
rect 8803 1173 8812 1207
rect 8760 1164 8812 1173
rect 9128 1207 9180 1216
rect 9128 1173 9137 1207
rect 9137 1173 9171 1207
rect 9171 1173 9180 1207
rect 9128 1164 9180 1173
rect 9496 1207 9548 1216
rect 9496 1173 9505 1207
rect 9505 1173 9539 1207
rect 9539 1173 9548 1207
rect 9496 1164 9548 1173
rect 9864 1207 9916 1216
rect 9864 1173 9873 1207
rect 9873 1173 9907 1207
rect 9907 1173 9916 1207
rect 9864 1164 9916 1173
rect 10232 1207 10284 1216
rect 10232 1173 10241 1207
rect 10241 1173 10275 1207
rect 10275 1173 10284 1207
rect 10232 1164 10284 1173
rect 10600 1207 10652 1216
rect 10600 1173 10609 1207
rect 10609 1173 10643 1207
rect 10643 1173 10652 1207
rect 10600 1164 10652 1173
rect 10968 1207 11020 1216
rect 10968 1173 10977 1207
rect 10977 1173 11011 1207
rect 11011 1173 11020 1207
rect 10968 1164 11020 1173
rect 11336 1207 11388 1216
rect 11336 1173 11345 1207
rect 11345 1173 11379 1207
rect 11379 1173 11388 1207
rect 11336 1164 11388 1173
rect 11704 1207 11756 1216
rect 11704 1173 11713 1207
rect 11713 1173 11747 1207
rect 11747 1173 11756 1207
rect 11704 1164 11756 1173
rect 12072 1207 12124 1216
rect 12072 1173 12081 1207
rect 12081 1173 12115 1207
rect 12115 1173 12124 1207
rect 12072 1164 12124 1173
rect 12808 1207 12860 1216
rect 12808 1173 12817 1207
rect 12817 1173 12851 1207
rect 12851 1173 12860 1207
rect 12808 1164 12860 1173
rect 13176 1207 13228 1216
rect 13176 1173 13185 1207
rect 13185 1173 13219 1207
rect 13219 1173 13228 1207
rect 13176 1164 13228 1173
rect 15660 1343 15712 1352
rect 15660 1309 15669 1343
rect 15669 1309 15703 1343
rect 15703 1309 15712 1343
rect 15660 1300 15712 1309
rect 15936 1343 15988 1352
rect 15936 1309 15945 1343
rect 15945 1309 15979 1343
rect 15979 1309 15988 1343
rect 15936 1300 15988 1309
rect 16028 1300 16080 1352
rect 16212 1343 16264 1352
rect 16212 1309 16221 1343
rect 16221 1309 16255 1343
rect 16255 1309 16264 1343
rect 16212 1300 16264 1309
rect 16580 1300 16632 1352
rect 16856 1343 16908 1352
rect 16856 1309 16865 1343
rect 16865 1309 16899 1343
rect 16899 1309 16908 1343
rect 16856 1300 16908 1309
rect 17132 1343 17184 1352
rect 17132 1309 17141 1343
rect 17141 1309 17175 1343
rect 17175 1309 17184 1343
rect 17132 1300 17184 1309
rect 17408 1343 17460 1352
rect 17408 1309 17417 1343
rect 17417 1309 17451 1343
rect 17451 1309 17460 1343
rect 17408 1300 17460 1309
rect 17684 1343 17736 1352
rect 17684 1309 17693 1343
rect 17693 1309 17727 1343
rect 17727 1309 17736 1343
rect 17684 1300 17736 1309
rect 13912 1207 13964 1216
rect 13912 1173 13921 1207
rect 13921 1173 13955 1207
rect 13955 1173 13964 1207
rect 13912 1164 13964 1173
rect 14280 1207 14332 1216
rect 14280 1173 14289 1207
rect 14289 1173 14323 1207
rect 14323 1173 14332 1207
rect 14280 1164 14332 1173
rect 14832 1207 14884 1216
rect 14832 1173 14841 1207
rect 14841 1173 14875 1207
rect 14875 1173 14884 1207
rect 14832 1164 14884 1173
rect 16764 1232 16816 1284
rect 18236 1343 18288 1352
rect 18236 1309 18245 1343
rect 18245 1309 18279 1343
rect 18279 1309 18288 1343
rect 18236 1300 18288 1309
rect 18512 1343 18564 1352
rect 18512 1309 18521 1343
rect 18521 1309 18555 1343
rect 18555 1309 18564 1343
rect 18512 1300 18564 1309
rect 19248 1368 19300 1420
rect 18420 1232 18472 1284
rect 17960 1164 18012 1216
rect 20444 1504 20496 1556
rect 24400 1504 24452 1556
rect 24676 1504 24728 1556
rect 26148 1504 26200 1556
rect 27620 1504 27672 1556
rect 28724 1504 28776 1556
rect 20168 1436 20220 1488
rect 20536 1368 20588 1420
rect 20628 1411 20680 1420
rect 20628 1377 20637 1411
rect 20637 1377 20671 1411
rect 20671 1377 20680 1411
rect 20628 1368 20680 1377
rect 21456 1436 21508 1488
rect 23388 1436 23440 1488
rect 28908 1436 28960 1488
rect 29828 1504 29880 1556
rect 30840 1504 30892 1556
rect 31300 1504 31352 1556
rect 32772 1504 32824 1556
rect 19156 1232 19208 1284
rect 19984 1300 20036 1352
rect 21088 1300 21140 1352
rect 22008 1343 22060 1352
rect 22008 1309 22017 1343
rect 22017 1309 22051 1343
rect 22051 1309 22060 1343
rect 22008 1300 22060 1309
rect 22284 1300 22336 1352
rect 19800 1232 19852 1284
rect 19064 1207 19116 1216
rect 19064 1173 19073 1207
rect 19073 1173 19107 1207
rect 19107 1173 19116 1207
rect 19064 1164 19116 1173
rect 23480 1300 23532 1352
rect 24032 1300 24084 1352
rect 24216 1300 24268 1352
rect 24768 1300 24820 1352
rect 25412 1368 25464 1420
rect 30472 1368 30524 1420
rect 30656 1368 30708 1420
rect 20076 1207 20128 1216
rect 20076 1173 20085 1207
rect 20085 1173 20119 1207
rect 20119 1173 20128 1207
rect 20076 1164 20128 1173
rect 21180 1207 21232 1216
rect 21180 1173 21189 1207
rect 21189 1173 21223 1207
rect 21223 1173 21232 1207
rect 21180 1164 21232 1173
rect 21548 1207 21600 1216
rect 21548 1173 21557 1207
rect 21557 1173 21591 1207
rect 21591 1173 21600 1207
rect 21548 1164 21600 1173
rect 21916 1164 21968 1216
rect 24860 1275 24912 1284
rect 24860 1241 24869 1275
rect 24869 1241 24903 1275
rect 24903 1241 24912 1275
rect 24860 1232 24912 1241
rect 26240 1300 26292 1352
rect 26516 1300 26568 1352
rect 27252 1300 27304 1352
rect 27528 1300 27580 1352
rect 27988 1300 28040 1352
rect 29000 1300 29052 1352
rect 30288 1300 30340 1352
rect 31024 1300 31076 1352
rect 31668 1436 31720 1488
rect 33140 1436 33192 1488
rect 34152 1504 34204 1556
rect 34980 1504 35032 1556
rect 34336 1436 34388 1488
rect 35900 1436 35952 1488
rect 36820 1504 36872 1556
rect 38292 1504 38344 1556
rect 39304 1504 39356 1556
rect 40776 1504 40828 1556
rect 41512 1504 41564 1556
rect 42800 1504 42852 1556
rect 45008 1547 45060 1556
rect 45008 1513 45017 1547
rect 45017 1513 45051 1547
rect 45051 1513 45060 1547
rect 45008 1504 45060 1513
rect 45744 1547 45796 1556
rect 45744 1513 45753 1547
rect 45753 1513 45787 1547
rect 45787 1513 45796 1547
rect 45744 1504 45796 1513
rect 37096 1436 37148 1488
rect 38844 1436 38896 1488
rect 32496 1368 32548 1420
rect 33600 1368 33652 1420
rect 33692 1368 33744 1420
rect 44088 1479 44140 1488
rect 44088 1445 44097 1479
rect 44097 1445 44131 1479
rect 44131 1445 44140 1479
rect 44088 1436 44140 1445
rect 44456 1479 44508 1488
rect 44456 1445 44465 1479
rect 44465 1445 44499 1479
rect 44499 1445 44508 1479
rect 44456 1436 44508 1445
rect 28080 1232 28132 1284
rect 30380 1275 30432 1284
rect 30380 1241 30389 1275
rect 30389 1241 30423 1275
rect 30423 1241 30432 1275
rect 30380 1232 30432 1241
rect 30472 1232 30524 1284
rect 32128 1300 32180 1352
rect 32956 1300 33008 1352
rect 33232 1300 33284 1352
rect 34888 1300 34940 1352
rect 37740 1300 37792 1352
rect 23020 1207 23072 1216
rect 23020 1173 23029 1207
rect 23029 1173 23063 1207
rect 23063 1173 23072 1207
rect 23020 1164 23072 1173
rect 23388 1207 23440 1216
rect 23388 1173 23397 1207
rect 23397 1173 23431 1207
rect 23431 1173 23440 1207
rect 23388 1164 23440 1173
rect 24124 1207 24176 1216
rect 24124 1173 24133 1207
rect 24133 1173 24167 1207
rect 24167 1173 24176 1207
rect 24124 1164 24176 1173
rect 24584 1207 24636 1216
rect 24584 1173 24593 1207
rect 24593 1173 24627 1207
rect 24627 1173 24636 1207
rect 24584 1164 24636 1173
rect 25044 1164 25096 1216
rect 25596 1164 25648 1216
rect 26516 1164 26568 1216
rect 27252 1164 27304 1216
rect 27988 1164 28040 1216
rect 30288 1164 30340 1216
rect 34796 1275 34848 1284
rect 34796 1241 34805 1275
rect 34805 1241 34839 1275
rect 34839 1241 34848 1275
rect 34796 1232 34848 1241
rect 35072 1232 35124 1284
rect 38108 1300 38160 1352
rect 39028 1343 39080 1352
rect 39028 1309 39037 1343
rect 39037 1309 39071 1343
rect 39071 1309 39080 1343
rect 39028 1300 39080 1309
rect 39488 1343 39540 1352
rect 39488 1309 39497 1343
rect 39497 1309 39531 1343
rect 39531 1309 39540 1343
rect 39488 1300 39540 1309
rect 40040 1300 40092 1352
rect 37464 1207 37516 1216
rect 37464 1173 37473 1207
rect 37473 1173 37507 1207
rect 37507 1173 37516 1207
rect 40224 1232 40276 1284
rect 41696 1343 41748 1352
rect 41696 1309 41705 1343
rect 41705 1309 41739 1343
rect 41739 1309 41748 1343
rect 41696 1300 41748 1309
rect 41880 1300 41932 1352
rect 41972 1232 42024 1284
rect 42340 1232 42392 1284
rect 43260 1343 43312 1352
rect 43260 1309 43269 1343
rect 43269 1309 43303 1343
rect 43303 1309 43312 1343
rect 43260 1300 43312 1309
rect 43536 1343 43588 1352
rect 43536 1309 43545 1343
rect 43545 1309 43579 1343
rect 43579 1309 43588 1343
rect 43536 1300 43588 1309
rect 43904 1343 43956 1352
rect 43904 1309 43913 1343
rect 43913 1309 43947 1343
rect 43947 1309 43956 1343
rect 43904 1300 43956 1309
rect 44272 1343 44324 1352
rect 44272 1309 44281 1343
rect 44281 1309 44315 1343
rect 44315 1309 44324 1343
rect 44272 1300 44324 1309
rect 44640 1343 44692 1352
rect 44640 1309 44649 1343
rect 44649 1309 44683 1343
rect 44683 1309 44692 1343
rect 44640 1300 44692 1309
rect 45192 1343 45244 1352
rect 45192 1309 45201 1343
rect 45201 1309 45235 1343
rect 45235 1309 45244 1343
rect 45192 1300 45244 1309
rect 45560 1343 45612 1352
rect 45560 1309 45569 1343
rect 45569 1309 45603 1343
rect 45603 1309 45612 1343
rect 45560 1300 45612 1309
rect 45928 1343 45980 1352
rect 45928 1309 45937 1343
rect 45937 1309 45971 1343
rect 45971 1309 45980 1343
rect 45928 1300 45980 1309
rect 46296 1343 46348 1352
rect 46296 1309 46305 1343
rect 46305 1309 46339 1343
rect 46339 1309 46348 1343
rect 46296 1300 46348 1309
rect 37464 1164 37516 1173
rect 39672 1207 39724 1216
rect 39672 1173 39681 1207
rect 39681 1173 39715 1207
rect 39715 1173 39724 1207
rect 39672 1164 39724 1173
rect 41144 1207 41196 1216
rect 41144 1173 41153 1207
rect 41153 1173 41187 1207
rect 41187 1173 41196 1207
rect 41144 1164 41196 1173
rect 41236 1164 41288 1216
rect 42708 1164 42760 1216
rect 42892 1207 42944 1216
rect 42892 1173 42901 1207
rect 42901 1173 42935 1207
rect 42935 1173 42944 1207
rect 42892 1164 42944 1173
rect 43168 1207 43220 1216
rect 43168 1173 43177 1207
rect 43177 1173 43211 1207
rect 43211 1173 43220 1207
rect 43168 1164 43220 1173
rect 43444 1207 43496 1216
rect 43444 1173 43453 1207
rect 43453 1173 43487 1207
rect 43487 1173 43496 1207
rect 43444 1164 43496 1173
rect 43720 1207 43772 1216
rect 43720 1173 43729 1207
rect 43729 1173 43763 1207
rect 43763 1173 43772 1207
rect 43720 1164 43772 1173
rect 43996 1232 44048 1284
rect 12380 1062 12432 1114
rect 12444 1062 12496 1114
rect 12508 1062 12560 1114
rect 12572 1062 12624 1114
rect 12636 1062 12688 1114
rect 23810 1062 23862 1114
rect 23874 1062 23926 1114
rect 23938 1062 23990 1114
rect 24002 1062 24054 1114
rect 24066 1062 24118 1114
rect 35240 1062 35292 1114
rect 35304 1062 35356 1114
rect 35368 1062 35420 1114
rect 35432 1062 35484 1114
rect 35496 1062 35548 1114
rect 46670 1062 46722 1114
rect 46734 1062 46786 1114
rect 46798 1062 46850 1114
rect 46862 1062 46914 1114
rect 46926 1062 46978 1114
rect 2136 960 2188 1012
rect 7288 960 7340 1012
rect 15108 960 15160 1012
rect 7932 892 7984 944
rect 3332 824 3384 876
rect 9772 824 9824 876
rect 5080 756 5132 808
rect 8668 756 8720 808
rect 2504 552 2556 604
rect 5540 552 5592 604
rect 1768 484 1820 536
rect 5724 484 5776 536
rect 5816 484 5868 536
rect 5448 416 5500 468
rect 6920 416 6972 468
rect 7656 688 7708 740
rect 11336 892 11388 944
rect 11704 892 11756 944
rect 17500 892 17552 944
rect 17224 824 17276 876
rect 18972 824 19024 876
rect 17224 688 17276 740
rect 18512 756 18564 808
rect 19156 756 19208 808
rect 19432 892 19484 944
rect 20536 824 20588 876
rect 21824 960 21876 1012
rect 30472 960 30524 1012
rect 31116 960 31168 1012
rect 41236 960 41288 1012
rect 44088 960 44140 1012
rect 24308 892 24360 944
rect 34796 892 34848 944
rect 35072 892 35124 944
rect 39672 892 39724 944
rect 28540 756 28592 808
rect 28356 688 28408 740
rect 29000 824 29052 876
rect 29276 756 29328 808
rect 30104 688 30156 740
rect 30840 688 30892 740
rect 31576 688 31628 740
rect 33968 688 34020 740
rect 37464 688 37516 740
rect 10232 620 10284 672
rect 32220 620 32272 672
rect 14740 552 14792 604
rect 8392 484 8444 536
rect 9864 484 9916 536
rect 32588 552 32640 604
rect 18236 484 18288 536
rect 18788 484 18840 536
rect 20536 484 20588 536
rect 42892 552 42944 604
rect 13912 416 13964 468
rect 27344 416 27396 468
rect 29368 416 29420 468
rect 41144 416 41196 468
rect 13636 348 13688 400
rect 14280 348 14332 400
rect 28172 348 28224 400
rect 28356 348 28408 400
rect 30564 348 30616 400
rect 30748 348 30800 400
rect 43444 552 43496 604
rect 43720 552 43772 604
rect 11244 280 11296 332
rect 14556 280 14608 332
rect 14832 280 14884 332
rect 20352 280 20404 332
rect 25688 280 25740 332
rect 12624 212 12676 264
rect 12808 212 12860 264
rect 27804 212 27856 264
rect 29920 144 29972 196
rect 30104 144 30156 196
rect 31024 144 31076 196
rect 13452 76 13504 128
rect 26792 76 26844 128
rect 40224 144 40276 196
<< metal2 >>
rect 1858 9840 1914 10000
rect 4066 9840 4122 10000
rect 6274 9840 6330 10000
rect 8482 9840 8538 10000
rect 10690 9840 10746 10000
rect 12898 9840 12954 10000
rect 15106 9840 15162 10000
rect 17314 9840 17370 10000
rect 19522 9840 19578 10000
rect 21730 9840 21786 10000
rect 23938 9840 23994 10000
rect 24044 9846 24256 9874
rect 1872 8634 1900 9840
rect 4080 8634 4108 9840
rect 6288 8634 6316 9840
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6380 8498 6408 8774
rect 6472 8566 6500 8774
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6564 8430 6592 8774
rect 8496 8634 8524 9840
rect 10704 8634 10732 9840
rect 12380 8732 12688 8741
rect 12380 8730 12386 8732
rect 12442 8730 12466 8732
rect 12522 8730 12546 8732
rect 12602 8730 12626 8732
rect 12682 8730 12688 8732
rect 12442 8678 12444 8730
rect 12624 8678 12626 8730
rect 12380 8676 12386 8678
rect 12442 8676 12466 8678
rect 12522 8676 12546 8678
rect 12602 8676 12626 8678
rect 12682 8676 12688 8678
rect 12380 8667 12688 8676
rect 12912 8634 12940 9840
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13004 8498 13032 8910
rect 15120 8634 15148 9840
rect 17328 8634 17356 9840
rect 19536 8634 19564 9840
rect 21744 8634 21772 9840
rect 23952 9738 23980 9840
rect 24044 9738 24072 9846
rect 23952 9710 24072 9738
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 22192 8968 22244 8974
rect 22192 8910 22244 8916
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6665 8188 6973 8197
rect 6665 8186 6671 8188
rect 6727 8186 6751 8188
rect 6807 8186 6831 8188
rect 6887 8186 6911 8188
rect 6967 8186 6973 8188
rect 6727 8134 6729 8186
rect 6909 8134 6911 8186
rect 6665 8132 6671 8134
rect 6727 8132 6751 8134
rect 6807 8132 6831 8134
rect 6887 8132 6911 8134
rect 6967 8132 6973 8134
rect 6665 8123 6973 8132
rect 12380 7644 12688 7653
rect 12380 7642 12386 7644
rect 12442 7642 12466 7644
rect 12522 7642 12546 7644
rect 12602 7642 12626 7644
rect 12682 7642 12688 7644
rect 12442 7590 12444 7642
rect 12624 7590 12626 7642
rect 12380 7588 12386 7590
rect 12442 7588 12466 7590
rect 12522 7588 12546 7590
rect 12602 7588 12626 7590
rect 12682 7588 12688 7590
rect 12380 7579 12688 7588
rect 6665 7100 6973 7109
rect 6665 7098 6671 7100
rect 6727 7098 6751 7100
rect 6807 7098 6831 7100
rect 6887 7098 6911 7100
rect 6967 7098 6973 7100
rect 6727 7046 6729 7098
rect 6909 7046 6911 7098
rect 6665 7044 6671 7046
rect 6727 7044 6751 7046
rect 6807 7044 6831 7046
rect 6887 7044 6911 7046
rect 6967 7044 6973 7046
rect 6665 7035 6973 7044
rect 12380 6556 12688 6565
rect 12380 6554 12386 6556
rect 12442 6554 12466 6556
rect 12522 6554 12546 6556
rect 12602 6554 12626 6556
rect 12682 6554 12688 6556
rect 12442 6502 12444 6554
rect 12624 6502 12626 6554
rect 12380 6500 12386 6502
rect 12442 6500 12466 6502
rect 12522 6500 12546 6502
rect 12602 6500 12626 6502
rect 12682 6500 12688 6502
rect 12380 6491 12688 6500
rect 6665 6012 6973 6021
rect 6665 6010 6671 6012
rect 6727 6010 6751 6012
rect 6807 6010 6831 6012
rect 6887 6010 6911 6012
rect 6967 6010 6973 6012
rect 6727 5958 6729 6010
rect 6909 5958 6911 6010
rect 6665 5956 6671 5958
rect 6727 5956 6751 5958
rect 6807 5956 6831 5958
rect 6887 5956 6911 5958
rect 6967 5956 6973 5958
rect 6665 5947 6973 5956
rect 12380 5468 12688 5477
rect 12380 5466 12386 5468
rect 12442 5466 12466 5468
rect 12522 5466 12546 5468
rect 12602 5466 12626 5468
rect 12682 5466 12688 5468
rect 12442 5414 12444 5466
rect 12624 5414 12626 5466
rect 12380 5412 12386 5414
rect 12442 5412 12466 5414
rect 12522 5412 12546 5414
rect 12602 5412 12626 5414
rect 12682 5412 12688 5414
rect 12380 5403 12688 5412
rect 6665 4924 6973 4933
rect 6665 4922 6671 4924
rect 6727 4922 6751 4924
rect 6807 4922 6831 4924
rect 6887 4922 6911 4924
rect 6967 4922 6973 4924
rect 6727 4870 6729 4922
rect 6909 4870 6911 4922
rect 6665 4868 6671 4870
rect 6727 4868 6751 4870
rect 6807 4868 6831 4870
rect 6887 4868 6911 4870
rect 6967 4868 6973 4870
rect 6665 4859 6973 4868
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 1124 1964 1176 1970
rect 1124 1906 1176 1912
rect 1136 160 1164 1906
rect 1584 1760 1636 1766
rect 1584 1702 1636 1708
rect 1596 1562 1624 1702
rect 1584 1556 1636 1562
rect 1584 1498 1636 1504
rect 2884 1358 2912 4150
rect 3988 2774 4016 4218
rect 6665 3836 6973 3845
rect 6665 3834 6671 3836
rect 6727 3834 6751 3836
rect 6807 3834 6831 3836
rect 6887 3834 6911 3836
rect 6967 3834 6973 3836
rect 6727 3782 6729 3834
rect 6909 3782 6911 3834
rect 6665 3780 6671 3782
rect 6727 3780 6751 3782
rect 6807 3780 6831 3782
rect 6887 3780 6911 3782
rect 6967 3780 6973 3782
rect 6665 3771 6973 3780
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 3988 2746 4108 2774
rect 3976 1964 4028 1970
rect 3976 1906 4028 1912
rect 1584 1352 1636 1358
rect 1584 1294 1636 1300
rect 1952 1352 2004 1358
rect 1952 1294 2004 1300
rect 2320 1352 2372 1358
rect 2320 1294 2372 1300
rect 2688 1352 2740 1358
rect 2688 1294 2740 1300
rect 2872 1352 2924 1358
rect 2872 1294 2924 1300
rect 3148 1352 3200 1358
rect 3148 1294 3200 1300
rect 3424 1352 3476 1358
rect 3424 1294 3476 1300
rect 1122 0 1178 160
rect 1490 82 1546 160
rect 1596 82 1624 1294
rect 1768 1216 1820 1222
rect 1768 1158 1820 1164
rect 1780 542 1808 1158
rect 1768 536 1820 542
rect 1768 478 1820 484
rect 1490 54 1624 82
rect 1858 82 1914 160
rect 1964 82 1992 1294
rect 2136 1216 2188 1222
rect 2136 1158 2188 1164
rect 2148 1018 2176 1158
rect 2136 1012 2188 1018
rect 2136 954 2188 960
rect 1858 54 1992 82
rect 2226 82 2282 160
rect 2332 82 2360 1294
rect 2504 1216 2556 1222
rect 2504 1158 2556 1164
rect 2516 610 2544 1158
rect 2504 604 2556 610
rect 2504 546 2556 552
rect 2226 54 2360 82
rect 2594 82 2650 160
rect 2700 82 2728 1294
rect 2964 1284 3016 1290
rect 2964 1226 3016 1232
rect 2976 160 3004 1226
rect 2594 54 2728 82
rect 1490 0 1546 54
rect 1858 0 1914 54
rect 2226 0 2282 54
rect 2594 0 2650 54
rect 2962 0 3018 160
rect 3160 82 3188 1294
rect 3332 1216 3384 1222
rect 3332 1158 3384 1164
rect 3344 882 3372 1158
rect 3332 876 3384 882
rect 3332 818 3384 824
rect 3330 82 3386 160
rect 3160 54 3386 82
rect 3436 82 3464 1294
rect 3698 82 3754 160
rect 3436 54 3754 82
rect 3988 82 4016 1906
rect 4080 1358 4108 2746
rect 4528 1964 4580 1970
rect 4528 1906 4580 1912
rect 4068 1352 4120 1358
rect 4068 1294 4120 1300
rect 4066 82 4122 160
rect 3988 54 4122 82
rect 3330 0 3386 54
rect 3698 0 3754 54
rect 4066 0 4122 54
rect 4434 82 4490 160
rect 4540 82 4568 1906
rect 4896 1352 4948 1358
rect 4896 1294 4948 1300
rect 5264 1352 5316 1358
rect 5264 1294 5316 1300
rect 4434 54 4568 82
rect 4802 82 4858 160
rect 4908 82 4936 1294
rect 5080 1216 5132 1222
rect 5080 1158 5132 1164
rect 5092 814 5120 1158
rect 5080 808 5132 814
rect 5080 750 5132 756
rect 4802 54 4936 82
rect 5170 82 5226 160
rect 5276 82 5304 1294
rect 5448 1216 5500 1222
rect 5448 1158 5500 1164
rect 5460 474 5488 1158
rect 5552 610 5580 3062
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5632 1352 5684 1358
rect 5632 1294 5684 1300
rect 5540 604 5592 610
rect 5540 546 5592 552
rect 5448 468 5500 474
rect 5448 410 5500 416
rect 5170 54 5304 82
rect 5538 82 5594 160
rect 5644 82 5672 1294
rect 5736 542 5764 2858
rect 6665 2748 6973 2757
rect 6665 2746 6671 2748
rect 6727 2746 6751 2748
rect 6807 2746 6831 2748
rect 6887 2746 6911 2748
rect 6967 2746 6973 2748
rect 6727 2694 6729 2746
rect 6909 2694 6911 2746
rect 6665 2692 6671 2694
rect 6727 2692 6751 2694
rect 6807 2692 6831 2694
rect 6887 2692 6911 2694
rect 6967 2692 6973 2694
rect 6665 2683 6973 2692
rect 6665 1660 6973 1669
rect 6665 1658 6671 1660
rect 6727 1658 6751 1660
rect 6807 1658 6831 1660
rect 6887 1658 6911 1660
rect 6967 1658 6973 1660
rect 6727 1606 6729 1658
rect 6909 1606 6911 1658
rect 6665 1604 6671 1606
rect 6727 1604 6751 1606
rect 6807 1604 6831 1606
rect 6887 1604 6911 1606
rect 6967 1604 6973 1606
rect 6665 1595 6973 1604
rect 7024 1358 7052 4490
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 12380 4380 12688 4389
rect 12380 4378 12386 4380
rect 12442 4378 12466 4380
rect 12522 4378 12546 4380
rect 12602 4378 12626 4380
rect 12682 4378 12688 4380
rect 12442 4326 12444 4378
rect 12624 4326 12626 4378
rect 12380 4324 12386 4326
rect 12442 4324 12466 4326
rect 12522 4324 12546 4326
rect 12602 4324 12626 4326
rect 12682 4324 12688 4326
rect 12380 4315 12688 4324
rect 15934 3632 15990 3641
rect 15934 3567 15990 3576
rect 13452 3528 13504 3534
rect 12070 3496 12126 3505
rect 13452 3470 13504 3476
rect 12070 3431 12126 3440
rect 12716 3460 12768 3466
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 8220 1562 8248 2518
rect 8666 2408 8722 2417
rect 8666 2343 8722 2352
rect 8208 1556 8260 1562
rect 8208 1498 8260 1504
rect 6000 1352 6052 1358
rect 6000 1294 6052 1300
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 6736 1352 6788 1358
rect 6736 1294 6788 1300
rect 7012 1352 7064 1358
rect 7012 1294 7064 1300
rect 7104 1352 7156 1358
rect 7104 1294 7156 1300
rect 7472 1352 7524 1358
rect 7472 1294 7524 1300
rect 7840 1352 7892 1358
rect 7840 1294 7892 1300
rect 8208 1352 8260 1358
rect 8208 1294 8260 1300
rect 8576 1352 8628 1358
rect 8576 1294 8628 1300
rect 5816 1216 5868 1222
rect 5816 1158 5868 1164
rect 5828 542 5856 1158
rect 5724 536 5776 542
rect 5724 478 5776 484
rect 5816 536 5868 542
rect 5816 478 5868 484
rect 5538 54 5672 82
rect 5906 82 5962 160
rect 6012 82 6040 1294
rect 5906 54 6040 82
rect 6274 82 6330 160
rect 6380 82 6408 1294
rect 6274 54 6408 82
rect 6642 82 6698 160
rect 6748 82 6776 1294
rect 6920 1216 6972 1222
rect 6920 1158 6972 1164
rect 6932 474 6960 1158
rect 6920 468 6972 474
rect 6920 410 6972 416
rect 6642 54 6776 82
rect 7010 82 7066 160
rect 7116 82 7144 1294
rect 7288 1216 7340 1222
rect 7288 1158 7340 1164
rect 7300 1018 7328 1158
rect 7288 1012 7340 1018
rect 7288 954 7340 960
rect 7010 54 7144 82
rect 7378 82 7434 160
rect 7484 82 7512 1294
rect 7656 1216 7708 1222
rect 7656 1158 7708 1164
rect 7668 746 7696 1158
rect 7656 740 7708 746
rect 7656 682 7708 688
rect 7378 54 7512 82
rect 7746 82 7802 160
rect 7852 82 7880 1294
rect 7932 1284 7984 1290
rect 7932 1226 7984 1232
rect 7944 950 7972 1226
rect 7932 944 7984 950
rect 7932 886 7984 892
rect 7746 54 7880 82
rect 8114 82 8170 160
rect 8220 82 8248 1294
rect 8392 1216 8444 1222
rect 8392 1158 8444 1164
rect 8404 542 8432 1158
rect 8392 536 8444 542
rect 8392 478 8444 484
rect 8114 54 8248 82
rect 8482 82 8538 160
rect 8588 82 8616 1294
rect 8680 814 8708 2343
rect 8772 1222 8800 3130
rect 9862 3088 9918 3097
rect 9862 3023 9918 3032
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 8944 1352 8996 1358
rect 8944 1294 8996 1300
rect 9312 1352 9364 1358
rect 9312 1294 9364 1300
rect 8760 1216 8812 1222
rect 8760 1158 8812 1164
rect 8668 808 8720 814
rect 8668 750 8720 756
rect 8482 54 8616 82
rect 8850 82 8906 160
rect 8956 82 8984 1294
rect 9128 1216 9180 1222
rect 9128 1158 9180 1164
rect 9140 377 9168 1158
rect 9126 368 9182 377
rect 9126 303 9182 312
rect 8850 54 8984 82
rect 9218 82 9274 160
rect 9324 82 9352 1294
rect 9496 1216 9548 1222
rect 9496 1158 9548 1164
rect 9508 513 9536 1158
rect 9494 504 9550 513
rect 9494 439 9550 448
rect 9600 160 9628 2790
rect 9692 1358 9720 2790
rect 9876 2774 9904 3023
rect 9784 2746 9904 2774
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 9784 882 9812 2746
rect 10048 1352 10100 1358
rect 10048 1294 10100 1300
rect 10416 1352 10468 1358
rect 10416 1294 10468 1300
rect 10784 1352 10836 1358
rect 10784 1294 10836 1300
rect 11152 1352 11204 1358
rect 11520 1352 11572 1358
rect 11152 1294 11204 1300
rect 11242 1320 11298 1329
rect 9864 1216 9916 1222
rect 9864 1158 9916 1164
rect 9772 876 9824 882
rect 9772 818 9824 824
rect 9876 542 9904 1158
rect 9864 536 9916 542
rect 9864 478 9916 484
rect 9218 54 9352 82
rect 4434 0 4490 54
rect 4802 0 4858 54
rect 5170 0 5226 54
rect 5538 0 5594 54
rect 5906 0 5962 54
rect 6274 0 6330 54
rect 6642 0 6698 54
rect 7010 0 7066 54
rect 7378 0 7434 54
rect 7746 0 7802 54
rect 8114 0 8170 54
rect 8482 0 8538 54
rect 8850 0 8906 54
rect 9218 0 9274 54
rect 9586 0 9642 160
rect 9954 82 10010 160
rect 10060 82 10088 1294
rect 10232 1216 10284 1222
rect 10232 1158 10284 1164
rect 10244 678 10272 1158
rect 10232 672 10284 678
rect 10232 614 10284 620
rect 9954 54 10088 82
rect 10322 82 10378 160
rect 10428 82 10456 1294
rect 10600 1216 10652 1222
rect 10600 1158 10652 1164
rect 10612 241 10640 1158
rect 10598 232 10654 241
rect 10598 167 10654 176
rect 10322 54 10456 82
rect 10690 82 10746 160
rect 10796 82 10824 1294
rect 10968 1216 11020 1222
rect 10968 1158 11020 1164
rect 10980 921 11008 1158
rect 10966 912 11022 921
rect 10966 847 11022 856
rect 10690 54 10824 82
rect 11058 82 11114 160
rect 11164 82 11192 1294
rect 11520 1294 11572 1300
rect 11888 1352 11940 1358
rect 11888 1294 11940 1300
rect 11242 1255 11298 1264
rect 11256 338 11284 1255
rect 11336 1216 11388 1222
rect 11336 1158 11388 1164
rect 11348 950 11376 1158
rect 11336 944 11388 950
rect 11336 886 11388 892
rect 11244 332 11296 338
rect 11244 274 11296 280
rect 11058 54 11192 82
rect 11426 82 11482 160
rect 11532 82 11560 1294
rect 11704 1216 11756 1222
rect 11704 1158 11756 1164
rect 11716 950 11744 1158
rect 11704 944 11756 950
rect 11704 886 11756 892
rect 11426 54 11560 82
rect 11794 82 11850 160
rect 11900 82 11928 1294
rect 12084 1222 12112 3431
rect 12716 3402 12768 3408
rect 12380 3292 12688 3301
rect 12380 3290 12386 3292
rect 12442 3290 12466 3292
rect 12522 3290 12546 3292
rect 12602 3290 12626 3292
rect 12682 3290 12688 3292
rect 12442 3238 12444 3290
rect 12624 3238 12626 3290
rect 12380 3236 12386 3238
rect 12442 3236 12466 3238
rect 12522 3236 12546 3238
rect 12602 3236 12626 3238
rect 12682 3236 12688 3238
rect 12380 3227 12688 3236
rect 12380 2204 12688 2213
rect 12380 2202 12386 2204
rect 12442 2202 12466 2204
rect 12522 2202 12546 2204
rect 12602 2202 12626 2204
rect 12682 2202 12688 2204
rect 12442 2150 12444 2202
rect 12624 2150 12626 2202
rect 12380 2148 12386 2150
rect 12442 2148 12466 2150
rect 12522 2148 12546 2150
rect 12602 2148 12626 2150
rect 12682 2148 12688 2150
rect 12380 2139 12688 2148
rect 12728 1562 12756 3402
rect 12716 1556 12768 1562
rect 12716 1498 12768 1504
rect 12256 1352 12308 1358
rect 12256 1294 12308 1300
rect 12624 1352 12676 1358
rect 12992 1352 13044 1358
rect 12676 1312 12756 1340
rect 12624 1294 12676 1300
rect 12072 1216 12124 1222
rect 12072 1158 12124 1164
rect 11794 54 11928 82
rect 12162 82 12218 160
rect 12268 82 12296 1294
rect 12380 1116 12688 1125
rect 12380 1114 12386 1116
rect 12442 1114 12466 1116
rect 12522 1114 12546 1116
rect 12602 1114 12626 1116
rect 12682 1114 12688 1116
rect 12442 1062 12444 1114
rect 12624 1062 12626 1114
rect 12380 1060 12386 1062
rect 12442 1060 12466 1062
rect 12522 1060 12546 1062
rect 12602 1060 12626 1062
rect 12682 1060 12688 1062
rect 12380 1051 12688 1060
rect 12622 640 12678 649
rect 12622 575 12678 584
rect 12636 270 12664 575
rect 12624 264 12676 270
rect 12624 206 12676 212
rect 12162 54 12296 82
rect 12530 82 12586 160
rect 12728 82 12756 1312
rect 12992 1294 13044 1300
rect 13360 1352 13412 1358
rect 13360 1294 13412 1300
rect 12808 1216 12860 1222
rect 12808 1158 12860 1164
rect 12820 270 12848 1158
rect 12808 264 12860 270
rect 12808 206 12860 212
rect 12530 54 12756 82
rect 12898 82 12954 160
rect 13004 82 13032 1294
rect 13176 1216 13228 1222
rect 13176 1158 13228 1164
rect 13188 1057 13216 1158
rect 13174 1048 13230 1057
rect 13174 983 13230 992
rect 12898 54 13032 82
rect 13266 82 13322 160
rect 13372 82 13400 1294
rect 13464 134 13492 3470
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 14002 2952 14058 2961
rect 13832 2910 14002 2938
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13648 406 13676 2246
rect 13832 1358 13860 2910
rect 14002 2887 14058 2896
rect 15108 2372 15160 2378
rect 15108 2314 15160 2320
rect 14556 1896 14608 1902
rect 14556 1838 14608 1844
rect 13728 1352 13780 1358
rect 13728 1294 13780 1300
rect 13820 1352 13872 1358
rect 13820 1294 13872 1300
rect 14096 1352 14148 1358
rect 14096 1294 14148 1300
rect 13636 400 13688 406
rect 13636 342 13688 348
rect 13266 54 13400 82
rect 13452 128 13504 134
rect 13452 70 13504 76
rect 13634 82 13690 160
rect 13740 82 13768 1294
rect 13912 1216 13964 1222
rect 13912 1158 13964 1164
rect 13924 474 13952 1158
rect 13912 468 13964 474
rect 13912 410 13964 416
rect 13634 54 13768 82
rect 14002 82 14058 160
rect 14108 82 14136 1294
rect 14280 1216 14332 1222
rect 14280 1158 14332 1164
rect 14292 406 14320 1158
rect 14280 400 14332 406
rect 14280 342 14332 348
rect 14568 338 14596 1838
rect 14738 1456 14794 1465
rect 15120 1426 15148 2314
rect 15212 2106 15240 3334
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 15200 2100 15252 2106
rect 15200 2042 15252 2048
rect 15396 1562 15424 2450
rect 15948 2106 15976 3567
rect 16486 2136 16542 2145
rect 15936 2100 15988 2106
rect 16960 2106 16988 4422
rect 17314 4040 17370 4049
rect 17314 3975 17370 3984
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 16486 2071 16488 2080
rect 15936 2042 15988 2048
rect 16540 2071 16542 2080
rect 16948 2100 17000 2106
rect 16488 2042 16540 2048
rect 16948 2042 17000 2048
rect 16578 2000 16634 2009
rect 15752 1964 15804 1970
rect 15752 1906 15804 1912
rect 16028 1964 16080 1970
rect 16028 1906 16080 1912
rect 16304 1964 16356 1970
rect 16578 1935 16634 1944
rect 16764 1964 16816 1970
rect 16304 1906 16356 1912
rect 15764 1562 15792 1906
rect 15384 1556 15436 1562
rect 15384 1498 15436 1504
rect 15752 1556 15804 1562
rect 15752 1498 15804 1504
rect 14738 1391 14794 1400
rect 15108 1420 15160 1426
rect 14648 1352 14700 1358
rect 14648 1294 14700 1300
rect 14556 332 14608 338
rect 14556 274 14608 280
rect 14002 54 14136 82
rect 14370 82 14426 160
rect 14660 82 14688 1294
rect 14752 610 14780 1391
rect 15108 1362 15160 1368
rect 16040 1358 16068 1906
rect 16210 1864 16266 1873
rect 16210 1799 16266 1808
rect 16224 1766 16252 1799
rect 16212 1760 16264 1766
rect 16212 1702 16264 1708
rect 16316 1562 16344 1906
rect 16304 1556 16356 1562
rect 16304 1498 16356 1504
rect 16592 1494 16620 1935
rect 16764 1906 16816 1912
rect 17040 1964 17092 1970
rect 17040 1906 17092 1912
rect 16580 1488 16632 1494
rect 16580 1430 16632 1436
rect 15016 1352 15068 1358
rect 15016 1294 15068 1300
rect 15384 1352 15436 1358
rect 15384 1294 15436 1300
rect 15660 1352 15712 1358
rect 15660 1294 15712 1300
rect 15936 1352 15988 1358
rect 15936 1294 15988 1300
rect 16028 1352 16080 1358
rect 16028 1294 16080 1300
rect 16212 1352 16264 1358
rect 16212 1294 16264 1300
rect 16580 1352 16632 1358
rect 16580 1294 16632 1300
rect 14832 1216 14884 1222
rect 14832 1158 14884 1164
rect 14740 604 14792 610
rect 14740 546 14792 552
rect 14844 338 14872 1158
rect 14832 332 14884 338
rect 14832 274 14884 280
rect 14370 54 14688 82
rect 14738 82 14794 160
rect 15028 82 15056 1294
rect 15106 1184 15162 1193
rect 15106 1119 15162 1128
rect 15120 1018 15148 1119
rect 15108 1012 15160 1018
rect 15108 954 15160 960
rect 14738 54 15056 82
rect 15106 82 15162 160
rect 15396 82 15424 1294
rect 15106 54 15424 82
rect 15474 82 15530 160
rect 15672 82 15700 1294
rect 15474 54 15700 82
rect 15842 82 15898 160
rect 15948 82 15976 1294
rect 16224 160 16252 1294
rect 16592 160 16620 1294
rect 16776 1290 16804 1906
rect 17052 1562 17080 1906
rect 17144 1834 17172 2790
rect 17328 2106 17356 3975
rect 17420 2650 17448 8434
rect 18095 8188 18403 8197
rect 18095 8186 18101 8188
rect 18157 8186 18181 8188
rect 18237 8186 18261 8188
rect 18317 8186 18341 8188
rect 18397 8186 18403 8188
rect 18157 8134 18159 8186
rect 18339 8134 18341 8186
rect 18095 8132 18101 8134
rect 18157 8132 18181 8134
rect 18237 8132 18261 8134
rect 18317 8132 18341 8134
rect 18397 8132 18403 8134
rect 18095 8123 18403 8132
rect 18095 7100 18403 7109
rect 18095 7098 18101 7100
rect 18157 7098 18181 7100
rect 18237 7098 18261 7100
rect 18317 7098 18341 7100
rect 18397 7098 18403 7100
rect 18157 7046 18159 7098
rect 18339 7046 18341 7098
rect 18095 7044 18101 7046
rect 18157 7044 18181 7046
rect 18237 7044 18261 7046
rect 18317 7044 18341 7046
rect 18397 7044 18403 7046
rect 18095 7035 18403 7044
rect 18095 6012 18403 6021
rect 18095 6010 18101 6012
rect 18157 6010 18181 6012
rect 18237 6010 18261 6012
rect 18317 6010 18341 6012
rect 18397 6010 18403 6012
rect 18157 5958 18159 6010
rect 18339 5958 18341 6010
rect 18095 5956 18101 5958
rect 18157 5956 18181 5958
rect 18237 5956 18261 5958
rect 18317 5956 18341 5958
rect 18397 5956 18403 5958
rect 18095 5947 18403 5956
rect 18095 4924 18403 4933
rect 18095 4922 18101 4924
rect 18157 4922 18181 4924
rect 18237 4922 18261 4924
rect 18317 4922 18341 4924
rect 18397 4922 18403 4924
rect 18157 4870 18159 4922
rect 18339 4870 18341 4922
rect 18095 4868 18101 4870
rect 18157 4868 18181 4870
rect 18237 4868 18261 4870
rect 18317 4868 18341 4870
rect 18397 4868 18403 4870
rect 18095 4859 18403 4868
rect 17774 4176 17830 4185
rect 17774 4111 17830 4120
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17316 2100 17368 2106
rect 17316 2042 17368 2048
rect 17224 2032 17276 2038
rect 17224 1974 17276 1980
rect 17132 1828 17184 1834
rect 17132 1770 17184 1776
rect 17236 1562 17264 1974
rect 17316 1964 17368 1970
rect 17316 1906 17368 1912
rect 17328 1562 17356 1906
rect 17512 1766 17540 2994
rect 17788 1970 17816 4111
rect 18095 3836 18403 3845
rect 18095 3834 18101 3836
rect 18157 3834 18181 3836
rect 18237 3834 18261 3836
rect 18317 3834 18341 3836
rect 18397 3834 18403 3836
rect 18157 3782 18159 3834
rect 18339 3782 18341 3834
rect 18095 3780 18101 3782
rect 18157 3780 18181 3782
rect 18237 3780 18261 3782
rect 18317 3780 18341 3782
rect 18397 3780 18403 3782
rect 18095 3771 18403 3780
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 18878 2816 18934 2825
rect 18095 2748 18403 2757
rect 18878 2751 18934 2760
rect 18095 2746 18101 2748
rect 18157 2746 18181 2748
rect 18237 2746 18261 2748
rect 18317 2746 18341 2748
rect 18397 2746 18403 2748
rect 18157 2694 18159 2746
rect 18339 2694 18341 2746
rect 18095 2692 18101 2694
rect 18157 2692 18181 2694
rect 18237 2692 18261 2694
rect 18317 2692 18341 2694
rect 18397 2692 18403 2694
rect 18095 2683 18403 2692
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 17972 2106 18000 2382
rect 18892 2106 18920 2751
rect 19352 2360 19380 2926
rect 19628 2650 19656 8434
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 19352 2332 19472 2360
rect 19338 2272 19394 2281
rect 19338 2207 19394 2216
rect 17960 2100 18012 2106
rect 17960 2042 18012 2048
rect 18880 2100 18932 2106
rect 18880 2042 18932 2048
rect 17776 1964 17828 1970
rect 17776 1906 17828 1912
rect 17960 1964 18012 1970
rect 17960 1906 18012 1912
rect 18696 1964 18748 1970
rect 18696 1906 18748 1912
rect 18880 1964 18932 1970
rect 18880 1906 18932 1912
rect 17684 1896 17736 1902
rect 17684 1838 17736 1844
rect 17500 1760 17552 1766
rect 17500 1702 17552 1708
rect 17696 1562 17724 1838
rect 17040 1556 17092 1562
rect 17040 1498 17092 1504
rect 17224 1556 17276 1562
rect 17224 1498 17276 1504
rect 17316 1556 17368 1562
rect 17316 1498 17368 1504
rect 17684 1556 17736 1562
rect 17684 1498 17736 1504
rect 16856 1352 16908 1358
rect 16856 1294 16908 1300
rect 17132 1352 17184 1358
rect 17408 1352 17460 1358
rect 17184 1312 17356 1340
rect 17132 1294 17184 1300
rect 16764 1284 16816 1290
rect 16764 1226 16816 1232
rect 15842 54 15976 82
rect 9954 0 10010 54
rect 10322 0 10378 54
rect 10690 0 10746 54
rect 11058 0 11114 54
rect 11426 0 11482 54
rect 11794 0 11850 54
rect 12162 0 12218 54
rect 12530 0 12586 54
rect 12898 0 12954 54
rect 13266 0 13322 54
rect 13634 0 13690 54
rect 14002 0 14058 54
rect 14370 0 14426 54
rect 14738 0 14794 54
rect 15106 0 15162 54
rect 15474 0 15530 54
rect 15842 0 15898 54
rect 16210 0 16266 160
rect 16578 0 16634 160
rect 16868 82 16896 1294
rect 17224 876 17276 882
rect 17224 818 17276 824
rect 17236 746 17264 818
rect 17224 740 17276 746
rect 17224 682 17276 688
rect 17328 160 17356 1312
rect 17408 1294 17460 1300
rect 17684 1352 17736 1358
rect 17736 1312 17816 1340
rect 17684 1294 17736 1300
rect 16946 82 17002 160
rect 16868 54 17002 82
rect 16946 0 17002 54
rect 17314 0 17370 160
rect 17420 82 17448 1294
rect 17498 1048 17554 1057
rect 17498 983 17554 992
rect 17512 950 17540 983
rect 17500 944 17552 950
rect 17500 886 17552 892
rect 17604 190 17724 218
rect 17604 82 17632 190
rect 17696 160 17724 190
rect 17420 54 17632 82
rect 17682 0 17738 160
rect 17788 82 17816 1312
rect 17972 1222 18000 1906
rect 18512 1760 18564 1766
rect 18512 1702 18564 1708
rect 18095 1660 18403 1669
rect 18095 1658 18101 1660
rect 18157 1658 18181 1660
rect 18237 1658 18261 1660
rect 18317 1658 18341 1660
rect 18397 1658 18403 1660
rect 18157 1606 18159 1658
rect 18339 1606 18341 1658
rect 18095 1604 18101 1606
rect 18157 1604 18181 1606
rect 18237 1604 18261 1606
rect 18317 1604 18341 1606
rect 18397 1604 18403 1606
rect 18095 1595 18403 1604
rect 18524 1601 18552 1702
rect 18510 1592 18566 1601
rect 18708 1562 18736 1906
rect 18510 1527 18566 1536
rect 18696 1556 18748 1562
rect 18696 1498 18748 1504
rect 18236 1352 18288 1358
rect 18236 1294 18288 1300
rect 18512 1352 18564 1358
rect 18892 1329 18920 1906
rect 19352 1902 19380 2207
rect 19444 2106 19472 2332
rect 19536 2122 19564 2586
rect 19996 2446 20024 3062
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 20088 2446 20116 2926
rect 20352 2916 20404 2922
rect 20352 2858 20404 2864
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20364 2446 20392 2858
rect 20640 2650 20668 2858
rect 21284 2650 21312 8366
rect 21362 3768 21418 3777
rect 21362 3703 21418 3712
rect 21376 2961 21404 3703
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21640 3120 21692 3126
rect 21640 3062 21692 3068
rect 21362 2952 21418 2961
rect 21362 2887 21418 2896
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 21548 2576 21600 2582
rect 20534 2544 20590 2553
rect 21548 2518 21600 2524
rect 20534 2479 20590 2488
rect 20628 2508 20680 2514
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 20352 2440 20404 2446
rect 20352 2382 20404 2388
rect 19892 2372 19944 2378
rect 19892 2314 19944 2320
rect 19432 2100 19484 2106
rect 19536 2094 19840 2122
rect 19432 2042 19484 2048
rect 19616 2032 19668 2038
rect 19616 1974 19668 1980
rect 19706 2000 19762 2009
rect 19432 1964 19484 1970
rect 19432 1906 19484 1912
rect 19524 1964 19576 1970
rect 19524 1906 19576 1912
rect 19340 1896 19392 1902
rect 19340 1838 19392 1844
rect 19156 1760 19208 1766
rect 18970 1728 19026 1737
rect 19156 1702 19208 1708
rect 18970 1663 19026 1672
rect 18512 1294 18564 1300
rect 18878 1320 18934 1329
rect 17960 1216 18012 1222
rect 17960 1158 18012 1164
rect 18248 542 18276 1294
rect 18420 1284 18472 1290
rect 18420 1226 18472 1232
rect 18236 536 18288 542
rect 18236 478 18288 484
rect 18432 160 18460 1226
rect 18524 814 18552 1294
rect 18878 1255 18934 1264
rect 18984 882 19012 1663
rect 19168 1290 19196 1702
rect 19248 1420 19300 1426
rect 19300 1380 19380 1408
rect 19248 1362 19300 1368
rect 19156 1284 19208 1290
rect 19156 1226 19208 1232
rect 19064 1216 19116 1222
rect 19064 1158 19116 1164
rect 18972 876 19024 882
rect 18972 818 19024 824
rect 18512 808 18564 814
rect 18512 750 18564 756
rect 18788 536 18840 542
rect 18788 478 18840 484
rect 18800 160 18828 478
rect 18050 82 18106 160
rect 17788 54 18106 82
rect 18050 0 18106 54
rect 18418 0 18474 160
rect 18786 0 18842 160
rect 19076 105 19104 1158
rect 19156 808 19208 814
rect 19156 750 19208 756
rect 19352 762 19380 1380
rect 19444 950 19472 1906
rect 19536 1562 19564 1906
rect 19524 1556 19576 1562
rect 19524 1498 19576 1504
rect 19432 944 19484 950
rect 19432 886 19484 892
rect 19628 785 19656 1974
rect 19706 1935 19762 1944
rect 19720 1902 19748 1935
rect 19708 1896 19760 1902
rect 19708 1838 19760 1844
rect 19812 1494 19840 2094
rect 19904 2009 19932 2314
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 19984 2100 20036 2106
rect 19984 2042 20036 2048
rect 20168 2100 20220 2106
rect 20168 2042 20220 2048
rect 19890 2000 19946 2009
rect 19890 1935 19946 1944
rect 19708 1488 19760 1494
rect 19708 1430 19760 1436
rect 19800 1488 19852 1494
rect 19800 1430 19852 1436
rect 19720 1329 19748 1430
rect 19996 1358 20024 2042
rect 20180 1494 20208 2042
rect 20258 2000 20314 2009
rect 20456 1970 20484 2246
rect 20548 2106 20576 2479
rect 20628 2450 20680 2456
rect 20536 2100 20588 2106
rect 20536 2042 20588 2048
rect 20258 1935 20260 1944
rect 20312 1935 20314 1944
rect 20352 1964 20404 1970
rect 20260 1906 20312 1912
rect 20352 1906 20404 1912
rect 20444 1964 20496 1970
rect 20444 1906 20496 1912
rect 20168 1488 20220 1494
rect 20168 1430 20220 1436
rect 19984 1352 20036 1358
rect 19706 1320 19762 1329
rect 19984 1294 20036 1300
rect 19706 1255 19762 1264
rect 19800 1284 19852 1290
rect 19852 1244 19932 1272
rect 19800 1226 19852 1232
rect 19614 776 19670 785
rect 19168 160 19196 750
rect 19352 734 19564 762
rect 19536 160 19564 734
rect 19614 711 19670 720
rect 19904 160 19932 1244
rect 20076 1216 20128 1222
rect 20128 1176 20300 1204
rect 20076 1158 20128 1164
rect 20272 160 20300 1176
rect 20364 338 20392 1906
rect 20444 1760 20496 1766
rect 20444 1702 20496 1708
rect 20456 1562 20484 1702
rect 20640 1578 20668 2450
rect 21560 2310 21588 2518
rect 21652 2446 21680 3062
rect 21640 2440 21692 2446
rect 21640 2382 21692 2388
rect 21744 2378 21772 3470
rect 22112 2650 22140 8434
rect 22204 2650 22232 8910
rect 22834 2952 22890 2961
rect 22834 2887 22890 2896
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22848 2446 22876 2887
rect 23492 2650 23520 8978
rect 23810 8732 24118 8741
rect 23810 8730 23816 8732
rect 23872 8730 23896 8732
rect 23952 8730 23976 8732
rect 24032 8730 24056 8732
rect 24112 8730 24118 8732
rect 23872 8678 23874 8730
rect 24054 8678 24056 8730
rect 23810 8676 23816 8678
rect 23872 8676 23896 8678
rect 23952 8676 23976 8678
rect 24032 8676 24056 8678
rect 24112 8676 24118 8678
rect 23810 8667 24118 8676
rect 24228 8634 24256 9846
rect 26146 9840 26202 10000
rect 28354 9840 28410 10000
rect 30562 9840 30618 10000
rect 32770 9840 32826 10000
rect 34978 9840 35034 10000
rect 37186 9840 37242 10000
rect 39394 9840 39450 10000
rect 41602 9840 41658 10000
rect 43810 9840 43866 10000
rect 46018 9840 46074 10000
rect 25320 8900 25372 8906
rect 25320 8842 25372 8848
rect 24216 8628 24268 8634
rect 24216 8570 24268 8576
rect 24308 8560 24360 8566
rect 24308 8502 24360 8508
rect 23810 7644 24118 7653
rect 23810 7642 23816 7644
rect 23872 7642 23896 7644
rect 23952 7642 23976 7644
rect 24032 7642 24056 7644
rect 24112 7642 24118 7644
rect 23872 7590 23874 7642
rect 24054 7590 24056 7642
rect 23810 7588 23816 7590
rect 23872 7588 23896 7590
rect 23952 7588 23976 7590
rect 24032 7588 24056 7590
rect 24112 7588 24118 7590
rect 23810 7579 24118 7588
rect 23810 6556 24118 6565
rect 23810 6554 23816 6556
rect 23872 6554 23896 6556
rect 23952 6554 23976 6556
rect 24032 6554 24056 6556
rect 24112 6554 24118 6556
rect 23872 6502 23874 6554
rect 24054 6502 24056 6554
rect 23810 6500 23816 6502
rect 23872 6500 23896 6502
rect 23952 6500 23976 6502
rect 24032 6500 24056 6502
rect 24112 6500 24118 6502
rect 23810 6491 24118 6500
rect 23810 5468 24118 5477
rect 23810 5466 23816 5468
rect 23872 5466 23896 5468
rect 23952 5466 23976 5468
rect 24032 5466 24056 5468
rect 24112 5466 24118 5468
rect 23872 5414 23874 5466
rect 24054 5414 24056 5466
rect 23810 5412 23816 5414
rect 23872 5412 23896 5414
rect 23952 5412 23976 5414
rect 24032 5412 24056 5414
rect 24112 5412 24118 5414
rect 23810 5403 24118 5412
rect 23810 4380 24118 4389
rect 23810 4378 23816 4380
rect 23872 4378 23896 4380
rect 23952 4378 23976 4380
rect 24032 4378 24056 4380
rect 24112 4378 24118 4380
rect 23872 4326 23874 4378
rect 24054 4326 24056 4378
rect 23810 4324 23816 4326
rect 23872 4324 23896 4326
rect 23952 4324 23976 4326
rect 24032 4324 24056 4326
rect 24112 4324 24118 4326
rect 23810 4315 24118 4324
rect 23810 3292 24118 3301
rect 23810 3290 23816 3292
rect 23872 3290 23896 3292
rect 23952 3290 23976 3292
rect 24032 3290 24056 3292
rect 24112 3290 24118 3292
rect 23872 3238 23874 3290
rect 24054 3238 24056 3290
rect 23810 3236 23816 3238
rect 23872 3236 23896 3238
rect 23952 3236 23976 3238
rect 24032 3236 24056 3238
rect 24112 3236 24118 3238
rect 23810 3227 24118 3236
rect 24320 2650 24348 8502
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 24308 2644 24360 2650
rect 24308 2586 24360 2592
rect 24688 2582 24716 8298
rect 24768 2848 24820 2854
rect 24768 2790 24820 2796
rect 24676 2576 24728 2582
rect 24676 2518 24728 2524
rect 22836 2440 22888 2446
rect 22836 2382 22888 2388
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 23572 2440 23624 2446
rect 24308 2440 24360 2446
rect 23572 2382 23624 2388
rect 23662 2408 23718 2417
rect 21732 2372 21784 2378
rect 21732 2314 21784 2320
rect 21088 2304 21140 2310
rect 21088 2246 21140 2252
rect 21548 2304 21600 2310
rect 22376 2304 22428 2310
rect 21548 2246 21600 2252
rect 21638 2272 21694 2281
rect 20812 1760 20864 1766
rect 20864 1720 21036 1748
rect 20812 1702 20864 1708
rect 20444 1556 20496 1562
rect 20444 1498 20496 1504
rect 20548 1550 20668 1578
rect 20548 1426 20576 1550
rect 20536 1420 20588 1426
rect 20536 1362 20588 1368
rect 20628 1420 20680 1426
rect 20628 1362 20680 1368
rect 20536 876 20588 882
rect 20536 818 20588 824
rect 20548 542 20576 818
rect 20536 536 20588 542
rect 20536 478 20588 484
rect 20352 332 20404 338
rect 20352 274 20404 280
rect 20640 160 20668 1362
rect 21008 160 21036 1720
rect 21100 1358 21128 2246
rect 22376 2246 22428 2252
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 21638 2207 21694 2216
rect 21652 1970 21680 2207
rect 22388 1970 22416 2246
rect 22572 1970 22600 2246
rect 21364 1964 21416 1970
rect 21364 1906 21416 1912
rect 21640 1964 21692 1970
rect 21640 1906 21692 1912
rect 22100 1964 22152 1970
rect 22100 1906 22152 1912
rect 22376 1964 22428 1970
rect 22376 1906 22428 1912
rect 22560 1964 22612 1970
rect 22560 1906 22612 1912
rect 21376 1465 21404 1906
rect 21824 1828 21876 1834
rect 21824 1770 21876 1776
rect 21456 1488 21508 1494
rect 21362 1456 21418 1465
rect 21456 1430 21508 1436
rect 21362 1391 21418 1400
rect 21088 1352 21140 1358
rect 21088 1294 21140 1300
rect 21180 1216 21232 1222
rect 21232 1176 21404 1204
rect 21180 1158 21232 1164
rect 21376 160 21404 1176
rect 21468 649 21496 1430
rect 21548 1216 21600 1222
rect 21548 1158 21600 1164
rect 21454 640 21510 649
rect 21454 575 21510 584
rect 19062 96 19118 105
rect 19062 31 19118 40
rect 19154 0 19210 160
rect 19522 0 19578 160
rect 19890 0 19946 160
rect 20258 0 20314 160
rect 20626 0 20682 160
rect 20994 0 21050 160
rect 21362 0 21418 160
rect 21560 82 21588 1158
rect 21836 1018 21864 1770
rect 21916 1760 21968 1766
rect 22112 1737 22140 1906
rect 22652 1760 22704 1766
rect 21916 1702 21968 1708
rect 22098 1728 22154 1737
rect 21928 1222 21956 1702
rect 22098 1663 22154 1672
rect 22480 1720 22652 1748
rect 22008 1352 22060 1358
rect 22284 1352 22336 1358
rect 22008 1294 22060 1300
rect 22112 1312 22284 1340
rect 21916 1216 21968 1222
rect 22020 1193 22048 1294
rect 21916 1158 21968 1164
rect 22006 1184 22062 1193
rect 22006 1119 22062 1128
rect 21824 1012 21876 1018
rect 21824 954 21876 960
rect 22112 160 22140 1312
rect 22284 1294 22336 1300
rect 22480 160 22508 1720
rect 22652 1702 22704 1708
rect 23400 1494 23428 2382
rect 23584 2106 23612 2382
rect 24308 2382 24360 2388
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 23662 2343 23718 2352
rect 23572 2100 23624 2106
rect 23572 2042 23624 2048
rect 23676 1970 23704 2343
rect 24216 2304 24268 2310
rect 24216 2246 24268 2252
rect 23810 2204 24118 2213
rect 23810 2202 23816 2204
rect 23872 2202 23896 2204
rect 23952 2202 23976 2204
rect 24032 2202 24056 2204
rect 24112 2202 24118 2204
rect 23872 2150 23874 2202
rect 24054 2150 24056 2202
rect 23810 2148 23816 2150
rect 23872 2148 23896 2150
rect 23952 2148 23976 2150
rect 24032 2148 24056 2150
rect 24112 2148 24118 2150
rect 23810 2139 24118 2148
rect 23664 1964 23716 1970
rect 23664 1906 23716 1912
rect 23480 1828 23532 1834
rect 23480 1770 23532 1776
rect 23388 1488 23440 1494
rect 23388 1430 23440 1436
rect 23492 1358 23520 1770
rect 23756 1760 23808 1766
rect 23584 1720 23756 1748
rect 23480 1352 23532 1358
rect 23480 1294 23532 1300
rect 23020 1216 23072 1222
rect 22848 1176 23020 1204
rect 22848 160 22876 1176
rect 23388 1216 23440 1222
rect 23020 1158 23072 1164
rect 23216 1176 23388 1204
rect 23216 160 23244 1176
rect 23388 1158 23440 1164
rect 23584 160 23612 1720
rect 23756 1702 23808 1708
rect 24032 1760 24084 1766
rect 24032 1702 24084 1708
rect 24044 1358 24072 1702
rect 24228 1358 24256 2246
rect 24320 2106 24348 2382
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 24398 2136 24454 2145
rect 24308 2100 24360 2106
rect 24398 2071 24454 2080
rect 24308 2042 24360 2048
rect 24412 1562 24440 2071
rect 24504 1970 24532 2246
rect 24492 1964 24544 1970
rect 24492 1906 24544 1912
rect 24596 1834 24624 2382
rect 24676 2100 24728 2106
rect 24676 2042 24728 2048
rect 24584 1828 24636 1834
rect 24584 1770 24636 1776
rect 24688 1714 24716 2042
rect 24780 1970 24808 2790
rect 24872 2650 24900 8434
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 25240 2774 25268 3334
rect 25148 2746 25268 2774
rect 24860 2644 24912 2650
rect 24860 2586 24912 2592
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 24952 2372 25004 2378
rect 24952 2314 25004 2320
rect 24768 1964 24820 1970
rect 24768 1906 24820 1912
rect 24964 1766 24992 2314
rect 25056 2106 25084 2382
rect 25044 2100 25096 2106
rect 25044 2042 25096 2048
rect 25148 1970 25176 2746
rect 25332 2650 25360 8842
rect 26160 8634 26188 9840
rect 28368 8634 28396 9840
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 28356 8628 28408 8634
rect 28356 8570 28408 8576
rect 26516 8492 26568 8498
rect 26516 8434 26568 8440
rect 28448 8492 28500 8498
rect 28448 8434 28500 8440
rect 26424 4548 26476 4554
rect 26424 4490 26476 4496
rect 25962 3088 26018 3097
rect 25962 3023 26018 3032
rect 26146 3088 26202 3097
rect 26146 3023 26202 3032
rect 25320 2644 25372 2650
rect 25320 2586 25372 2592
rect 25976 2446 26004 3023
rect 26160 2825 26188 3023
rect 26146 2816 26202 2825
rect 26146 2751 26202 2760
rect 25872 2440 25924 2446
rect 25872 2382 25924 2388
rect 25964 2440 26016 2446
rect 25964 2382 26016 2388
rect 25884 2106 25912 2382
rect 25872 2100 25924 2106
rect 25872 2042 25924 2048
rect 26436 1970 26464 4490
rect 26528 2650 26556 8434
rect 27436 4276 27488 4282
rect 27436 4218 27488 4224
rect 26516 2644 26568 2650
rect 26516 2586 26568 2592
rect 27344 2440 27396 2446
rect 26606 2408 26662 2417
rect 27344 2382 27396 2388
rect 26606 2343 26662 2352
rect 26976 2372 27028 2378
rect 26516 2304 26568 2310
rect 26516 2246 26568 2252
rect 25136 1964 25188 1970
rect 25136 1906 25188 1912
rect 25412 1964 25464 1970
rect 25412 1906 25464 1912
rect 25688 1964 25740 1970
rect 25688 1906 25740 1912
rect 26424 1964 26476 1970
rect 26424 1906 26476 1912
rect 24860 1760 24912 1766
rect 24688 1686 24808 1714
rect 24860 1702 24912 1708
rect 24952 1760 25004 1766
rect 24952 1702 25004 1708
rect 24400 1556 24452 1562
rect 24400 1498 24452 1504
rect 24676 1556 24728 1562
rect 24676 1498 24728 1504
rect 24032 1352 24084 1358
rect 24032 1294 24084 1300
rect 24216 1352 24268 1358
rect 24216 1294 24268 1300
rect 24306 1320 24362 1329
rect 24306 1255 24362 1264
rect 24124 1216 24176 1222
rect 24176 1176 24256 1204
rect 24124 1158 24176 1164
rect 23810 1116 24118 1125
rect 23810 1114 23816 1116
rect 23872 1114 23896 1116
rect 23952 1114 23976 1116
rect 24032 1114 24056 1116
rect 24112 1114 24118 1116
rect 23872 1062 23874 1114
rect 24054 1062 24056 1114
rect 23810 1060 23816 1062
rect 23872 1060 23896 1062
rect 23952 1060 23976 1062
rect 24032 1060 24056 1062
rect 24112 1060 24118 1062
rect 23810 1051 24118 1060
rect 23952 190 24072 218
rect 23952 160 23980 190
rect 21730 82 21786 160
rect 21560 54 21786 82
rect 21730 0 21786 54
rect 22098 0 22154 160
rect 22466 0 22522 160
rect 22834 0 22890 160
rect 23202 0 23258 160
rect 23570 0 23626 160
rect 23938 0 23994 160
rect 24044 82 24072 190
rect 24228 82 24256 1176
rect 24320 950 24348 1255
rect 24584 1216 24636 1222
rect 24584 1158 24636 1164
rect 24308 944 24360 950
rect 24308 886 24360 892
rect 24044 54 24256 82
rect 24306 82 24362 160
rect 24596 82 24624 1158
rect 24688 160 24716 1498
rect 24780 1358 24808 1686
rect 24768 1352 24820 1358
rect 24768 1294 24820 1300
rect 24872 1290 24900 1702
rect 25424 1426 25452 1906
rect 25412 1420 25464 1426
rect 25412 1362 25464 1368
rect 24860 1284 24912 1290
rect 24860 1226 24912 1232
rect 25044 1216 25096 1222
rect 25596 1216 25648 1222
rect 25044 1158 25096 1164
rect 25424 1176 25596 1204
rect 25056 160 25084 1158
rect 25424 160 25452 1176
rect 25596 1158 25648 1164
rect 25700 338 25728 1906
rect 26056 1760 26108 1766
rect 26056 1702 26108 1708
rect 26240 1760 26292 1766
rect 26240 1702 26292 1708
rect 25688 332 25740 338
rect 25688 274 25740 280
rect 24306 54 24624 82
rect 24306 0 24362 54
rect 24674 0 24730 160
rect 25042 0 25098 160
rect 25410 0 25466 160
rect 25778 82 25834 160
rect 26068 82 26096 1702
rect 26148 1556 26200 1562
rect 26148 1498 26200 1504
rect 26160 160 26188 1498
rect 26252 1358 26280 1702
rect 26528 1358 26556 2246
rect 26620 1902 26648 2343
rect 26976 2314 27028 2320
rect 26988 2106 27016 2314
rect 27160 2304 27212 2310
rect 27160 2246 27212 2252
rect 27172 2106 27200 2246
rect 26976 2100 27028 2106
rect 26976 2042 27028 2048
rect 27160 2100 27212 2106
rect 27160 2042 27212 2048
rect 26884 1964 26936 1970
rect 27252 1964 27304 1970
rect 26936 1924 27252 1952
rect 26884 1906 26936 1912
rect 27252 1906 27304 1912
rect 26608 1896 26660 1902
rect 26608 1838 26660 1844
rect 26792 1828 26844 1834
rect 26792 1770 26844 1776
rect 26240 1352 26292 1358
rect 26240 1294 26292 1300
rect 26516 1352 26568 1358
rect 26516 1294 26568 1300
rect 26516 1216 26568 1222
rect 26516 1158 26568 1164
rect 26528 160 26556 1158
rect 25778 54 26096 82
rect 25778 0 25834 54
rect 26146 0 26202 160
rect 26514 0 26570 160
rect 26804 134 26832 1770
rect 27252 1760 27304 1766
rect 27252 1702 27304 1708
rect 27264 1358 27292 1702
rect 27252 1352 27304 1358
rect 27252 1294 27304 1300
rect 27252 1216 27304 1222
rect 27172 1176 27252 1204
rect 26792 128 26844 134
rect 26792 70 26844 76
rect 26882 82 26938 160
rect 27172 82 27200 1176
rect 27252 1158 27304 1164
rect 27356 474 27384 2382
rect 27448 1970 27476 4218
rect 27712 4208 27764 4214
rect 27712 4150 27764 4156
rect 27724 1970 27752 4150
rect 28262 3768 28318 3777
rect 28262 3703 28318 3712
rect 28172 3188 28224 3194
rect 28172 3130 28224 3136
rect 27804 2440 27856 2446
rect 27804 2382 27856 2388
rect 27436 1964 27488 1970
rect 27436 1906 27488 1912
rect 27712 1964 27764 1970
rect 27712 1906 27764 1912
rect 27528 1760 27580 1766
rect 27528 1702 27580 1708
rect 27540 1358 27568 1702
rect 27620 1556 27672 1562
rect 27620 1498 27672 1504
rect 27528 1352 27580 1358
rect 27528 1294 27580 1300
rect 27632 1204 27660 1498
rect 27540 1176 27660 1204
rect 27344 468 27396 474
rect 27344 410 27396 416
rect 26882 54 27200 82
rect 27250 82 27306 160
rect 27540 82 27568 1176
rect 27816 270 27844 2382
rect 28080 2304 28132 2310
rect 28080 2246 28132 2252
rect 28184 2258 28212 3130
rect 28276 2446 28304 3703
rect 28460 2650 28488 8434
rect 28448 2644 28500 2650
rect 28448 2586 28500 2592
rect 28908 2644 28960 2650
rect 28908 2586 28960 2592
rect 28264 2440 28316 2446
rect 28264 2382 28316 2388
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 27988 1760 28040 1766
rect 27988 1702 28040 1708
rect 28000 1358 28028 1702
rect 27988 1352 28040 1358
rect 27988 1294 28040 1300
rect 28092 1290 28120 2246
rect 28184 2230 28304 2258
rect 28276 1970 28304 2230
rect 28172 1964 28224 1970
rect 28172 1906 28224 1912
rect 28264 1964 28316 1970
rect 28264 1906 28316 1912
rect 28080 1284 28132 1290
rect 28080 1226 28132 1232
rect 27988 1216 28040 1222
rect 27908 1176 27988 1204
rect 27804 264 27856 270
rect 27804 206 27856 212
rect 27250 54 27568 82
rect 27618 82 27674 160
rect 27908 82 27936 1176
rect 27988 1158 28040 1164
rect 28184 406 28212 1906
rect 28264 1760 28316 1766
rect 28264 1702 28316 1708
rect 28172 400 28224 406
rect 28172 342 28224 348
rect 28000 190 28120 218
rect 28000 160 28028 190
rect 27618 54 27936 82
rect 26882 0 26938 54
rect 27250 0 27306 54
rect 27618 0 27674 54
rect 27986 0 28042 160
rect 28092 82 28120 190
rect 28276 82 28304 1702
rect 28552 814 28580 2382
rect 28920 2106 28948 2586
rect 29000 2304 29052 2310
rect 29000 2246 29052 2252
rect 28908 2100 28960 2106
rect 28908 2042 28960 2048
rect 28644 1562 28764 1578
rect 28644 1556 28776 1562
rect 28644 1550 28724 1556
rect 28540 808 28592 814
rect 28540 750 28592 756
rect 28356 740 28408 746
rect 28356 682 28408 688
rect 28368 406 28396 682
rect 28356 400 28408 406
rect 28356 342 28408 348
rect 28092 54 28304 82
rect 28354 82 28410 160
rect 28644 82 28672 1550
rect 28724 1498 28776 1504
rect 28908 1488 28960 1494
rect 28908 1430 28960 1436
rect 28354 54 28672 82
rect 28722 82 28778 160
rect 28920 82 28948 1430
rect 29012 1358 29040 2246
rect 29196 2106 29224 8774
rect 30576 8634 30604 9840
rect 32784 8634 32812 9840
rect 34992 8634 35020 9840
rect 35240 8732 35548 8741
rect 35240 8730 35246 8732
rect 35302 8730 35326 8732
rect 35382 8730 35406 8732
rect 35462 8730 35486 8732
rect 35542 8730 35548 8732
rect 35302 8678 35304 8730
rect 35484 8678 35486 8730
rect 35240 8676 35246 8678
rect 35302 8676 35326 8678
rect 35382 8676 35406 8678
rect 35462 8676 35486 8678
rect 35542 8676 35548 8678
rect 35240 8667 35548 8676
rect 37200 8634 37228 9840
rect 39408 8634 39436 9840
rect 41616 8634 41644 9840
rect 43824 8634 43852 9840
rect 46032 8634 46060 9840
rect 46670 8732 46978 8741
rect 46670 8730 46676 8732
rect 46732 8730 46756 8732
rect 46812 8730 46836 8732
rect 46892 8730 46916 8732
rect 46972 8730 46978 8732
rect 46732 8678 46734 8730
rect 46914 8678 46916 8730
rect 46670 8676 46676 8678
rect 46732 8676 46756 8678
rect 46812 8676 46836 8678
rect 46892 8676 46916 8678
rect 46972 8676 46978 8678
rect 46670 8667 46978 8676
rect 30564 8628 30616 8634
rect 30564 8570 30616 8576
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 34980 8628 35032 8634
rect 34980 8570 35032 8576
rect 37188 8628 37240 8634
rect 37188 8570 37240 8576
rect 39396 8628 39448 8634
rect 39396 8570 39448 8576
rect 41604 8628 41656 8634
rect 41604 8570 41656 8576
rect 43812 8628 43864 8634
rect 43812 8570 43864 8576
rect 46020 8628 46072 8634
rect 46020 8570 46072 8576
rect 30656 8492 30708 8498
rect 30656 8434 30708 8440
rect 33140 8492 33192 8498
rect 33140 8434 33192 8440
rect 35072 8492 35124 8498
rect 35072 8434 35124 8440
rect 37372 8492 37424 8498
rect 37372 8434 37424 8440
rect 41696 8492 41748 8498
rect 41696 8434 41748 8440
rect 45008 8492 45060 8498
rect 45008 8434 45060 8440
rect 46112 8492 46164 8498
rect 46112 8434 46164 8440
rect 29525 8188 29833 8197
rect 29525 8186 29531 8188
rect 29587 8186 29611 8188
rect 29667 8186 29691 8188
rect 29747 8186 29771 8188
rect 29827 8186 29833 8188
rect 29587 8134 29589 8186
rect 29769 8134 29771 8186
rect 29525 8132 29531 8134
rect 29587 8132 29611 8134
rect 29667 8132 29691 8134
rect 29747 8132 29771 8134
rect 29827 8132 29833 8134
rect 29525 8123 29833 8132
rect 29525 7100 29833 7109
rect 29525 7098 29531 7100
rect 29587 7098 29611 7100
rect 29667 7098 29691 7100
rect 29747 7098 29771 7100
rect 29827 7098 29833 7100
rect 29587 7046 29589 7098
rect 29769 7046 29771 7098
rect 29525 7044 29531 7046
rect 29587 7044 29611 7046
rect 29667 7044 29691 7046
rect 29747 7044 29771 7046
rect 29827 7044 29833 7046
rect 29525 7035 29833 7044
rect 30668 6914 30696 8434
rect 30668 6886 30880 6914
rect 29525 6012 29833 6021
rect 29525 6010 29531 6012
rect 29587 6010 29611 6012
rect 29667 6010 29691 6012
rect 29747 6010 29771 6012
rect 29827 6010 29833 6012
rect 29587 5958 29589 6010
rect 29769 5958 29771 6010
rect 29525 5956 29531 5958
rect 29587 5956 29611 5958
rect 29667 5956 29691 5958
rect 29747 5956 29771 5958
rect 29827 5956 29833 5958
rect 29525 5947 29833 5956
rect 29525 4924 29833 4933
rect 29525 4922 29531 4924
rect 29587 4922 29611 4924
rect 29667 4922 29691 4924
rect 29747 4922 29771 4924
rect 29827 4922 29833 4924
rect 29587 4870 29589 4922
rect 29769 4870 29771 4922
rect 29525 4868 29531 4870
rect 29587 4868 29611 4870
rect 29667 4868 29691 4870
rect 29747 4868 29771 4870
rect 29827 4868 29833 4870
rect 29525 4859 29833 4868
rect 29525 3836 29833 3845
rect 29525 3834 29531 3836
rect 29587 3834 29611 3836
rect 29667 3834 29691 3836
rect 29747 3834 29771 3836
rect 29827 3834 29833 3836
rect 29587 3782 29589 3834
rect 29769 3782 29771 3834
rect 29525 3780 29531 3782
rect 29587 3780 29611 3782
rect 29667 3780 29691 3782
rect 29747 3780 29771 3782
rect 29827 3780 29833 3782
rect 29525 3771 29833 3780
rect 30562 3496 30618 3505
rect 29368 3460 29420 3466
rect 30562 3431 30618 3440
rect 29368 3402 29420 3408
rect 29184 2100 29236 2106
rect 29184 2042 29236 2048
rect 29380 2038 29408 3402
rect 30576 2774 30604 3431
rect 29525 2748 29833 2757
rect 29525 2746 29531 2748
rect 29587 2746 29611 2748
rect 29667 2746 29691 2748
rect 29747 2746 29771 2748
rect 29827 2746 29833 2748
rect 29587 2694 29589 2746
rect 29769 2694 29771 2746
rect 29525 2692 29531 2694
rect 29587 2692 29611 2694
rect 29667 2692 29691 2694
rect 29747 2692 29771 2694
rect 29827 2692 29833 2694
rect 29525 2683 29833 2692
rect 30484 2746 30604 2774
rect 30852 2774 30880 6886
rect 31116 3120 31168 3126
rect 31116 3062 31168 3068
rect 30852 2746 31064 2774
rect 30012 2440 30064 2446
rect 30012 2382 30064 2388
rect 30104 2440 30156 2446
rect 30104 2382 30156 2388
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 30024 2106 30052 2382
rect 30012 2100 30064 2106
rect 30012 2042 30064 2048
rect 29368 2032 29420 2038
rect 29368 1974 29420 1980
rect 29276 1964 29328 1970
rect 29276 1906 29328 1912
rect 29644 1964 29696 1970
rect 29644 1906 29696 1912
rect 29092 1760 29144 1766
rect 29092 1702 29144 1708
rect 29000 1352 29052 1358
rect 29000 1294 29052 1300
rect 29000 876 29052 882
rect 29000 818 29052 824
rect 29012 785 29040 818
rect 28998 776 29054 785
rect 28998 711 29054 720
rect 29104 160 29132 1702
rect 29288 814 29316 1906
rect 29368 1828 29420 1834
rect 29368 1770 29420 1776
rect 29276 808 29328 814
rect 29276 750 29328 756
rect 29380 474 29408 1770
rect 29656 1748 29684 1906
rect 29656 1720 29960 1748
rect 29525 1660 29833 1669
rect 29525 1658 29531 1660
rect 29587 1658 29611 1660
rect 29667 1658 29691 1660
rect 29747 1658 29771 1660
rect 29827 1658 29833 1660
rect 29587 1606 29589 1658
rect 29769 1606 29771 1658
rect 29525 1604 29531 1606
rect 29587 1604 29611 1606
rect 29667 1604 29691 1606
rect 29747 1604 29771 1606
rect 29827 1604 29833 1606
rect 29525 1595 29833 1604
rect 29828 1556 29880 1562
rect 29828 1498 29880 1504
rect 29368 468 29420 474
rect 29368 410 29420 416
rect 29840 218 29868 1498
rect 29472 190 29592 218
rect 29472 160 29500 190
rect 28722 54 28948 82
rect 28354 0 28410 54
rect 28722 0 28778 54
rect 29090 0 29146 160
rect 29458 0 29514 160
rect 29564 82 29592 190
rect 29748 190 29868 218
rect 29932 202 29960 1720
rect 30116 746 30144 2382
rect 30392 2281 30420 2382
rect 30378 2272 30434 2281
rect 30378 2207 30434 2216
rect 30484 1970 30512 2746
rect 30932 2644 30984 2650
rect 30932 2586 30984 2592
rect 30840 2508 30892 2514
rect 30840 2450 30892 2456
rect 30748 2440 30800 2446
rect 30576 2400 30748 2428
rect 30472 1964 30524 1970
rect 30472 1906 30524 1912
rect 30380 1828 30432 1834
rect 30380 1770 30432 1776
rect 30288 1760 30340 1766
rect 30288 1702 30340 1708
rect 30300 1358 30328 1702
rect 30288 1352 30340 1358
rect 30288 1294 30340 1300
rect 30392 1290 30420 1770
rect 30470 1592 30526 1601
rect 30470 1527 30526 1536
rect 30484 1426 30512 1527
rect 30472 1420 30524 1426
rect 30472 1362 30524 1368
rect 30380 1284 30432 1290
rect 30380 1226 30432 1232
rect 30472 1284 30524 1290
rect 30472 1226 30524 1232
rect 30288 1216 30340 1222
rect 30288 1158 30340 1164
rect 30104 740 30156 746
rect 30104 682 30156 688
rect 29920 196 29972 202
rect 29748 82 29776 190
rect 29564 54 29776 82
rect 29826 82 29882 160
rect 29920 138 29972 144
rect 30104 196 30156 202
rect 30104 138 30156 144
rect 30116 82 30144 138
rect 29826 54 30144 82
rect 30194 82 30250 160
rect 30300 82 30328 1158
rect 30484 1018 30512 1226
rect 30472 1012 30524 1018
rect 30472 954 30524 960
rect 30576 406 30604 2400
rect 30748 2382 30800 2388
rect 30656 2304 30708 2310
rect 30656 2246 30708 2252
rect 30668 1426 30696 2246
rect 30748 1964 30800 1970
rect 30748 1906 30800 1912
rect 30656 1420 30708 1426
rect 30656 1362 30708 1368
rect 30760 406 30788 1906
rect 30852 1562 30880 2450
rect 30944 2106 30972 2586
rect 31036 2582 31064 2746
rect 31024 2576 31076 2582
rect 31024 2518 31076 2524
rect 31024 2372 31076 2378
rect 31024 2314 31076 2320
rect 30932 2100 30984 2106
rect 30932 2042 30984 2048
rect 30932 1760 30984 1766
rect 31036 1737 31064 2314
rect 30932 1702 30984 1708
rect 31022 1728 31078 1737
rect 30840 1556 30892 1562
rect 30840 1498 30892 1504
rect 30840 740 30892 746
rect 30840 682 30892 688
rect 30564 400 30616 406
rect 30564 342 30616 348
rect 30748 400 30800 406
rect 30748 342 30800 348
rect 30194 54 30328 82
rect 30562 82 30618 160
rect 30852 82 30880 682
rect 30944 160 30972 1702
rect 31022 1663 31078 1672
rect 31024 1352 31076 1358
rect 31024 1294 31076 1300
rect 31036 202 31064 1294
rect 31128 1018 31156 3062
rect 32128 2848 32180 2854
rect 32128 2790 32180 2796
rect 31208 2576 31260 2582
rect 31208 2518 31260 2524
rect 31220 2038 31248 2518
rect 31484 2440 31536 2446
rect 31484 2382 31536 2388
rect 31208 2032 31260 2038
rect 31208 1974 31260 1980
rect 31300 1556 31352 1562
rect 31300 1498 31352 1504
rect 31116 1012 31168 1018
rect 31116 954 31168 960
rect 31024 196 31076 202
rect 30562 54 30880 82
rect 29826 0 29882 54
rect 30194 0 30250 54
rect 30562 0 30618 54
rect 30930 0 30986 160
rect 31312 160 31340 1498
rect 31496 1193 31524 2382
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 31588 1970 31616 2246
rect 31576 1964 31628 1970
rect 31576 1906 31628 1912
rect 32140 1902 32168 2790
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 32494 2136 32550 2145
rect 32494 2071 32550 2080
rect 32312 1964 32364 1970
rect 32312 1906 32364 1912
rect 32128 1896 32180 1902
rect 32324 1850 32352 1906
rect 32508 1902 32536 2071
rect 32588 1964 32640 1970
rect 32588 1906 32640 1912
rect 32128 1838 32180 1844
rect 31668 1828 31720 1834
rect 31668 1770 31720 1776
rect 32232 1822 32352 1850
rect 32496 1896 32548 1902
rect 32496 1838 32548 1844
rect 31680 1578 31708 1770
rect 32128 1760 32180 1766
rect 32128 1702 32180 1708
rect 31588 1550 31708 1578
rect 31482 1184 31538 1193
rect 31482 1119 31538 1128
rect 31588 746 31616 1550
rect 31668 1488 31720 1494
rect 31668 1430 31720 1436
rect 31576 740 31628 746
rect 31576 682 31628 688
rect 31680 160 31708 1430
rect 32140 1358 32168 1702
rect 32128 1352 32180 1358
rect 32128 1294 32180 1300
rect 32232 678 32260 1822
rect 32496 1760 32548 1766
rect 32496 1702 32548 1708
rect 32508 1544 32536 1702
rect 32324 1516 32536 1544
rect 32220 672 32272 678
rect 32220 614 32272 620
rect 31024 138 31076 144
rect 31298 0 31354 160
rect 31666 0 31722 160
rect 32034 82 32090 160
rect 32324 82 32352 1516
rect 32496 1420 32548 1426
rect 32496 1362 32548 1368
rect 32508 241 32536 1362
rect 32600 610 32628 1906
rect 32772 1556 32824 1562
rect 32692 1516 32772 1544
rect 32588 604 32640 610
rect 32588 546 32640 552
rect 32494 232 32550 241
rect 32494 167 32550 176
rect 32034 54 32352 82
rect 32402 82 32458 160
rect 32692 82 32720 1516
rect 32772 1498 32824 1504
rect 32876 785 32904 2382
rect 33152 2310 33180 8434
rect 34794 3088 34850 3097
rect 33968 3052 34020 3058
rect 34850 3046 34928 3074
rect 34794 3023 34850 3032
rect 33968 2994 34020 3000
rect 33324 2440 33376 2446
rect 33324 2382 33376 2388
rect 32956 2304 33008 2310
rect 32956 2246 33008 2252
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 32968 1358 32996 2246
rect 33336 2106 33364 2382
rect 33324 2100 33376 2106
rect 33324 2042 33376 2048
rect 33336 1970 33456 1986
rect 33336 1964 33468 1970
rect 33336 1958 33416 1964
rect 33232 1760 33284 1766
rect 33232 1702 33284 1708
rect 33140 1488 33192 1494
rect 33060 1448 33140 1476
rect 32956 1352 33008 1358
rect 32956 1294 33008 1300
rect 32862 776 32918 785
rect 32862 711 32918 720
rect 32402 54 32720 82
rect 32770 82 32826 160
rect 33060 82 33088 1448
rect 33140 1430 33192 1436
rect 33244 1358 33272 1702
rect 33232 1352 33284 1358
rect 33232 1294 33284 1300
rect 33336 921 33364 1958
rect 33416 1906 33468 1912
rect 33784 1896 33836 1902
rect 33612 1844 33784 1850
rect 33612 1838 33836 1844
rect 33416 1828 33468 1834
rect 33416 1770 33468 1776
rect 33612 1822 33824 1838
rect 33322 912 33378 921
rect 33322 847 33378 856
rect 32770 54 33088 82
rect 33138 82 33194 160
rect 33428 82 33456 1770
rect 33612 1426 33640 1822
rect 33784 1760 33836 1766
rect 33784 1702 33836 1708
rect 33690 1592 33746 1601
rect 33690 1527 33746 1536
rect 33704 1426 33732 1527
rect 33600 1420 33652 1426
rect 33600 1362 33652 1368
rect 33692 1420 33744 1426
rect 33692 1362 33744 1368
rect 33138 54 33456 82
rect 33506 82 33562 160
rect 33796 82 33824 1702
rect 33980 746 34008 2994
rect 34612 1760 34664 1766
rect 34612 1702 34664 1708
rect 34152 1556 34204 1562
rect 34152 1498 34204 1504
rect 33968 740 34020 746
rect 33968 682 34020 688
rect 33506 54 33824 82
rect 33874 82 33930 160
rect 34164 82 34192 1498
rect 34336 1488 34388 1494
rect 34256 1448 34336 1476
rect 34256 160 34284 1448
rect 34336 1430 34388 1436
rect 34624 160 34652 1702
rect 34900 1358 34928 3046
rect 35084 2650 35112 8434
rect 35240 7644 35548 7653
rect 35240 7642 35246 7644
rect 35302 7642 35326 7644
rect 35382 7642 35406 7644
rect 35462 7642 35486 7644
rect 35542 7642 35548 7644
rect 35302 7590 35304 7642
rect 35484 7590 35486 7642
rect 35240 7588 35246 7590
rect 35302 7588 35326 7590
rect 35382 7588 35406 7590
rect 35462 7588 35486 7590
rect 35542 7588 35548 7590
rect 35240 7579 35548 7588
rect 35240 6556 35548 6565
rect 35240 6554 35246 6556
rect 35302 6554 35326 6556
rect 35382 6554 35406 6556
rect 35462 6554 35486 6556
rect 35542 6554 35548 6556
rect 35302 6502 35304 6554
rect 35484 6502 35486 6554
rect 35240 6500 35246 6502
rect 35302 6500 35326 6502
rect 35382 6500 35406 6502
rect 35462 6500 35486 6502
rect 35542 6500 35548 6502
rect 35240 6491 35548 6500
rect 35240 5468 35548 5477
rect 35240 5466 35246 5468
rect 35302 5466 35326 5468
rect 35382 5466 35406 5468
rect 35462 5466 35486 5468
rect 35542 5466 35548 5468
rect 35302 5414 35304 5466
rect 35484 5414 35486 5466
rect 35240 5412 35246 5414
rect 35302 5412 35326 5414
rect 35382 5412 35406 5414
rect 35462 5412 35486 5414
rect 35542 5412 35548 5414
rect 35240 5403 35548 5412
rect 35240 4380 35548 4389
rect 35240 4378 35246 4380
rect 35302 4378 35326 4380
rect 35382 4378 35406 4380
rect 35462 4378 35486 4380
rect 35542 4378 35548 4380
rect 35302 4326 35304 4378
rect 35484 4326 35486 4378
rect 35240 4324 35246 4326
rect 35302 4324 35326 4326
rect 35382 4324 35406 4326
rect 35462 4324 35486 4326
rect 35542 4324 35548 4326
rect 35240 4315 35548 4324
rect 36266 4040 36322 4049
rect 36266 3975 36322 3984
rect 35240 3292 35548 3301
rect 35240 3290 35246 3292
rect 35302 3290 35326 3292
rect 35382 3290 35406 3292
rect 35462 3290 35486 3292
rect 35542 3290 35548 3292
rect 35302 3238 35304 3290
rect 35484 3238 35486 3290
rect 35240 3236 35246 3238
rect 35302 3236 35326 3238
rect 35382 3236 35406 3238
rect 35462 3236 35486 3238
rect 35542 3236 35548 3238
rect 35240 3227 35548 3236
rect 35072 2644 35124 2650
rect 35072 2586 35124 2592
rect 36084 2508 36136 2514
rect 36084 2450 36136 2456
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 35240 2204 35548 2213
rect 35240 2202 35246 2204
rect 35302 2202 35326 2204
rect 35382 2202 35406 2204
rect 35462 2202 35486 2204
rect 35542 2202 35548 2204
rect 35302 2150 35304 2202
rect 35484 2150 35486 2202
rect 35240 2148 35246 2150
rect 35302 2148 35326 2150
rect 35382 2148 35406 2150
rect 35462 2148 35486 2150
rect 35542 2148 35548 2150
rect 35240 2139 35548 2148
rect 35912 2106 35940 2382
rect 35900 2100 35952 2106
rect 35900 2042 35952 2048
rect 35532 2032 35584 2038
rect 35716 2032 35768 2038
rect 35584 1992 35716 2020
rect 35532 1974 35584 1980
rect 35716 1974 35768 1980
rect 36096 1873 36124 2450
rect 36280 1970 36308 3975
rect 37384 2650 37412 8434
rect 40955 8188 41263 8197
rect 40955 8186 40961 8188
rect 41017 8186 41041 8188
rect 41097 8186 41121 8188
rect 41177 8186 41201 8188
rect 41257 8186 41263 8188
rect 41017 8134 41019 8186
rect 41199 8134 41201 8186
rect 40955 8132 40961 8134
rect 41017 8132 41041 8134
rect 41097 8132 41121 8134
rect 41177 8132 41201 8134
rect 41257 8132 41263 8134
rect 40955 8123 41263 8132
rect 40955 7100 41263 7109
rect 40955 7098 40961 7100
rect 41017 7098 41041 7100
rect 41097 7098 41121 7100
rect 41177 7098 41201 7100
rect 41257 7098 41263 7100
rect 41017 7046 41019 7098
rect 41199 7046 41201 7098
rect 40955 7044 40961 7046
rect 41017 7044 41041 7046
rect 41097 7044 41121 7046
rect 41177 7044 41201 7046
rect 41257 7044 41263 7046
rect 40955 7035 41263 7044
rect 40955 6012 41263 6021
rect 40955 6010 40961 6012
rect 41017 6010 41041 6012
rect 41097 6010 41121 6012
rect 41177 6010 41201 6012
rect 41257 6010 41263 6012
rect 41017 5958 41019 6010
rect 41199 5958 41201 6010
rect 40955 5956 40961 5958
rect 41017 5956 41041 5958
rect 41097 5956 41121 5958
rect 41177 5956 41201 5958
rect 41257 5956 41263 5958
rect 40955 5947 41263 5956
rect 40955 4924 41263 4933
rect 40955 4922 40961 4924
rect 41017 4922 41041 4924
rect 41097 4922 41121 4924
rect 41177 4922 41201 4924
rect 41257 4922 41263 4924
rect 41017 4870 41019 4922
rect 41199 4870 41201 4922
rect 40955 4868 40961 4870
rect 41017 4868 41041 4870
rect 41097 4868 41121 4870
rect 41177 4868 41201 4870
rect 41257 4868 41263 4870
rect 40955 4859 41263 4868
rect 38108 4480 38160 4486
rect 38108 4422 38160 4428
rect 37832 2916 37884 2922
rect 37832 2858 37884 2864
rect 37844 2774 37872 2858
rect 37752 2746 37872 2774
rect 37372 2644 37424 2650
rect 37372 2586 37424 2592
rect 36268 1964 36320 1970
rect 36268 1906 36320 1912
rect 37372 1964 37424 1970
rect 37372 1906 37424 1912
rect 36082 1864 36138 1873
rect 35992 1828 36044 1834
rect 36082 1799 36138 1808
rect 37280 1828 37332 1834
rect 35992 1770 36044 1776
rect 37280 1770 37332 1776
rect 34980 1556 35032 1562
rect 34980 1498 35032 1504
rect 34888 1352 34940 1358
rect 34888 1294 34940 1300
rect 34796 1284 34848 1290
rect 34796 1226 34848 1232
rect 34808 950 34836 1226
rect 34796 944 34848 950
rect 34796 886 34848 892
rect 34992 160 35020 1498
rect 35900 1488 35952 1494
rect 35636 1448 35900 1476
rect 35072 1284 35124 1290
rect 35072 1226 35124 1232
rect 35084 950 35112 1226
rect 35240 1116 35548 1125
rect 35240 1114 35246 1116
rect 35302 1114 35326 1116
rect 35382 1114 35406 1116
rect 35462 1114 35486 1116
rect 35542 1114 35548 1116
rect 35302 1062 35304 1114
rect 35484 1062 35486 1114
rect 35240 1060 35246 1062
rect 35302 1060 35326 1062
rect 35382 1060 35406 1062
rect 35462 1060 35486 1062
rect 35542 1060 35548 1062
rect 35240 1051 35548 1060
rect 35072 944 35124 950
rect 35072 886 35124 892
rect 33874 54 34192 82
rect 32034 0 32090 54
rect 32402 0 32458 54
rect 32770 0 32826 54
rect 33138 0 33194 54
rect 33506 0 33562 54
rect 33874 0 33930 54
rect 34242 0 34298 160
rect 34610 0 34666 160
rect 34978 0 35034 160
rect 35346 82 35402 160
rect 35636 82 35664 1448
rect 35900 1430 35952 1436
rect 36004 1340 36032 1770
rect 36084 1760 36136 1766
rect 36084 1702 36136 1708
rect 35820 1312 36032 1340
rect 35346 54 35664 82
rect 35714 82 35770 160
rect 35820 82 35848 1312
rect 36096 160 36124 1702
rect 36820 1556 36872 1562
rect 36740 1516 36820 1544
rect 35714 54 35848 82
rect 35346 0 35402 54
rect 35714 0 35770 54
rect 36082 0 36138 160
rect 36450 82 36506 160
rect 36740 82 36768 1516
rect 36820 1498 36872 1504
rect 37096 1488 37148 1494
rect 37292 1442 37320 1770
rect 37384 1465 37412 1906
rect 37096 1430 37148 1436
rect 36450 54 36768 82
rect 36818 82 36874 160
rect 37108 82 37136 1430
rect 37200 1414 37320 1442
rect 37370 1456 37426 1465
rect 37200 160 37228 1414
rect 37370 1391 37426 1400
rect 37752 1358 37780 2746
rect 38016 2304 38068 2310
rect 37844 2264 38016 2292
rect 37740 1352 37792 1358
rect 37740 1294 37792 1300
rect 37464 1216 37516 1222
rect 37464 1158 37516 1164
rect 37476 746 37504 1158
rect 37464 740 37516 746
rect 37464 682 37516 688
rect 36818 54 37136 82
rect 36450 0 36506 54
rect 36818 0 36874 54
rect 37186 0 37242 160
rect 37554 82 37610 160
rect 37844 82 37872 2264
rect 38016 2246 38068 2252
rect 38120 1358 38148 4422
rect 41602 4176 41658 4185
rect 41602 4111 41658 4120
rect 40955 3836 41263 3845
rect 40955 3834 40961 3836
rect 41017 3834 41041 3836
rect 41097 3834 41121 3836
rect 41177 3834 41201 3836
rect 41257 3834 41263 3836
rect 41017 3782 41019 3834
rect 41199 3782 41201 3834
rect 40955 3780 40961 3782
rect 41017 3780 41041 3782
rect 41097 3780 41121 3782
rect 41177 3780 41201 3782
rect 41257 3780 41263 3782
rect 40955 3771 41263 3780
rect 38934 3632 38990 3641
rect 38990 3590 39068 3618
rect 38934 3567 38990 3576
rect 38568 2848 38620 2854
rect 38568 2790 38620 2796
rect 38198 2000 38254 2009
rect 38198 1935 38200 1944
rect 38252 1935 38254 1944
rect 38200 1906 38252 1912
rect 38580 1902 38608 2790
rect 38658 2544 38714 2553
rect 38714 2502 38792 2530
rect 38658 2479 38714 2488
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 38672 2106 38700 2246
rect 38660 2100 38712 2106
rect 38660 2042 38712 2048
rect 38764 1970 38792 2502
rect 38752 1964 38804 1970
rect 38752 1906 38804 1912
rect 38568 1896 38620 1902
rect 38212 1834 38424 1850
rect 38568 1838 38620 1844
rect 38200 1828 38424 1834
rect 38252 1822 38424 1828
rect 38200 1770 38252 1776
rect 38396 1766 38424 1822
rect 38476 1828 38528 1834
rect 38476 1770 38528 1776
rect 38384 1760 38436 1766
rect 38488 1737 38516 1770
rect 38936 1760 38988 1766
rect 38384 1702 38436 1708
rect 38474 1728 38530 1737
rect 38936 1702 38988 1708
rect 38474 1663 38530 1672
rect 38292 1556 38344 1562
rect 38212 1516 38292 1544
rect 38108 1352 38160 1358
rect 38108 1294 38160 1300
rect 37554 54 37872 82
rect 37922 82 37978 160
rect 38212 82 38240 1516
rect 38292 1498 38344 1504
rect 38844 1488 38896 1494
rect 38580 1448 38844 1476
rect 37922 54 38240 82
rect 38290 82 38346 160
rect 38580 82 38608 1448
rect 38844 1430 38896 1436
rect 38290 54 38608 82
rect 38658 82 38714 160
rect 38948 82 38976 1702
rect 39040 1358 39068 3590
rect 40955 2748 41263 2757
rect 40955 2746 40961 2748
rect 41017 2746 41041 2748
rect 41097 2746 41121 2748
rect 41177 2746 41201 2748
rect 41257 2746 41263 2748
rect 41017 2694 41019 2746
rect 41199 2694 41201 2746
rect 40955 2692 40961 2694
rect 41017 2692 41041 2694
rect 41097 2692 41121 2694
rect 41177 2692 41201 2694
rect 41257 2692 41263 2694
rect 40955 2683 41263 2692
rect 41512 2576 41564 2582
rect 41512 2518 41564 2524
rect 39118 2408 39174 2417
rect 39118 2343 39174 2352
rect 39132 1766 39160 2343
rect 40512 1970 40632 1986
rect 40132 1964 40184 1970
rect 40132 1906 40184 1912
rect 40512 1964 40644 1970
rect 40512 1958 40592 1964
rect 39120 1760 39172 1766
rect 39120 1702 39172 1708
rect 39304 1556 39356 1562
rect 39304 1498 39356 1504
rect 39028 1352 39080 1358
rect 39028 1294 39080 1300
rect 38658 54 38976 82
rect 39026 82 39082 160
rect 39316 82 39344 1498
rect 39488 1352 39540 1358
rect 39488 1294 39540 1300
rect 40040 1352 40092 1358
rect 40040 1294 40092 1300
rect 39026 54 39344 82
rect 39394 82 39450 160
rect 39500 82 39528 1294
rect 39672 1216 39724 1222
rect 39672 1158 39724 1164
rect 39684 950 39712 1158
rect 39672 944 39724 950
rect 39672 886 39724 892
rect 39394 54 39528 82
rect 39762 82 39818 160
rect 40052 82 40080 1294
rect 40144 160 40172 1906
rect 40224 1284 40276 1290
rect 40224 1226 40276 1232
rect 40236 202 40264 1226
rect 40224 196 40276 202
rect 39762 54 40080 82
rect 37554 0 37610 54
rect 37922 0 37978 54
rect 38290 0 38346 54
rect 38658 0 38714 54
rect 39026 0 39082 54
rect 39394 0 39450 54
rect 39762 0 39818 54
rect 40130 0 40186 160
rect 40512 160 40540 1958
rect 40592 1906 40644 1912
rect 41052 1964 41104 1970
rect 41052 1906 41104 1912
rect 41328 1964 41380 1970
rect 41328 1906 41380 1912
rect 41064 1850 41092 1906
rect 40776 1828 40828 1834
rect 40776 1770 40828 1776
rect 40880 1822 41092 1850
rect 40788 1562 40816 1770
rect 40776 1556 40828 1562
rect 40776 1498 40828 1504
rect 40880 160 40908 1822
rect 40955 1660 41263 1669
rect 40955 1658 40961 1660
rect 41017 1658 41041 1660
rect 41097 1658 41121 1660
rect 41177 1658 41201 1660
rect 41257 1658 41263 1660
rect 41017 1606 41019 1658
rect 41199 1606 41201 1658
rect 40955 1604 40961 1606
rect 41017 1604 41041 1606
rect 41097 1604 41121 1606
rect 41177 1604 41201 1606
rect 41257 1604 41263 1606
rect 40955 1595 41263 1604
rect 41144 1216 41196 1222
rect 41144 1158 41196 1164
rect 41236 1216 41288 1222
rect 41236 1158 41288 1164
rect 41156 474 41184 1158
rect 41248 1018 41276 1158
rect 41236 1012 41288 1018
rect 41236 954 41288 960
rect 41144 468 41196 474
rect 41144 410 41196 416
rect 40224 138 40276 144
rect 40498 0 40554 160
rect 40866 0 40922 160
rect 41234 82 41290 160
rect 41340 82 41368 1906
rect 41524 1562 41552 2518
rect 41512 1556 41564 1562
rect 41512 1498 41564 1504
rect 41616 1340 41644 4111
rect 41708 2650 41736 8434
rect 44732 8424 44784 8430
rect 44732 8366 44784 8372
rect 44744 2650 44772 8366
rect 45020 2650 45048 8434
rect 46124 2650 46152 8434
rect 46670 7644 46978 7653
rect 46670 7642 46676 7644
rect 46732 7642 46756 7644
rect 46812 7642 46836 7644
rect 46892 7642 46916 7644
rect 46972 7642 46978 7644
rect 46732 7590 46734 7642
rect 46914 7590 46916 7642
rect 46670 7588 46676 7590
rect 46732 7588 46756 7590
rect 46812 7588 46836 7590
rect 46892 7588 46916 7590
rect 46972 7588 46978 7590
rect 46670 7579 46978 7588
rect 46670 6556 46978 6565
rect 46670 6554 46676 6556
rect 46732 6554 46756 6556
rect 46812 6554 46836 6556
rect 46892 6554 46916 6556
rect 46972 6554 46978 6556
rect 46732 6502 46734 6554
rect 46914 6502 46916 6554
rect 46670 6500 46676 6502
rect 46732 6500 46756 6502
rect 46812 6500 46836 6502
rect 46892 6500 46916 6502
rect 46972 6500 46978 6502
rect 46670 6491 46978 6500
rect 46670 5468 46978 5477
rect 46670 5466 46676 5468
rect 46732 5466 46756 5468
rect 46812 5466 46836 5468
rect 46892 5466 46916 5468
rect 46972 5466 46978 5468
rect 46732 5414 46734 5466
rect 46914 5414 46916 5466
rect 46670 5412 46676 5414
rect 46732 5412 46756 5414
rect 46812 5412 46836 5414
rect 46892 5412 46916 5414
rect 46972 5412 46978 5414
rect 46670 5403 46978 5412
rect 46670 4380 46978 4389
rect 46670 4378 46676 4380
rect 46732 4378 46756 4380
rect 46812 4378 46836 4380
rect 46892 4378 46916 4380
rect 46972 4378 46978 4380
rect 46732 4326 46734 4378
rect 46914 4326 46916 4378
rect 46670 4324 46676 4326
rect 46732 4324 46756 4326
rect 46812 4324 46836 4326
rect 46892 4324 46916 4326
rect 46972 4324 46978 4326
rect 46670 4315 46978 4324
rect 46670 3292 46978 3301
rect 46670 3290 46676 3292
rect 46732 3290 46756 3292
rect 46812 3290 46836 3292
rect 46892 3290 46916 3292
rect 46972 3290 46978 3292
rect 46732 3238 46734 3290
rect 46914 3238 46916 3290
rect 46670 3236 46676 3238
rect 46732 3236 46756 3238
rect 46812 3236 46836 3238
rect 46892 3236 46916 3238
rect 46972 3236 46978 3238
rect 46670 3227 46978 3236
rect 41696 2644 41748 2650
rect 41696 2586 41748 2592
rect 44732 2644 44784 2650
rect 44732 2586 44784 2592
rect 45008 2644 45060 2650
rect 45008 2586 45060 2592
rect 46112 2644 46164 2650
rect 46112 2586 46164 2592
rect 44456 2576 44508 2582
rect 44456 2518 44508 2524
rect 42248 2440 42300 2446
rect 42248 2382 42300 2388
rect 42260 2106 42288 2382
rect 42800 2372 42852 2378
rect 42800 2314 42852 2320
rect 42248 2100 42300 2106
rect 42248 2042 42300 2048
rect 42812 1562 42840 2314
rect 43996 1964 44048 1970
rect 43996 1906 44048 1912
rect 42800 1556 42852 1562
rect 42800 1498 42852 1504
rect 41696 1352 41748 1358
rect 41616 1312 41696 1340
rect 41696 1294 41748 1300
rect 41880 1352 41932 1358
rect 43260 1352 43312 1358
rect 41880 1294 41932 1300
rect 43166 1320 43222 1329
rect 41234 54 41368 82
rect 41602 82 41658 160
rect 41892 82 41920 1294
rect 41972 1284 42024 1290
rect 41972 1226 42024 1232
rect 42340 1284 42392 1290
rect 43260 1294 43312 1300
rect 43536 1352 43588 1358
rect 43536 1294 43588 1300
rect 43904 1352 43956 1358
rect 43904 1294 43956 1300
rect 43166 1255 43222 1264
rect 42340 1226 42392 1232
rect 41984 160 42012 1226
rect 42352 160 42380 1226
rect 43180 1222 43208 1255
rect 42708 1216 42760 1222
rect 42708 1158 42760 1164
rect 42892 1216 42944 1222
rect 42892 1158 42944 1164
rect 43168 1216 43220 1222
rect 43168 1158 43220 1164
rect 42720 160 42748 1158
rect 42904 610 42932 1158
rect 42892 604 42944 610
rect 42892 546 42944 552
rect 41602 54 41920 82
rect 41234 0 41290 54
rect 41602 0 41658 54
rect 41970 0 42026 160
rect 42338 0 42394 160
rect 42706 0 42762 160
rect 43074 82 43130 160
rect 43272 82 43300 1294
rect 43444 1216 43496 1222
rect 43444 1158 43496 1164
rect 43456 610 43484 1158
rect 43444 604 43496 610
rect 43444 546 43496 552
rect 43074 54 43300 82
rect 43442 82 43498 160
rect 43548 82 43576 1294
rect 43720 1216 43772 1222
rect 43720 1158 43772 1164
rect 43732 610 43760 1158
rect 43720 604 43772 610
rect 43720 546 43772 552
rect 43442 54 43576 82
rect 43810 82 43866 160
rect 43916 82 43944 1294
rect 44008 1290 44036 1906
rect 44468 1494 44496 2518
rect 44548 2440 44600 2446
rect 44548 2382 44600 2388
rect 45192 2440 45244 2446
rect 45192 2382 45244 2388
rect 45836 2440 45888 2446
rect 45836 2382 45888 2388
rect 44560 2106 44588 2382
rect 45204 2106 45232 2382
rect 45848 2106 45876 2382
rect 46670 2204 46978 2213
rect 46670 2202 46676 2204
rect 46732 2202 46756 2204
rect 46812 2202 46836 2204
rect 46892 2202 46916 2204
rect 46972 2202 46978 2204
rect 46732 2150 46734 2202
rect 46914 2150 46916 2202
rect 46670 2148 46676 2150
rect 46732 2148 46756 2150
rect 46812 2148 46836 2150
rect 46892 2148 46916 2150
rect 46972 2148 46978 2150
rect 46670 2139 46978 2148
rect 44548 2100 44600 2106
rect 44548 2042 44600 2048
rect 45192 2100 45244 2106
rect 45192 2042 45244 2048
rect 45836 2100 45888 2106
rect 45836 2042 45888 2048
rect 45008 2032 45060 2038
rect 45008 1974 45060 1980
rect 45020 1562 45048 1974
rect 46480 1964 46532 1970
rect 46480 1906 46532 1912
rect 45744 1896 45796 1902
rect 45744 1838 45796 1844
rect 45756 1562 45784 1838
rect 45008 1556 45060 1562
rect 45008 1498 45060 1504
rect 45744 1556 45796 1562
rect 45744 1498 45796 1504
rect 44088 1488 44140 1494
rect 44088 1430 44140 1436
rect 44456 1488 44508 1494
rect 44456 1430 44508 1436
rect 43996 1284 44048 1290
rect 43996 1226 44048 1232
rect 44100 1018 44128 1430
rect 44272 1352 44324 1358
rect 44640 1352 44692 1358
rect 44272 1294 44324 1300
rect 44560 1312 44640 1340
rect 44088 1012 44140 1018
rect 44088 954 44140 960
rect 43810 54 43944 82
rect 44178 82 44234 160
rect 44284 82 44312 1294
rect 44560 160 44588 1312
rect 44640 1294 44692 1300
rect 45192 1352 45244 1358
rect 45192 1294 45244 1300
rect 45560 1352 45612 1358
rect 45560 1294 45612 1300
rect 45928 1352 45980 1358
rect 45928 1294 45980 1300
rect 46296 1352 46348 1358
rect 46296 1294 46348 1300
rect 44178 54 44312 82
rect 43074 0 43130 54
rect 43442 0 43498 54
rect 43810 0 43866 54
rect 44178 0 44234 54
rect 44546 0 44602 160
rect 44914 82 44970 160
rect 45204 82 45232 1294
rect 45296 190 45416 218
rect 45296 160 45324 190
rect 44914 54 45232 82
rect 44914 0 44970 54
rect 45282 0 45338 160
rect 45388 82 45416 190
rect 45572 82 45600 1294
rect 45388 54 45600 82
rect 45650 82 45706 160
rect 45940 82 45968 1294
rect 45650 54 45968 82
rect 46018 82 46074 160
rect 46308 82 46336 1294
rect 46018 54 46336 82
rect 46386 82 46442 160
rect 46492 82 46520 1906
rect 46572 1896 46624 1902
rect 46572 1838 46624 1844
rect 46386 54 46520 82
rect 46584 82 46612 1838
rect 46670 1116 46978 1125
rect 46670 1114 46676 1116
rect 46732 1114 46756 1116
rect 46812 1114 46836 1116
rect 46892 1114 46916 1116
rect 46972 1114 46978 1116
rect 46732 1062 46734 1114
rect 46914 1062 46916 1114
rect 46670 1060 46676 1062
rect 46732 1060 46756 1062
rect 46812 1060 46836 1062
rect 46892 1060 46916 1062
rect 46972 1060 46978 1062
rect 46670 1051 46978 1060
rect 46754 82 46810 160
rect 46584 54 46810 82
rect 45650 0 45706 54
rect 46018 0 46074 54
rect 46386 0 46442 54
rect 46754 0 46810 54
<< via2 >>
rect 12386 8730 12442 8732
rect 12466 8730 12522 8732
rect 12546 8730 12602 8732
rect 12626 8730 12682 8732
rect 12386 8678 12432 8730
rect 12432 8678 12442 8730
rect 12466 8678 12496 8730
rect 12496 8678 12508 8730
rect 12508 8678 12522 8730
rect 12546 8678 12560 8730
rect 12560 8678 12572 8730
rect 12572 8678 12602 8730
rect 12626 8678 12636 8730
rect 12636 8678 12682 8730
rect 12386 8676 12442 8678
rect 12466 8676 12522 8678
rect 12546 8676 12602 8678
rect 12626 8676 12682 8678
rect 6671 8186 6727 8188
rect 6751 8186 6807 8188
rect 6831 8186 6887 8188
rect 6911 8186 6967 8188
rect 6671 8134 6717 8186
rect 6717 8134 6727 8186
rect 6751 8134 6781 8186
rect 6781 8134 6793 8186
rect 6793 8134 6807 8186
rect 6831 8134 6845 8186
rect 6845 8134 6857 8186
rect 6857 8134 6887 8186
rect 6911 8134 6921 8186
rect 6921 8134 6967 8186
rect 6671 8132 6727 8134
rect 6751 8132 6807 8134
rect 6831 8132 6887 8134
rect 6911 8132 6967 8134
rect 12386 7642 12442 7644
rect 12466 7642 12522 7644
rect 12546 7642 12602 7644
rect 12626 7642 12682 7644
rect 12386 7590 12432 7642
rect 12432 7590 12442 7642
rect 12466 7590 12496 7642
rect 12496 7590 12508 7642
rect 12508 7590 12522 7642
rect 12546 7590 12560 7642
rect 12560 7590 12572 7642
rect 12572 7590 12602 7642
rect 12626 7590 12636 7642
rect 12636 7590 12682 7642
rect 12386 7588 12442 7590
rect 12466 7588 12522 7590
rect 12546 7588 12602 7590
rect 12626 7588 12682 7590
rect 6671 7098 6727 7100
rect 6751 7098 6807 7100
rect 6831 7098 6887 7100
rect 6911 7098 6967 7100
rect 6671 7046 6717 7098
rect 6717 7046 6727 7098
rect 6751 7046 6781 7098
rect 6781 7046 6793 7098
rect 6793 7046 6807 7098
rect 6831 7046 6845 7098
rect 6845 7046 6857 7098
rect 6857 7046 6887 7098
rect 6911 7046 6921 7098
rect 6921 7046 6967 7098
rect 6671 7044 6727 7046
rect 6751 7044 6807 7046
rect 6831 7044 6887 7046
rect 6911 7044 6967 7046
rect 12386 6554 12442 6556
rect 12466 6554 12522 6556
rect 12546 6554 12602 6556
rect 12626 6554 12682 6556
rect 12386 6502 12432 6554
rect 12432 6502 12442 6554
rect 12466 6502 12496 6554
rect 12496 6502 12508 6554
rect 12508 6502 12522 6554
rect 12546 6502 12560 6554
rect 12560 6502 12572 6554
rect 12572 6502 12602 6554
rect 12626 6502 12636 6554
rect 12636 6502 12682 6554
rect 12386 6500 12442 6502
rect 12466 6500 12522 6502
rect 12546 6500 12602 6502
rect 12626 6500 12682 6502
rect 6671 6010 6727 6012
rect 6751 6010 6807 6012
rect 6831 6010 6887 6012
rect 6911 6010 6967 6012
rect 6671 5958 6717 6010
rect 6717 5958 6727 6010
rect 6751 5958 6781 6010
rect 6781 5958 6793 6010
rect 6793 5958 6807 6010
rect 6831 5958 6845 6010
rect 6845 5958 6857 6010
rect 6857 5958 6887 6010
rect 6911 5958 6921 6010
rect 6921 5958 6967 6010
rect 6671 5956 6727 5958
rect 6751 5956 6807 5958
rect 6831 5956 6887 5958
rect 6911 5956 6967 5958
rect 12386 5466 12442 5468
rect 12466 5466 12522 5468
rect 12546 5466 12602 5468
rect 12626 5466 12682 5468
rect 12386 5414 12432 5466
rect 12432 5414 12442 5466
rect 12466 5414 12496 5466
rect 12496 5414 12508 5466
rect 12508 5414 12522 5466
rect 12546 5414 12560 5466
rect 12560 5414 12572 5466
rect 12572 5414 12602 5466
rect 12626 5414 12636 5466
rect 12636 5414 12682 5466
rect 12386 5412 12442 5414
rect 12466 5412 12522 5414
rect 12546 5412 12602 5414
rect 12626 5412 12682 5414
rect 6671 4922 6727 4924
rect 6751 4922 6807 4924
rect 6831 4922 6887 4924
rect 6911 4922 6967 4924
rect 6671 4870 6717 4922
rect 6717 4870 6727 4922
rect 6751 4870 6781 4922
rect 6781 4870 6793 4922
rect 6793 4870 6807 4922
rect 6831 4870 6845 4922
rect 6845 4870 6857 4922
rect 6857 4870 6887 4922
rect 6911 4870 6921 4922
rect 6921 4870 6967 4922
rect 6671 4868 6727 4870
rect 6751 4868 6807 4870
rect 6831 4868 6887 4870
rect 6911 4868 6967 4870
rect 6671 3834 6727 3836
rect 6751 3834 6807 3836
rect 6831 3834 6887 3836
rect 6911 3834 6967 3836
rect 6671 3782 6717 3834
rect 6717 3782 6727 3834
rect 6751 3782 6781 3834
rect 6781 3782 6793 3834
rect 6793 3782 6807 3834
rect 6831 3782 6845 3834
rect 6845 3782 6857 3834
rect 6857 3782 6887 3834
rect 6911 3782 6921 3834
rect 6921 3782 6967 3834
rect 6671 3780 6727 3782
rect 6751 3780 6807 3782
rect 6831 3780 6887 3782
rect 6911 3780 6967 3782
rect 6671 2746 6727 2748
rect 6751 2746 6807 2748
rect 6831 2746 6887 2748
rect 6911 2746 6967 2748
rect 6671 2694 6717 2746
rect 6717 2694 6727 2746
rect 6751 2694 6781 2746
rect 6781 2694 6793 2746
rect 6793 2694 6807 2746
rect 6831 2694 6845 2746
rect 6845 2694 6857 2746
rect 6857 2694 6887 2746
rect 6911 2694 6921 2746
rect 6921 2694 6967 2746
rect 6671 2692 6727 2694
rect 6751 2692 6807 2694
rect 6831 2692 6887 2694
rect 6911 2692 6967 2694
rect 6671 1658 6727 1660
rect 6751 1658 6807 1660
rect 6831 1658 6887 1660
rect 6911 1658 6967 1660
rect 6671 1606 6717 1658
rect 6717 1606 6727 1658
rect 6751 1606 6781 1658
rect 6781 1606 6793 1658
rect 6793 1606 6807 1658
rect 6831 1606 6845 1658
rect 6845 1606 6857 1658
rect 6857 1606 6887 1658
rect 6911 1606 6921 1658
rect 6921 1606 6967 1658
rect 6671 1604 6727 1606
rect 6751 1604 6807 1606
rect 6831 1604 6887 1606
rect 6911 1604 6967 1606
rect 12386 4378 12442 4380
rect 12466 4378 12522 4380
rect 12546 4378 12602 4380
rect 12626 4378 12682 4380
rect 12386 4326 12432 4378
rect 12432 4326 12442 4378
rect 12466 4326 12496 4378
rect 12496 4326 12508 4378
rect 12508 4326 12522 4378
rect 12546 4326 12560 4378
rect 12560 4326 12572 4378
rect 12572 4326 12602 4378
rect 12626 4326 12636 4378
rect 12636 4326 12682 4378
rect 12386 4324 12442 4326
rect 12466 4324 12522 4326
rect 12546 4324 12602 4326
rect 12626 4324 12682 4326
rect 15934 3576 15990 3632
rect 12070 3440 12126 3496
rect 8666 2352 8722 2408
rect 9862 3032 9918 3088
rect 9126 312 9182 368
rect 9494 448 9550 504
rect 10598 176 10654 232
rect 10966 856 11022 912
rect 11242 1264 11298 1320
rect 12386 3290 12442 3292
rect 12466 3290 12522 3292
rect 12546 3290 12602 3292
rect 12626 3290 12682 3292
rect 12386 3238 12432 3290
rect 12432 3238 12442 3290
rect 12466 3238 12496 3290
rect 12496 3238 12508 3290
rect 12508 3238 12522 3290
rect 12546 3238 12560 3290
rect 12560 3238 12572 3290
rect 12572 3238 12602 3290
rect 12626 3238 12636 3290
rect 12636 3238 12682 3290
rect 12386 3236 12442 3238
rect 12466 3236 12522 3238
rect 12546 3236 12602 3238
rect 12626 3236 12682 3238
rect 12386 2202 12442 2204
rect 12466 2202 12522 2204
rect 12546 2202 12602 2204
rect 12626 2202 12682 2204
rect 12386 2150 12432 2202
rect 12432 2150 12442 2202
rect 12466 2150 12496 2202
rect 12496 2150 12508 2202
rect 12508 2150 12522 2202
rect 12546 2150 12560 2202
rect 12560 2150 12572 2202
rect 12572 2150 12602 2202
rect 12626 2150 12636 2202
rect 12636 2150 12682 2202
rect 12386 2148 12442 2150
rect 12466 2148 12522 2150
rect 12546 2148 12602 2150
rect 12626 2148 12682 2150
rect 12386 1114 12442 1116
rect 12466 1114 12522 1116
rect 12546 1114 12602 1116
rect 12626 1114 12682 1116
rect 12386 1062 12432 1114
rect 12432 1062 12442 1114
rect 12466 1062 12496 1114
rect 12496 1062 12508 1114
rect 12508 1062 12522 1114
rect 12546 1062 12560 1114
rect 12560 1062 12572 1114
rect 12572 1062 12602 1114
rect 12626 1062 12636 1114
rect 12636 1062 12682 1114
rect 12386 1060 12442 1062
rect 12466 1060 12522 1062
rect 12546 1060 12602 1062
rect 12626 1060 12682 1062
rect 12622 584 12678 640
rect 13174 992 13230 1048
rect 14002 2896 14058 2952
rect 14738 1400 14794 1456
rect 16486 2100 16542 2136
rect 17314 3984 17370 4040
rect 16486 2080 16488 2100
rect 16488 2080 16540 2100
rect 16540 2080 16542 2100
rect 16578 1944 16634 2000
rect 16210 1808 16266 1864
rect 15106 1128 15162 1184
rect 18101 8186 18157 8188
rect 18181 8186 18237 8188
rect 18261 8186 18317 8188
rect 18341 8186 18397 8188
rect 18101 8134 18147 8186
rect 18147 8134 18157 8186
rect 18181 8134 18211 8186
rect 18211 8134 18223 8186
rect 18223 8134 18237 8186
rect 18261 8134 18275 8186
rect 18275 8134 18287 8186
rect 18287 8134 18317 8186
rect 18341 8134 18351 8186
rect 18351 8134 18397 8186
rect 18101 8132 18157 8134
rect 18181 8132 18237 8134
rect 18261 8132 18317 8134
rect 18341 8132 18397 8134
rect 18101 7098 18157 7100
rect 18181 7098 18237 7100
rect 18261 7098 18317 7100
rect 18341 7098 18397 7100
rect 18101 7046 18147 7098
rect 18147 7046 18157 7098
rect 18181 7046 18211 7098
rect 18211 7046 18223 7098
rect 18223 7046 18237 7098
rect 18261 7046 18275 7098
rect 18275 7046 18287 7098
rect 18287 7046 18317 7098
rect 18341 7046 18351 7098
rect 18351 7046 18397 7098
rect 18101 7044 18157 7046
rect 18181 7044 18237 7046
rect 18261 7044 18317 7046
rect 18341 7044 18397 7046
rect 18101 6010 18157 6012
rect 18181 6010 18237 6012
rect 18261 6010 18317 6012
rect 18341 6010 18397 6012
rect 18101 5958 18147 6010
rect 18147 5958 18157 6010
rect 18181 5958 18211 6010
rect 18211 5958 18223 6010
rect 18223 5958 18237 6010
rect 18261 5958 18275 6010
rect 18275 5958 18287 6010
rect 18287 5958 18317 6010
rect 18341 5958 18351 6010
rect 18351 5958 18397 6010
rect 18101 5956 18157 5958
rect 18181 5956 18237 5958
rect 18261 5956 18317 5958
rect 18341 5956 18397 5958
rect 18101 4922 18157 4924
rect 18181 4922 18237 4924
rect 18261 4922 18317 4924
rect 18341 4922 18397 4924
rect 18101 4870 18147 4922
rect 18147 4870 18157 4922
rect 18181 4870 18211 4922
rect 18211 4870 18223 4922
rect 18223 4870 18237 4922
rect 18261 4870 18275 4922
rect 18275 4870 18287 4922
rect 18287 4870 18317 4922
rect 18341 4870 18351 4922
rect 18351 4870 18397 4922
rect 18101 4868 18157 4870
rect 18181 4868 18237 4870
rect 18261 4868 18317 4870
rect 18341 4868 18397 4870
rect 17774 4120 17830 4176
rect 18101 3834 18157 3836
rect 18181 3834 18237 3836
rect 18261 3834 18317 3836
rect 18341 3834 18397 3836
rect 18101 3782 18147 3834
rect 18147 3782 18157 3834
rect 18181 3782 18211 3834
rect 18211 3782 18223 3834
rect 18223 3782 18237 3834
rect 18261 3782 18275 3834
rect 18275 3782 18287 3834
rect 18287 3782 18317 3834
rect 18341 3782 18351 3834
rect 18351 3782 18397 3834
rect 18101 3780 18157 3782
rect 18181 3780 18237 3782
rect 18261 3780 18317 3782
rect 18341 3780 18397 3782
rect 18878 2760 18934 2816
rect 18101 2746 18157 2748
rect 18181 2746 18237 2748
rect 18261 2746 18317 2748
rect 18341 2746 18397 2748
rect 18101 2694 18147 2746
rect 18147 2694 18157 2746
rect 18181 2694 18211 2746
rect 18211 2694 18223 2746
rect 18223 2694 18237 2746
rect 18261 2694 18275 2746
rect 18275 2694 18287 2746
rect 18287 2694 18317 2746
rect 18341 2694 18351 2746
rect 18351 2694 18397 2746
rect 18101 2692 18157 2694
rect 18181 2692 18237 2694
rect 18261 2692 18317 2694
rect 18341 2692 18397 2694
rect 19338 2216 19394 2272
rect 17498 992 17554 1048
rect 18101 1658 18157 1660
rect 18181 1658 18237 1660
rect 18261 1658 18317 1660
rect 18341 1658 18397 1660
rect 18101 1606 18147 1658
rect 18147 1606 18157 1658
rect 18181 1606 18211 1658
rect 18211 1606 18223 1658
rect 18223 1606 18237 1658
rect 18261 1606 18275 1658
rect 18275 1606 18287 1658
rect 18287 1606 18317 1658
rect 18341 1606 18351 1658
rect 18351 1606 18397 1658
rect 18101 1604 18157 1606
rect 18181 1604 18237 1606
rect 18261 1604 18317 1606
rect 18341 1604 18397 1606
rect 18510 1536 18566 1592
rect 21362 3712 21418 3768
rect 21362 2896 21418 2952
rect 20534 2488 20590 2544
rect 18970 1672 19026 1728
rect 18878 1264 18934 1320
rect 19706 1944 19762 2000
rect 19890 1944 19946 2000
rect 20258 1964 20314 2000
rect 20258 1944 20260 1964
rect 20260 1944 20312 1964
rect 20312 1944 20314 1964
rect 19706 1264 19762 1320
rect 19614 720 19670 776
rect 22834 2896 22890 2952
rect 23816 8730 23872 8732
rect 23896 8730 23952 8732
rect 23976 8730 24032 8732
rect 24056 8730 24112 8732
rect 23816 8678 23862 8730
rect 23862 8678 23872 8730
rect 23896 8678 23926 8730
rect 23926 8678 23938 8730
rect 23938 8678 23952 8730
rect 23976 8678 23990 8730
rect 23990 8678 24002 8730
rect 24002 8678 24032 8730
rect 24056 8678 24066 8730
rect 24066 8678 24112 8730
rect 23816 8676 23872 8678
rect 23896 8676 23952 8678
rect 23976 8676 24032 8678
rect 24056 8676 24112 8678
rect 23816 7642 23872 7644
rect 23896 7642 23952 7644
rect 23976 7642 24032 7644
rect 24056 7642 24112 7644
rect 23816 7590 23862 7642
rect 23862 7590 23872 7642
rect 23896 7590 23926 7642
rect 23926 7590 23938 7642
rect 23938 7590 23952 7642
rect 23976 7590 23990 7642
rect 23990 7590 24002 7642
rect 24002 7590 24032 7642
rect 24056 7590 24066 7642
rect 24066 7590 24112 7642
rect 23816 7588 23872 7590
rect 23896 7588 23952 7590
rect 23976 7588 24032 7590
rect 24056 7588 24112 7590
rect 23816 6554 23872 6556
rect 23896 6554 23952 6556
rect 23976 6554 24032 6556
rect 24056 6554 24112 6556
rect 23816 6502 23862 6554
rect 23862 6502 23872 6554
rect 23896 6502 23926 6554
rect 23926 6502 23938 6554
rect 23938 6502 23952 6554
rect 23976 6502 23990 6554
rect 23990 6502 24002 6554
rect 24002 6502 24032 6554
rect 24056 6502 24066 6554
rect 24066 6502 24112 6554
rect 23816 6500 23872 6502
rect 23896 6500 23952 6502
rect 23976 6500 24032 6502
rect 24056 6500 24112 6502
rect 23816 5466 23872 5468
rect 23896 5466 23952 5468
rect 23976 5466 24032 5468
rect 24056 5466 24112 5468
rect 23816 5414 23862 5466
rect 23862 5414 23872 5466
rect 23896 5414 23926 5466
rect 23926 5414 23938 5466
rect 23938 5414 23952 5466
rect 23976 5414 23990 5466
rect 23990 5414 24002 5466
rect 24002 5414 24032 5466
rect 24056 5414 24066 5466
rect 24066 5414 24112 5466
rect 23816 5412 23872 5414
rect 23896 5412 23952 5414
rect 23976 5412 24032 5414
rect 24056 5412 24112 5414
rect 23816 4378 23872 4380
rect 23896 4378 23952 4380
rect 23976 4378 24032 4380
rect 24056 4378 24112 4380
rect 23816 4326 23862 4378
rect 23862 4326 23872 4378
rect 23896 4326 23926 4378
rect 23926 4326 23938 4378
rect 23938 4326 23952 4378
rect 23976 4326 23990 4378
rect 23990 4326 24002 4378
rect 24002 4326 24032 4378
rect 24056 4326 24066 4378
rect 24066 4326 24112 4378
rect 23816 4324 23872 4326
rect 23896 4324 23952 4326
rect 23976 4324 24032 4326
rect 24056 4324 24112 4326
rect 23816 3290 23872 3292
rect 23896 3290 23952 3292
rect 23976 3290 24032 3292
rect 24056 3290 24112 3292
rect 23816 3238 23862 3290
rect 23862 3238 23872 3290
rect 23896 3238 23926 3290
rect 23926 3238 23938 3290
rect 23938 3238 23952 3290
rect 23976 3238 23990 3290
rect 23990 3238 24002 3290
rect 24002 3238 24032 3290
rect 24056 3238 24066 3290
rect 24066 3238 24112 3290
rect 23816 3236 23872 3238
rect 23896 3236 23952 3238
rect 23976 3236 24032 3238
rect 24056 3236 24112 3238
rect 21638 2216 21694 2272
rect 21362 1400 21418 1456
rect 21454 584 21510 640
rect 19062 40 19118 96
rect 22098 1672 22154 1728
rect 22006 1128 22062 1184
rect 23662 2352 23718 2408
rect 23816 2202 23872 2204
rect 23896 2202 23952 2204
rect 23976 2202 24032 2204
rect 24056 2202 24112 2204
rect 23816 2150 23862 2202
rect 23862 2150 23872 2202
rect 23896 2150 23926 2202
rect 23926 2150 23938 2202
rect 23938 2150 23952 2202
rect 23976 2150 23990 2202
rect 23990 2150 24002 2202
rect 24002 2150 24032 2202
rect 24056 2150 24066 2202
rect 24066 2150 24112 2202
rect 23816 2148 23872 2150
rect 23896 2148 23952 2150
rect 23976 2148 24032 2150
rect 24056 2148 24112 2150
rect 24398 2080 24454 2136
rect 25962 3032 26018 3088
rect 26146 3032 26202 3088
rect 26146 2760 26202 2816
rect 26606 2352 26662 2408
rect 24306 1264 24362 1320
rect 23816 1114 23872 1116
rect 23896 1114 23952 1116
rect 23976 1114 24032 1116
rect 24056 1114 24112 1116
rect 23816 1062 23862 1114
rect 23862 1062 23872 1114
rect 23896 1062 23926 1114
rect 23926 1062 23938 1114
rect 23938 1062 23952 1114
rect 23976 1062 23990 1114
rect 23990 1062 24002 1114
rect 24002 1062 24032 1114
rect 24056 1062 24066 1114
rect 24066 1062 24112 1114
rect 23816 1060 23872 1062
rect 23896 1060 23952 1062
rect 23976 1060 24032 1062
rect 24056 1060 24112 1062
rect 28262 3712 28318 3768
rect 35246 8730 35302 8732
rect 35326 8730 35382 8732
rect 35406 8730 35462 8732
rect 35486 8730 35542 8732
rect 35246 8678 35292 8730
rect 35292 8678 35302 8730
rect 35326 8678 35356 8730
rect 35356 8678 35368 8730
rect 35368 8678 35382 8730
rect 35406 8678 35420 8730
rect 35420 8678 35432 8730
rect 35432 8678 35462 8730
rect 35486 8678 35496 8730
rect 35496 8678 35542 8730
rect 35246 8676 35302 8678
rect 35326 8676 35382 8678
rect 35406 8676 35462 8678
rect 35486 8676 35542 8678
rect 46676 8730 46732 8732
rect 46756 8730 46812 8732
rect 46836 8730 46892 8732
rect 46916 8730 46972 8732
rect 46676 8678 46722 8730
rect 46722 8678 46732 8730
rect 46756 8678 46786 8730
rect 46786 8678 46798 8730
rect 46798 8678 46812 8730
rect 46836 8678 46850 8730
rect 46850 8678 46862 8730
rect 46862 8678 46892 8730
rect 46916 8678 46926 8730
rect 46926 8678 46972 8730
rect 46676 8676 46732 8678
rect 46756 8676 46812 8678
rect 46836 8676 46892 8678
rect 46916 8676 46972 8678
rect 29531 8186 29587 8188
rect 29611 8186 29667 8188
rect 29691 8186 29747 8188
rect 29771 8186 29827 8188
rect 29531 8134 29577 8186
rect 29577 8134 29587 8186
rect 29611 8134 29641 8186
rect 29641 8134 29653 8186
rect 29653 8134 29667 8186
rect 29691 8134 29705 8186
rect 29705 8134 29717 8186
rect 29717 8134 29747 8186
rect 29771 8134 29781 8186
rect 29781 8134 29827 8186
rect 29531 8132 29587 8134
rect 29611 8132 29667 8134
rect 29691 8132 29747 8134
rect 29771 8132 29827 8134
rect 29531 7098 29587 7100
rect 29611 7098 29667 7100
rect 29691 7098 29747 7100
rect 29771 7098 29827 7100
rect 29531 7046 29577 7098
rect 29577 7046 29587 7098
rect 29611 7046 29641 7098
rect 29641 7046 29653 7098
rect 29653 7046 29667 7098
rect 29691 7046 29705 7098
rect 29705 7046 29717 7098
rect 29717 7046 29747 7098
rect 29771 7046 29781 7098
rect 29781 7046 29827 7098
rect 29531 7044 29587 7046
rect 29611 7044 29667 7046
rect 29691 7044 29747 7046
rect 29771 7044 29827 7046
rect 29531 6010 29587 6012
rect 29611 6010 29667 6012
rect 29691 6010 29747 6012
rect 29771 6010 29827 6012
rect 29531 5958 29577 6010
rect 29577 5958 29587 6010
rect 29611 5958 29641 6010
rect 29641 5958 29653 6010
rect 29653 5958 29667 6010
rect 29691 5958 29705 6010
rect 29705 5958 29717 6010
rect 29717 5958 29747 6010
rect 29771 5958 29781 6010
rect 29781 5958 29827 6010
rect 29531 5956 29587 5958
rect 29611 5956 29667 5958
rect 29691 5956 29747 5958
rect 29771 5956 29827 5958
rect 29531 4922 29587 4924
rect 29611 4922 29667 4924
rect 29691 4922 29747 4924
rect 29771 4922 29827 4924
rect 29531 4870 29577 4922
rect 29577 4870 29587 4922
rect 29611 4870 29641 4922
rect 29641 4870 29653 4922
rect 29653 4870 29667 4922
rect 29691 4870 29705 4922
rect 29705 4870 29717 4922
rect 29717 4870 29747 4922
rect 29771 4870 29781 4922
rect 29781 4870 29827 4922
rect 29531 4868 29587 4870
rect 29611 4868 29667 4870
rect 29691 4868 29747 4870
rect 29771 4868 29827 4870
rect 29531 3834 29587 3836
rect 29611 3834 29667 3836
rect 29691 3834 29747 3836
rect 29771 3834 29827 3836
rect 29531 3782 29577 3834
rect 29577 3782 29587 3834
rect 29611 3782 29641 3834
rect 29641 3782 29653 3834
rect 29653 3782 29667 3834
rect 29691 3782 29705 3834
rect 29705 3782 29717 3834
rect 29717 3782 29747 3834
rect 29771 3782 29781 3834
rect 29781 3782 29827 3834
rect 29531 3780 29587 3782
rect 29611 3780 29667 3782
rect 29691 3780 29747 3782
rect 29771 3780 29827 3782
rect 30562 3440 30618 3496
rect 29531 2746 29587 2748
rect 29611 2746 29667 2748
rect 29691 2746 29747 2748
rect 29771 2746 29827 2748
rect 29531 2694 29577 2746
rect 29577 2694 29587 2746
rect 29611 2694 29641 2746
rect 29641 2694 29653 2746
rect 29653 2694 29667 2746
rect 29691 2694 29705 2746
rect 29705 2694 29717 2746
rect 29717 2694 29747 2746
rect 29771 2694 29781 2746
rect 29781 2694 29827 2746
rect 29531 2692 29587 2694
rect 29611 2692 29667 2694
rect 29691 2692 29747 2694
rect 29771 2692 29827 2694
rect 28998 720 29054 776
rect 29531 1658 29587 1660
rect 29611 1658 29667 1660
rect 29691 1658 29747 1660
rect 29771 1658 29827 1660
rect 29531 1606 29577 1658
rect 29577 1606 29587 1658
rect 29611 1606 29641 1658
rect 29641 1606 29653 1658
rect 29653 1606 29667 1658
rect 29691 1606 29705 1658
rect 29705 1606 29717 1658
rect 29717 1606 29747 1658
rect 29771 1606 29781 1658
rect 29781 1606 29827 1658
rect 29531 1604 29587 1606
rect 29611 1604 29667 1606
rect 29691 1604 29747 1606
rect 29771 1604 29827 1606
rect 30378 2216 30434 2272
rect 30470 1536 30526 1592
rect 31022 1672 31078 1728
rect 32494 2080 32550 2136
rect 31482 1128 31538 1184
rect 32494 176 32550 232
rect 34794 3032 34850 3088
rect 32862 720 32918 776
rect 33322 856 33378 912
rect 33690 1536 33746 1592
rect 35246 7642 35302 7644
rect 35326 7642 35382 7644
rect 35406 7642 35462 7644
rect 35486 7642 35542 7644
rect 35246 7590 35292 7642
rect 35292 7590 35302 7642
rect 35326 7590 35356 7642
rect 35356 7590 35368 7642
rect 35368 7590 35382 7642
rect 35406 7590 35420 7642
rect 35420 7590 35432 7642
rect 35432 7590 35462 7642
rect 35486 7590 35496 7642
rect 35496 7590 35542 7642
rect 35246 7588 35302 7590
rect 35326 7588 35382 7590
rect 35406 7588 35462 7590
rect 35486 7588 35542 7590
rect 35246 6554 35302 6556
rect 35326 6554 35382 6556
rect 35406 6554 35462 6556
rect 35486 6554 35542 6556
rect 35246 6502 35292 6554
rect 35292 6502 35302 6554
rect 35326 6502 35356 6554
rect 35356 6502 35368 6554
rect 35368 6502 35382 6554
rect 35406 6502 35420 6554
rect 35420 6502 35432 6554
rect 35432 6502 35462 6554
rect 35486 6502 35496 6554
rect 35496 6502 35542 6554
rect 35246 6500 35302 6502
rect 35326 6500 35382 6502
rect 35406 6500 35462 6502
rect 35486 6500 35542 6502
rect 35246 5466 35302 5468
rect 35326 5466 35382 5468
rect 35406 5466 35462 5468
rect 35486 5466 35542 5468
rect 35246 5414 35292 5466
rect 35292 5414 35302 5466
rect 35326 5414 35356 5466
rect 35356 5414 35368 5466
rect 35368 5414 35382 5466
rect 35406 5414 35420 5466
rect 35420 5414 35432 5466
rect 35432 5414 35462 5466
rect 35486 5414 35496 5466
rect 35496 5414 35542 5466
rect 35246 5412 35302 5414
rect 35326 5412 35382 5414
rect 35406 5412 35462 5414
rect 35486 5412 35542 5414
rect 35246 4378 35302 4380
rect 35326 4378 35382 4380
rect 35406 4378 35462 4380
rect 35486 4378 35542 4380
rect 35246 4326 35292 4378
rect 35292 4326 35302 4378
rect 35326 4326 35356 4378
rect 35356 4326 35368 4378
rect 35368 4326 35382 4378
rect 35406 4326 35420 4378
rect 35420 4326 35432 4378
rect 35432 4326 35462 4378
rect 35486 4326 35496 4378
rect 35496 4326 35542 4378
rect 35246 4324 35302 4326
rect 35326 4324 35382 4326
rect 35406 4324 35462 4326
rect 35486 4324 35542 4326
rect 36266 3984 36322 4040
rect 35246 3290 35302 3292
rect 35326 3290 35382 3292
rect 35406 3290 35462 3292
rect 35486 3290 35542 3292
rect 35246 3238 35292 3290
rect 35292 3238 35302 3290
rect 35326 3238 35356 3290
rect 35356 3238 35368 3290
rect 35368 3238 35382 3290
rect 35406 3238 35420 3290
rect 35420 3238 35432 3290
rect 35432 3238 35462 3290
rect 35486 3238 35496 3290
rect 35496 3238 35542 3290
rect 35246 3236 35302 3238
rect 35326 3236 35382 3238
rect 35406 3236 35462 3238
rect 35486 3236 35542 3238
rect 35246 2202 35302 2204
rect 35326 2202 35382 2204
rect 35406 2202 35462 2204
rect 35486 2202 35542 2204
rect 35246 2150 35292 2202
rect 35292 2150 35302 2202
rect 35326 2150 35356 2202
rect 35356 2150 35368 2202
rect 35368 2150 35382 2202
rect 35406 2150 35420 2202
rect 35420 2150 35432 2202
rect 35432 2150 35462 2202
rect 35486 2150 35496 2202
rect 35496 2150 35542 2202
rect 35246 2148 35302 2150
rect 35326 2148 35382 2150
rect 35406 2148 35462 2150
rect 35486 2148 35542 2150
rect 40961 8186 41017 8188
rect 41041 8186 41097 8188
rect 41121 8186 41177 8188
rect 41201 8186 41257 8188
rect 40961 8134 41007 8186
rect 41007 8134 41017 8186
rect 41041 8134 41071 8186
rect 41071 8134 41083 8186
rect 41083 8134 41097 8186
rect 41121 8134 41135 8186
rect 41135 8134 41147 8186
rect 41147 8134 41177 8186
rect 41201 8134 41211 8186
rect 41211 8134 41257 8186
rect 40961 8132 41017 8134
rect 41041 8132 41097 8134
rect 41121 8132 41177 8134
rect 41201 8132 41257 8134
rect 40961 7098 41017 7100
rect 41041 7098 41097 7100
rect 41121 7098 41177 7100
rect 41201 7098 41257 7100
rect 40961 7046 41007 7098
rect 41007 7046 41017 7098
rect 41041 7046 41071 7098
rect 41071 7046 41083 7098
rect 41083 7046 41097 7098
rect 41121 7046 41135 7098
rect 41135 7046 41147 7098
rect 41147 7046 41177 7098
rect 41201 7046 41211 7098
rect 41211 7046 41257 7098
rect 40961 7044 41017 7046
rect 41041 7044 41097 7046
rect 41121 7044 41177 7046
rect 41201 7044 41257 7046
rect 40961 6010 41017 6012
rect 41041 6010 41097 6012
rect 41121 6010 41177 6012
rect 41201 6010 41257 6012
rect 40961 5958 41007 6010
rect 41007 5958 41017 6010
rect 41041 5958 41071 6010
rect 41071 5958 41083 6010
rect 41083 5958 41097 6010
rect 41121 5958 41135 6010
rect 41135 5958 41147 6010
rect 41147 5958 41177 6010
rect 41201 5958 41211 6010
rect 41211 5958 41257 6010
rect 40961 5956 41017 5958
rect 41041 5956 41097 5958
rect 41121 5956 41177 5958
rect 41201 5956 41257 5958
rect 40961 4922 41017 4924
rect 41041 4922 41097 4924
rect 41121 4922 41177 4924
rect 41201 4922 41257 4924
rect 40961 4870 41007 4922
rect 41007 4870 41017 4922
rect 41041 4870 41071 4922
rect 41071 4870 41083 4922
rect 41083 4870 41097 4922
rect 41121 4870 41135 4922
rect 41135 4870 41147 4922
rect 41147 4870 41177 4922
rect 41201 4870 41211 4922
rect 41211 4870 41257 4922
rect 40961 4868 41017 4870
rect 41041 4868 41097 4870
rect 41121 4868 41177 4870
rect 41201 4868 41257 4870
rect 36082 1808 36138 1864
rect 35246 1114 35302 1116
rect 35326 1114 35382 1116
rect 35406 1114 35462 1116
rect 35486 1114 35542 1116
rect 35246 1062 35292 1114
rect 35292 1062 35302 1114
rect 35326 1062 35356 1114
rect 35356 1062 35368 1114
rect 35368 1062 35382 1114
rect 35406 1062 35420 1114
rect 35420 1062 35432 1114
rect 35432 1062 35462 1114
rect 35486 1062 35496 1114
rect 35496 1062 35542 1114
rect 35246 1060 35302 1062
rect 35326 1060 35382 1062
rect 35406 1060 35462 1062
rect 35486 1060 35542 1062
rect 37370 1400 37426 1456
rect 41602 4120 41658 4176
rect 40961 3834 41017 3836
rect 41041 3834 41097 3836
rect 41121 3834 41177 3836
rect 41201 3834 41257 3836
rect 40961 3782 41007 3834
rect 41007 3782 41017 3834
rect 41041 3782 41071 3834
rect 41071 3782 41083 3834
rect 41083 3782 41097 3834
rect 41121 3782 41135 3834
rect 41135 3782 41147 3834
rect 41147 3782 41177 3834
rect 41201 3782 41211 3834
rect 41211 3782 41257 3834
rect 40961 3780 41017 3782
rect 41041 3780 41097 3782
rect 41121 3780 41177 3782
rect 41201 3780 41257 3782
rect 38934 3576 38990 3632
rect 38198 1964 38254 2000
rect 38198 1944 38200 1964
rect 38200 1944 38252 1964
rect 38252 1944 38254 1964
rect 38658 2488 38714 2544
rect 38474 1672 38530 1728
rect 40961 2746 41017 2748
rect 41041 2746 41097 2748
rect 41121 2746 41177 2748
rect 41201 2746 41257 2748
rect 40961 2694 41007 2746
rect 41007 2694 41017 2746
rect 41041 2694 41071 2746
rect 41071 2694 41083 2746
rect 41083 2694 41097 2746
rect 41121 2694 41135 2746
rect 41135 2694 41147 2746
rect 41147 2694 41177 2746
rect 41201 2694 41211 2746
rect 41211 2694 41257 2746
rect 40961 2692 41017 2694
rect 41041 2692 41097 2694
rect 41121 2692 41177 2694
rect 41201 2692 41257 2694
rect 39118 2352 39174 2408
rect 40961 1658 41017 1660
rect 41041 1658 41097 1660
rect 41121 1658 41177 1660
rect 41201 1658 41257 1660
rect 40961 1606 41007 1658
rect 41007 1606 41017 1658
rect 41041 1606 41071 1658
rect 41071 1606 41083 1658
rect 41083 1606 41097 1658
rect 41121 1606 41135 1658
rect 41135 1606 41147 1658
rect 41147 1606 41177 1658
rect 41201 1606 41211 1658
rect 41211 1606 41257 1658
rect 40961 1604 41017 1606
rect 41041 1604 41097 1606
rect 41121 1604 41177 1606
rect 41201 1604 41257 1606
rect 46676 7642 46732 7644
rect 46756 7642 46812 7644
rect 46836 7642 46892 7644
rect 46916 7642 46972 7644
rect 46676 7590 46722 7642
rect 46722 7590 46732 7642
rect 46756 7590 46786 7642
rect 46786 7590 46798 7642
rect 46798 7590 46812 7642
rect 46836 7590 46850 7642
rect 46850 7590 46862 7642
rect 46862 7590 46892 7642
rect 46916 7590 46926 7642
rect 46926 7590 46972 7642
rect 46676 7588 46732 7590
rect 46756 7588 46812 7590
rect 46836 7588 46892 7590
rect 46916 7588 46972 7590
rect 46676 6554 46732 6556
rect 46756 6554 46812 6556
rect 46836 6554 46892 6556
rect 46916 6554 46972 6556
rect 46676 6502 46722 6554
rect 46722 6502 46732 6554
rect 46756 6502 46786 6554
rect 46786 6502 46798 6554
rect 46798 6502 46812 6554
rect 46836 6502 46850 6554
rect 46850 6502 46862 6554
rect 46862 6502 46892 6554
rect 46916 6502 46926 6554
rect 46926 6502 46972 6554
rect 46676 6500 46732 6502
rect 46756 6500 46812 6502
rect 46836 6500 46892 6502
rect 46916 6500 46972 6502
rect 46676 5466 46732 5468
rect 46756 5466 46812 5468
rect 46836 5466 46892 5468
rect 46916 5466 46972 5468
rect 46676 5414 46722 5466
rect 46722 5414 46732 5466
rect 46756 5414 46786 5466
rect 46786 5414 46798 5466
rect 46798 5414 46812 5466
rect 46836 5414 46850 5466
rect 46850 5414 46862 5466
rect 46862 5414 46892 5466
rect 46916 5414 46926 5466
rect 46926 5414 46972 5466
rect 46676 5412 46732 5414
rect 46756 5412 46812 5414
rect 46836 5412 46892 5414
rect 46916 5412 46972 5414
rect 46676 4378 46732 4380
rect 46756 4378 46812 4380
rect 46836 4378 46892 4380
rect 46916 4378 46972 4380
rect 46676 4326 46722 4378
rect 46722 4326 46732 4378
rect 46756 4326 46786 4378
rect 46786 4326 46798 4378
rect 46798 4326 46812 4378
rect 46836 4326 46850 4378
rect 46850 4326 46862 4378
rect 46862 4326 46892 4378
rect 46916 4326 46926 4378
rect 46926 4326 46972 4378
rect 46676 4324 46732 4326
rect 46756 4324 46812 4326
rect 46836 4324 46892 4326
rect 46916 4324 46972 4326
rect 46676 3290 46732 3292
rect 46756 3290 46812 3292
rect 46836 3290 46892 3292
rect 46916 3290 46972 3292
rect 46676 3238 46722 3290
rect 46722 3238 46732 3290
rect 46756 3238 46786 3290
rect 46786 3238 46798 3290
rect 46798 3238 46812 3290
rect 46836 3238 46850 3290
rect 46850 3238 46862 3290
rect 46862 3238 46892 3290
rect 46916 3238 46926 3290
rect 46926 3238 46972 3290
rect 46676 3236 46732 3238
rect 46756 3236 46812 3238
rect 46836 3236 46892 3238
rect 46916 3236 46972 3238
rect 43166 1264 43222 1320
rect 46676 2202 46732 2204
rect 46756 2202 46812 2204
rect 46836 2202 46892 2204
rect 46916 2202 46972 2204
rect 46676 2150 46722 2202
rect 46722 2150 46732 2202
rect 46756 2150 46786 2202
rect 46786 2150 46798 2202
rect 46798 2150 46812 2202
rect 46836 2150 46850 2202
rect 46850 2150 46862 2202
rect 46862 2150 46892 2202
rect 46916 2150 46926 2202
rect 46926 2150 46972 2202
rect 46676 2148 46732 2150
rect 46756 2148 46812 2150
rect 46836 2148 46892 2150
rect 46916 2148 46972 2150
rect 46676 1114 46732 1116
rect 46756 1114 46812 1116
rect 46836 1114 46892 1116
rect 46916 1114 46972 1116
rect 46676 1062 46722 1114
rect 46722 1062 46732 1114
rect 46756 1062 46786 1114
rect 46786 1062 46798 1114
rect 46798 1062 46812 1114
rect 46836 1062 46850 1114
rect 46850 1062 46862 1114
rect 46862 1062 46892 1114
rect 46916 1062 46926 1114
rect 46926 1062 46972 1114
rect 46676 1060 46732 1062
rect 46756 1060 46812 1062
rect 46836 1060 46892 1062
rect 46916 1060 46972 1062
<< metal3 >>
rect 12376 8736 12692 8737
rect 12376 8672 12382 8736
rect 12446 8672 12462 8736
rect 12526 8672 12542 8736
rect 12606 8672 12622 8736
rect 12686 8672 12692 8736
rect 12376 8671 12692 8672
rect 23806 8736 24122 8737
rect 23806 8672 23812 8736
rect 23876 8672 23892 8736
rect 23956 8672 23972 8736
rect 24036 8672 24052 8736
rect 24116 8672 24122 8736
rect 23806 8671 24122 8672
rect 35236 8736 35552 8737
rect 35236 8672 35242 8736
rect 35306 8672 35322 8736
rect 35386 8672 35402 8736
rect 35466 8672 35482 8736
rect 35546 8672 35552 8736
rect 35236 8671 35552 8672
rect 46666 8736 46982 8737
rect 46666 8672 46672 8736
rect 46736 8672 46752 8736
rect 46816 8672 46832 8736
rect 46896 8672 46912 8736
rect 46976 8672 46982 8736
rect 46666 8671 46982 8672
rect 6661 8192 6977 8193
rect 6661 8128 6667 8192
rect 6731 8128 6747 8192
rect 6811 8128 6827 8192
rect 6891 8128 6907 8192
rect 6971 8128 6977 8192
rect 6661 8127 6977 8128
rect 18091 8192 18407 8193
rect 18091 8128 18097 8192
rect 18161 8128 18177 8192
rect 18241 8128 18257 8192
rect 18321 8128 18337 8192
rect 18401 8128 18407 8192
rect 18091 8127 18407 8128
rect 29521 8192 29837 8193
rect 29521 8128 29527 8192
rect 29591 8128 29607 8192
rect 29671 8128 29687 8192
rect 29751 8128 29767 8192
rect 29831 8128 29837 8192
rect 29521 8127 29837 8128
rect 40951 8192 41267 8193
rect 40951 8128 40957 8192
rect 41021 8128 41037 8192
rect 41101 8128 41117 8192
rect 41181 8128 41197 8192
rect 41261 8128 41267 8192
rect 40951 8127 41267 8128
rect 12376 7648 12692 7649
rect 12376 7584 12382 7648
rect 12446 7584 12462 7648
rect 12526 7584 12542 7648
rect 12606 7584 12622 7648
rect 12686 7584 12692 7648
rect 12376 7583 12692 7584
rect 23806 7648 24122 7649
rect 23806 7584 23812 7648
rect 23876 7584 23892 7648
rect 23956 7584 23972 7648
rect 24036 7584 24052 7648
rect 24116 7584 24122 7648
rect 23806 7583 24122 7584
rect 35236 7648 35552 7649
rect 35236 7584 35242 7648
rect 35306 7584 35322 7648
rect 35386 7584 35402 7648
rect 35466 7584 35482 7648
rect 35546 7584 35552 7648
rect 35236 7583 35552 7584
rect 46666 7648 46982 7649
rect 46666 7584 46672 7648
rect 46736 7584 46752 7648
rect 46816 7584 46832 7648
rect 46896 7584 46912 7648
rect 46976 7584 46982 7648
rect 46666 7583 46982 7584
rect 6661 7104 6977 7105
rect 6661 7040 6667 7104
rect 6731 7040 6747 7104
rect 6811 7040 6827 7104
rect 6891 7040 6907 7104
rect 6971 7040 6977 7104
rect 6661 7039 6977 7040
rect 18091 7104 18407 7105
rect 18091 7040 18097 7104
rect 18161 7040 18177 7104
rect 18241 7040 18257 7104
rect 18321 7040 18337 7104
rect 18401 7040 18407 7104
rect 18091 7039 18407 7040
rect 29521 7104 29837 7105
rect 29521 7040 29527 7104
rect 29591 7040 29607 7104
rect 29671 7040 29687 7104
rect 29751 7040 29767 7104
rect 29831 7040 29837 7104
rect 29521 7039 29837 7040
rect 40951 7104 41267 7105
rect 40951 7040 40957 7104
rect 41021 7040 41037 7104
rect 41101 7040 41117 7104
rect 41181 7040 41197 7104
rect 41261 7040 41267 7104
rect 40951 7039 41267 7040
rect 12376 6560 12692 6561
rect 12376 6496 12382 6560
rect 12446 6496 12462 6560
rect 12526 6496 12542 6560
rect 12606 6496 12622 6560
rect 12686 6496 12692 6560
rect 12376 6495 12692 6496
rect 23806 6560 24122 6561
rect 23806 6496 23812 6560
rect 23876 6496 23892 6560
rect 23956 6496 23972 6560
rect 24036 6496 24052 6560
rect 24116 6496 24122 6560
rect 23806 6495 24122 6496
rect 35236 6560 35552 6561
rect 35236 6496 35242 6560
rect 35306 6496 35322 6560
rect 35386 6496 35402 6560
rect 35466 6496 35482 6560
rect 35546 6496 35552 6560
rect 35236 6495 35552 6496
rect 46666 6560 46982 6561
rect 46666 6496 46672 6560
rect 46736 6496 46752 6560
rect 46816 6496 46832 6560
rect 46896 6496 46912 6560
rect 46976 6496 46982 6560
rect 46666 6495 46982 6496
rect 6661 6016 6977 6017
rect 6661 5952 6667 6016
rect 6731 5952 6747 6016
rect 6811 5952 6827 6016
rect 6891 5952 6907 6016
rect 6971 5952 6977 6016
rect 6661 5951 6977 5952
rect 18091 6016 18407 6017
rect 18091 5952 18097 6016
rect 18161 5952 18177 6016
rect 18241 5952 18257 6016
rect 18321 5952 18337 6016
rect 18401 5952 18407 6016
rect 18091 5951 18407 5952
rect 29521 6016 29837 6017
rect 29521 5952 29527 6016
rect 29591 5952 29607 6016
rect 29671 5952 29687 6016
rect 29751 5952 29767 6016
rect 29831 5952 29837 6016
rect 29521 5951 29837 5952
rect 40951 6016 41267 6017
rect 40951 5952 40957 6016
rect 41021 5952 41037 6016
rect 41101 5952 41117 6016
rect 41181 5952 41197 6016
rect 41261 5952 41267 6016
rect 40951 5951 41267 5952
rect 12376 5472 12692 5473
rect 12376 5408 12382 5472
rect 12446 5408 12462 5472
rect 12526 5408 12542 5472
rect 12606 5408 12622 5472
rect 12686 5408 12692 5472
rect 12376 5407 12692 5408
rect 23806 5472 24122 5473
rect 23806 5408 23812 5472
rect 23876 5408 23892 5472
rect 23956 5408 23972 5472
rect 24036 5408 24052 5472
rect 24116 5408 24122 5472
rect 23806 5407 24122 5408
rect 35236 5472 35552 5473
rect 35236 5408 35242 5472
rect 35306 5408 35322 5472
rect 35386 5408 35402 5472
rect 35466 5408 35482 5472
rect 35546 5408 35552 5472
rect 35236 5407 35552 5408
rect 46666 5472 46982 5473
rect 46666 5408 46672 5472
rect 46736 5408 46752 5472
rect 46816 5408 46832 5472
rect 46896 5408 46912 5472
rect 46976 5408 46982 5472
rect 46666 5407 46982 5408
rect 6661 4928 6977 4929
rect 6661 4864 6667 4928
rect 6731 4864 6747 4928
rect 6811 4864 6827 4928
rect 6891 4864 6907 4928
rect 6971 4864 6977 4928
rect 6661 4863 6977 4864
rect 18091 4928 18407 4929
rect 18091 4864 18097 4928
rect 18161 4864 18177 4928
rect 18241 4864 18257 4928
rect 18321 4864 18337 4928
rect 18401 4864 18407 4928
rect 18091 4863 18407 4864
rect 29521 4928 29837 4929
rect 29521 4864 29527 4928
rect 29591 4864 29607 4928
rect 29671 4864 29687 4928
rect 29751 4864 29767 4928
rect 29831 4864 29837 4928
rect 29521 4863 29837 4864
rect 40951 4928 41267 4929
rect 40951 4864 40957 4928
rect 41021 4864 41037 4928
rect 41101 4864 41117 4928
rect 41181 4864 41197 4928
rect 41261 4864 41267 4928
rect 40951 4863 41267 4864
rect 12376 4384 12692 4385
rect 12376 4320 12382 4384
rect 12446 4320 12462 4384
rect 12526 4320 12542 4384
rect 12606 4320 12622 4384
rect 12686 4320 12692 4384
rect 12376 4319 12692 4320
rect 23806 4384 24122 4385
rect 23806 4320 23812 4384
rect 23876 4320 23892 4384
rect 23956 4320 23972 4384
rect 24036 4320 24052 4384
rect 24116 4320 24122 4384
rect 23806 4319 24122 4320
rect 35236 4384 35552 4385
rect 35236 4320 35242 4384
rect 35306 4320 35322 4384
rect 35386 4320 35402 4384
rect 35466 4320 35482 4384
rect 35546 4320 35552 4384
rect 35236 4319 35552 4320
rect 46666 4384 46982 4385
rect 46666 4320 46672 4384
rect 46736 4320 46752 4384
rect 46816 4320 46832 4384
rect 46896 4320 46912 4384
rect 46976 4320 46982 4384
rect 46666 4319 46982 4320
rect 17769 4178 17835 4181
rect 41597 4178 41663 4181
rect 17769 4176 41663 4178
rect 17769 4120 17774 4176
rect 17830 4120 41602 4176
rect 41658 4120 41663 4176
rect 17769 4118 41663 4120
rect 17769 4115 17835 4118
rect 41597 4115 41663 4118
rect 17309 4042 17375 4045
rect 36261 4042 36327 4045
rect 17309 4040 36327 4042
rect 17309 3984 17314 4040
rect 17370 3984 36266 4040
rect 36322 3984 36327 4040
rect 17309 3982 36327 3984
rect 17309 3979 17375 3982
rect 36261 3979 36327 3982
rect 6661 3840 6977 3841
rect 6661 3776 6667 3840
rect 6731 3776 6747 3840
rect 6811 3776 6827 3840
rect 6891 3776 6907 3840
rect 6971 3776 6977 3840
rect 6661 3775 6977 3776
rect 18091 3840 18407 3841
rect 18091 3776 18097 3840
rect 18161 3776 18177 3840
rect 18241 3776 18257 3840
rect 18321 3776 18337 3840
rect 18401 3776 18407 3840
rect 18091 3775 18407 3776
rect 29521 3840 29837 3841
rect 29521 3776 29527 3840
rect 29591 3776 29607 3840
rect 29671 3776 29687 3840
rect 29751 3776 29767 3840
rect 29831 3776 29837 3840
rect 29521 3775 29837 3776
rect 40951 3840 41267 3841
rect 40951 3776 40957 3840
rect 41021 3776 41037 3840
rect 41101 3776 41117 3840
rect 41181 3776 41197 3840
rect 41261 3776 41267 3840
rect 40951 3775 41267 3776
rect 21357 3770 21423 3773
rect 28257 3770 28323 3773
rect 21357 3768 28323 3770
rect 21357 3712 21362 3768
rect 21418 3712 28262 3768
rect 28318 3712 28323 3768
rect 21357 3710 28323 3712
rect 21357 3707 21423 3710
rect 28257 3707 28323 3710
rect 15929 3634 15995 3637
rect 38929 3634 38995 3637
rect 15929 3632 38995 3634
rect 15929 3576 15934 3632
rect 15990 3576 38934 3632
rect 38990 3576 38995 3632
rect 15929 3574 38995 3576
rect 15929 3571 15995 3574
rect 38929 3571 38995 3574
rect 12065 3498 12131 3501
rect 30557 3498 30623 3501
rect 12065 3496 30623 3498
rect 12065 3440 12070 3496
rect 12126 3440 30562 3496
rect 30618 3440 30623 3496
rect 12065 3438 30623 3440
rect 12065 3435 12131 3438
rect 30557 3435 30623 3438
rect 12376 3296 12692 3297
rect 12376 3232 12382 3296
rect 12446 3232 12462 3296
rect 12526 3232 12542 3296
rect 12606 3232 12622 3296
rect 12686 3232 12692 3296
rect 12376 3231 12692 3232
rect 23806 3296 24122 3297
rect 23806 3232 23812 3296
rect 23876 3232 23892 3296
rect 23956 3232 23972 3296
rect 24036 3232 24052 3296
rect 24116 3232 24122 3296
rect 23806 3231 24122 3232
rect 35236 3296 35552 3297
rect 35236 3232 35242 3296
rect 35306 3232 35322 3296
rect 35386 3232 35402 3296
rect 35466 3232 35482 3296
rect 35546 3232 35552 3296
rect 35236 3231 35552 3232
rect 46666 3296 46982 3297
rect 46666 3232 46672 3296
rect 46736 3232 46752 3296
rect 46816 3232 46832 3296
rect 46896 3232 46912 3296
rect 46976 3232 46982 3296
rect 46666 3231 46982 3232
rect 9857 3090 9923 3093
rect 25957 3090 26023 3093
rect 9857 3088 26023 3090
rect 9857 3032 9862 3088
rect 9918 3032 25962 3088
rect 26018 3032 26023 3088
rect 9857 3030 26023 3032
rect 9857 3027 9923 3030
rect 25957 3027 26023 3030
rect 26141 3090 26207 3093
rect 34789 3090 34855 3093
rect 26141 3088 34855 3090
rect 26141 3032 26146 3088
rect 26202 3032 34794 3088
rect 34850 3032 34855 3088
rect 26141 3030 34855 3032
rect 26141 3027 26207 3030
rect 34789 3027 34855 3030
rect 13997 2954 14063 2957
rect 21357 2954 21423 2957
rect 13997 2952 21423 2954
rect 13997 2896 14002 2952
rect 14058 2896 21362 2952
rect 21418 2896 21423 2952
rect 13997 2894 21423 2896
rect 13997 2891 14063 2894
rect 21357 2891 21423 2894
rect 22829 2954 22895 2957
rect 30230 2954 30236 2956
rect 22829 2952 30236 2954
rect 22829 2896 22834 2952
rect 22890 2896 30236 2952
rect 22829 2894 30236 2896
rect 22829 2891 22895 2894
rect 30230 2892 30236 2894
rect 30300 2892 30306 2956
rect 18873 2818 18939 2821
rect 26141 2818 26207 2821
rect 18873 2816 26207 2818
rect 18873 2760 18878 2816
rect 18934 2760 26146 2816
rect 26202 2760 26207 2816
rect 18873 2758 26207 2760
rect 18873 2755 18939 2758
rect 26141 2755 26207 2758
rect 6661 2752 6977 2753
rect 6661 2688 6667 2752
rect 6731 2688 6747 2752
rect 6811 2688 6827 2752
rect 6891 2688 6907 2752
rect 6971 2688 6977 2752
rect 6661 2687 6977 2688
rect 18091 2752 18407 2753
rect 18091 2688 18097 2752
rect 18161 2688 18177 2752
rect 18241 2688 18257 2752
rect 18321 2688 18337 2752
rect 18401 2688 18407 2752
rect 18091 2687 18407 2688
rect 29521 2752 29837 2753
rect 29521 2688 29527 2752
rect 29591 2688 29607 2752
rect 29671 2688 29687 2752
rect 29751 2688 29767 2752
rect 29831 2688 29837 2752
rect 29521 2687 29837 2688
rect 40951 2752 41267 2753
rect 40951 2688 40957 2752
rect 41021 2688 41037 2752
rect 41101 2688 41117 2752
rect 41181 2688 41197 2752
rect 41261 2688 41267 2752
rect 40951 2687 41267 2688
rect 20529 2546 20595 2549
rect 38653 2546 38719 2549
rect 20529 2544 38719 2546
rect 20529 2488 20534 2544
rect 20590 2488 38658 2544
rect 38714 2488 38719 2544
rect 20529 2486 38719 2488
rect 20529 2483 20595 2486
rect 38653 2483 38719 2486
rect 8661 2410 8727 2413
rect 23657 2410 23723 2413
rect 8661 2408 23723 2410
rect 8661 2352 8666 2408
rect 8722 2352 23662 2408
rect 23718 2352 23723 2408
rect 8661 2350 23723 2352
rect 8661 2347 8727 2350
rect 23657 2347 23723 2350
rect 26601 2410 26667 2413
rect 39113 2410 39179 2413
rect 26601 2408 39179 2410
rect 26601 2352 26606 2408
rect 26662 2352 39118 2408
rect 39174 2352 39179 2408
rect 26601 2350 39179 2352
rect 26601 2347 26667 2350
rect 39113 2347 39179 2350
rect 19333 2274 19399 2277
rect 21633 2274 21699 2277
rect 19333 2272 21699 2274
rect 19333 2216 19338 2272
rect 19394 2216 21638 2272
rect 21694 2216 21699 2272
rect 19333 2214 21699 2216
rect 19333 2211 19399 2214
rect 21633 2211 21699 2214
rect 30373 2276 30439 2277
rect 30373 2272 30420 2276
rect 30484 2274 30490 2276
rect 30373 2216 30378 2272
rect 30373 2212 30420 2216
rect 30484 2214 30530 2274
rect 30484 2212 30490 2214
rect 30373 2211 30439 2212
rect 12376 2208 12692 2209
rect 12376 2144 12382 2208
rect 12446 2144 12462 2208
rect 12526 2144 12542 2208
rect 12606 2144 12622 2208
rect 12686 2144 12692 2208
rect 12376 2143 12692 2144
rect 23806 2208 24122 2209
rect 23806 2144 23812 2208
rect 23876 2144 23892 2208
rect 23956 2144 23972 2208
rect 24036 2144 24052 2208
rect 24116 2144 24122 2208
rect 23806 2143 24122 2144
rect 35236 2208 35552 2209
rect 35236 2144 35242 2208
rect 35306 2144 35322 2208
rect 35386 2144 35402 2208
rect 35466 2144 35482 2208
rect 35546 2144 35552 2208
rect 35236 2143 35552 2144
rect 46666 2208 46982 2209
rect 46666 2144 46672 2208
rect 46736 2144 46752 2208
rect 46816 2144 46832 2208
rect 46896 2144 46912 2208
rect 46976 2144 46982 2208
rect 46666 2143 46982 2144
rect 16481 2138 16547 2141
rect 24393 2138 24459 2141
rect 32489 2138 32555 2141
rect 16481 2136 22110 2138
rect 16481 2080 16486 2136
rect 16542 2080 22110 2136
rect 16481 2078 22110 2080
rect 16481 2075 16547 2078
rect 16573 2002 16639 2005
rect 19701 2002 19767 2005
rect 16573 2000 19767 2002
rect 16573 1944 16578 2000
rect 16634 1944 19706 2000
rect 19762 1944 19767 2000
rect 16573 1942 19767 1944
rect 16573 1939 16639 1942
rect 19701 1939 19767 1942
rect 19885 2002 19951 2005
rect 20253 2002 20319 2005
rect 19885 2000 20319 2002
rect 19885 1944 19890 2000
rect 19946 1944 20258 2000
rect 20314 1944 20319 2000
rect 19885 1942 20319 1944
rect 22050 2002 22110 2078
rect 24393 2136 32555 2138
rect 24393 2080 24398 2136
rect 24454 2080 32494 2136
rect 32550 2080 32555 2136
rect 24393 2078 32555 2080
rect 24393 2075 24459 2078
rect 32489 2075 32555 2078
rect 38193 2002 38259 2005
rect 22050 2000 38259 2002
rect 22050 1944 38198 2000
rect 38254 1944 38259 2000
rect 22050 1942 38259 1944
rect 19885 1939 19951 1942
rect 20253 1939 20319 1942
rect 38193 1939 38259 1942
rect 16205 1866 16271 1869
rect 36077 1866 36143 1869
rect 16205 1864 36143 1866
rect 16205 1808 16210 1864
rect 16266 1808 36082 1864
rect 36138 1808 36143 1864
rect 16205 1806 36143 1808
rect 16205 1803 16271 1806
rect 36077 1803 36143 1806
rect 18965 1730 19031 1733
rect 22093 1730 22159 1733
rect 18965 1728 22159 1730
rect 18965 1672 18970 1728
rect 19026 1672 22098 1728
rect 22154 1672 22159 1728
rect 18965 1670 22159 1672
rect 18965 1667 19031 1670
rect 22093 1667 22159 1670
rect 31017 1730 31083 1733
rect 38469 1730 38535 1733
rect 31017 1728 38535 1730
rect 31017 1672 31022 1728
rect 31078 1672 38474 1728
rect 38530 1672 38535 1728
rect 31017 1670 38535 1672
rect 31017 1667 31083 1670
rect 38469 1667 38535 1670
rect 6661 1664 6977 1665
rect 6661 1600 6667 1664
rect 6731 1600 6747 1664
rect 6811 1600 6827 1664
rect 6891 1600 6907 1664
rect 6971 1600 6977 1664
rect 6661 1599 6977 1600
rect 18091 1664 18407 1665
rect 18091 1600 18097 1664
rect 18161 1600 18177 1664
rect 18241 1600 18257 1664
rect 18321 1600 18337 1664
rect 18401 1600 18407 1664
rect 18091 1599 18407 1600
rect 29521 1664 29837 1665
rect 29521 1600 29527 1664
rect 29591 1600 29607 1664
rect 29671 1600 29687 1664
rect 29751 1600 29767 1664
rect 29831 1600 29837 1664
rect 29521 1599 29837 1600
rect 40951 1664 41267 1665
rect 40951 1600 40957 1664
rect 41021 1600 41037 1664
rect 41101 1600 41117 1664
rect 41181 1600 41197 1664
rect 41261 1600 41267 1664
rect 40951 1599 41267 1600
rect 18505 1594 18571 1597
rect 30465 1594 30531 1597
rect 33685 1594 33751 1597
rect 18505 1592 22110 1594
rect 18505 1536 18510 1592
rect 18566 1536 22110 1592
rect 18505 1534 22110 1536
rect 18505 1531 18571 1534
rect 14733 1458 14799 1461
rect 21357 1458 21423 1461
rect 14733 1456 21423 1458
rect 14733 1400 14738 1456
rect 14794 1400 21362 1456
rect 21418 1400 21423 1456
rect 14733 1398 21423 1400
rect 22050 1458 22110 1534
rect 30465 1592 33751 1594
rect 30465 1536 30470 1592
rect 30526 1536 33690 1592
rect 33746 1536 33751 1592
rect 30465 1534 33751 1536
rect 30465 1531 30531 1534
rect 33685 1531 33751 1534
rect 37365 1458 37431 1461
rect 22050 1456 37431 1458
rect 22050 1400 37370 1456
rect 37426 1400 37431 1456
rect 22050 1398 37431 1400
rect 14733 1395 14799 1398
rect 21357 1395 21423 1398
rect 37365 1395 37431 1398
rect 11237 1322 11303 1325
rect 18873 1322 18939 1325
rect 11237 1320 18939 1322
rect 11237 1264 11242 1320
rect 11298 1264 18878 1320
rect 18934 1264 18939 1320
rect 11237 1262 18939 1264
rect 11237 1259 11303 1262
rect 18873 1259 18939 1262
rect 19701 1322 19767 1325
rect 24301 1322 24367 1325
rect 19701 1320 24367 1322
rect 19701 1264 19706 1320
rect 19762 1264 24306 1320
rect 24362 1264 24367 1320
rect 19701 1262 24367 1264
rect 19701 1259 19767 1262
rect 24301 1259 24367 1262
rect 30230 1260 30236 1324
rect 30300 1322 30306 1324
rect 43161 1322 43227 1325
rect 30300 1320 43227 1322
rect 30300 1264 43166 1320
rect 43222 1264 43227 1320
rect 30300 1262 43227 1264
rect 30300 1260 30306 1262
rect 43161 1259 43227 1262
rect 15101 1186 15167 1189
rect 22001 1186 22067 1189
rect 31477 1186 31543 1189
rect 15101 1184 22067 1186
rect 15101 1128 15106 1184
rect 15162 1128 22006 1184
rect 22062 1128 22067 1184
rect 15101 1126 22067 1128
rect 15101 1123 15167 1126
rect 22001 1123 22067 1126
rect 26742 1184 31543 1186
rect 26742 1128 31482 1184
rect 31538 1128 31543 1184
rect 26742 1126 31543 1128
rect 12376 1120 12692 1121
rect 12376 1056 12382 1120
rect 12446 1056 12462 1120
rect 12526 1056 12542 1120
rect 12606 1056 12622 1120
rect 12686 1056 12692 1120
rect 12376 1055 12692 1056
rect 23806 1120 24122 1121
rect 23806 1056 23812 1120
rect 23876 1056 23892 1120
rect 23956 1056 23972 1120
rect 24036 1056 24052 1120
rect 24116 1056 24122 1120
rect 23806 1055 24122 1056
rect 13169 1050 13235 1053
rect 17493 1050 17559 1053
rect 13169 1048 17559 1050
rect 13169 992 13174 1048
rect 13230 992 17498 1048
rect 17554 992 17559 1048
rect 13169 990 17559 992
rect 13169 987 13235 990
rect 17493 987 17559 990
rect 10961 914 11027 917
rect 26742 914 26802 1126
rect 31477 1123 31543 1126
rect 35236 1120 35552 1121
rect 35236 1056 35242 1120
rect 35306 1056 35322 1120
rect 35386 1056 35402 1120
rect 35466 1056 35482 1120
rect 35546 1056 35552 1120
rect 35236 1055 35552 1056
rect 46666 1120 46982 1121
rect 46666 1056 46672 1120
rect 46736 1056 46752 1120
rect 46816 1056 46832 1120
rect 46896 1056 46912 1120
rect 46976 1056 46982 1120
rect 46666 1055 46982 1056
rect 33317 914 33383 917
rect 10961 912 26802 914
rect 10961 856 10966 912
rect 11022 856 26802 912
rect 10961 854 26802 856
rect 29134 912 33383 914
rect 29134 856 33322 912
rect 33378 856 33383 912
rect 29134 854 33383 856
rect 10961 851 11027 854
rect 19609 778 19675 781
rect 28993 778 29059 781
rect 19609 776 29059 778
rect 19609 720 19614 776
rect 19670 720 28998 776
rect 29054 720 29059 776
rect 19609 718 29059 720
rect 19609 715 19675 718
rect 28993 715 29059 718
rect 12617 642 12683 645
rect 21449 642 21515 645
rect 12617 640 21515 642
rect 12617 584 12622 640
rect 12678 584 21454 640
rect 21510 584 21515 640
rect 12617 582 21515 584
rect 12617 579 12683 582
rect 21449 579 21515 582
rect 9489 506 9555 509
rect 29134 506 29194 854
rect 33317 851 33383 854
rect 32857 778 32923 781
rect 9489 504 29194 506
rect 9489 448 9494 504
rect 9550 448 29194 504
rect 9489 446 29194 448
rect 31710 776 32923 778
rect 31710 720 32862 776
rect 32918 720 32923 776
rect 31710 718 32923 720
rect 9489 443 9555 446
rect 9121 370 9187 373
rect 31710 370 31770 718
rect 32857 715 32923 718
rect 9121 368 31770 370
rect 9121 312 9126 368
rect 9182 312 31770 368
rect 9121 310 31770 312
rect 9121 307 9187 310
rect 10593 234 10659 237
rect 30414 234 30420 236
rect 10593 232 30420 234
rect 10593 176 10598 232
rect 10654 176 30420 232
rect 10593 174 30420 176
rect 10593 171 10659 174
rect 30414 172 30420 174
rect 30484 172 30490 236
rect 32489 234 32555 237
rect 31710 232 32555 234
rect 31710 176 32494 232
rect 32550 176 32555 232
rect 31710 174 32555 176
rect 19057 98 19123 101
rect 31710 98 31770 174
rect 32489 171 32555 174
rect 19057 96 31770 98
rect 19057 40 19062 96
rect 19118 40 31770 96
rect 19057 38 31770 40
rect 19057 35 19123 38
<< via3 >>
rect 12382 8732 12446 8736
rect 12382 8676 12386 8732
rect 12386 8676 12442 8732
rect 12442 8676 12446 8732
rect 12382 8672 12446 8676
rect 12462 8732 12526 8736
rect 12462 8676 12466 8732
rect 12466 8676 12522 8732
rect 12522 8676 12526 8732
rect 12462 8672 12526 8676
rect 12542 8732 12606 8736
rect 12542 8676 12546 8732
rect 12546 8676 12602 8732
rect 12602 8676 12606 8732
rect 12542 8672 12606 8676
rect 12622 8732 12686 8736
rect 12622 8676 12626 8732
rect 12626 8676 12682 8732
rect 12682 8676 12686 8732
rect 12622 8672 12686 8676
rect 23812 8732 23876 8736
rect 23812 8676 23816 8732
rect 23816 8676 23872 8732
rect 23872 8676 23876 8732
rect 23812 8672 23876 8676
rect 23892 8732 23956 8736
rect 23892 8676 23896 8732
rect 23896 8676 23952 8732
rect 23952 8676 23956 8732
rect 23892 8672 23956 8676
rect 23972 8732 24036 8736
rect 23972 8676 23976 8732
rect 23976 8676 24032 8732
rect 24032 8676 24036 8732
rect 23972 8672 24036 8676
rect 24052 8732 24116 8736
rect 24052 8676 24056 8732
rect 24056 8676 24112 8732
rect 24112 8676 24116 8732
rect 24052 8672 24116 8676
rect 35242 8732 35306 8736
rect 35242 8676 35246 8732
rect 35246 8676 35302 8732
rect 35302 8676 35306 8732
rect 35242 8672 35306 8676
rect 35322 8732 35386 8736
rect 35322 8676 35326 8732
rect 35326 8676 35382 8732
rect 35382 8676 35386 8732
rect 35322 8672 35386 8676
rect 35402 8732 35466 8736
rect 35402 8676 35406 8732
rect 35406 8676 35462 8732
rect 35462 8676 35466 8732
rect 35402 8672 35466 8676
rect 35482 8732 35546 8736
rect 35482 8676 35486 8732
rect 35486 8676 35542 8732
rect 35542 8676 35546 8732
rect 35482 8672 35546 8676
rect 46672 8732 46736 8736
rect 46672 8676 46676 8732
rect 46676 8676 46732 8732
rect 46732 8676 46736 8732
rect 46672 8672 46736 8676
rect 46752 8732 46816 8736
rect 46752 8676 46756 8732
rect 46756 8676 46812 8732
rect 46812 8676 46816 8732
rect 46752 8672 46816 8676
rect 46832 8732 46896 8736
rect 46832 8676 46836 8732
rect 46836 8676 46892 8732
rect 46892 8676 46896 8732
rect 46832 8672 46896 8676
rect 46912 8732 46976 8736
rect 46912 8676 46916 8732
rect 46916 8676 46972 8732
rect 46972 8676 46976 8732
rect 46912 8672 46976 8676
rect 6667 8188 6731 8192
rect 6667 8132 6671 8188
rect 6671 8132 6727 8188
rect 6727 8132 6731 8188
rect 6667 8128 6731 8132
rect 6747 8188 6811 8192
rect 6747 8132 6751 8188
rect 6751 8132 6807 8188
rect 6807 8132 6811 8188
rect 6747 8128 6811 8132
rect 6827 8188 6891 8192
rect 6827 8132 6831 8188
rect 6831 8132 6887 8188
rect 6887 8132 6891 8188
rect 6827 8128 6891 8132
rect 6907 8188 6971 8192
rect 6907 8132 6911 8188
rect 6911 8132 6967 8188
rect 6967 8132 6971 8188
rect 6907 8128 6971 8132
rect 18097 8188 18161 8192
rect 18097 8132 18101 8188
rect 18101 8132 18157 8188
rect 18157 8132 18161 8188
rect 18097 8128 18161 8132
rect 18177 8188 18241 8192
rect 18177 8132 18181 8188
rect 18181 8132 18237 8188
rect 18237 8132 18241 8188
rect 18177 8128 18241 8132
rect 18257 8188 18321 8192
rect 18257 8132 18261 8188
rect 18261 8132 18317 8188
rect 18317 8132 18321 8188
rect 18257 8128 18321 8132
rect 18337 8188 18401 8192
rect 18337 8132 18341 8188
rect 18341 8132 18397 8188
rect 18397 8132 18401 8188
rect 18337 8128 18401 8132
rect 29527 8188 29591 8192
rect 29527 8132 29531 8188
rect 29531 8132 29587 8188
rect 29587 8132 29591 8188
rect 29527 8128 29591 8132
rect 29607 8188 29671 8192
rect 29607 8132 29611 8188
rect 29611 8132 29667 8188
rect 29667 8132 29671 8188
rect 29607 8128 29671 8132
rect 29687 8188 29751 8192
rect 29687 8132 29691 8188
rect 29691 8132 29747 8188
rect 29747 8132 29751 8188
rect 29687 8128 29751 8132
rect 29767 8188 29831 8192
rect 29767 8132 29771 8188
rect 29771 8132 29827 8188
rect 29827 8132 29831 8188
rect 29767 8128 29831 8132
rect 40957 8188 41021 8192
rect 40957 8132 40961 8188
rect 40961 8132 41017 8188
rect 41017 8132 41021 8188
rect 40957 8128 41021 8132
rect 41037 8188 41101 8192
rect 41037 8132 41041 8188
rect 41041 8132 41097 8188
rect 41097 8132 41101 8188
rect 41037 8128 41101 8132
rect 41117 8188 41181 8192
rect 41117 8132 41121 8188
rect 41121 8132 41177 8188
rect 41177 8132 41181 8188
rect 41117 8128 41181 8132
rect 41197 8188 41261 8192
rect 41197 8132 41201 8188
rect 41201 8132 41257 8188
rect 41257 8132 41261 8188
rect 41197 8128 41261 8132
rect 12382 7644 12446 7648
rect 12382 7588 12386 7644
rect 12386 7588 12442 7644
rect 12442 7588 12446 7644
rect 12382 7584 12446 7588
rect 12462 7644 12526 7648
rect 12462 7588 12466 7644
rect 12466 7588 12522 7644
rect 12522 7588 12526 7644
rect 12462 7584 12526 7588
rect 12542 7644 12606 7648
rect 12542 7588 12546 7644
rect 12546 7588 12602 7644
rect 12602 7588 12606 7644
rect 12542 7584 12606 7588
rect 12622 7644 12686 7648
rect 12622 7588 12626 7644
rect 12626 7588 12682 7644
rect 12682 7588 12686 7644
rect 12622 7584 12686 7588
rect 23812 7644 23876 7648
rect 23812 7588 23816 7644
rect 23816 7588 23872 7644
rect 23872 7588 23876 7644
rect 23812 7584 23876 7588
rect 23892 7644 23956 7648
rect 23892 7588 23896 7644
rect 23896 7588 23952 7644
rect 23952 7588 23956 7644
rect 23892 7584 23956 7588
rect 23972 7644 24036 7648
rect 23972 7588 23976 7644
rect 23976 7588 24032 7644
rect 24032 7588 24036 7644
rect 23972 7584 24036 7588
rect 24052 7644 24116 7648
rect 24052 7588 24056 7644
rect 24056 7588 24112 7644
rect 24112 7588 24116 7644
rect 24052 7584 24116 7588
rect 35242 7644 35306 7648
rect 35242 7588 35246 7644
rect 35246 7588 35302 7644
rect 35302 7588 35306 7644
rect 35242 7584 35306 7588
rect 35322 7644 35386 7648
rect 35322 7588 35326 7644
rect 35326 7588 35382 7644
rect 35382 7588 35386 7644
rect 35322 7584 35386 7588
rect 35402 7644 35466 7648
rect 35402 7588 35406 7644
rect 35406 7588 35462 7644
rect 35462 7588 35466 7644
rect 35402 7584 35466 7588
rect 35482 7644 35546 7648
rect 35482 7588 35486 7644
rect 35486 7588 35542 7644
rect 35542 7588 35546 7644
rect 35482 7584 35546 7588
rect 46672 7644 46736 7648
rect 46672 7588 46676 7644
rect 46676 7588 46732 7644
rect 46732 7588 46736 7644
rect 46672 7584 46736 7588
rect 46752 7644 46816 7648
rect 46752 7588 46756 7644
rect 46756 7588 46812 7644
rect 46812 7588 46816 7644
rect 46752 7584 46816 7588
rect 46832 7644 46896 7648
rect 46832 7588 46836 7644
rect 46836 7588 46892 7644
rect 46892 7588 46896 7644
rect 46832 7584 46896 7588
rect 46912 7644 46976 7648
rect 46912 7588 46916 7644
rect 46916 7588 46972 7644
rect 46972 7588 46976 7644
rect 46912 7584 46976 7588
rect 6667 7100 6731 7104
rect 6667 7044 6671 7100
rect 6671 7044 6727 7100
rect 6727 7044 6731 7100
rect 6667 7040 6731 7044
rect 6747 7100 6811 7104
rect 6747 7044 6751 7100
rect 6751 7044 6807 7100
rect 6807 7044 6811 7100
rect 6747 7040 6811 7044
rect 6827 7100 6891 7104
rect 6827 7044 6831 7100
rect 6831 7044 6887 7100
rect 6887 7044 6891 7100
rect 6827 7040 6891 7044
rect 6907 7100 6971 7104
rect 6907 7044 6911 7100
rect 6911 7044 6967 7100
rect 6967 7044 6971 7100
rect 6907 7040 6971 7044
rect 18097 7100 18161 7104
rect 18097 7044 18101 7100
rect 18101 7044 18157 7100
rect 18157 7044 18161 7100
rect 18097 7040 18161 7044
rect 18177 7100 18241 7104
rect 18177 7044 18181 7100
rect 18181 7044 18237 7100
rect 18237 7044 18241 7100
rect 18177 7040 18241 7044
rect 18257 7100 18321 7104
rect 18257 7044 18261 7100
rect 18261 7044 18317 7100
rect 18317 7044 18321 7100
rect 18257 7040 18321 7044
rect 18337 7100 18401 7104
rect 18337 7044 18341 7100
rect 18341 7044 18397 7100
rect 18397 7044 18401 7100
rect 18337 7040 18401 7044
rect 29527 7100 29591 7104
rect 29527 7044 29531 7100
rect 29531 7044 29587 7100
rect 29587 7044 29591 7100
rect 29527 7040 29591 7044
rect 29607 7100 29671 7104
rect 29607 7044 29611 7100
rect 29611 7044 29667 7100
rect 29667 7044 29671 7100
rect 29607 7040 29671 7044
rect 29687 7100 29751 7104
rect 29687 7044 29691 7100
rect 29691 7044 29747 7100
rect 29747 7044 29751 7100
rect 29687 7040 29751 7044
rect 29767 7100 29831 7104
rect 29767 7044 29771 7100
rect 29771 7044 29827 7100
rect 29827 7044 29831 7100
rect 29767 7040 29831 7044
rect 40957 7100 41021 7104
rect 40957 7044 40961 7100
rect 40961 7044 41017 7100
rect 41017 7044 41021 7100
rect 40957 7040 41021 7044
rect 41037 7100 41101 7104
rect 41037 7044 41041 7100
rect 41041 7044 41097 7100
rect 41097 7044 41101 7100
rect 41037 7040 41101 7044
rect 41117 7100 41181 7104
rect 41117 7044 41121 7100
rect 41121 7044 41177 7100
rect 41177 7044 41181 7100
rect 41117 7040 41181 7044
rect 41197 7100 41261 7104
rect 41197 7044 41201 7100
rect 41201 7044 41257 7100
rect 41257 7044 41261 7100
rect 41197 7040 41261 7044
rect 12382 6556 12446 6560
rect 12382 6500 12386 6556
rect 12386 6500 12442 6556
rect 12442 6500 12446 6556
rect 12382 6496 12446 6500
rect 12462 6556 12526 6560
rect 12462 6500 12466 6556
rect 12466 6500 12522 6556
rect 12522 6500 12526 6556
rect 12462 6496 12526 6500
rect 12542 6556 12606 6560
rect 12542 6500 12546 6556
rect 12546 6500 12602 6556
rect 12602 6500 12606 6556
rect 12542 6496 12606 6500
rect 12622 6556 12686 6560
rect 12622 6500 12626 6556
rect 12626 6500 12682 6556
rect 12682 6500 12686 6556
rect 12622 6496 12686 6500
rect 23812 6556 23876 6560
rect 23812 6500 23816 6556
rect 23816 6500 23872 6556
rect 23872 6500 23876 6556
rect 23812 6496 23876 6500
rect 23892 6556 23956 6560
rect 23892 6500 23896 6556
rect 23896 6500 23952 6556
rect 23952 6500 23956 6556
rect 23892 6496 23956 6500
rect 23972 6556 24036 6560
rect 23972 6500 23976 6556
rect 23976 6500 24032 6556
rect 24032 6500 24036 6556
rect 23972 6496 24036 6500
rect 24052 6556 24116 6560
rect 24052 6500 24056 6556
rect 24056 6500 24112 6556
rect 24112 6500 24116 6556
rect 24052 6496 24116 6500
rect 35242 6556 35306 6560
rect 35242 6500 35246 6556
rect 35246 6500 35302 6556
rect 35302 6500 35306 6556
rect 35242 6496 35306 6500
rect 35322 6556 35386 6560
rect 35322 6500 35326 6556
rect 35326 6500 35382 6556
rect 35382 6500 35386 6556
rect 35322 6496 35386 6500
rect 35402 6556 35466 6560
rect 35402 6500 35406 6556
rect 35406 6500 35462 6556
rect 35462 6500 35466 6556
rect 35402 6496 35466 6500
rect 35482 6556 35546 6560
rect 35482 6500 35486 6556
rect 35486 6500 35542 6556
rect 35542 6500 35546 6556
rect 35482 6496 35546 6500
rect 46672 6556 46736 6560
rect 46672 6500 46676 6556
rect 46676 6500 46732 6556
rect 46732 6500 46736 6556
rect 46672 6496 46736 6500
rect 46752 6556 46816 6560
rect 46752 6500 46756 6556
rect 46756 6500 46812 6556
rect 46812 6500 46816 6556
rect 46752 6496 46816 6500
rect 46832 6556 46896 6560
rect 46832 6500 46836 6556
rect 46836 6500 46892 6556
rect 46892 6500 46896 6556
rect 46832 6496 46896 6500
rect 46912 6556 46976 6560
rect 46912 6500 46916 6556
rect 46916 6500 46972 6556
rect 46972 6500 46976 6556
rect 46912 6496 46976 6500
rect 6667 6012 6731 6016
rect 6667 5956 6671 6012
rect 6671 5956 6727 6012
rect 6727 5956 6731 6012
rect 6667 5952 6731 5956
rect 6747 6012 6811 6016
rect 6747 5956 6751 6012
rect 6751 5956 6807 6012
rect 6807 5956 6811 6012
rect 6747 5952 6811 5956
rect 6827 6012 6891 6016
rect 6827 5956 6831 6012
rect 6831 5956 6887 6012
rect 6887 5956 6891 6012
rect 6827 5952 6891 5956
rect 6907 6012 6971 6016
rect 6907 5956 6911 6012
rect 6911 5956 6967 6012
rect 6967 5956 6971 6012
rect 6907 5952 6971 5956
rect 18097 6012 18161 6016
rect 18097 5956 18101 6012
rect 18101 5956 18157 6012
rect 18157 5956 18161 6012
rect 18097 5952 18161 5956
rect 18177 6012 18241 6016
rect 18177 5956 18181 6012
rect 18181 5956 18237 6012
rect 18237 5956 18241 6012
rect 18177 5952 18241 5956
rect 18257 6012 18321 6016
rect 18257 5956 18261 6012
rect 18261 5956 18317 6012
rect 18317 5956 18321 6012
rect 18257 5952 18321 5956
rect 18337 6012 18401 6016
rect 18337 5956 18341 6012
rect 18341 5956 18397 6012
rect 18397 5956 18401 6012
rect 18337 5952 18401 5956
rect 29527 6012 29591 6016
rect 29527 5956 29531 6012
rect 29531 5956 29587 6012
rect 29587 5956 29591 6012
rect 29527 5952 29591 5956
rect 29607 6012 29671 6016
rect 29607 5956 29611 6012
rect 29611 5956 29667 6012
rect 29667 5956 29671 6012
rect 29607 5952 29671 5956
rect 29687 6012 29751 6016
rect 29687 5956 29691 6012
rect 29691 5956 29747 6012
rect 29747 5956 29751 6012
rect 29687 5952 29751 5956
rect 29767 6012 29831 6016
rect 29767 5956 29771 6012
rect 29771 5956 29827 6012
rect 29827 5956 29831 6012
rect 29767 5952 29831 5956
rect 40957 6012 41021 6016
rect 40957 5956 40961 6012
rect 40961 5956 41017 6012
rect 41017 5956 41021 6012
rect 40957 5952 41021 5956
rect 41037 6012 41101 6016
rect 41037 5956 41041 6012
rect 41041 5956 41097 6012
rect 41097 5956 41101 6012
rect 41037 5952 41101 5956
rect 41117 6012 41181 6016
rect 41117 5956 41121 6012
rect 41121 5956 41177 6012
rect 41177 5956 41181 6012
rect 41117 5952 41181 5956
rect 41197 6012 41261 6016
rect 41197 5956 41201 6012
rect 41201 5956 41257 6012
rect 41257 5956 41261 6012
rect 41197 5952 41261 5956
rect 12382 5468 12446 5472
rect 12382 5412 12386 5468
rect 12386 5412 12442 5468
rect 12442 5412 12446 5468
rect 12382 5408 12446 5412
rect 12462 5468 12526 5472
rect 12462 5412 12466 5468
rect 12466 5412 12522 5468
rect 12522 5412 12526 5468
rect 12462 5408 12526 5412
rect 12542 5468 12606 5472
rect 12542 5412 12546 5468
rect 12546 5412 12602 5468
rect 12602 5412 12606 5468
rect 12542 5408 12606 5412
rect 12622 5468 12686 5472
rect 12622 5412 12626 5468
rect 12626 5412 12682 5468
rect 12682 5412 12686 5468
rect 12622 5408 12686 5412
rect 23812 5468 23876 5472
rect 23812 5412 23816 5468
rect 23816 5412 23872 5468
rect 23872 5412 23876 5468
rect 23812 5408 23876 5412
rect 23892 5468 23956 5472
rect 23892 5412 23896 5468
rect 23896 5412 23952 5468
rect 23952 5412 23956 5468
rect 23892 5408 23956 5412
rect 23972 5468 24036 5472
rect 23972 5412 23976 5468
rect 23976 5412 24032 5468
rect 24032 5412 24036 5468
rect 23972 5408 24036 5412
rect 24052 5468 24116 5472
rect 24052 5412 24056 5468
rect 24056 5412 24112 5468
rect 24112 5412 24116 5468
rect 24052 5408 24116 5412
rect 35242 5468 35306 5472
rect 35242 5412 35246 5468
rect 35246 5412 35302 5468
rect 35302 5412 35306 5468
rect 35242 5408 35306 5412
rect 35322 5468 35386 5472
rect 35322 5412 35326 5468
rect 35326 5412 35382 5468
rect 35382 5412 35386 5468
rect 35322 5408 35386 5412
rect 35402 5468 35466 5472
rect 35402 5412 35406 5468
rect 35406 5412 35462 5468
rect 35462 5412 35466 5468
rect 35402 5408 35466 5412
rect 35482 5468 35546 5472
rect 35482 5412 35486 5468
rect 35486 5412 35542 5468
rect 35542 5412 35546 5468
rect 35482 5408 35546 5412
rect 46672 5468 46736 5472
rect 46672 5412 46676 5468
rect 46676 5412 46732 5468
rect 46732 5412 46736 5468
rect 46672 5408 46736 5412
rect 46752 5468 46816 5472
rect 46752 5412 46756 5468
rect 46756 5412 46812 5468
rect 46812 5412 46816 5468
rect 46752 5408 46816 5412
rect 46832 5468 46896 5472
rect 46832 5412 46836 5468
rect 46836 5412 46892 5468
rect 46892 5412 46896 5468
rect 46832 5408 46896 5412
rect 46912 5468 46976 5472
rect 46912 5412 46916 5468
rect 46916 5412 46972 5468
rect 46972 5412 46976 5468
rect 46912 5408 46976 5412
rect 6667 4924 6731 4928
rect 6667 4868 6671 4924
rect 6671 4868 6727 4924
rect 6727 4868 6731 4924
rect 6667 4864 6731 4868
rect 6747 4924 6811 4928
rect 6747 4868 6751 4924
rect 6751 4868 6807 4924
rect 6807 4868 6811 4924
rect 6747 4864 6811 4868
rect 6827 4924 6891 4928
rect 6827 4868 6831 4924
rect 6831 4868 6887 4924
rect 6887 4868 6891 4924
rect 6827 4864 6891 4868
rect 6907 4924 6971 4928
rect 6907 4868 6911 4924
rect 6911 4868 6967 4924
rect 6967 4868 6971 4924
rect 6907 4864 6971 4868
rect 18097 4924 18161 4928
rect 18097 4868 18101 4924
rect 18101 4868 18157 4924
rect 18157 4868 18161 4924
rect 18097 4864 18161 4868
rect 18177 4924 18241 4928
rect 18177 4868 18181 4924
rect 18181 4868 18237 4924
rect 18237 4868 18241 4924
rect 18177 4864 18241 4868
rect 18257 4924 18321 4928
rect 18257 4868 18261 4924
rect 18261 4868 18317 4924
rect 18317 4868 18321 4924
rect 18257 4864 18321 4868
rect 18337 4924 18401 4928
rect 18337 4868 18341 4924
rect 18341 4868 18397 4924
rect 18397 4868 18401 4924
rect 18337 4864 18401 4868
rect 29527 4924 29591 4928
rect 29527 4868 29531 4924
rect 29531 4868 29587 4924
rect 29587 4868 29591 4924
rect 29527 4864 29591 4868
rect 29607 4924 29671 4928
rect 29607 4868 29611 4924
rect 29611 4868 29667 4924
rect 29667 4868 29671 4924
rect 29607 4864 29671 4868
rect 29687 4924 29751 4928
rect 29687 4868 29691 4924
rect 29691 4868 29747 4924
rect 29747 4868 29751 4924
rect 29687 4864 29751 4868
rect 29767 4924 29831 4928
rect 29767 4868 29771 4924
rect 29771 4868 29827 4924
rect 29827 4868 29831 4924
rect 29767 4864 29831 4868
rect 40957 4924 41021 4928
rect 40957 4868 40961 4924
rect 40961 4868 41017 4924
rect 41017 4868 41021 4924
rect 40957 4864 41021 4868
rect 41037 4924 41101 4928
rect 41037 4868 41041 4924
rect 41041 4868 41097 4924
rect 41097 4868 41101 4924
rect 41037 4864 41101 4868
rect 41117 4924 41181 4928
rect 41117 4868 41121 4924
rect 41121 4868 41177 4924
rect 41177 4868 41181 4924
rect 41117 4864 41181 4868
rect 41197 4924 41261 4928
rect 41197 4868 41201 4924
rect 41201 4868 41257 4924
rect 41257 4868 41261 4924
rect 41197 4864 41261 4868
rect 12382 4380 12446 4384
rect 12382 4324 12386 4380
rect 12386 4324 12442 4380
rect 12442 4324 12446 4380
rect 12382 4320 12446 4324
rect 12462 4380 12526 4384
rect 12462 4324 12466 4380
rect 12466 4324 12522 4380
rect 12522 4324 12526 4380
rect 12462 4320 12526 4324
rect 12542 4380 12606 4384
rect 12542 4324 12546 4380
rect 12546 4324 12602 4380
rect 12602 4324 12606 4380
rect 12542 4320 12606 4324
rect 12622 4380 12686 4384
rect 12622 4324 12626 4380
rect 12626 4324 12682 4380
rect 12682 4324 12686 4380
rect 12622 4320 12686 4324
rect 23812 4380 23876 4384
rect 23812 4324 23816 4380
rect 23816 4324 23872 4380
rect 23872 4324 23876 4380
rect 23812 4320 23876 4324
rect 23892 4380 23956 4384
rect 23892 4324 23896 4380
rect 23896 4324 23952 4380
rect 23952 4324 23956 4380
rect 23892 4320 23956 4324
rect 23972 4380 24036 4384
rect 23972 4324 23976 4380
rect 23976 4324 24032 4380
rect 24032 4324 24036 4380
rect 23972 4320 24036 4324
rect 24052 4380 24116 4384
rect 24052 4324 24056 4380
rect 24056 4324 24112 4380
rect 24112 4324 24116 4380
rect 24052 4320 24116 4324
rect 35242 4380 35306 4384
rect 35242 4324 35246 4380
rect 35246 4324 35302 4380
rect 35302 4324 35306 4380
rect 35242 4320 35306 4324
rect 35322 4380 35386 4384
rect 35322 4324 35326 4380
rect 35326 4324 35382 4380
rect 35382 4324 35386 4380
rect 35322 4320 35386 4324
rect 35402 4380 35466 4384
rect 35402 4324 35406 4380
rect 35406 4324 35462 4380
rect 35462 4324 35466 4380
rect 35402 4320 35466 4324
rect 35482 4380 35546 4384
rect 35482 4324 35486 4380
rect 35486 4324 35542 4380
rect 35542 4324 35546 4380
rect 35482 4320 35546 4324
rect 46672 4380 46736 4384
rect 46672 4324 46676 4380
rect 46676 4324 46732 4380
rect 46732 4324 46736 4380
rect 46672 4320 46736 4324
rect 46752 4380 46816 4384
rect 46752 4324 46756 4380
rect 46756 4324 46812 4380
rect 46812 4324 46816 4380
rect 46752 4320 46816 4324
rect 46832 4380 46896 4384
rect 46832 4324 46836 4380
rect 46836 4324 46892 4380
rect 46892 4324 46896 4380
rect 46832 4320 46896 4324
rect 46912 4380 46976 4384
rect 46912 4324 46916 4380
rect 46916 4324 46972 4380
rect 46972 4324 46976 4380
rect 46912 4320 46976 4324
rect 6667 3836 6731 3840
rect 6667 3780 6671 3836
rect 6671 3780 6727 3836
rect 6727 3780 6731 3836
rect 6667 3776 6731 3780
rect 6747 3836 6811 3840
rect 6747 3780 6751 3836
rect 6751 3780 6807 3836
rect 6807 3780 6811 3836
rect 6747 3776 6811 3780
rect 6827 3836 6891 3840
rect 6827 3780 6831 3836
rect 6831 3780 6887 3836
rect 6887 3780 6891 3836
rect 6827 3776 6891 3780
rect 6907 3836 6971 3840
rect 6907 3780 6911 3836
rect 6911 3780 6967 3836
rect 6967 3780 6971 3836
rect 6907 3776 6971 3780
rect 18097 3836 18161 3840
rect 18097 3780 18101 3836
rect 18101 3780 18157 3836
rect 18157 3780 18161 3836
rect 18097 3776 18161 3780
rect 18177 3836 18241 3840
rect 18177 3780 18181 3836
rect 18181 3780 18237 3836
rect 18237 3780 18241 3836
rect 18177 3776 18241 3780
rect 18257 3836 18321 3840
rect 18257 3780 18261 3836
rect 18261 3780 18317 3836
rect 18317 3780 18321 3836
rect 18257 3776 18321 3780
rect 18337 3836 18401 3840
rect 18337 3780 18341 3836
rect 18341 3780 18397 3836
rect 18397 3780 18401 3836
rect 18337 3776 18401 3780
rect 29527 3836 29591 3840
rect 29527 3780 29531 3836
rect 29531 3780 29587 3836
rect 29587 3780 29591 3836
rect 29527 3776 29591 3780
rect 29607 3836 29671 3840
rect 29607 3780 29611 3836
rect 29611 3780 29667 3836
rect 29667 3780 29671 3836
rect 29607 3776 29671 3780
rect 29687 3836 29751 3840
rect 29687 3780 29691 3836
rect 29691 3780 29747 3836
rect 29747 3780 29751 3836
rect 29687 3776 29751 3780
rect 29767 3836 29831 3840
rect 29767 3780 29771 3836
rect 29771 3780 29827 3836
rect 29827 3780 29831 3836
rect 29767 3776 29831 3780
rect 40957 3836 41021 3840
rect 40957 3780 40961 3836
rect 40961 3780 41017 3836
rect 41017 3780 41021 3836
rect 40957 3776 41021 3780
rect 41037 3836 41101 3840
rect 41037 3780 41041 3836
rect 41041 3780 41097 3836
rect 41097 3780 41101 3836
rect 41037 3776 41101 3780
rect 41117 3836 41181 3840
rect 41117 3780 41121 3836
rect 41121 3780 41177 3836
rect 41177 3780 41181 3836
rect 41117 3776 41181 3780
rect 41197 3836 41261 3840
rect 41197 3780 41201 3836
rect 41201 3780 41257 3836
rect 41257 3780 41261 3836
rect 41197 3776 41261 3780
rect 12382 3292 12446 3296
rect 12382 3236 12386 3292
rect 12386 3236 12442 3292
rect 12442 3236 12446 3292
rect 12382 3232 12446 3236
rect 12462 3292 12526 3296
rect 12462 3236 12466 3292
rect 12466 3236 12522 3292
rect 12522 3236 12526 3292
rect 12462 3232 12526 3236
rect 12542 3292 12606 3296
rect 12542 3236 12546 3292
rect 12546 3236 12602 3292
rect 12602 3236 12606 3292
rect 12542 3232 12606 3236
rect 12622 3292 12686 3296
rect 12622 3236 12626 3292
rect 12626 3236 12682 3292
rect 12682 3236 12686 3292
rect 12622 3232 12686 3236
rect 23812 3292 23876 3296
rect 23812 3236 23816 3292
rect 23816 3236 23872 3292
rect 23872 3236 23876 3292
rect 23812 3232 23876 3236
rect 23892 3292 23956 3296
rect 23892 3236 23896 3292
rect 23896 3236 23952 3292
rect 23952 3236 23956 3292
rect 23892 3232 23956 3236
rect 23972 3292 24036 3296
rect 23972 3236 23976 3292
rect 23976 3236 24032 3292
rect 24032 3236 24036 3292
rect 23972 3232 24036 3236
rect 24052 3292 24116 3296
rect 24052 3236 24056 3292
rect 24056 3236 24112 3292
rect 24112 3236 24116 3292
rect 24052 3232 24116 3236
rect 35242 3292 35306 3296
rect 35242 3236 35246 3292
rect 35246 3236 35302 3292
rect 35302 3236 35306 3292
rect 35242 3232 35306 3236
rect 35322 3292 35386 3296
rect 35322 3236 35326 3292
rect 35326 3236 35382 3292
rect 35382 3236 35386 3292
rect 35322 3232 35386 3236
rect 35402 3292 35466 3296
rect 35402 3236 35406 3292
rect 35406 3236 35462 3292
rect 35462 3236 35466 3292
rect 35402 3232 35466 3236
rect 35482 3292 35546 3296
rect 35482 3236 35486 3292
rect 35486 3236 35542 3292
rect 35542 3236 35546 3292
rect 35482 3232 35546 3236
rect 46672 3292 46736 3296
rect 46672 3236 46676 3292
rect 46676 3236 46732 3292
rect 46732 3236 46736 3292
rect 46672 3232 46736 3236
rect 46752 3292 46816 3296
rect 46752 3236 46756 3292
rect 46756 3236 46812 3292
rect 46812 3236 46816 3292
rect 46752 3232 46816 3236
rect 46832 3292 46896 3296
rect 46832 3236 46836 3292
rect 46836 3236 46892 3292
rect 46892 3236 46896 3292
rect 46832 3232 46896 3236
rect 46912 3292 46976 3296
rect 46912 3236 46916 3292
rect 46916 3236 46972 3292
rect 46972 3236 46976 3292
rect 46912 3232 46976 3236
rect 30236 2892 30300 2956
rect 6667 2748 6731 2752
rect 6667 2692 6671 2748
rect 6671 2692 6727 2748
rect 6727 2692 6731 2748
rect 6667 2688 6731 2692
rect 6747 2748 6811 2752
rect 6747 2692 6751 2748
rect 6751 2692 6807 2748
rect 6807 2692 6811 2748
rect 6747 2688 6811 2692
rect 6827 2748 6891 2752
rect 6827 2692 6831 2748
rect 6831 2692 6887 2748
rect 6887 2692 6891 2748
rect 6827 2688 6891 2692
rect 6907 2748 6971 2752
rect 6907 2692 6911 2748
rect 6911 2692 6967 2748
rect 6967 2692 6971 2748
rect 6907 2688 6971 2692
rect 18097 2748 18161 2752
rect 18097 2692 18101 2748
rect 18101 2692 18157 2748
rect 18157 2692 18161 2748
rect 18097 2688 18161 2692
rect 18177 2748 18241 2752
rect 18177 2692 18181 2748
rect 18181 2692 18237 2748
rect 18237 2692 18241 2748
rect 18177 2688 18241 2692
rect 18257 2748 18321 2752
rect 18257 2692 18261 2748
rect 18261 2692 18317 2748
rect 18317 2692 18321 2748
rect 18257 2688 18321 2692
rect 18337 2748 18401 2752
rect 18337 2692 18341 2748
rect 18341 2692 18397 2748
rect 18397 2692 18401 2748
rect 18337 2688 18401 2692
rect 29527 2748 29591 2752
rect 29527 2692 29531 2748
rect 29531 2692 29587 2748
rect 29587 2692 29591 2748
rect 29527 2688 29591 2692
rect 29607 2748 29671 2752
rect 29607 2692 29611 2748
rect 29611 2692 29667 2748
rect 29667 2692 29671 2748
rect 29607 2688 29671 2692
rect 29687 2748 29751 2752
rect 29687 2692 29691 2748
rect 29691 2692 29747 2748
rect 29747 2692 29751 2748
rect 29687 2688 29751 2692
rect 29767 2748 29831 2752
rect 29767 2692 29771 2748
rect 29771 2692 29827 2748
rect 29827 2692 29831 2748
rect 29767 2688 29831 2692
rect 40957 2748 41021 2752
rect 40957 2692 40961 2748
rect 40961 2692 41017 2748
rect 41017 2692 41021 2748
rect 40957 2688 41021 2692
rect 41037 2748 41101 2752
rect 41037 2692 41041 2748
rect 41041 2692 41097 2748
rect 41097 2692 41101 2748
rect 41037 2688 41101 2692
rect 41117 2748 41181 2752
rect 41117 2692 41121 2748
rect 41121 2692 41177 2748
rect 41177 2692 41181 2748
rect 41117 2688 41181 2692
rect 41197 2748 41261 2752
rect 41197 2692 41201 2748
rect 41201 2692 41257 2748
rect 41257 2692 41261 2748
rect 41197 2688 41261 2692
rect 30420 2272 30484 2276
rect 30420 2216 30434 2272
rect 30434 2216 30484 2272
rect 30420 2212 30484 2216
rect 12382 2204 12446 2208
rect 12382 2148 12386 2204
rect 12386 2148 12442 2204
rect 12442 2148 12446 2204
rect 12382 2144 12446 2148
rect 12462 2204 12526 2208
rect 12462 2148 12466 2204
rect 12466 2148 12522 2204
rect 12522 2148 12526 2204
rect 12462 2144 12526 2148
rect 12542 2204 12606 2208
rect 12542 2148 12546 2204
rect 12546 2148 12602 2204
rect 12602 2148 12606 2204
rect 12542 2144 12606 2148
rect 12622 2204 12686 2208
rect 12622 2148 12626 2204
rect 12626 2148 12682 2204
rect 12682 2148 12686 2204
rect 12622 2144 12686 2148
rect 23812 2204 23876 2208
rect 23812 2148 23816 2204
rect 23816 2148 23872 2204
rect 23872 2148 23876 2204
rect 23812 2144 23876 2148
rect 23892 2204 23956 2208
rect 23892 2148 23896 2204
rect 23896 2148 23952 2204
rect 23952 2148 23956 2204
rect 23892 2144 23956 2148
rect 23972 2204 24036 2208
rect 23972 2148 23976 2204
rect 23976 2148 24032 2204
rect 24032 2148 24036 2204
rect 23972 2144 24036 2148
rect 24052 2204 24116 2208
rect 24052 2148 24056 2204
rect 24056 2148 24112 2204
rect 24112 2148 24116 2204
rect 24052 2144 24116 2148
rect 35242 2204 35306 2208
rect 35242 2148 35246 2204
rect 35246 2148 35302 2204
rect 35302 2148 35306 2204
rect 35242 2144 35306 2148
rect 35322 2204 35386 2208
rect 35322 2148 35326 2204
rect 35326 2148 35382 2204
rect 35382 2148 35386 2204
rect 35322 2144 35386 2148
rect 35402 2204 35466 2208
rect 35402 2148 35406 2204
rect 35406 2148 35462 2204
rect 35462 2148 35466 2204
rect 35402 2144 35466 2148
rect 35482 2204 35546 2208
rect 35482 2148 35486 2204
rect 35486 2148 35542 2204
rect 35542 2148 35546 2204
rect 35482 2144 35546 2148
rect 46672 2204 46736 2208
rect 46672 2148 46676 2204
rect 46676 2148 46732 2204
rect 46732 2148 46736 2204
rect 46672 2144 46736 2148
rect 46752 2204 46816 2208
rect 46752 2148 46756 2204
rect 46756 2148 46812 2204
rect 46812 2148 46816 2204
rect 46752 2144 46816 2148
rect 46832 2204 46896 2208
rect 46832 2148 46836 2204
rect 46836 2148 46892 2204
rect 46892 2148 46896 2204
rect 46832 2144 46896 2148
rect 46912 2204 46976 2208
rect 46912 2148 46916 2204
rect 46916 2148 46972 2204
rect 46972 2148 46976 2204
rect 46912 2144 46976 2148
rect 6667 1660 6731 1664
rect 6667 1604 6671 1660
rect 6671 1604 6727 1660
rect 6727 1604 6731 1660
rect 6667 1600 6731 1604
rect 6747 1660 6811 1664
rect 6747 1604 6751 1660
rect 6751 1604 6807 1660
rect 6807 1604 6811 1660
rect 6747 1600 6811 1604
rect 6827 1660 6891 1664
rect 6827 1604 6831 1660
rect 6831 1604 6887 1660
rect 6887 1604 6891 1660
rect 6827 1600 6891 1604
rect 6907 1660 6971 1664
rect 6907 1604 6911 1660
rect 6911 1604 6967 1660
rect 6967 1604 6971 1660
rect 6907 1600 6971 1604
rect 18097 1660 18161 1664
rect 18097 1604 18101 1660
rect 18101 1604 18157 1660
rect 18157 1604 18161 1660
rect 18097 1600 18161 1604
rect 18177 1660 18241 1664
rect 18177 1604 18181 1660
rect 18181 1604 18237 1660
rect 18237 1604 18241 1660
rect 18177 1600 18241 1604
rect 18257 1660 18321 1664
rect 18257 1604 18261 1660
rect 18261 1604 18317 1660
rect 18317 1604 18321 1660
rect 18257 1600 18321 1604
rect 18337 1660 18401 1664
rect 18337 1604 18341 1660
rect 18341 1604 18397 1660
rect 18397 1604 18401 1660
rect 18337 1600 18401 1604
rect 29527 1660 29591 1664
rect 29527 1604 29531 1660
rect 29531 1604 29587 1660
rect 29587 1604 29591 1660
rect 29527 1600 29591 1604
rect 29607 1660 29671 1664
rect 29607 1604 29611 1660
rect 29611 1604 29667 1660
rect 29667 1604 29671 1660
rect 29607 1600 29671 1604
rect 29687 1660 29751 1664
rect 29687 1604 29691 1660
rect 29691 1604 29747 1660
rect 29747 1604 29751 1660
rect 29687 1600 29751 1604
rect 29767 1660 29831 1664
rect 29767 1604 29771 1660
rect 29771 1604 29827 1660
rect 29827 1604 29831 1660
rect 29767 1600 29831 1604
rect 40957 1660 41021 1664
rect 40957 1604 40961 1660
rect 40961 1604 41017 1660
rect 41017 1604 41021 1660
rect 40957 1600 41021 1604
rect 41037 1660 41101 1664
rect 41037 1604 41041 1660
rect 41041 1604 41097 1660
rect 41097 1604 41101 1660
rect 41037 1600 41101 1604
rect 41117 1660 41181 1664
rect 41117 1604 41121 1660
rect 41121 1604 41177 1660
rect 41177 1604 41181 1660
rect 41117 1600 41181 1604
rect 41197 1660 41261 1664
rect 41197 1604 41201 1660
rect 41201 1604 41257 1660
rect 41257 1604 41261 1660
rect 41197 1600 41261 1604
rect 30236 1260 30300 1324
rect 12382 1116 12446 1120
rect 12382 1060 12386 1116
rect 12386 1060 12442 1116
rect 12442 1060 12446 1116
rect 12382 1056 12446 1060
rect 12462 1116 12526 1120
rect 12462 1060 12466 1116
rect 12466 1060 12522 1116
rect 12522 1060 12526 1116
rect 12462 1056 12526 1060
rect 12542 1116 12606 1120
rect 12542 1060 12546 1116
rect 12546 1060 12602 1116
rect 12602 1060 12606 1116
rect 12542 1056 12606 1060
rect 12622 1116 12686 1120
rect 12622 1060 12626 1116
rect 12626 1060 12682 1116
rect 12682 1060 12686 1116
rect 12622 1056 12686 1060
rect 23812 1116 23876 1120
rect 23812 1060 23816 1116
rect 23816 1060 23872 1116
rect 23872 1060 23876 1116
rect 23812 1056 23876 1060
rect 23892 1116 23956 1120
rect 23892 1060 23896 1116
rect 23896 1060 23952 1116
rect 23952 1060 23956 1116
rect 23892 1056 23956 1060
rect 23972 1116 24036 1120
rect 23972 1060 23976 1116
rect 23976 1060 24032 1116
rect 24032 1060 24036 1116
rect 23972 1056 24036 1060
rect 24052 1116 24116 1120
rect 24052 1060 24056 1116
rect 24056 1060 24112 1116
rect 24112 1060 24116 1116
rect 24052 1056 24116 1060
rect 35242 1116 35306 1120
rect 35242 1060 35246 1116
rect 35246 1060 35302 1116
rect 35302 1060 35306 1116
rect 35242 1056 35306 1060
rect 35322 1116 35386 1120
rect 35322 1060 35326 1116
rect 35326 1060 35382 1116
rect 35382 1060 35386 1116
rect 35322 1056 35386 1060
rect 35402 1116 35466 1120
rect 35402 1060 35406 1116
rect 35406 1060 35462 1116
rect 35462 1060 35466 1116
rect 35402 1056 35466 1060
rect 35482 1116 35546 1120
rect 35482 1060 35486 1116
rect 35486 1060 35542 1116
rect 35542 1060 35546 1116
rect 35482 1056 35546 1060
rect 46672 1116 46736 1120
rect 46672 1060 46676 1116
rect 46676 1060 46732 1116
rect 46732 1060 46736 1116
rect 46672 1056 46736 1060
rect 46752 1116 46816 1120
rect 46752 1060 46756 1116
rect 46756 1060 46812 1116
rect 46812 1060 46816 1116
rect 46752 1056 46816 1060
rect 46832 1116 46896 1120
rect 46832 1060 46836 1116
rect 46836 1060 46892 1116
rect 46892 1060 46896 1116
rect 46832 1056 46896 1060
rect 46912 1116 46976 1120
rect 46912 1060 46916 1116
rect 46916 1060 46972 1116
rect 46972 1060 46976 1116
rect 46912 1056 46976 1060
rect 30420 172 30484 236
<< metal4 >>
rect 6659 8192 6979 8752
rect 6659 8128 6667 8192
rect 6731 8128 6747 8192
rect 6811 8128 6827 8192
rect 6891 8128 6907 8192
rect 6971 8128 6979 8192
rect 6659 7104 6979 8128
rect 6659 7040 6667 7104
rect 6731 7040 6747 7104
rect 6811 7040 6827 7104
rect 6891 7040 6907 7104
rect 6971 7040 6979 7104
rect 6659 6016 6979 7040
rect 6659 5952 6667 6016
rect 6731 5952 6747 6016
rect 6811 5952 6827 6016
rect 6891 5952 6907 6016
rect 6971 5952 6979 6016
rect 6659 4928 6979 5952
rect 6659 4864 6667 4928
rect 6731 4864 6747 4928
rect 6811 4864 6827 4928
rect 6891 4864 6907 4928
rect 6971 4864 6979 4928
rect 6659 3840 6979 4864
rect 6659 3776 6667 3840
rect 6731 3776 6747 3840
rect 6811 3776 6827 3840
rect 6891 3776 6907 3840
rect 6971 3776 6979 3840
rect 6659 2752 6979 3776
rect 6659 2688 6667 2752
rect 6731 2688 6747 2752
rect 6811 2688 6827 2752
rect 6891 2688 6907 2752
rect 6971 2688 6979 2752
rect 6659 1664 6979 2688
rect 6659 1600 6667 1664
rect 6731 1600 6747 1664
rect 6811 1600 6827 1664
rect 6891 1600 6907 1664
rect 6971 1600 6979 1664
rect 6659 1040 6979 1600
rect 12374 8736 12694 8752
rect 12374 8672 12382 8736
rect 12446 8672 12462 8736
rect 12526 8672 12542 8736
rect 12606 8672 12622 8736
rect 12686 8672 12694 8736
rect 12374 7648 12694 8672
rect 12374 7584 12382 7648
rect 12446 7584 12462 7648
rect 12526 7584 12542 7648
rect 12606 7584 12622 7648
rect 12686 7584 12694 7648
rect 12374 6560 12694 7584
rect 12374 6496 12382 6560
rect 12446 6496 12462 6560
rect 12526 6496 12542 6560
rect 12606 6496 12622 6560
rect 12686 6496 12694 6560
rect 12374 5472 12694 6496
rect 12374 5408 12382 5472
rect 12446 5408 12462 5472
rect 12526 5408 12542 5472
rect 12606 5408 12622 5472
rect 12686 5408 12694 5472
rect 12374 4384 12694 5408
rect 12374 4320 12382 4384
rect 12446 4320 12462 4384
rect 12526 4320 12542 4384
rect 12606 4320 12622 4384
rect 12686 4320 12694 4384
rect 12374 3296 12694 4320
rect 12374 3232 12382 3296
rect 12446 3232 12462 3296
rect 12526 3232 12542 3296
rect 12606 3232 12622 3296
rect 12686 3232 12694 3296
rect 12374 2208 12694 3232
rect 12374 2144 12382 2208
rect 12446 2144 12462 2208
rect 12526 2144 12542 2208
rect 12606 2144 12622 2208
rect 12686 2144 12694 2208
rect 12374 1120 12694 2144
rect 12374 1056 12382 1120
rect 12446 1056 12462 1120
rect 12526 1056 12542 1120
rect 12606 1056 12622 1120
rect 12686 1056 12694 1120
rect 12374 1040 12694 1056
rect 18089 8192 18409 8752
rect 18089 8128 18097 8192
rect 18161 8128 18177 8192
rect 18241 8128 18257 8192
rect 18321 8128 18337 8192
rect 18401 8128 18409 8192
rect 18089 7104 18409 8128
rect 18089 7040 18097 7104
rect 18161 7040 18177 7104
rect 18241 7040 18257 7104
rect 18321 7040 18337 7104
rect 18401 7040 18409 7104
rect 18089 6016 18409 7040
rect 18089 5952 18097 6016
rect 18161 5952 18177 6016
rect 18241 5952 18257 6016
rect 18321 5952 18337 6016
rect 18401 5952 18409 6016
rect 18089 4928 18409 5952
rect 18089 4864 18097 4928
rect 18161 4864 18177 4928
rect 18241 4864 18257 4928
rect 18321 4864 18337 4928
rect 18401 4864 18409 4928
rect 18089 3840 18409 4864
rect 18089 3776 18097 3840
rect 18161 3776 18177 3840
rect 18241 3776 18257 3840
rect 18321 3776 18337 3840
rect 18401 3776 18409 3840
rect 18089 2752 18409 3776
rect 18089 2688 18097 2752
rect 18161 2688 18177 2752
rect 18241 2688 18257 2752
rect 18321 2688 18337 2752
rect 18401 2688 18409 2752
rect 18089 1664 18409 2688
rect 18089 1600 18097 1664
rect 18161 1600 18177 1664
rect 18241 1600 18257 1664
rect 18321 1600 18337 1664
rect 18401 1600 18409 1664
rect 18089 1040 18409 1600
rect 23804 8736 24124 8752
rect 23804 8672 23812 8736
rect 23876 8672 23892 8736
rect 23956 8672 23972 8736
rect 24036 8672 24052 8736
rect 24116 8672 24124 8736
rect 23804 7648 24124 8672
rect 23804 7584 23812 7648
rect 23876 7584 23892 7648
rect 23956 7584 23972 7648
rect 24036 7584 24052 7648
rect 24116 7584 24124 7648
rect 23804 6560 24124 7584
rect 23804 6496 23812 6560
rect 23876 6496 23892 6560
rect 23956 6496 23972 6560
rect 24036 6496 24052 6560
rect 24116 6496 24124 6560
rect 23804 5472 24124 6496
rect 23804 5408 23812 5472
rect 23876 5408 23892 5472
rect 23956 5408 23972 5472
rect 24036 5408 24052 5472
rect 24116 5408 24124 5472
rect 23804 4384 24124 5408
rect 23804 4320 23812 4384
rect 23876 4320 23892 4384
rect 23956 4320 23972 4384
rect 24036 4320 24052 4384
rect 24116 4320 24124 4384
rect 23804 3296 24124 4320
rect 23804 3232 23812 3296
rect 23876 3232 23892 3296
rect 23956 3232 23972 3296
rect 24036 3232 24052 3296
rect 24116 3232 24124 3296
rect 23804 2208 24124 3232
rect 23804 2144 23812 2208
rect 23876 2144 23892 2208
rect 23956 2144 23972 2208
rect 24036 2144 24052 2208
rect 24116 2144 24124 2208
rect 23804 1120 24124 2144
rect 23804 1056 23812 1120
rect 23876 1056 23892 1120
rect 23956 1056 23972 1120
rect 24036 1056 24052 1120
rect 24116 1056 24124 1120
rect 23804 1040 24124 1056
rect 29519 8192 29839 8752
rect 29519 8128 29527 8192
rect 29591 8128 29607 8192
rect 29671 8128 29687 8192
rect 29751 8128 29767 8192
rect 29831 8128 29839 8192
rect 29519 7104 29839 8128
rect 29519 7040 29527 7104
rect 29591 7040 29607 7104
rect 29671 7040 29687 7104
rect 29751 7040 29767 7104
rect 29831 7040 29839 7104
rect 29519 6016 29839 7040
rect 29519 5952 29527 6016
rect 29591 5952 29607 6016
rect 29671 5952 29687 6016
rect 29751 5952 29767 6016
rect 29831 5952 29839 6016
rect 29519 4928 29839 5952
rect 29519 4864 29527 4928
rect 29591 4864 29607 4928
rect 29671 4864 29687 4928
rect 29751 4864 29767 4928
rect 29831 4864 29839 4928
rect 29519 3840 29839 4864
rect 29519 3776 29527 3840
rect 29591 3776 29607 3840
rect 29671 3776 29687 3840
rect 29751 3776 29767 3840
rect 29831 3776 29839 3840
rect 29519 2752 29839 3776
rect 35234 8736 35554 8752
rect 35234 8672 35242 8736
rect 35306 8672 35322 8736
rect 35386 8672 35402 8736
rect 35466 8672 35482 8736
rect 35546 8672 35554 8736
rect 35234 7648 35554 8672
rect 35234 7584 35242 7648
rect 35306 7584 35322 7648
rect 35386 7584 35402 7648
rect 35466 7584 35482 7648
rect 35546 7584 35554 7648
rect 35234 6560 35554 7584
rect 35234 6496 35242 6560
rect 35306 6496 35322 6560
rect 35386 6496 35402 6560
rect 35466 6496 35482 6560
rect 35546 6496 35554 6560
rect 35234 5472 35554 6496
rect 35234 5408 35242 5472
rect 35306 5408 35322 5472
rect 35386 5408 35402 5472
rect 35466 5408 35482 5472
rect 35546 5408 35554 5472
rect 35234 4384 35554 5408
rect 35234 4320 35242 4384
rect 35306 4320 35322 4384
rect 35386 4320 35402 4384
rect 35466 4320 35482 4384
rect 35546 4320 35554 4384
rect 35234 3296 35554 4320
rect 35234 3232 35242 3296
rect 35306 3232 35322 3296
rect 35386 3232 35402 3296
rect 35466 3232 35482 3296
rect 35546 3232 35554 3296
rect 30235 2956 30301 2957
rect 30235 2892 30236 2956
rect 30300 2892 30301 2956
rect 30235 2891 30301 2892
rect 29519 2688 29527 2752
rect 29591 2688 29607 2752
rect 29671 2688 29687 2752
rect 29751 2688 29767 2752
rect 29831 2688 29839 2752
rect 29519 1664 29839 2688
rect 29519 1600 29527 1664
rect 29591 1600 29607 1664
rect 29671 1600 29687 1664
rect 29751 1600 29767 1664
rect 29831 1600 29839 1664
rect 29519 1040 29839 1600
rect 30238 1325 30298 2891
rect 30419 2276 30485 2277
rect 30419 2212 30420 2276
rect 30484 2212 30485 2276
rect 30419 2211 30485 2212
rect 30235 1324 30301 1325
rect 30235 1260 30236 1324
rect 30300 1260 30301 1324
rect 30235 1259 30301 1260
rect 30422 237 30482 2211
rect 35234 2208 35554 3232
rect 35234 2144 35242 2208
rect 35306 2144 35322 2208
rect 35386 2144 35402 2208
rect 35466 2144 35482 2208
rect 35546 2144 35554 2208
rect 35234 1120 35554 2144
rect 35234 1056 35242 1120
rect 35306 1056 35322 1120
rect 35386 1056 35402 1120
rect 35466 1056 35482 1120
rect 35546 1056 35554 1120
rect 35234 1040 35554 1056
rect 40949 8192 41269 8752
rect 40949 8128 40957 8192
rect 41021 8128 41037 8192
rect 41101 8128 41117 8192
rect 41181 8128 41197 8192
rect 41261 8128 41269 8192
rect 40949 7104 41269 8128
rect 40949 7040 40957 7104
rect 41021 7040 41037 7104
rect 41101 7040 41117 7104
rect 41181 7040 41197 7104
rect 41261 7040 41269 7104
rect 40949 6016 41269 7040
rect 40949 5952 40957 6016
rect 41021 5952 41037 6016
rect 41101 5952 41117 6016
rect 41181 5952 41197 6016
rect 41261 5952 41269 6016
rect 40949 4928 41269 5952
rect 40949 4864 40957 4928
rect 41021 4864 41037 4928
rect 41101 4864 41117 4928
rect 41181 4864 41197 4928
rect 41261 4864 41269 4928
rect 40949 3840 41269 4864
rect 40949 3776 40957 3840
rect 41021 3776 41037 3840
rect 41101 3776 41117 3840
rect 41181 3776 41197 3840
rect 41261 3776 41269 3840
rect 40949 2752 41269 3776
rect 40949 2688 40957 2752
rect 41021 2688 41037 2752
rect 41101 2688 41117 2752
rect 41181 2688 41197 2752
rect 41261 2688 41269 2752
rect 40949 1664 41269 2688
rect 40949 1600 40957 1664
rect 41021 1600 41037 1664
rect 41101 1600 41117 1664
rect 41181 1600 41197 1664
rect 41261 1600 41269 1664
rect 40949 1040 41269 1600
rect 46664 8736 46984 8752
rect 46664 8672 46672 8736
rect 46736 8672 46752 8736
rect 46816 8672 46832 8736
rect 46896 8672 46912 8736
rect 46976 8672 46984 8736
rect 46664 7648 46984 8672
rect 46664 7584 46672 7648
rect 46736 7584 46752 7648
rect 46816 7584 46832 7648
rect 46896 7584 46912 7648
rect 46976 7584 46984 7648
rect 46664 6560 46984 7584
rect 46664 6496 46672 6560
rect 46736 6496 46752 6560
rect 46816 6496 46832 6560
rect 46896 6496 46912 6560
rect 46976 6496 46984 6560
rect 46664 5472 46984 6496
rect 46664 5408 46672 5472
rect 46736 5408 46752 5472
rect 46816 5408 46832 5472
rect 46896 5408 46912 5472
rect 46976 5408 46984 5472
rect 46664 4384 46984 5408
rect 46664 4320 46672 4384
rect 46736 4320 46752 4384
rect 46816 4320 46832 4384
rect 46896 4320 46912 4384
rect 46976 4320 46984 4384
rect 46664 3296 46984 4320
rect 46664 3232 46672 3296
rect 46736 3232 46752 3296
rect 46816 3232 46832 3296
rect 46896 3232 46912 3296
rect 46976 3232 46984 3296
rect 46664 2208 46984 3232
rect 46664 2144 46672 2208
rect 46736 2144 46752 2208
rect 46816 2144 46832 2208
rect 46896 2144 46912 2208
rect 46976 2144 46984 2208
rect 46664 1120 46984 2144
rect 46664 1056 46672 1120
rect 46736 1056 46752 1120
rect 46816 1056 46832 1120
rect 46896 1056 46912 1120
rect 46976 1056 46984 1120
rect 46664 1040 46984 1056
rect 30419 236 30485 237
rect 30419 172 30420 236
rect 30484 172 30485 236
rect 30419 171 30485 172
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37444 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_8 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1840 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_12
timestamp 1688980957
transform 1 0 2208 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_16
timestamp 1688980957
transform 1 0 2576 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_20
timestamp 1688980957
transform 1 0 2944 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_39
timestamp 1688980957
transform 1 0 4692 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_44
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_48
timestamp 1688980957
transform 1 0 5520 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_52
timestamp 1688980957
transform 1 0 5888 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_60
timestamp 1688980957
transform 1 0 6624 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_64
timestamp 1688980957
transform 1 0 6992 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_68
timestamp 1688980957
transform 1 0 7360 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_72
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_76
timestamp 1688980957
transform 1 0 8096 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_80
timestamp 1688980957
transform 1 0 8464 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_88
timestamp 1688980957
transform 1 0 9200 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_92
timestamp 1688980957
transform 1 0 9568 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_96
timestamp 1688980957
transform 1 0 9936 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_100
timestamp 1688980957
transform 1 0 10304 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_104
timestamp 1688980957
transform 1 0 10672 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_108
timestamp 1688980957
transform 1 0 11040 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_116
timestamp 1688980957
transform 1 0 11776 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_120
timestamp 1688980957
transform 1 0 12144 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_124
timestamp 1688980957
transform 1 0 12512 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_128
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_132
timestamp 1688980957
transform 1 0 13248 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_136
timestamp 1688980957
transform 1 0 13616 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_144
timestamp 1688980957
transform 1 0 14352 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_148
timestamp 1688980957
transform 1 0 14720 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_152
timestamp 1688980957
transform 1 0 15088 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_203
timestamp 1688980957
transform 1 0 19780 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_214
timestamp 1688980957
transform 1 0 20792 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_234
timestamp 1688980957
transform 1 0 22632 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_246
timestamp 1688980957
transform 1 0 23736 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_271
timestamp 1688980957
transform 1 0 26036 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_299
timestamp 1688980957
transform 1 0 28612 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_315
timestamp 1688980957
transform 1 0 30084 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1688980957
transform 1 0 31924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34316 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_397
timestamp 1688980957
transform 1 0 37628 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_436
timestamp 1688980957
transform 1 0 41216 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_464
timestamp 1688980957
transform 1 0 43792 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_468
timestamp 1688980957
transform 1 0 44160 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_472
timestamp 1688980957
transform 1 0 44528 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_480
timestamp 1688980957
transform 1 0 45264 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_484
timestamp 1688980957
transform 1 0 45632 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_488
timestamp 1688980957
transform 1 0 46000 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_492
timestamp 1688980957
transform 1 0 46368 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_18
timestamp 1688980957
transform 1 0 2760 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_30
timestamp 1688980957
transform 1 0 3864 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_36
timestamp 1688980957
transform 1 0 4416 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_40
timestamp 1688980957
transform 1 0 4784 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_52 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5888 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_149 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_157
timestamp 1688980957
transform 1 0 15548 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_216
timestamp 1688980957
transform 1 0 20976 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_236
timestamp 1688980957
transform 1 0 22816 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_248
timestamp 1688980957
transform 1 0 23920 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_258
timestamp 1688980957
transform 1 0 24840 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_268
timestamp 1688980957
transform 1 0 25760 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_296
timestamp 1688980957
transform 1 0 28336 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_301
timestamp 1688980957
transform 1 0 28796 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_312
timestamp 1688980957
transform 1 0 29808 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_323
timestamp 1688980957
transform 1 0 30820 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_343
timestamp 1688980957
transform 1 0 32660 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_352
timestamp 1688980957
transform 1 0 33488 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_366
timestamp 1688980957
transform 1 0 34776 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_372
timestamp 1688980957
transform 1 0 35328 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_377
timestamp 1688980957
transform 1 0 35788 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_387
timestamp 1688980957
transform 1 0 36708 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_399
timestamp 1688980957
transform 1 0 37812 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_407
timestamp 1688980957
transform 1 0 38548 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_415
timestamp 1688980957
transform 1 0 39284 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_427
timestamp 1688980957
transform 1 0 40388 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_440
timestamp 1688980957
transform 1 0 41584 0 -1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_452
timestamp 1688980957
transform 1 0 42688 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_464
timestamp 1688980957
transform 1 0 43792 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_476
timestamp 1688980957
transform 1 0 44896 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_487
timestamp 1688980957
transform 1 0 45908 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_184
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_202
timestamp 1688980957
transform 1 0 19688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_216
timestamp 1688980957
transform 1 0 20976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_220
timestamp 1688980957
transform 1 0 21344 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_224
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_231
timestamp 1688980957
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_243
timestamp 1688980957
transform 1 0 23460 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 1688980957
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_271
timestamp 1688980957
transform 1 0 26036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_275
timestamp 1688980957
transform 1 0 26404 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_279
timestamp 1688980957
transform 1 0 26772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_286
timestamp 1688980957
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_299
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_303
timestamp 1688980957
transform 1 0 28980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_318
timestamp 1688980957
transform 1 0 30360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_331
timestamp 1688980957
transform 1 0 31556 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_340
timestamp 1688980957
transform 1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_346
timestamp 1688980957
transform 1 0 32936 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_351
timestamp 1688980957
transform 1 0 33396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_371
timestamp 1688980957
transform 1 0 35236 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_375
timestamp 1688980957
transform 1 0 35604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_387
timestamp 1688980957
transform 1 0 36708 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_395
timestamp 1688980957
transform 1 0 37444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_402
timestamp 1688980957
transform 1 0 38088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_409
timestamp 1688980957
transform 1 0 38732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_417
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_448
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_460
timestamp 1688980957
transform 1 0 43424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 1688980957
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_480
timestamp 1688980957
transform 1 0 45264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_487
timestamp 1688980957
transform 1 0 45908 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_493
timestamp 1688980957
transform 1 0 46460 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_473
timestamp 1688980957
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_485
timestamp 1688980957
transform 1 0 45724 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_493
timestamp 1688980957
transform 1 0 46460 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1688980957
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_477
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_489
timestamp 1688980957
transform 1 0 46092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_493
timestamp 1688980957
transform 1 0 46460 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_473
timestamp 1688980957
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_485
timestamp 1688980957
transform 1 0 45724 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_493
timestamp 1688980957
transform 1 0 46460 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_469
timestamp 1688980957
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 1688980957
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_489
timestamp 1688980957
transform 1 0 46092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_493
timestamp 1688980957
transform 1 0 46460 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_473
timestamp 1688980957
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_485
timestamp 1688980957
transform 1 0 45724 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_493
timestamp 1688980957
transform 1 0 46460 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 1688980957
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_477
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_489
timestamp 1688980957
transform 1 0 46092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_493
timestamp 1688980957
transform 1 0 46460 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_473
timestamp 1688980957
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_485
timestamp 1688980957
transform 1 0 45724 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_493
timestamp 1688980957
transform 1 0 46460 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_469
timestamp 1688980957
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 1688980957
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_477
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_489
timestamp 1688980957
transform 1 0 46092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_493
timestamp 1688980957
transform 1 0 46460 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_461
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_473
timestamp 1688980957
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_485
timestamp 1688980957
transform 1 0 45724 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_493
timestamp 1688980957
transform 1 0 46460 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_469
timestamp 1688980957
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 1688980957
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_477
timestamp 1688980957
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_489
timestamp 1688980957
transform 1 0 46092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_493
timestamp 1688980957
transform 1 0 46460 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_13
timestamp 1688980957
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_25
timestamp 1688980957
transform 1 0 3404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_37
timestamp 1688980957
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_49
timestamp 1688980957
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_61
timestamp 1688980957
transform 1 0 6716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_73
timestamp 1688980957
transform 1 0 7820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_89
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_101
timestamp 1688980957
transform 1 0 10396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 1688980957
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_133
timestamp 1688980957
transform 1 0 13340 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_139
timestamp 1688980957
transform 1 0 13892 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_157
timestamp 1688980957
transform 1 0 15548 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 1688980957
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_197
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_229
timestamp 1688980957
transform 1 0 22172 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_241
timestamp 1688980957
transform 1 0 23276 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_257
timestamp 1688980957
transform 1 0 24748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_269
timestamp 1688980957
transform 1 0 25852 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_277
timestamp 1688980957
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_301
timestamp 1688980957
transform 1 0 28796 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_307
timestamp 1688980957
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_309
timestamp 1688980957
transform 1 0 29532 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_325
timestamp 1688980957
transform 1 0 31004 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_333
timestamp 1688980957
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_365
timestamp 1688980957
transform 1 0 34684 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 1688980957
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 1688980957
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_399
timestamp 1688980957
transform 1 0 37812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_411
timestamp 1688980957
transform 1 0 38916 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_419
timestamp 1688980957
transform 1 0 39652 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_425
timestamp 1688980957
transform 1 0 40204 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_437
timestamp 1688980957
transform 1 0 41308 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_445
timestamp 1688980957
transform 1 0 42044 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_461
timestamp 1688980957
transform 1 0 43516 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_469
timestamp 1688980957
transform 1 0 44252 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_475
timestamp 1688980957
transform 1 0 44804 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_477
timestamp 1688980957
transform 1 0 44988 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_493
timestamp 1688980957
transform 1 0 46460 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40940 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 43516 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 43884 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 44252 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 44620 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44988 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 45356 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 45724 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 46092 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 46276 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 46000 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 40480 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 40756 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 41032 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 41308 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 42412 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 41400 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 42688 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 42964 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 43240 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 1564 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 1932 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 2300 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 5612 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 6716 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 7084 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1688980957
transform 1 0 7820 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 8188 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 2668 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 3128 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 3404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 4140 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 4508 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 5244 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 12236 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 12604 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 12972 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 13340 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 9292 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1688980957
transform 1 0 9660 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform 1 0 10028 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1688980957
transform 1 0 10396 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 10764 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1688980957
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1688980957
transform 1 0 11868 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 14444 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform 1 0 17480 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform 1 0 18032 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform 1 0 18584 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform 1 0 14812 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform 1 0 15456 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1688980957
transform 1 0 16008 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1688980957
transform 1 0 16928 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1688980957
transform 1 0 39468 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28888 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__00_
timestamp 1688980957
transform 1 0 23000 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__01_
timestamp 1688980957
transform 1 0 24012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__02_
timestamp 1688980957
transform 1 0 24564 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__03_
timestamp 1688980957
transform 1 0 24932 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__04_
timestamp 1688980957
transform 1 0 26220 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__05_
timestamp 1688980957
transform 1 0 25760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__06_
timestamp 1688980957
transform 1 0 27232 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__07_
timestamp 1688980957
transform 1 0 27508 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__08_
timestamp 1688980957
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__09_
timestamp 1688980957
transform 1 0 20056 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__10_
timestamp 1688980957
transform 1 0 21160 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__11_
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__12_
timestamp 1688980957
transform 1 0 21436 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__13_
timestamp 1688980957
transform 1 0 21896 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__14_
timestamp 1688980957
transform 1 0 22172 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__15_
timestamp 1688980957
transform 1 0 23184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__16_
timestamp 1688980957
transform 1 0 27784 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__17_
timestamp 1688980957
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__18_
timestamp 1688980957
transform 1 0 30452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__19_
timestamp 1688980957
transform 1 0 32108 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__20_
timestamp 1688980957
transform 1 0 32384 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__21_
timestamp 1688980957
transform 1 0 33212 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__22_
timestamp 1688980957
transform 1 0 32660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__23_
timestamp 1688980957
transform 1 0 28060 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__24_
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__25_
timestamp 1688980957
transform 1 0 28336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__26_
timestamp 1688980957
transform 1 0 29256 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__27_
timestamp 1688980957
transform 1 0 29532 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__28_
timestamp 1688980957
transform 1 0 30268 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__29_
timestamp 1688980957
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__30_
timestamp 1688980957
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__31_
timestamp 1688980957
transform 1 0 31280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__32_
timestamp 1688980957
transform 1 0 19504 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__33_
timestamp 1688980957
transform 1 0 19504 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__34_
timestamp 1688980957
transform 1 0 16284 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__35_
timestamp 1688980957
transform 1 0 16008 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__36_
timestamp 1688980957
transform 1 0 15732 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__37_
timestamp 1688980957
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__38_
timestamp 1688980957
transform 1 0 20332 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__39_
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__40_
timestamp 1688980957
transform 1 0 18676 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__41_
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__42_
timestamp 1688980957
transform 1 0 18400 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__43_
timestamp 1688980957
transform 1 0 18124 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__44_
timestamp 1688980957
transform 1 0 17848 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__45_
timestamp 1688980957
transform 1 0 17296 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__46_
timestamp 1688980957
transform 1 0 17020 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__47_
timestamp 1688980957
transform 1 0 16744 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__48_
timestamp 1688980957
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__49_
timestamp 1688980957
transform 1 0 18952 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__50_
timestamp 1688980957
transform 1 0 20148 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__51_
timestamp 1688980957
transform 1 0 19780 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 26036 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output76 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1688980957
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1688980957
transform 1 0 32844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1688980957
transform 1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1688980957
transform 1 0 39836 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1688980957
transform 1 0 41676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1688980957
transform 1 0 43884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1688980957
transform 1 0 46092 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1688980957
transform 1 0 12972 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 14996 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1688980957
transform 1 0 17388 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1688980957
transform 1 0 19596 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1688980957
transform 1 0 19872 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 20240 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform 1 0 20608 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1688980957
transform 1 0 20976 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 24748 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1688980957
transform 1 0 25300 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1688980957
transform 1 0 25668 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform 1 0 25852 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 26220 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1688980957
transform 1 0 26956 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1688980957
transform 1 0 27324 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 27692 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1688980957
transform 1 0 21344 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 22080 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1688980957
transform 1 0 22448 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1688980957
transform 1 0 22816 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 23184 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1688980957
transform 1 0 23552 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1688980957
transform 1 0 23920 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1688980957
transform 1 0 28244 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 32108 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 32660 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1688980957
transform 1 0 32844 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 33212 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform 1 0 33764 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1688980957
transform 1 0 34132 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1688980957
transform 1 0 28428 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform 1 0 28796 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 29532 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1688980957
transform 1 0 29900 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 30268 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 30820 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform 1 0 31372 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1688980957
transform 1 0 31556 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 31004 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 33580 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 37996 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1688980957
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output133
timestamp 1688980957
transform 1 0 38916 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output134
timestamp 1688980957
transform 1 0 39836 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 38732 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 40388 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 34684 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform 1 0 35236 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1688980957
transform 1 0 35420 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 35788 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 36340 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 37260 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 36156 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 37812 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 38364 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 46828 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 46828 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 46828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 46828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 46828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 46828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 46828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 46828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 46828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 46828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 46828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 46828 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 46828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 46828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 26956 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform 1 0 24288 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform 1 0 25208 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform 1 0 26496 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform 1 0 23276 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 17572 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform 1 0 19228 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 25484 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 30544 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 34500 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 35880 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 45080 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 42412 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 45356 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 45632 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 23552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 19872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 22080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 26496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 28704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 31004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 33120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 35328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 44528 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 45632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 44896 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 37168 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 44896 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 39762 0 39818 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 43442 0 43498 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 43810 0 43866 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 44178 0 44234 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 44546 0 44602 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 44914 0 44970 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 45282 0 45338 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 45650 0 45706 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 46018 0 46074 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 46386 0 46442 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 46754 0 46810 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 40130 0 40186 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 40498 0 40554 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 40866 0 40922 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 41234 0 41290 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 41602 0 41658 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 41970 0 42026 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 42338 0 42394 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 42706 0 42762 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 43074 0 43130 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 4066 9840 4122 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 26146 9840 26202 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 28354 9840 28410 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 30562 9840 30618 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 32770 9840 32826 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 34978 9840 35034 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 37186 9840 37242 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 39394 9840 39450 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 41602 9840 41658 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 43810 9840 43866 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 46018 9840 46074 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 6274 9840 6330 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 8482 9840 8538 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 10690 9840 10746 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 12898 9840 12954 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 15106 9840 15162 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 17314 9840 17370 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 19522 9840 19578 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 21730 9840 21786 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 23938 9840 23994 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 1122 0 1178 160 0 FreeSans 224 90 0 0 N1END[0]
port 40 nsew signal input
flabel metal2 s 1490 0 1546 160 0 FreeSans 224 90 0 0 N1END[1]
port 41 nsew signal input
flabel metal2 s 1858 0 1914 160 0 FreeSans 224 90 0 0 N1END[2]
port 42 nsew signal input
flabel metal2 s 2226 0 2282 160 0 FreeSans 224 90 0 0 N1END[3]
port 43 nsew signal input
flabel metal2 s 5538 0 5594 160 0 FreeSans 224 90 0 0 N2END[0]
port 44 nsew signal input
flabel metal2 s 5906 0 5962 160 0 FreeSans 224 90 0 0 N2END[1]
port 45 nsew signal input
flabel metal2 s 6274 0 6330 160 0 FreeSans 224 90 0 0 N2END[2]
port 46 nsew signal input
flabel metal2 s 6642 0 6698 160 0 FreeSans 224 90 0 0 N2END[3]
port 47 nsew signal input
flabel metal2 s 7010 0 7066 160 0 FreeSans 224 90 0 0 N2END[4]
port 48 nsew signal input
flabel metal2 s 7378 0 7434 160 0 FreeSans 224 90 0 0 N2END[5]
port 49 nsew signal input
flabel metal2 s 7746 0 7802 160 0 FreeSans 224 90 0 0 N2END[6]
port 50 nsew signal input
flabel metal2 s 8114 0 8170 160 0 FreeSans 224 90 0 0 N2END[7]
port 51 nsew signal input
flabel metal2 s 2594 0 2650 160 0 FreeSans 224 90 0 0 N2MID[0]
port 52 nsew signal input
flabel metal2 s 2962 0 3018 160 0 FreeSans 224 90 0 0 N2MID[1]
port 53 nsew signal input
flabel metal2 s 3330 0 3386 160 0 FreeSans 224 90 0 0 N2MID[2]
port 54 nsew signal input
flabel metal2 s 3698 0 3754 160 0 FreeSans 224 90 0 0 N2MID[3]
port 55 nsew signal input
flabel metal2 s 4066 0 4122 160 0 FreeSans 224 90 0 0 N2MID[4]
port 56 nsew signal input
flabel metal2 s 4434 0 4490 160 0 FreeSans 224 90 0 0 N2MID[5]
port 57 nsew signal input
flabel metal2 s 4802 0 4858 160 0 FreeSans 224 90 0 0 N2MID[6]
port 58 nsew signal input
flabel metal2 s 5170 0 5226 160 0 FreeSans 224 90 0 0 N2MID[7]
port 59 nsew signal input
flabel metal2 s 8482 0 8538 160 0 FreeSans 224 90 0 0 N4END[0]
port 60 nsew signal input
flabel metal2 s 12162 0 12218 160 0 FreeSans 224 90 0 0 N4END[10]
port 61 nsew signal input
flabel metal2 s 12530 0 12586 160 0 FreeSans 224 90 0 0 N4END[11]
port 62 nsew signal input
flabel metal2 s 12898 0 12954 160 0 FreeSans 224 90 0 0 N4END[12]
port 63 nsew signal input
flabel metal2 s 13266 0 13322 160 0 FreeSans 224 90 0 0 N4END[13]
port 64 nsew signal input
flabel metal2 s 13634 0 13690 160 0 FreeSans 224 90 0 0 N4END[14]
port 65 nsew signal input
flabel metal2 s 14002 0 14058 160 0 FreeSans 224 90 0 0 N4END[15]
port 66 nsew signal input
flabel metal2 s 8850 0 8906 160 0 FreeSans 224 90 0 0 N4END[1]
port 67 nsew signal input
flabel metal2 s 9218 0 9274 160 0 FreeSans 224 90 0 0 N4END[2]
port 68 nsew signal input
flabel metal2 s 9586 0 9642 160 0 FreeSans 224 90 0 0 N4END[3]
port 69 nsew signal input
flabel metal2 s 9954 0 10010 160 0 FreeSans 224 90 0 0 N4END[4]
port 70 nsew signal input
flabel metal2 s 10322 0 10378 160 0 FreeSans 224 90 0 0 N4END[5]
port 71 nsew signal input
flabel metal2 s 10690 0 10746 160 0 FreeSans 224 90 0 0 N4END[6]
port 72 nsew signal input
flabel metal2 s 11058 0 11114 160 0 FreeSans 224 90 0 0 N4END[7]
port 73 nsew signal input
flabel metal2 s 11426 0 11482 160 0 FreeSans 224 90 0 0 N4END[8]
port 74 nsew signal input
flabel metal2 s 11794 0 11850 160 0 FreeSans 224 90 0 0 N4END[9]
port 75 nsew signal input
flabel metal2 s 14370 0 14426 160 0 FreeSans 224 90 0 0 NN4END[0]
port 76 nsew signal input
flabel metal2 s 18050 0 18106 160 0 FreeSans 224 90 0 0 NN4END[10]
port 77 nsew signal input
flabel metal2 s 18418 0 18474 160 0 FreeSans 224 90 0 0 NN4END[11]
port 78 nsew signal input
flabel metal2 s 18786 0 18842 160 0 FreeSans 224 90 0 0 NN4END[12]
port 79 nsew signal input
flabel metal2 s 19154 0 19210 160 0 FreeSans 224 90 0 0 NN4END[13]
port 80 nsew signal input
flabel metal2 s 19522 0 19578 160 0 FreeSans 224 90 0 0 NN4END[14]
port 81 nsew signal input
flabel metal2 s 19890 0 19946 160 0 FreeSans 224 90 0 0 NN4END[15]
port 82 nsew signal input
flabel metal2 s 14738 0 14794 160 0 FreeSans 224 90 0 0 NN4END[1]
port 83 nsew signal input
flabel metal2 s 15106 0 15162 160 0 FreeSans 224 90 0 0 NN4END[2]
port 84 nsew signal input
flabel metal2 s 15474 0 15530 160 0 FreeSans 224 90 0 0 NN4END[3]
port 85 nsew signal input
flabel metal2 s 15842 0 15898 160 0 FreeSans 224 90 0 0 NN4END[4]
port 86 nsew signal input
flabel metal2 s 16210 0 16266 160 0 FreeSans 224 90 0 0 NN4END[5]
port 87 nsew signal input
flabel metal2 s 16578 0 16634 160 0 FreeSans 224 90 0 0 NN4END[6]
port 88 nsew signal input
flabel metal2 s 16946 0 17002 160 0 FreeSans 224 90 0 0 NN4END[7]
port 89 nsew signal input
flabel metal2 s 17314 0 17370 160 0 FreeSans 224 90 0 0 NN4END[8]
port 90 nsew signal input
flabel metal2 s 17682 0 17738 160 0 FreeSans 224 90 0 0 NN4END[9]
port 91 nsew signal input
flabel metal2 s 20258 0 20314 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 92 nsew signal tristate
flabel metal2 s 20626 0 20682 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 93 nsew signal tristate
flabel metal2 s 20994 0 21050 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 94 nsew signal tristate
flabel metal2 s 21362 0 21418 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 95 nsew signal tristate
flabel metal2 s 24674 0 24730 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 96 nsew signal tristate
flabel metal2 s 25042 0 25098 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 97 nsew signal tristate
flabel metal2 s 25410 0 25466 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 98 nsew signal tristate
flabel metal2 s 25778 0 25834 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 99 nsew signal tristate
flabel metal2 s 26146 0 26202 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 100 nsew signal tristate
flabel metal2 s 26514 0 26570 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 101 nsew signal tristate
flabel metal2 s 26882 0 26938 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 102 nsew signal tristate
flabel metal2 s 27250 0 27306 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 103 nsew signal tristate
flabel metal2 s 21730 0 21786 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 104 nsew signal tristate
flabel metal2 s 22098 0 22154 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 105 nsew signal tristate
flabel metal2 s 22466 0 22522 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 106 nsew signal tristate
flabel metal2 s 22834 0 22890 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 107 nsew signal tristate
flabel metal2 s 23202 0 23258 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 108 nsew signal tristate
flabel metal2 s 23570 0 23626 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 109 nsew signal tristate
flabel metal2 s 23938 0 23994 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 110 nsew signal tristate
flabel metal2 s 24306 0 24362 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 111 nsew signal tristate
flabel metal2 s 27618 0 27674 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 112 nsew signal tristate
flabel metal2 s 31298 0 31354 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 113 nsew signal tristate
flabel metal2 s 31666 0 31722 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 114 nsew signal tristate
flabel metal2 s 32034 0 32090 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 115 nsew signal tristate
flabel metal2 s 32402 0 32458 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 116 nsew signal tristate
flabel metal2 s 32770 0 32826 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 117 nsew signal tristate
flabel metal2 s 33138 0 33194 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 118 nsew signal tristate
flabel metal2 s 27986 0 28042 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 119 nsew signal tristate
flabel metal2 s 28354 0 28410 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 120 nsew signal tristate
flabel metal2 s 28722 0 28778 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 121 nsew signal tristate
flabel metal2 s 29090 0 29146 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 122 nsew signal tristate
flabel metal2 s 29458 0 29514 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 123 nsew signal tristate
flabel metal2 s 29826 0 29882 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 124 nsew signal tristate
flabel metal2 s 30194 0 30250 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 125 nsew signal tristate
flabel metal2 s 30562 0 30618 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 126 nsew signal tristate
flabel metal2 s 30930 0 30986 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 127 nsew signal tristate
flabel metal2 s 33506 0 33562 160 0 FreeSans 224 90 0 0 SS4BEG[0]
port 128 nsew signal tristate
flabel metal2 s 37186 0 37242 160 0 FreeSans 224 90 0 0 SS4BEG[10]
port 129 nsew signal tristate
flabel metal2 s 37554 0 37610 160 0 FreeSans 224 90 0 0 SS4BEG[11]
port 130 nsew signal tristate
flabel metal2 s 37922 0 37978 160 0 FreeSans 224 90 0 0 SS4BEG[12]
port 131 nsew signal tristate
flabel metal2 s 38290 0 38346 160 0 FreeSans 224 90 0 0 SS4BEG[13]
port 132 nsew signal tristate
flabel metal2 s 38658 0 38714 160 0 FreeSans 224 90 0 0 SS4BEG[14]
port 133 nsew signal tristate
flabel metal2 s 39026 0 39082 160 0 FreeSans 224 90 0 0 SS4BEG[15]
port 134 nsew signal tristate
flabel metal2 s 33874 0 33930 160 0 FreeSans 224 90 0 0 SS4BEG[1]
port 135 nsew signal tristate
flabel metal2 s 34242 0 34298 160 0 FreeSans 224 90 0 0 SS4BEG[2]
port 136 nsew signal tristate
flabel metal2 s 34610 0 34666 160 0 FreeSans 224 90 0 0 SS4BEG[3]
port 137 nsew signal tristate
flabel metal2 s 34978 0 35034 160 0 FreeSans 224 90 0 0 SS4BEG[4]
port 138 nsew signal tristate
flabel metal2 s 35346 0 35402 160 0 FreeSans 224 90 0 0 SS4BEG[5]
port 139 nsew signal tristate
flabel metal2 s 35714 0 35770 160 0 FreeSans 224 90 0 0 SS4BEG[6]
port 140 nsew signal tristate
flabel metal2 s 36082 0 36138 160 0 FreeSans 224 90 0 0 SS4BEG[7]
port 141 nsew signal tristate
flabel metal2 s 36450 0 36506 160 0 FreeSans 224 90 0 0 SS4BEG[8]
port 142 nsew signal tristate
flabel metal2 s 36818 0 36874 160 0 FreeSans 224 90 0 0 SS4BEG[9]
port 143 nsew signal tristate
flabel metal2 s 39394 0 39450 160 0 FreeSans 224 90 0 0 UserCLK
port 144 nsew signal input
flabel metal2 s 1858 9840 1914 10000 0 FreeSans 224 90 0 0 UserCLKo
port 145 nsew signal tristate
flabel metal4 s 6659 1040 6979 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 18089 1040 18409 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 29519 1040 29839 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 40949 1040 41269 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 12374 1040 12694 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 23804 1040 24124 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 35234 1040 35554 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 46664 1040 46984 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
rlabel metal1 23966 8160 23966 8160 0 vccd1
rlabel via1 24044 8704 24044 8704 0 vssd1
rlabel metal2 39935 68 39935 68 0 FrameStrobe[0]
rlabel metal2 43523 68 43523 68 0 FrameStrobe[10]
rlabel metal2 43891 68 43891 68 0 FrameStrobe[11]
rlabel metal2 44259 68 44259 68 0 FrameStrobe[12]
rlabel metal2 44574 704 44574 704 0 FrameStrobe[13]
rlabel metal2 45087 68 45087 68 0 FrameStrobe[14]
rlabel metal2 45310 143 45310 143 0 FrameStrobe[15]
rlabel metal2 45823 68 45823 68 0 FrameStrobe[16]
rlabel metal2 46191 68 46191 68 0 FrameStrobe[17]
rlabel metal2 46467 68 46467 68 0 FrameStrobe[18]
rlabel metal2 46683 68 46683 68 0 FrameStrobe[19]
rlabel metal2 40158 1010 40158 1010 0 FrameStrobe[1]
rlabel metal2 40526 1027 40526 1027 0 FrameStrobe[2]
rlabel metal2 40894 959 40894 959 0 FrameStrobe[3]
rlabel metal2 41315 68 41315 68 0 FrameStrobe[4]
rlabel metal2 41775 68 41775 68 0 FrameStrobe[5]
rlabel metal2 41998 670 41998 670 0 FrameStrobe[6]
rlabel metal2 42366 670 42366 670 0 FrameStrobe[7]
rlabel metal2 42734 636 42734 636 0 FrameStrobe[8]
rlabel metal2 43201 68 43201 68 0 FrameStrobe[9]
rlabel metal2 4094 9224 4094 9224 0 FrameStrobe_O[0]
rlabel metal2 26174 9224 26174 9224 0 FrameStrobe_O[10]
rlabel metal1 28520 8602 28520 8602 0 FrameStrobe_O[11]
rlabel metal1 30728 8602 30728 8602 0 FrameStrobe_O[12]
rlabel metal1 32936 8602 32936 8602 0 FrameStrobe_O[13]
rlabel metal1 35144 8602 35144 8602 0 FrameStrobe_O[14]
rlabel metal2 37214 9224 37214 9224 0 FrameStrobe_O[15]
rlabel metal1 39744 8602 39744 8602 0 FrameStrobe_O[16]
rlabel metal1 41768 8602 41768 8602 0 FrameStrobe_O[17]
rlabel metal1 43976 8602 43976 8602 0 FrameStrobe_O[18]
rlabel metal1 46184 8602 46184 8602 0 FrameStrobe_O[19]
rlabel metal1 6440 8602 6440 8602 0 FrameStrobe_O[1]
rlabel metal1 8832 8602 8832 8602 0 FrameStrobe_O[2]
rlabel metal1 10856 8602 10856 8602 0 FrameStrobe_O[3]
rlabel metal1 13064 8602 13064 8602 0 FrameStrobe_O[4]
rlabel metal2 15134 9224 15134 9224 0 FrameStrobe_O[5]
rlabel metal1 17480 8602 17480 8602 0 FrameStrobe_O[6]
rlabel metal1 19688 8602 19688 8602 0 FrameStrobe_O[7]
rlabel metal1 21896 8602 21896 8602 0 FrameStrobe_O[8]
rlabel metal1 24426 8602 24426 8602 0 FrameStrobe_O[9]
rlabel metal2 27002 2210 27002 2210 0 FrameStrobe_O_i\[0\]
rlabel metal1 26726 2448 26726 2448 0 FrameStrobe_O_i\[10\]
rlabel metal1 30314 2074 30314 2074 0 FrameStrobe_O_i\[11\]
rlabel metal1 31947 2278 31947 2278 0 FrameStrobe_O_i\[12\]
rlabel metal1 33948 2074 33948 2074 0 FrameStrobe_O_i\[13\]
rlabel metal2 35926 2244 35926 2244 0 FrameStrobe_O_i\[14\]
rlabel metal1 37812 2414 37812 2414 0 FrameStrobe_O_i\[15\]
rlabel metal1 44850 2074 44850 2074 0 FrameStrobe_O_i\[16\]
rlabel metal1 42366 2074 42366 2074 0 FrameStrobe_O_i\[17\]
rlabel metal1 45310 2074 45310 2074 0 FrameStrobe_O_i\[18\]
rlabel metal1 45770 2074 45770 2074 0 FrameStrobe_O_i\[19\]
rlabel metal2 24334 2244 24334 2244 0 FrameStrobe_O_i\[1\]
rlabel metal1 24932 1802 24932 1802 0 FrameStrobe_O_i\[2\]
rlabel metal1 26220 2074 26220 2074 0 FrameStrobe_O_i\[3\]
rlabel metal1 23460 2074 23460 2074 0 FrameStrobe_O_i\[4\]
rlabel metal1 21298 2414 21298 2414 0 FrameStrobe_O_i\[5\]
rlabel metal1 17802 2074 17802 2074 0 FrameStrobe_O_i\[6\]
rlabel metal2 19458 2210 19458 2210 0 FrameStrobe_O_i\[7\]
rlabel metal1 22494 2414 22494 2414 0 FrameStrobe_O_i\[8\]
rlabel metal1 25300 2074 25300 2074 0 FrameStrobe_O_i\[9\]
rlabel metal2 1150 1010 1150 1010 0 N1END[0]
rlabel metal2 1571 68 1571 68 0 N1END[1]
rlabel metal2 1939 68 1939 68 0 N1END[2]
rlabel metal2 2307 68 2307 68 0 N1END[3]
rlabel metal2 5619 68 5619 68 0 N2END[0]
rlabel metal2 5987 68 5987 68 0 N2END[1]
rlabel metal2 6355 68 6355 68 0 N2END[2]
rlabel metal2 6723 68 6723 68 0 N2END[3]
rlabel metal2 7091 68 7091 68 0 N2END[4]
rlabel metal2 7459 68 7459 68 0 N2END[5]
rlabel metal2 7827 68 7827 68 0 N2END[6]
rlabel metal2 8195 68 8195 68 0 N2END[7]
rlabel metal2 2675 68 2675 68 0 N2MID[0]
rlabel metal2 2990 670 2990 670 0 N2MID[1]
rlabel metal2 3259 68 3259 68 0 N2MID[2]
rlabel metal2 3581 68 3581 68 0 N2MID[3]
rlabel metal2 4041 68 4041 68 0 N2MID[4]
rlabel metal2 4515 68 4515 68 0 N2MID[5]
rlabel metal2 4883 68 4883 68 0 N2MID[6]
rlabel metal2 5251 68 5251 68 0 N2MID[7]
rlabel metal2 8563 68 8563 68 0 N4END[0]
rlabel metal2 12243 68 12243 68 0 N4END[10]
rlabel metal2 12657 68 12657 68 0 N4END[11]
rlabel metal2 12979 68 12979 68 0 N4END[12]
rlabel metal2 13347 68 13347 68 0 N4END[13]
rlabel metal2 13715 68 13715 68 0 N4END[14]
rlabel metal2 14083 68 14083 68 0 N4END[15]
rlabel metal2 8931 68 8931 68 0 N4END[1]
rlabel metal2 9299 68 9299 68 0 N4END[2]
rlabel metal1 9660 2822 9660 2822 0 N4END[3]
rlabel metal2 10035 68 10035 68 0 N4END[4]
rlabel metal2 10403 68 10403 68 0 N4END[5]
rlabel metal2 10771 68 10771 68 0 N4END[6]
rlabel metal2 11139 68 11139 68 0 N4END[7]
rlabel metal2 11507 68 11507 68 0 N4END[8]
rlabel metal2 11875 68 11875 68 0 N4END[9]
rlabel metal2 14543 68 14543 68 0 NN4END[0]
rlabel metal2 17933 68 17933 68 0 NN4END[10]
rlabel metal2 18446 670 18446 670 0 NN4END[11]
rlabel metal2 18814 296 18814 296 0 NN4END[12]
rlabel metal2 19182 432 19182 432 0 NN4END[13]
rlabel metal2 19550 415 19550 415 0 NN4END[14]
rlabel metal2 19918 670 19918 670 0 NN4END[15]
rlabel metal2 14911 68 14911 68 0 NN4END[1]
rlabel metal2 15279 68 15279 68 0 NN4END[2]
rlabel metal2 15601 68 15601 68 0 NN4END[3]
rlabel metal2 15923 68 15923 68 0 NN4END[4]
rlabel metal2 16238 704 16238 704 0 NN4END[5]
rlabel metal2 16606 704 16606 704 0 NN4END[6]
rlabel metal2 16921 68 16921 68 0 NN4END[7]
rlabel metal2 17342 704 17342 704 0 NN4END[8]
rlabel metal2 17710 143 17710 143 0 NN4END[9]
rlabel metal2 20286 636 20286 636 0 S1BEG[0]
rlabel metal2 20654 738 20654 738 0 S1BEG[1]
rlabel metal2 21022 908 21022 908 0 S1BEG[2]
rlabel metal2 21390 636 21390 636 0 S1BEG[3]
rlabel metal2 24702 806 24702 806 0 S2BEG[0]
rlabel metal2 25070 636 25070 636 0 S2BEG[1]
rlabel metal2 25438 636 25438 636 0 S2BEG[2]
rlabel metal2 25951 68 25951 68 0 S2BEG[3]
rlabel metal2 26174 806 26174 806 0 S2BEG[4]
rlabel metal2 26542 636 26542 636 0 S2BEG[5]
rlabel metal2 27055 68 27055 68 0 S2BEG[6]
rlabel metal2 27423 68 27423 68 0 S2BEG[7]
rlabel metal2 21659 68 21659 68 0 S2BEGb[0]
rlabel metal2 22126 704 22126 704 0 S2BEGb[1]
rlabel metal2 22494 908 22494 908 0 S2BEGb[2]
rlabel metal2 22862 636 22862 636 0 S2BEGb[3]
rlabel metal2 23230 636 23230 636 0 S2BEGb[4]
rlabel metal2 23598 908 23598 908 0 S2BEGb[5]
rlabel metal2 23966 143 23966 143 0 S2BEGb[6]
rlabel metal2 24479 68 24479 68 0 S2BEGb[7]
rlabel metal2 27791 68 27791 68 0 S4BEG[0]
rlabel metal2 31326 806 31326 806 0 S4BEG[10]
rlabel metal2 31694 772 31694 772 0 S4BEG[11]
rlabel metal2 32207 68 32207 68 0 S4BEG[12]
rlabel metal2 32575 68 32575 68 0 S4BEG[13]
rlabel metal2 32943 68 32943 68 0 S4BEG[14]
rlabel metal2 33311 68 33311 68 0 S4BEG[15]
rlabel metal2 28014 143 28014 143 0 S4BEG[1]
rlabel metal2 28527 68 28527 68 0 S4BEG[2]
rlabel metal2 28849 68 28849 68 0 S4BEG[3]
rlabel metal2 29118 908 29118 908 0 S4BEG[4]
rlabel metal2 29486 143 29486 143 0 S4BEG[5]
rlabel metal2 29999 68 29999 68 0 S4BEG[6]
rlabel metal2 30275 68 30275 68 0 S4BEG[7]
rlabel metal2 30735 68 30735 68 0 S4BEG[8]
rlabel metal2 30958 908 30958 908 0 S4BEG[9]
rlabel metal2 33679 68 33679 68 0 SS4BEG[0]
rlabel metal2 37214 755 37214 755 0 SS4BEG[10]
rlabel metal2 37727 68 37727 68 0 SS4BEG[11]
rlabel metal2 38095 68 38095 68 0 SS4BEG[12]
rlabel metal2 38463 68 38463 68 0 SS4BEG[13]
rlabel metal2 38831 68 38831 68 0 SS4BEG[14]
rlabel metal2 39199 68 39199 68 0 SS4BEG[15]
rlabel metal2 34047 68 34047 68 0 SS4BEG[1]
rlabel metal2 34270 772 34270 772 0 SS4BEG[2]
rlabel metal2 34638 908 34638 908 0 SS4BEG[3]
rlabel metal2 35006 806 35006 806 0 SS4BEG[4]
rlabel metal2 35519 68 35519 68 0 SS4BEG[5]
rlabel metal2 35795 68 35795 68 0 SS4BEG[6]
rlabel metal2 36110 908 36110 908 0 SS4BEG[7]
rlabel metal2 36623 68 36623 68 0 SS4BEG[8]
rlabel metal2 36991 68 36991 68 0 SS4BEG[9]
rlabel metal2 39475 68 39475 68 0 UserCLK
rlabel metal1 2024 8602 2024 8602 0 UserCLKo
rlabel metal2 41170 816 41170 816 0 net1
rlabel metal1 45586 1972 45586 1972 0 net10
rlabel metal1 25714 1292 25714 1292 0 net100
rlabel metal1 25898 1972 25898 1972 0 net101
rlabel metal1 26312 1326 26312 1326 0 net102
rlabel metal1 26772 1326 26772 1326 0 net103
rlabel metal1 27324 1326 27324 1326 0 net104
rlabel metal1 27692 1326 27692 1326 0 net105
rlabel metal1 21252 1326 21252 1326 0 net106
rlabel metal1 22218 1360 22218 1360 0 net107
rlabel metal1 21206 2040 21206 2040 0 net108
rlabel metal1 22862 1292 22862 1292 0 net109
rlabel metal1 45954 1938 45954 1938 0 net11
rlabel metal2 21942 1462 21942 1462 0 net110
rlabel metal1 22862 2040 22862 2040 0 net111
rlabel metal1 23736 1326 23736 1326 0 net112
rlabel metal1 24334 1326 24334 1326 0 net113
rlabel metal1 28152 1326 28152 1326 0 net114
rlabel metal1 32062 1258 32062 1258 0 net115
rlabel metal1 32476 1326 32476 1326 0 net116
rlabel metal1 32890 1972 32890 1972 0 net117
rlabel metal1 33304 1326 33304 1326 0 net118
rlabel metal1 33442 1258 33442 1258 0 net119
rlabel metal1 28106 2482 28106 2482 0 net12
rlabel metal1 28520 2074 28520 2074 0 net120
rlabel metal1 28474 1972 28474 1972 0 net121
rlabel metal1 28520 1258 28520 1258 0 net122
rlabel metal1 29348 1326 29348 1326 0 net123
rlabel metal1 29946 2006 29946 2006 0 net124
rlabel metal2 30406 1530 30406 1530 0 net125
rlabel metal1 30636 1326 30636 1326 0 net126
rlabel metal1 31510 1360 31510 1360 0 net127
rlabel metal2 31602 2108 31602 2108 0 net128
rlabel metal1 31188 2006 31188 2006 0 net129
rlabel metal1 40802 1462 40802 1462 0 net13
rlabel metal1 33718 1904 33718 1904 0 net130
rlabel via2 16514 2091 16514 2091 0 net131
rlabel metal2 16238 1785 16238 1785 0 net132
rlabel metal2 39008 3604 39008 3604 0 net133
rlabel metal1 29256 2890 29256 2890 0 net134
rlabel metal2 20562 2295 20562 2295 0 net135
rlabel metal2 40250 714 40250 714 0 net136
rlabel metal2 34822 1088 34822 1088 0 net137
rlabel metal3 22540 2788 22540 2788 0 net138
rlabel metal2 19090 629 19090 629 0 net139
rlabel metal1 41262 1836 41262 1836 0 net14
rlabel metal2 19642 1377 19642 1377 0 net140
rlabel metal1 36478 1224 36478 1224 0 net141
rlabel metal2 18538 1649 18538 1649 0 net142
rlabel metal1 17434 2074 17434 2074 0 net143
rlabel metal1 25760 3026 25760 3026 0 net144
rlabel metal1 27554 4454 27554 4454 0 net145
rlabel metal2 6578 8602 6578 8602 0 net146
rlabel metal2 39146 2057 39146 2057 0 net15
rlabel metal1 26404 3094 26404 3094 0 net16
rlabel metal2 41630 2737 41630 2737 0 net17
rlabel metal2 42918 884 42918 884 0 net18
rlabel metal2 43194 1241 43194 1241 0 net19
rlabel metal1 43746 408 43746 408 0 net2
rlabel metal1 43470 442 43470 442 0 net20
rlabel metal2 1610 1632 1610 1632 0 net21
rlabel metal2 1794 850 1794 850 0 net22
rlabel metal2 2162 1088 2162 1088 0 net23
rlabel metal2 2530 884 2530 884 0 net24
rlabel metal2 12650 425 12650 425 0 net25
rlabel metal1 20010 2584 20010 2584 0 net26
rlabel metal2 17250 782 17250 782 0 net27
rlabel metal2 14582 1088 14582 1088 0 net28
rlabel metal2 15134 1071 15134 1071 0 net29
rlabel metal1 43010 510 43010 510 0 net3
rlabel metal2 14766 1003 14766 1003 0 net30
rlabel metal1 13662 1326 13662 1326 0 net31
rlabel metal2 13662 1326 13662 1326 0 net32
rlabel metal1 15318 4182 15318 4182 0 net33
rlabel metal2 4002 3505 4002 3505 0 net34
rlabel metal3 17940 3060 17940 3060 0 net35
rlabel metal1 16744 4522 16744 4522 0 net36
rlabel metal1 20240 3366 20240 3366 0 net37
rlabel metal1 20976 2822 20976 2822 0 net38
rlabel metal2 5106 986 5106 986 0 net39
rlabel metal2 44482 2006 44482 2006 0 net4
rlabel metal1 17618 3502 17618 3502 0 net40
rlabel metal1 18492 3162 18492 3162 0 net41
rlabel metal1 21068 3434 21068 3434 0 net42
rlabel metal2 12834 714 12834 714 0 net43
rlabel metal2 28566 1598 28566 1598 0 net44
rlabel metal2 13938 2924 13938 2924 0 net45
rlabel metal2 13938 816 13938 816 0 net46
rlabel metal2 14306 782 14306 782 0 net47
rlabel metal2 32890 1581 32890 1581 0 net48
rlabel metal2 33350 1428 33350 1428 0 net49
rlabel metal1 43838 1530 43838 1530 0 net5
rlabel metal1 17250 544 17250 544 0 net50
rlabel metal2 32246 1241 32246 1241 0 net51
rlabel metal2 10626 697 10626 697 0 net52
rlabel metal2 10994 1037 10994 1037 0 net53
rlabel metal1 17342 748 17342 748 0 net54
rlabel metal2 30130 1564 30130 1564 0 net55
rlabel metal3 21344 3468 21344 3468 0 net56
rlabel metal1 14490 1224 14490 1224 0 net57
rlabel metal1 17618 1530 17618 1530 0 net58
rlabel metal1 17894 1190 17894 1190 0 net59
rlabel metal2 45034 1768 45034 1768 0 net6
rlabel metal1 18906 1292 18906 1292 0 net60
rlabel metal1 18538 1530 18538 1530 0 net61
rlabel metal1 19550 1360 19550 1360 0 net62
rlabel metal2 19550 1734 19550 1734 0 net63
rlabel metal2 14858 748 14858 748 0 net64
rlabel metal1 15318 1530 15318 1530 0 net65
rlabel metal1 15640 1530 15640 1530 0 net66
rlabel metal1 15778 1224 15778 1224 0 net67
rlabel metal1 16192 1530 16192 1530 0 net68
rlabel metal1 16560 1190 16560 1190 0 net69
rlabel metal1 44620 1190 44620 1190 0 net7
rlabel metal1 16882 1530 16882 1530 0 net70
rlabel metal1 17158 1462 17158 1462 0 net71
rlabel metal2 17250 1768 17250 1768 0 net72
rlabel metal1 39698 850 39698 850 0 net73
rlabel metal1 6486 8840 6486 8840 0 net74
rlabel metal1 26358 8466 26358 8466 0 net75
rlabel metal1 28612 2618 28612 2618 0 net76
rlabel metal2 30774 6900 30774 6900 0 net77
rlabel metal1 33028 8466 33028 8466 0 net78
rlabel metal1 35236 2618 35236 2618 0 net79
rlabel metal1 45310 1904 45310 1904 0 net8
rlabel metal1 37490 2618 37490 2618 0 net80
rlabel metal1 42320 8398 42320 8398 0 net81
rlabel metal1 41906 2618 41906 2618 0 net82
rlabel metal1 44482 8466 44482 8466 0 net83
rlabel metal1 45908 2618 45908 2618 0 net84
rlabel metal1 6394 8908 6394 8908 0 net85
rlabel metal1 8970 8500 8970 8500 0 net86
rlabel metal1 10810 8398 10810 8398 0 net87
rlabel metal2 13018 8704 13018 8704 0 net88
rlabel metal1 18929 8398 18929 8398 0 net89
rlabel metal2 44022 1598 44022 1598 0 net9
rlabel metal1 17618 2618 17618 2618 0 net90
rlabel metal1 19780 2618 19780 2618 0 net91
rlabel metal1 21988 8466 21988 8466 0 net92
rlabel metal1 24656 8466 24656 8466 0 net93
rlabel metal1 19872 1326 19872 1326 0 net94
rlabel metal1 20148 1258 20148 1258 0 net95
rlabel metal1 20562 1938 20562 1938 0 net96
rlabel metal1 20516 1326 20516 1326 0 net97
rlabel metal2 24886 1496 24886 1496 0 net98
rlabel metal1 25346 1360 25346 1360 0 net99
<< properties >>
string FIXED_BBOX 0 0 48000 10000
<< end >>
