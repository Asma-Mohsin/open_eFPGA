magic
tech sky130A
magscale 1 2
timestamp 1733308812
<< viali >>
rect 4997 7497 5031 7531
rect 5549 7497 5583 7531
rect 6377 7497 6411 7531
rect 7021 7497 7055 7531
rect 7573 7497 7607 7531
rect 8125 7497 8159 7531
rect 8677 7497 8711 7531
rect 9873 7497 9907 7531
rect 10977 7497 11011 7531
rect 11805 7497 11839 7531
rect 12173 7497 12207 7531
rect 12725 7497 12759 7531
rect 13277 7497 13311 7531
rect 13829 7497 13863 7531
rect 14749 7497 14783 7531
rect 15301 7497 15335 7531
rect 15853 7497 15887 7531
rect 16405 7497 16439 7531
rect 17325 7497 17359 7531
rect 17877 7497 17911 7531
rect 18429 7497 18463 7531
rect 20821 7497 20855 7531
rect 22569 7497 22603 7531
rect 23397 7497 23431 7531
rect 23765 7497 23799 7531
rect 25237 7497 25271 7531
rect 25973 7497 26007 7531
rect 27813 7497 27847 7531
rect 31401 7497 31435 7531
rect 31953 7497 31987 7531
rect 33425 7497 33459 7531
rect 33701 7497 33735 7531
rect 34161 7497 34195 7531
rect 34897 7497 34931 7531
rect 35449 7497 35483 7531
rect 36553 7497 36587 7531
rect 38025 7497 38059 7531
rect 40049 7497 40083 7531
rect 41245 7497 41279 7531
rect 5273 7429 5307 7463
rect 6745 7429 6779 7463
rect 7849 7429 7883 7463
rect 8401 7429 8435 7463
rect 11253 7429 11287 7463
rect 15025 7429 15059 7463
rect 20361 7429 20395 7463
rect 36461 7429 36495 7463
rect 40509 7429 40543 7463
rect 4721 7361 4755 7395
rect 5825 7361 5859 7395
rect 6561 7361 6595 7395
rect 7297 7361 7331 7395
rect 9137 7361 9171 7395
rect 9505 7361 9539 7395
rect 10149 7361 10183 7395
rect 10701 7361 10735 7395
rect 12449 7361 12483 7395
rect 13001 7361 13035 7395
rect 13553 7361 13587 7395
rect 14289 7361 14323 7395
rect 14473 7361 14507 7395
rect 15577 7361 15611 7395
rect 16129 7361 16163 7395
rect 16865 7361 16899 7395
rect 17049 7361 17083 7395
rect 17601 7361 17635 7395
rect 18153 7361 18187 7395
rect 18705 7361 18739 7395
rect 19441 7361 19475 7395
rect 19993 7361 20027 7395
rect 20637 7361 20671 7395
rect 20913 7361 20947 7395
rect 21373 7361 21407 7395
rect 21649 7361 21683 7395
rect 22017 7361 22051 7395
rect 22293 7361 22327 7395
rect 22385 7361 22419 7395
rect 22845 7361 22879 7395
rect 23121 7361 23155 7395
rect 23213 7361 23247 7395
rect 23673 7361 23707 7395
rect 23949 7361 23983 7395
rect 24225 7361 24259 7395
rect 24409 7361 24443 7395
rect 24869 7361 24903 7395
rect 24961 7361 24995 7395
rect 25421 7361 25455 7395
rect 25697 7361 25731 7395
rect 25789 7361 25823 7395
rect 26249 7361 26283 7395
rect 26525 7361 26559 7395
rect 26801 7361 26835 7395
rect 27169 7361 27203 7395
rect 27445 7361 27479 7395
rect 27721 7361 27755 7395
rect 27997 7361 28031 7395
rect 28273 7361 28307 7395
rect 28549 7361 28583 7395
rect 28825 7361 28859 7395
rect 29101 7361 29135 7395
rect 29377 7361 29411 7395
rect 29745 7361 29779 7395
rect 30021 7361 30055 7395
rect 30297 7361 30331 7395
rect 30573 7361 30607 7395
rect 30665 7361 30699 7395
rect 30941 7361 30975 7395
rect 31217 7361 31251 7395
rect 31493 7361 31527 7395
rect 31769 7361 31803 7395
rect 32137 7361 32171 7395
rect 32413 7361 32447 7395
rect 32689 7361 32723 7395
rect 32965 7361 32999 7395
rect 33241 7361 33275 7395
rect 33517 7361 33551 7395
rect 34069 7361 34103 7395
rect 34805 7361 34839 7395
rect 35357 7361 35391 7395
rect 35909 7361 35943 7395
rect 37105 7361 37139 7395
rect 37381 7361 37415 7395
rect 37933 7361 37967 7395
rect 38485 7361 38519 7395
rect 39037 7361 39071 7395
rect 39681 7361 39715 7395
rect 39957 7361 39991 7395
rect 41153 7361 41187 7395
rect 41429 7361 41463 7395
rect 6101 7225 6135 7259
rect 8953 7225 8987 7259
rect 10517 7225 10551 7259
rect 14105 7225 14139 7259
rect 21189 7225 21223 7259
rect 22661 7225 22695 7259
rect 24593 7225 24627 7259
rect 24685 7225 24719 7259
rect 25513 7225 25547 7259
rect 26985 7225 27019 7259
rect 28089 7225 28123 7259
rect 29193 7225 29227 7259
rect 33149 7225 33183 7259
rect 16681 7157 16715 7191
rect 18797 7157 18831 7191
rect 19533 7157 19567 7191
rect 21097 7157 21131 7191
rect 21465 7157 21499 7191
rect 21833 7157 21867 7191
rect 22109 7157 22143 7191
rect 22937 7157 22971 7191
rect 23489 7157 23523 7191
rect 24041 7157 24075 7191
rect 25145 7157 25179 7191
rect 26065 7157 26099 7191
rect 26341 7157 26375 7191
rect 26617 7157 26651 7191
rect 27261 7157 27295 7191
rect 27537 7157 27571 7191
rect 28365 7157 28399 7191
rect 28641 7157 28675 7191
rect 28917 7157 28951 7191
rect 29561 7157 29595 7191
rect 29837 7157 29871 7191
rect 30113 7157 30147 7191
rect 30389 7157 30423 7191
rect 30849 7157 30883 7191
rect 31125 7157 31159 7191
rect 31677 7157 31711 7191
rect 32321 7157 32355 7191
rect 32597 7157 32631 7191
rect 32873 7157 32907 7191
rect 36001 7157 36035 7191
rect 36921 7157 36955 7191
rect 37473 7157 37507 7191
rect 38761 7157 38795 7191
rect 39129 7157 39163 7191
rect 39497 7157 39531 7191
rect 40601 7157 40635 7191
rect 40969 7157 41003 7191
rect 5181 6953 5215 6987
rect 5733 6953 5767 6987
rect 6837 6953 6871 6987
rect 13093 6953 13127 6987
rect 13645 6953 13679 6987
rect 14565 6953 14599 6987
rect 18889 6953 18923 6987
rect 26433 6953 26467 6987
rect 21741 6885 21775 6919
rect 7573 6817 7607 6851
rect 8125 6817 8159 6851
rect 8677 6817 8711 6851
rect 9597 6817 9631 6851
rect 10517 6817 10551 6851
rect 11069 6817 11103 6851
rect 11621 6817 11655 6851
rect 12725 6817 12759 6851
rect 15301 6817 15335 6851
rect 15853 6817 15887 6851
rect 16405 6817 16439 6851
rect 16957 6817 16991 6851
rect 17509 6817 17543 6851
rect 18061 6817 18095 6851
rect 18613 6817 18647 6851
rect 35725 6817 35759 6851
rect 36277 6817 36311 6851
rect 37933 6817 37967 6851
rect 40785 6817 40819 6851
rect 6193 6749 6227 6783
rect 6745 6749 6779 6783
rect 7849 6749 7883 6783
rect 9303 6749 9337 6783
rect 12265 6749 12299 6783
rect 14289 6749 14323 6783
rect 15577 6749 15611 6783
rect 19073 6749 19107 6783
rect 19349 6749 19383 6783
rect 19625 6749 19659 6783
rect 19901 6749 19935 6783
rect 20177 6749 20211 6783
rect 20453 6749 20487 6783
rect 20729 6749 20763 6783
rect 21005 6749 21039 6783
rect 21281 6749 21315 6783
rect 21557 6749 21591 6783
rect 22845 6749 22879 6783
rect 23029 6749 23063 6783
rect 24869 6749 24903 6783
rect 25145 6749 25179 6783
rect 25421 6749 25455 6783
rect 26249 6749 26283 6783
rect 26525 6749 26559 6783
rect 26801 6749 26835 6783
rect 27169 6749 27203 6783
rect 27537 6749 27571 6783
rect 27905 6749 27939 6783
rect 28273 6749 28307 6783
rect 28733 6749 28767 6783
rect 29193 6749 29227 6783
rect 29653 6749 29687 6783
rect 30021 6749 30055 6783
rect 30297 6749 30331 6783
rect 31217 6749 31251 6783
rect 32597 6749 32631 6783
rect 33149 6749 33183 6783
rect 33425 6749 33459 6783
rect 33885 6749 33919 6783
rect 34161 6749 34195 6783
rect 34253 6749 34287 6783
rect 34897 6749 34931 6783
rect 35173 6749 35207 6783
rect 39313 6749 39347 6783
rect 39957 6749 39991 6783
rect 40509 6749 40543 6783
rect 5089 6681 5123 6715
rect 5641 6681 5675 6715
rect 7297 6681 7331 6715
rect 8401 6681 8435 6715
rect 10241 6681 10275 6715
rect 10793 6681 10827 6715
rect 11345 6681 11379 6715
rect 11897 6681 11931 6715
rect 12449 6681 12483 6715
rect 13001 6681 13035 6715
rect 13553 6681 13587 6715
rect 14473 6681 14507 6715
rect 15025 6681 15059 6715
rect 16129 6681 16163 6715
rect 16681 6681 16715 6715
rect 17233 6681 17267 6715
rect 17785 6681 17819 6715
rect 18337 6681 18371 6715
rect 35449 6681 35483 6715
rect 36001 6681 36035 6715
rect 36553 6681 36587 6715
rect 37105 6681 37139 6715
rect 37657 6681 37691 6715
rect 38209 6681 38243 6715
rect 38761 6681 38795 6715
rect 6285 6613 6319 6647
rect 14105 6613 14139 6647
rect 19533 6613 19567 6647
rect 19809 6613 19843 6647
rect 20085 6613 20119 6647
rect 20361 6613 20395 6647
rect 20637 6613 20671 6647
rect 20913 6613 20947 6647
rect 21189 6613 21223 6647
rect 21465 6613 21499 6647
rect 22661 6613 22695 6647
rect 23213 6613 23247 6647
rect 25053 6613 25087 6647
rect 25329 6613 25363 6647
rect 25605 6613 25639 6647
rect 26709 6613 26743 6647
rect 26985 6613 27019 6647
rect 27353 6613 27387 6647
rect 27721 6613 27755 6647
rect 28089 6613 28123 6647
rect 28457 6613 28491 6647
rect 28917 6613 28951 6647
rect 29377 6613 29411 6647
rect 29837 6613 29871 6647
rect 30205 6613 30239 6647
rect 30481 6613 30515 6647
rect 31401 6613 31435 6647
rect 32413 6613 32447 6647
rect 33333 6613 33367 6647
rect 33609 6613 33643 6647
rect 33701 6613 33735 6647
rect 33977 6613 34011 6647
rect 34437 6613 34471 6647
rect 34989 6613 35023 6647
rect 36645 6613 36679 6647
rect 37197 6613 37231 6647
rect 38301 6613 38335 6647
rect 38853 6613 38887 6647
rect 39405 6613 39439 6647
rect 40049 6613 40083 6647
rect 6009 6409 6043 6443
rect 7849 6409 7883 6443
rect 8677 6409 8711 6443
rect 9229 6409 9263 6443
rect 9781 6409 9815 6443
rect 11529 6409 11563 6443
rect 11989 6409 12023 6443
rect 13829 6409 13863 6443
rect 14289 6409 14323 6443
rect 14657 6409 14691 6443
rect 15301 6409 15335 6443
rect 15669 6409 15703 6443
rect 16129 6409 16163 6443
rect 17601 6409 17635 6443
rect 18061 6409 18095 6443
rect 18337 6409 18371 6443
rect 18613 6409 18647 6443
rect 18981 6409 19015 6443
rect 22477 6409 22511 6443
rect 37289 6409 37323 6443
rect 9689 6341 9723 6375
rect 10241 6341 10275 6375
rect 5917 6273 5951 6307
rect 6193 6273 6227 6307
rect 8033 6273 8067 6307
rect 8585 6273 8619 6307
rect 9137 6273 9171 6307
rect 11069 6273 11103 6307
rect 11713 6273 11747 6307
rect 11897 6273 11931 6307
rect 14013 6273 14047 6307
rect 14197 6273 14231 6307
rect 14841 6273 14875 6307
rect 15485 6273 15519 6307
rect 15853 6273 15887 6307
rect 16313 6273 16347 6307
rect 16865 6273 16899 6307
rect 17233 6273 17267 6307
rect 17509 6273 17543 6307
rect 17785 6273 17819 6307
rect 18245 6273 18279 6307
rect 18521 6273 18555 6307
rect 18797 6273 18831 6307
rect 19165 6273 19199 6307
rect 20453 6273 20487 6307
rect 21833 6273 21867 6307
rect 22293 6273 22327 6307
rect 22753 6273 22787 6307
rect 25789 6273 25823 6307
rect 34253 6273 34287 6307
rect 37473 6273 37507 6307
rect 37749 6273 37783 6307
rect 5733 6137 5767 6171
rect 10885 6137 10919 6171
rect 16681 6137 16715 6171
rect 17325 6137 17359 6171
rect 37565 6137 37599 6171
rect 10333 6069 10367 6103
rect 20637 6069 20671 6103
rect 22017 6069 22051 6103
rect 22937 6069 22971 6103
rect 25973 6069 26007 6103
rect 34069 6069 34103 6103
rect 13001 5865 13035 5899
rect 12817 5661 12851 5695
rect 20821 5185 20855 5219
rect 21005 4981 21039 5015
rect 18889 3145 18923 3179
rect 18705 3009 18739 3043
rect 22937 3009 22971 3043
rect 25053 3009 25087 3043
rect 23121 2873 23155 2907
rect 25237 2805 25271 2839
rect 3985 2601 4019 2635
rect 11989 2601 12023 2635
rect 18337 2601 18371 2635
rect 20453 2601 20487 2635
rect 22569 2601 22603 2635
rect 24685 2601 24719 2635
rect 33149 2601 33183 2635
rect 34713 2601 34747 2635
rect 36829 2601 36863 2635
rect 37841 2601 37875 2635
rect 39497 2601 39531 2635
rect 41613 2601 41647 2635
rect 43361 2601 43395 2635
rect 16221 2533 16255 2567
rect 16865 2533 16899 2567
rect 29101 2533 29135 2567
rect 35265 2533 35299 2567
rect 37381 2533 37415 2567
rect 6653 2465 6687 2499
rect 8033 2465 8067 2499
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 6377 2397 6411 2431
rect 7757 2397 7791 2431
rect 9873 2397 9907 2431
rect 12173 2397 12207 2431
rect 14289 2397 14323 2431
rect 16405 2397 16439 2431
rect 16681 2397 16715 2431
rect 18521 2397 18555 2431
rect 20637 2397 20671 2431
rect 22753 2397 22787 2431
rect 24869 2397 24903 2431
rect 27169 2397 27203 2431
rect 28917 2397 28951 2431
rect 31033 2397 31067 2431
rect 33333 2397 33367 2431
rect 34897 2397 34931 2431
rect 35449 2397 35483 2431
rect 37013 2397 37047 2431
rect 37565 2397 37599 2431
rect 38025 2397 38059 2431
rect 39681 2397 39715 2431
rect 41797 2397 41831 2431
rect 43545 2397 43579 2431
rect 3893 2329 3927 2363
rect 14657 2329 14691 2363
rect 14841 2329 14875 2363
rect 10057 2261 10091 2295
rect 14105 2261 14139 2295
rect 26985 2261 27019 2295
rect 31217 2261 31251 2295
<< metal1 >>
rect 16390 8508 16396 8560
rect 16448 8548 16454 8560
rect 32582 8548 32588 8560
rect 16448 8520 32588 8548
rect 16448 8508 16454 8520
rect 32582 8508 32588 8520
rect 32640 8508 32646 8560
rect 15838 8440 15844 8492
rect 15896 8480 15902 8492
rect 33502 8480 33508 8492
rect 15896 8452 33508 8480
rect 15896 8440 15902 8452
rect 33502 8440 33508 8452
rect 33560 8440 33566 8492
rect 15470 8372 15476 8424
rect 15528 8412 15534 8424
rect 33686 8412 33692 8424
rect 15528 8384 33692 8412
rect 15528 8372 15534 8384
rect 33686 8372 33692 8384
rect 33744 8372 33750 8424
rect 13354 8304 13360 8356
rect 13412 8344 13418 8356
rect 36170 8344 36176 8356
rect 13412 8316 36176 8344
rect 13412 8304 13418 8316
rect 36170 8304 36176 8316
rect 36228 8304 36234 8356
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 14274 8276 14280 8288
rect 13872 8248 14280 8276
rect 13872 8236 13878 8248
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 25314 8236 25320 8288
rect 25372 8276 25378 8288
rect 25958 8276 25964 8288
rect 25372 8248 25964 8276
rect 25372 8236 25378 8248
rect 25958 8236 25964 8248
rect 26016 8236 26022 8288
rect 28810 8236 28816 8288
rect 28868 8276 28874 8288
rect 29730 8276 29736 8288
rect 28868 8248 29736 8276
rect 28868 8236 28874 8248
rect 29730 8236 29736 8248
rect 29788 8236 29794 8288
rect 29914 8236 29920 8288
rect 29972 8276 29978 8288
rect 30742 8276 30748 8288
rect 29972 8248 30748 8276
rect 29972 8236 29978 8248
rect 30742 8236 30748 8248
rect 30800 8236 30806 8288
rect 9646 8180 16344 8208
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 9646 8072 9674 8180
rect 16316 8152 16344 8180
rect 23198 8168 23204 8220
rect 23256 8208 23262 8220
rect 23256 8180 31524 8208
rect 23256 8168 23262 8180
rect 12434 8100 12440 8152
rect 12492 8140 12498 8152
rect 16114 8140 16120 8152
rect 12492 8112 16120 8140
rect 12492 8100 12498 8112
rect 16114 8100 16120 8112
rect 16172 8100 16178 8152
rect 16298 8100 16304 8152
rect 16356 8100 16362 8152
rect 19426 8100 19432 8152
rect 19484 8140 19490 8152
rect 19484 8112 29132 8140
rect 19484 8100 19490 8112
rect 7800 8044 9674 8072
rect 7800 8032 7806 8044
rect 13630 8032 13636 8084
rect 13688 8072 13694 8084
rect 22094 8072 22100 8084
rect 13688 8044 22100 8072
rect 13688 8032 13694 8044
rect 22094 8032 22100 8044
rect 22152 8032 22158 8084
rect 29104 8072 29132 8112
rect 29178 8100 29184 8152
rect 29236 8140 29242 8152
rect 30282 8140 30288 8152
rect 29236 8112 30288 8140
rect 29236 8100 29242 8112
rect 30282 8100 30288 8112
rect 30340 8100 30346 8152
rect 31202 8072 31208 8084
rect 29104 8044 31208 8072
rect 31202 8032 31208 8044
rect 31260 8032 31266 8084
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 11790 8004 11796 8016
rect 11112 7976 11796 8004
rect 11112 7964 11118 7976
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 12158 7964 12164 8016
rect 12216 8004 12222 8016
rect 20714 8004 20720 8016
rect 12216 7976 20720 8004
rect 12216 7964 12222 7976
rect 20714 7964 20720 7976
rect 20772 7964 20778 8016
rect 23290 7964 23296 8016
rect 23348 8004 23354 8016
rect 30650 8004 30656 8016
rect 23348 7976 30656 8004
rect 23348 7964 23354 7976
rect 30650 7964 30656 7976
rect 30708 7964 30714 8016
rect 31496 7948 31524 8180
rect 14090 7896 14096 7948
rect 14148 7936 14154 7948
rect 25314 7936 25320 7948
rect 14148 7908 25320 7936
rect 14148 7896 14154 7908
rect 25314 7896 25320 7908
rect 25372 7896 25378 7948
rect 26786 7896 26792 7948
rect 26844 7936 26850 7948
rect 31386 7936 31392 7948
rect 26844 7908 31392 7936
rect 26844 7896 26850 7908
rect 31386 7896 31392 7908
rect 31444 7896 31450 7948
rect 31478 7896 31484 7948
rect 31536 7896 31542 7948
rect 20346 7868 20352 7880
rect 13648 7840 20352 7868
rect 8386 7760 8392 7812
rect 8444 7800 8450 7812
rect 13648 7800 13676 7840
rect 20346 7828 20352 7840
rect 20404 7828 20410 7880
rect 26878 7828 26884 7880
rect 26936 7868 26942 7880
rect 32674 7868 32680 7880
rect 26936 7840 32680 7868
rect 26936 7828 26942 7840
rect 32674 7828 32680 7840
rect 32732 7828 32738 7880
rect 8444 7772 13676 7800
rect 8444 7760 8450 7772
rect 16298 7760 16304 7812
rect 16356 7800 16362 7812
rect 22922 7800 22928 7812
rect 16356 7772 22928 7800
rect 16356 7760 16362 7772
rect 22922 7760 22928 7772
rect 22980 7760 22986 7812
rect 27430 7760 27436 7812
rect 27488 7800 27494 7812
rect 28534 7800 28540 7812
rect 27488 7772 28540 7800
rect 27488 7760 27494 7772
rect 28534 7760 28540 7772
rect 28592 7760 28598 7812
rect 6730 7692 6736 7744
rect 6788 7732 6794 7744
rect 21082 7732 21088 7744
rect 6788 7704 21088 7732
rect 6788 7692 6794 7704
rect 21082 7692 21088 7704
rect 21140 7692 21146 7744
rect 27246 7692 27252 7744
rect 27304 7732 27310 7744
rect 28442 7732 28448 7744
rect 27304 7704 28448 7732
rect 27304 7692 27310 7704
rect 28442 7692 28448 7704
rect 28500 7692 28506 7744
rect 1104 7642 44040 7664
rect 1104 7590 11644 7642
rect 11696 7590 11708 7642
rect 11760 7590 11772 7642
rect 11824 7590 11836 7642
rect 11888 7590 11900 7642
rect 11952 7590 22338 7642
rect 22390 7590 22402 7642
rect 22454 7590 22466 7642
rect 22518 7590 22530 7642
rect 22582 7590 22594 7642
rect 22646 7590 33032 7642
rect 33084 7590 33096 7642
rect 33148 7590 33160 7642
rect 33212 7590 33224 7642
rect 33276 7590 33288 7642
rect 33340 7590 43726 7642
rect 43778 7590 43790 7642
rect 43842 7590 43854 7642
rect 43906 7590 43918 7642
rect 43970 7590 43982 7642
rect 44034 7590 44040 7642
rect 1104 7568 44040 7590
rect 4985 7531 5043 7537
rect 4985 7497 4997 7531
rect 5031 7528 5043 7531
rect 5442 7528 5448 7540
rect 5031 7500 5448 7528
rect 5031 7497 5043 7500
rect 4985 7491 5043 7497
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 5537 7531 5595 7537
rect 5537 7497 5549 7531
rect 5583 7528 5595 7531
rect 5994 7528 6000 7540
rect 5583 7500 6000 7528
rect 5583 7497 5595 7500
rect 5537 7491 5595 7497
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 6365 7531 6423 7537
rect 6365 7497 6377 7531
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 7009 7531 7067 7537
rect 7009 7497 7021 7531
rect 7055 7528 7067 7531
rect 7374 7528 7380 7540
rect 7055 7500 7380 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 5261 7463 5319 7469
rect 5261 7429 5273 7463
rect 5307 7460 5319 7463
rect 6380 7460 6408 7491
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 7561 7531 7619 7537
rect 7561 7497 7573 7531
rect 7607 7528 7619 7531
rect 7926 7528 7932 7540
rect 7607 7500 7932 7528
rect 7607 7497 7619 7500
rect 7561 7491 7619 7497
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 8113 7531 8171 7537
rect 8113 7497 8125 7531
rect 8159 7528 8171 7531
rect 8478 7528 8484 7540
rect 8159 7500 8484 7528
rect 8159 7497 8171 7500
rect 8113 7491 8171 7497
rect 8478 7488 8484 7500
rect 8536 7488 8542 7540
rect 8665 7531 8723 7537
rect 8665 7497 8677 7531
rect 8711 7528 8723 7531
rect 9030 7528 9036 7540
rect 8711 7500 9036 7528
rect 8711 7497 8723 7500
rect 8665 7491 8723 7497
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 9861 7531 9919 7537
rect 9861 7497 9873 7531
rect 9907 7528 9919 7531
rect 10686 7528 10692 7540
rect 9907 7500 10692 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 10965 7531 11023 7537
rect 10965 7497 10977 7531
rect 11011 7528 11023 7531
rect 11054 7528 11060 7540
rect 11011 7500 11060 7528
rect 11011 7497 11023 7500
rect 10965 7491 11023 7497
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 11793 7531 11851 7537
rect 11793 7528 11805 7531
rect 11164 7500 11805 7528
rect 5307 7432 6408 7460
rect 5307 7429 5319 7432
rect 5261 7423 5319 7429
rect 6730 7420 6736 7472
rect 6788 7420 6794 7472
rect 7837 7463 7895 7469
rect 7837 7429 7849 7463
rect 7883 7429 7895 7463
rect 7837 7423 7895 7429
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7392 4767 7395
rect 5534 7392 5540 7404
rect 4755 7364 5540 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 5810 7352 5816 7404
rect 5868 7352 5874 7404
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6564 7324 6592 7355
rect 7282 7352 7288 7404
rect 7340 7352 7346 7404
rect 7852 7392 7880 7423
rect 8386 7420 8392 7472
rect 8444 7420 8450 7472
rect 10042 7460 10048 7472
rect 9048 7432 10048 7460
rect 9048 7392 9076 7432
rect 10042 7420 10048 7432
rect 10100 7420 10106 7472
rect 7852 7364 9076 7392
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 9493 7395 9551 7401
rect 9493 7361 9505 7395
rect 9539 7392 9551 7395
rect 10137 7395 10195 7401
rect 10137 7392 10149 7395
rect 9539 7364 10149 7392
rect 9539 7361 9551 7364
rect 9493 7355 9551 7361
rect 10137 7361 10149 7364
rect 10183 7392 10195 7395
rect 10594 7392 10600 7404
rect 10183 7364 10600 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 6730 7324 6736 7336
rect 6564 7296 6736 7324
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 9140 7324 9168 7355
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 10689 7395 10747 7401
rect 10689 7361 10701 7395
rect 10735 7392 10747 7395
rect 11164 7392 11192 7500
rect 11793 7497 11805 7500
rect 11839 7528 11851 7531
rect 12066 7528 12072 7540
rect 11839 7500 12072 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 12066 7488 12072 7500
rect 12124 7488 12130 7540
rect 12158 7488 12164 7540
rect 12216 7488 12222 7540
rect 12713 7531 12771 7537
rect 12713 7497 12725 7531
rect 12759 7528 12771 7531
rect 13170 7528 13176 7540
rect 12759 7500 13176 7528
rect 12759 7497 12771 7500
rect 12713 7491 12771 7497
rect 13170 7488 13176 7500
rect 13228 7488 13234 7540
rect 13265 7531 13323 7537
rect 13265 7497 13277 7531
rect 13311 7528 13323 7531
rect 13722 7528 13728 7540
rect 13311 7500 13728 7528
rect 13311 7497 13323 7500
rect 13265 7491 13323 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 13814 7488 13820 7540
rect 13872 7488 13878 7540
rect 14737 7531 14795 7537
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 15102 7528 15108 7540
rect 14783 7500 15108 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 15102 7488 15108 7500
rect 15160 7488 15166 7540
rect 15289 7531 15347 7537
rect 15289 7497 15301 7531
rect 15335 7528 15347 7531
rect 15654 7528 15660 7540
rect 15335 7500 15660 7528
rect 15335 7497 15347 7500
rect 15289 7491 15347 7497
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 15841 7531 15899 7537
rect 15841 7497 15853 7531
rect 15887 7528 15899 7531
rect 16206 7528 16212 7540
rect 15887 7500 16212 7528
rect 15887 7497 15899 7500
rect 15841 7491 15899 7497
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 16393 7531 16451 7537
rect 16393 7497 16405 7531
rect 16439 7528 16451 7531
rect 16758 7528 16764 7540
rect 16439 7500 16764 7528
rect 16439 7497 16451 7500
rect 16393 7491 16451 7497
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 17310 7488 17316 7540
rect 17368 7488 17374 7540
rect 17862 7488 17868 7540
rect 17920 7488 17926 7540
rect 18414 7488 18420 7540
rect 18472 7488 18478 7540
rect 20809 7531 20867 7537
rect 20809 7497 20821 7531
rect 20855 7497 20867 7531
rect 20809 7491 20867 7497
rect 11241 7463 11299 7469
rect 11241 7429 11253 7463
rect 11287 7460 11299 7463
rect 12176 7460 12204 7488
rect 11287 7432 12204 7460
rect 11287 7429 11299 7432
rect 11241 7423 11299 7429
rect 14642 7420 14648 7472
rect 14700 7460 14706 7472
rect 15013 7463 15071 7469
rect 15013 7460 15025 7463
rect 14700 7432 15025 7460
rect 14700 7420 14706 7432
rect 15013 7429 15025 7432
rect 15059 7429 15071 7463
rect 15013 7423 15071 7429
rect 19150 7420 19156 7472
rect 19208 7460 19214 7472
rect 20349 7463 20407 7469
rect 20349 7460 20361 7463
rect 19208 7432 20361 7460
rect 19208 7420 19214 7432
rect 20349 7429 20361 7432
rect 20395 7429 20407 7463
rect 20824 7460 20852 7491
rect 21082 7488 21088 7540
rect 21140 7528 21146 7540
rect 22557 7531 22615 7537
rect 22557 7528 22569 7531
rect 21140 7500 22569 7528
rect 21140 7488 21146 7500
rect 22557 7497 22569 7500
rect 22603 7497 22615 7531
rect 22557 7491 22615 7497
rect 22922 7488 22928 7540
rect 22980 7528 22986 7540
rect 23385 7531 23443 7537
rect 23385 7528 23397 7531
rect 22980 7500 23397 7528
rect 22980 7488 22986 7500
rect 23385 7497 23397 7500
rect 23431 7497 23443 7531
rect 23385 7491 23443 7497
rect 23753 7531 23811 7537
rect 23753 7497 23765 7531
rect 23799 7497 23811 7531
rect 25225 7531 25283 7537
rect 25225 7528 25237 7531
rect 23753 7491 23811 7497
rect 24412 7500 25237 7528
rect 20990 7460 20996 7472
rect 20824 7432 20996 7460
rect 20349 7423 20407 7429
rect 20990 7420 20996 7432
rect 21048 7420 21054 7472
rect 23768 7460 23796 7491
rect 22388 7432 23796 7460
rect 10735 7364 11192 7392
rect 10735 7361 10747 7364
rect 10689 7355 10747 7361
rect 12434 7352 12440 7404
rect 12492 7352 12498 7404
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7392 13047 7395
rect 13262 7392 13268 7404
rect 13035 7364 13268 7392
rect 13035 7361 13047 7364
rect 12989 7355 13047 7361
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7392 13599 7395
rect 14182 7392 14188 7404
rect 13587 7364 14188 7392
rect 13587 7361 13599 7364
rect 13541 7355 13599 7361
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 14274 7352 14280 7404
rect 14332 7352 14338 7404
rect 14458 7352 14464 7404
rect 14516 7352 14522 7404
rect 15562 7352 15568 7404
rect 15620 7352 15626 7404
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7392 16175 7395
rect 16574 7392 16580 7404
rect 16163 7364 16580 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17310 7392 17316 7404
rect 17083 7364 17316 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 16868 7324 16896 7355
rect 17310 7352 17316 7364
rect 17368 7352 17374 7404
rect 17589 7395 17647 7401
rect 17589 7361 17601 7395
rect 17635 7392 17647 7395
rect 17862 7392 17868 7404
rect 17635 7364 17868 7392
rect 17635 7361 17647 7364
rect 17589 7355 17647 7361
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7392 18199 7395
rect 18598 7392 18604 7404
rect 18187 7364 18604 7392
rect 18187 7361 18199 7364
rect 18141 7355 18199 7361
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7392 18751 7395
rect 18966 7392 18972 7404
rect 18739 7364 18972 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 18966 7352 18972 7364
rect 19024 7352 19030 7404
rect 19429 7395 19487 7401
rect 19429 7361 19441 7395
rect 19475 7361 19487 7395
rect 19429 7355 19487 7361
rect 17678 7324 17684 7336
rect 9140 7296 11652 7324
rect 6089 7259 6147 7265
rect 6089 7225 6101 7259
rect 6135 7256 6147 7259
rect 6546 7256 6552 7268
rect 6135 7228 6552 7256
rect 6135 7225 6147 7228
rect 6089 7219 6147 7225
rect 6546 7216 6552 7228
rect 6604 7216 6610 7268
rect 8941 7259 8999 7265
rect 8941 7225 8953 7259
rect 8987 7256 8999 7259
rect 9674 7256 9680 7268
rect 8987 7228 9680 7256
rect 8987 7225 8999 7228
rect 8941 7219 8999 7225
rect 9674 7216 9680 7228
rect 9732 7216 9738 7268
rect 10505 7259 10563 7265
rect 10505 7225 10517 7259
rect 10551 7256 10563 7259
rect 11238 7256 11244 7268
rect 10551 7228 11244 7256
rect 10551 7225 10563 7228
rect 10505 7219 10563 7225
rect 11238 7216 11244 7228
rect 11296 7216 11302 7268
rect 11624 7256 11652 7296
rect 11900 7296 16804 7324
rect 16868 7296 17684 7324
rect 11900 7256 11928 7296
rect 11624 7228 11928 7256
rect 12066 7216 12072 7268
rect 12124 7216 12130 7268
rect 12250 7216 12256 7268
rect 12308 7256 12314 7268
rect 13630 7256 13636 7268
rect 12308 7228 13636 7256
rect 12308 7216 12314 7228
rect 13630 7216 13636 7228
rect 13688 7216 13694 7268
rect 14093 7259 14151 7265
rect 14093 7225 14105 7259
rect 14139 7256 14151 7259
rect 14642 7256 14648 7268
rect 14139 7228 14648 7256
rect 14139 7225 14151 7228
rect 14093 7219 14151 7225
rect 14642 7216 14648 7228
rect 14700 7216 14706 7268
rect 16776 7256 16804 7296
rect 17678 7284 17684 7296
rect 17736 7284 17742 7336
rect 19444 7324 19472 7355
rect 19978 7352 19984 7404
rect 20036 7352 20042 7404
rect 20625 7395 20683 7401
rect 20625 7361 20637 7395
rect 20671 7392 20683 7395
rect 20806 7392 20812 7404
rect 20671 7364 20812 7392
rect 20671 7361 20683 7364
rect 20625 7355 20683 7361
rect 20806 7352 20812 7364
rect 20864 7352 20870 7404
rect 20901 7395 20959 7401
rect 20901 7361 20913 7395
rect 20947 7392 20959 7395
rect 21174 7392 21180 7404
rect 20947 7364 21180 7392
rect 20947 7361 20959 7364
rect 20901 7355 20959 7361
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 21358 7352 21364 7404
rect 21416 7352 21422 7404
rect 21634 7352 21640 7404
rect 21692 7352 21698 7404
rect 22002 7352 22008 7404
rect 22060 7352 22066 7404
rect 22278 7352 22284 7404
rect 22336 7352 22342 7404
rect 22388 7401 22416 7432
rect 22373 7395 22431 7401
rect 22373 7361 22385 7395
rect 22419 7361 22431 7395
rect 22373 7355 22431 7361
rect 22830 7352 22836 7404
rect 22888 7352 22894 7404
rect 23106 7352 23112 7404
rect 23164 7352 23170 7404
rect 23201 7395 23259 7401
rect 23201 7361 23213 7395
rect 23247 7361 23259 7395
rect 23201 7355 23259 7361
rect 23216 7324 23244 7355
rect 23382 7352 23388 7404
rect 23440 7392 23446 7404
rect 23661 7395 23719 7401
rect 23661 7392 23673 7395
rect 23440 7364 23673 7392
rect 23440 7352 23446 7364
rect 23661 7361 23673 7364
rect 23707 7361 23719 7395
rect 23661 7355 23719 7361
rect 23934 7352 23940 7404
rect 23992 7352 23998 7404
rect 24210 7352 24216 7404
rect 24268 7352 24274 7404
rect 24412 7401 24440 7500
rect 25225 7497 25237 7500
rect 25271 7497 25283 7531
rect 25225 7491 25283 7497
rect 25314 7488 25320 7540
rect 25372 7528 25378 7540
rect 25961 7531 26019 7537
rect 25961 7528 25973 7531
rect 25372 7500 25973 7528
rect 25372 7488 25378 7500
rect 25961 7497 25973 7500
rect 26007 7497 26019 7531
rect 25961 7491 26019 7497
rect 26142 7488 26148 7540
rect 26200 7528 26206 7540
rect 26200 7500 26924 7528
rect 26200 7488 26206 7500
rect 24670 7420 24676 7472
rect 24728 7460 24734 7472
rect 24728 7432 25084 7460
rect 24728 7420 24734 7432
rect 24397 7395 24455 7401
rect 24397 7361 24409 7395
rect 24443 7361 24455 7395
rect 24397 7355 24455 7361
rect 24486 7352 24492 7404
rect 24544 7392 24550 7404
rect 24857 7395 24915 7401
rect 24857 7392 24869 7395
rect 24544 7364 24869 7392
rect 24544 7352 24550 7364
rect 24857 7361 24869 7364
rect 24903 7361 24915 7395
rect 24857 7355 24915 7361
rect 24949 7395 25007 7401
rect 24949 7361 24961 7395
rect 24995 7361 25007 7395
rect 25056 7392 25084 7432
rect 25498 7420 25504 7472
rect 25556 7460 25562 7472
rect 25556 7432 25820 7460
rect 25556 7420 25562 7432
rect 25792 7401 25820 7432
rect 25866 7420 25872 7472
rect 25924 7460 25930 7472
rect 25924 7432 26832 7460
rect 25924 7420 25930 7432
rect 25409 7395 25467 7401
rect 25409 7392 25421 7395
rect 25056 7364 25421 7392
rect 24949 7355 25007 7361
rect 25409 7361 25421 7364
rect 25455 7361 25467 7395
rect 25409 7355 25467 7361
rect 25685 7395 25743 7401
rect 25685 7361 25697 7395
rect 25731 7361 25743 7395
rect 25685 7355 25743 7361
rect 25777 7395 25835 7401
rect 25777 7361 25789 7395
rect 25823 7361 25835 7395
rect 25777 7355 25835 7361
rect 24964 7324 24992 7355
rect 19444 7296 23152 7324
rect 23216 7296 24716 7324
rect 24964 7296 25544 7324
rect 23124 7268 23152 7296
rect 16776 7228 19656 7256
rect 12084 7188 12112 7216
rect 16298 7188 16304 7200
rect 12084 7160 16304 7188
rect 16298 7148 16304 7160
rect 16356 7148 16362 7200
rect 16669 7191 16727 7197
rect 16669 7157 16681 7191
rect 16715 7188 16727 7191
rect 17402 7188 17408 7200
rect 16715 7160 17408 7188
rect 16715 7157 16727 7160
rect 16669 7151 16727 7157
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 18782 7148 18788 7200
rect 18840 7148 18846 7200
rect 19242 7148 19248 7200
rect 19300 7188 19306 7200
rect 19521 7191 19579 7197
rect 19521 7188 19533 7191
rect 19300 7160 19533 7188
rect 19300 7148 19306 7160
rect 19521 7157 19533 7160
rect 19567 7157 19579 7191
rect 19628 7188 19656 7228
rect 20530 7216 20536 7268
rect 20588 7256 20594 7268
rect 21177 7259 21235 7265
rect 21177 7256 21189 7259
rect 20588 7228 21189 7256
rect 20588 7216 20594 7228
rect 21177 7225 21189 7228
rect 21223 7225 21235 7259
rect 21177 7219 21235 7225
rect 21910 7216 21916 7268
rect 21968 7256 21974 7268
rect 22649 7259 22707 7265
rect 22649 7256 22661 7259
rect 21968 7228 22661 7256
rect 21968 7216 21974 7228
rect 22649 7225 22661 7228
rect 22695 7225 22707 7259
rect 22649 7219 22707 7225
rect 23106 7216 23112 7268
rect 23164 7216 23170 7268
rect 24578 7216 24584 7268
rect 24636 7216 24642 7268
rect 24688 7265 24716 7296
rect 24673 7259 24731 7265
rect 24673 7225 24685 7259
rect 24719 7225 24731 7259
rect 24673 7219 24731 7225
rect 24762 7216 24768 7268
rect 24820 7256 24826 7268
rect 25516 7265 25544 7296
rect 25501 7259 25559 7265
rect 24820 7228 25268 7256
rect 24820 7216 24826 7228
rect 21085 7191 21143 7197
rect 21085 7188 21097 7191
rect 19628 7160 21097 7188
rect 19521 7151 19579 7157
rect 21085 7157 21097 7160
rect 21131 7157 21143 7191
rect 21085 7151 21143 7157
rect 21450 7148 21456 7200
rect 21508 7148 21514 7200
rect 21818 7148 21824 7200
rect 21876 7148 21882 7200
rect 22094 7148 22100 7200
rect 22152 7148 22158 7200
rect 22922 7148 22928 7200
rect 22980 7148 22986 7200
rect 23474 7148 23480 7200
rect 23532 7148 23538 7200
rect 24026 7148 24032 7200
rect 24084 7148 24090 7200
rect 25130 7148 25136 7200
rect 25188 7148 25194 7200
rect 25240 7188 25268 7228
rect 25501 7225 25513 7259
rect 25547 7225 25559 7259
rect 25501 7219 25559 7225
rect 25700 7188 25728 7355
rect 25958 7352 25964 7404
rect 26016 7392 26022 7404
rect 26804 7401 26832 7432
rect 26237 7395 26295 7401
rect 26237 7392 26249 7395
rect 26016 7364 26249 7392
rect 26016 7352 26022 7364
rect 26237 7361 26249 7364
rect 26283 7361 26295 7395
rect 26237 7355 26295 7361
rect 26513 7395 26571 7401
rect 26513 7361 26525 7395
rect 26559 7361 26571 7395
rect 26513 7355 26571 7361
rect 26789 7395 26847 7401
rect 26789 7361 26801 7395
rect 26835 7361 26847 7395
rect 26896 7392 26924 7500
rect 27062 7488 27068 7540
rect 27120 7528 27126 7540
rect 27801 7531 27859 7537
rect 27801 7528 27813 7531
rect 27120 7500 27813 7528
rect 27120 7488 27126 7500
rect 27801 7497 27813 7500
rect 27847 7497 27859 7531
rect 27801 7491 27859 7497
rect 28350 7488 28356 7540
rect 28408 7528 28414 7540
rect 28408 7500 29408 7528
rect 28408 7488 28414 7500
rect 26970 7420 26976 7472
rect 27028 7460 27034 7472
rect 27028 7432 27752 7460
rect 27028 7420 27034 7432
rect 27724 7401 27752 7432
rect 27890 7420 27896 7472
rect 27948 7460 27954 7472
rect 27948 7432 28856 7460
rect 27948 7420 27954 7432
rect 27157 7395 27215 7401
rect 27157 7392 27169 7395
rect 26896 7364 27169 7392
rect 26789 7355 26847 7361
rect 27157 7361 27169 7364
rect 27203 7361 27215 7395
rect 27157 7355 27215 7361
rect 27433 7395 27491 7401
rect 27433 7361 27445 7395
rect 27479 7361 27491 7395
rect 27433 7355 27491 7361
rect 27709 7395 27767 7401
rect 27709 7361 27721 7395
rect 27755 7361 27767 7395
rect 27709 7355 27767 7361
rect 27985 7395 28043 7401
rect 27985 7361 27997 7395
rect 28031 7361 28043 7395
rect 27985 7355 28043 7361
rect 28261 7395 28319 7401
rect 28261 7361 28273 7395
rect 28307 7392 28319 7395
rect 28442 7392 28448 7404
rect 28307 7364 28448 7392
rect 28307 7361 28319 7364
rect 28261 7355 28319 7361
rect 25866 7284 25872 7336
rect 25924 7324 25930 7336
rect 26528 7324 26556 7355
rect 25924 7296 26556 7324
rect 25924 7284 25930 7296
rect 26694 7284 26700 7336
rect 26752 7324 26758 7336
rect 27448 7324 27476 7355
rect 26752 7296 27476 7324
rect 26752 7284 26758 7296
rect 27522 7284 27528 7336
rect 27580 7324 27586 7336
rect 28000 7324 28028 7355
rect 28442 7352 28448 7364
rect 28500 7352 28506 7404
rect 28534 7352 28540 7404
rect 28592 7352 28598 7404
rect 28828 7401 28856 7432
rect 29380 7401 29408 7500
rect 29454 7488 29460 7540
rect 29512 7528 29518 7540
rect 29512 7500 30420 7528
rect 29512 7488 29518 7500
rect 28813 7395 28871 7401
rect 28813 7361 28825 7395
rect 28859 7361 28871 7395
rect 28813 7355 28871 7361
rect 29089 7395 29147 7401
rect 29089 7361 29101 7395
rect 29135 7361 29147 7395
rect 29089 7355 29147 7361
rect 29365 7395 29423 7401
rect 29365 7361 29377 7395
rect 29411 7361 29423 7395
rect 29365 7355 29423 7361
rect 27580 7296 28028 7324
rect 27580 7284 27586 7296
rect 28350 7284 28356 7336
rect 28408 7324 28414 7336
rect 29104 7324 29132 7355
rect 29730 7352 29736 7404
rect 29788 7352 29794 7404
rect 30009 7395 30067 7401
rect 30009 7361 30021 7395
rect 30055 7361 30067 7395
rect 30009 7355 30067 7361
rect 28408 7296 29132 7324
rect 28408 7284 28414 7296
rect 26973 7259 27031 7265
rect 26973 7256 26985 7259
rect 25884 7228 26985 7256
rect 25884 7200 25912 7228
rect 26973 7225 26985 7228
rect 27019 7225 27031 7259
rect 26973 7219 27031 7225
rect 27430 7216 27436 7268
rect 27488 7256 27494 7268
rect 28077 7259 28135 7265
rect 28077 7256 28089 7259
rect 27488 7228 28089 7256
rect 27488 7216 27494 7228
rect 28077 7225 28089 7228
rect 28123 7225 28135 7259
rect 28077 7219 28135 7225
rect 28810 7216 28816 7268
rect 28868 7256 28874 7268
rect 29181 7259 29239 7265
rect 29181 7256 29193 7259
rect 28868 7228 29193 7256
rect 28868 7216 28874 7228
rect 29181 7225 29193 7228
rect 29227 7225 29239 7259
rect 30024 7256 30052 7355
rect 30282 7352 30288 7404
rect 30340 7352 30346 7404
rect 30392 7392 30420 7500
rect 30466 7488 30472 7540
rect 30524 7528 30530 7540
rect 30524 7500 31248 7528
rect 30524 7488 30530 7500
rect 30561 7395 30619 7401
rect 30561 7392 30573 7395
rect 30392 7364 30573 7392
rect 30561 7361 30573 7364
rect 30607 7361 30619 7395
rect 30561 7355 30619 7361
rect 30653 7395 30711 7401
rect 30653 7361 30665 7395
rect 30699 7392 30711 7395
rect 30742 7392 30748 7404
rect 30699 7364 30748 7392
rect 30699 7361 30711 7364
rect 30653 7355 30711 7361
rect 30742 7352 30748 7364
rect 30800 7352 30806 7404
rect 31220 7401 31248 7500
rect 31386 7488 31392 7540
rect 31444 7488 31450 7540
rect 31478 7488 31484 7540
rect 31536 7528 31542 7540
rect 31941 7531 31999 7537
rect 31941 7528 31953 7531
rect 31536 7500 31953 7528
rect 31536 7488 31542 7500
rect 31941 7497 31953 7500
rect 31987 7497 31999 7531
rect 31941 7491 31999 7497
rect 32490 7488 32496 7540
rect 32548 7528 32554 7540
rect 33413 7531 33471 7537
rect 32548 7500 33272 7528
rect 32548 7488 32554 7500
rect 31294 7420 31300 7472
rect 31352 7460 31358 7472
rect 31352 7432 32168 7460
rect 31352 7420 31358 7432
rect 30929 7395 30987 7401
rect 30929 7361 30941 7395
rect 30975 7361 30987 7395
rect 30929 7355 30987 7361
rect 31205 7395 31263 7401
rect 31205 7361 31217 7395
rect 31251 7361 31263 7395
rect 31205 7355 31263 7361
rect 30190 7284 30196 7336
rect 30248 7324 30254 7336
rect 30944 7324 30972 7355
rect 31478 7352 31484 7404
rect 31536 7352 31542 7404
rect 32140 7401 32168 7432
rect 32214 7420 32220 7472
rect 32272 7460 32278 7472
rect 32272 7432 32996 7460
rect 32272 7420 32278 7432
rect 32968 7401 32996 7432
rect 33244 7401 33272 7500
rect 33413 7497 33425 7531
rect 33459 7528 33471 7531
rect 33502 7528 33508 7540
rect 33459 7500 33508 7528
rect 33459 7497 33471 7500
rect 33413 7491 33471 7497
rect 33502 7488 33508 7500
rect 33560 7488 33566 7540
rect 33686 7488 33692 7540
rect 33744 7488 33750 7540
rect 33870 7488 33876 7540
rect 33928 7528 33934 7540
rect 34149 7531 34207 7537
rect 34149 7528 34161 7531
rect 33928 7500 34161 7528
rect 33928 7488 33934 7500
rect 34149 7497 34161 7500
rect 34195 7497 34207 7531
rect 34149 7491 34207 7497
rect 34606 7488 34612 7540
rect 34664 7528 34670 7540
rect 34885 7531 34943 7537
rect 34885 7528 34897 7531
rect 34664 7500 34897 7528
rect 34664 7488 34670 7500
rect 34885 7497 34897 7500
rect 34931 7497 34943 7531
rect 34885 7491 34943 7497
rect 35437 7531 35495 7537
rect 35437 7497 35449 7531
rect 35483 7497 35495 7531
rect 35437 7491 35495 7497
rect 34698 7420 34704 7472
rect 34756 7460 34762 7472
rect 35452 7460 35480 7491
rect 35710 7488 35716 7540
rect 35768 7528 35774 7540
rect 36541 7531 36599 7537
rect 36541 7528 36553 7531
rect 35768 7500 36553 7528
rect 35768 7488 35774 7500
rect 36541 7497 36553 7500
rect 36587 7497 36599 7531
rect 36541 7491 36599 7497
rect 37090 7488 37096 7540
rect 37148 7528 37154 7540
rect 38013 7531 38071 7537
rect 38013 7528 38025 7531
rect 37148 7500 38025 7528
rect 37148 7488 37154 7500
rect 38013 7497 38025 7500
rect 38059 7497 38071 7531
rect 38013 7491 38071 7497
rect 39114 7488 39120 7540
rect 39172 7528 39178 7540
rect 40037 7531 40095 7537
rect 40037 7528 40049 7531
rect 39172 7500 40049 7528
rect 39172 7488 39178 7500
rect 40037 7497 40049 7500
rect 40083 7497 40095 7531
rect 41233 7531 41291 7537
rect 41233 7528 41245 7531
rect 40037 7491 40095 7497
rect 40512 7500 41245 7528
rect 34756 7432 35480 7460
rect 34756 7420 34762 7432
rect 36170 7420 36176 7472
rect 36228 7460 36234 7472
rect 36449 7463 36507 7469
rect 36449 7460 36461 7463
rect 36228 7432 36461 7460
rect 36228 7420 36234 7432
rect 36449 7429 36461 7432
rect 36495 7429 36507 7463
rect 36449 7423 36507 7429
rect 36814 7420 36820 7472
rect 36872 7460 36878 7472
rect 40512 7469 40540 7500
rect 41233 7497 41245 7500
rect 41279 7497 41291 7531
rect 41233 7491 41291 7497
rect 40497 7463 40555 7469
rect 36872 7432 38516 7460
rect 36872 7420 36878 7432
rect 31757 7395 31815 7401
rect 31757 7361 31769 7395
rect 31803 7361 31815 7395
rect 31757 7355 31815 7361
rect 32125 7395 32183 7401
rect 32125 7361 32137 7395
rect 32171 7361 32183 7395
rect 32125 7355 32183 7361
rect 32401 7395 32459 7401
rect 32677 7396 32735 7401
rect 32401 7361 32413 7395
rect 32447 7361 32459 7395
rect 32600 7395 32735 7396
rect 32600 7392 32689 7395
rect 32401 7355 32459 7361
rect 32508 7368 32689 7392
rect 32508 7364 32628 7368
rect 30248 7296 30972 7324
rect 30248 7284 30254 7296
rect 31018 7284 31024 7336
rect 31076 7324 31082 7336
rect 31772 7324 31800 7355
rect 31076 7296 31800 7324
rect 31076 7284 31082 7296
rect 31846 7284 31852 7336
rect 31904 7324 31910 7336
rect 32416 7324 32444 7355
rect 31904 7296 32444 7324
rect 31904 7284 31910 7296
rect 29181 7219 29239 7225
rect 29288 7228 30052 7256
rect 25240 7160 25728 7188
rect 25866 7148 25872 7200
rect 25924 7148 25930 7200
rect 26050 7148 26056 7200
rect 26108 7148 26114 7200
rect 26142 7148 26148 7200
rect 26200 7188 26206 7200
rect 26329 7191 26387 7197
rect 26329 7188 26341 7191
rect 26200 7160 26341 7188
rect 26200 7148 26206 7160
rect 26329 7157 26341 7160
rect 26375 7157 26387 7191
rect 26329 7151 26387 7157
rect 26602 7148 26608 7200
rect 26660 7148 26666 7200
rect 27246 7148 27252 7200
rect 27304 7148 27310 7200
rect 27522 7148 27528 7200
rect 27580 7148 27586 7200
rect 28350 7148 28356 7200
rect 28408 7148 28414 7200
rect 28626 7148 28632 7200
rect 28684 7148 28690 7200
rect 28902 7148 28908 7200
rect 28960 7148 28966 7200
rect 29086 7148 29092 7200
rect 29144 7188 29150 7200
rect 29288 7188 29316 7228
rect 30558 7216 30564 7268
rect 30616 7256 30622 7268
rect 31478 7256 31484 7268
rect 30616 7228 31484 7256
rect 30616 7216 30622 7228
rect 31478 7216 31484 7228
rect 31536 7216 31542 7268
rect 31938 7216 31944 7268
rect 31996 7256 32002 7268
rect 32508 7256 32536 7364
rect 32677 7361 32689 7368
rect 32723 7361 32735 7395
rect 32677 7355 32735 7361
rect 32953 7395 33011 7401
rect 32953 7361 32965 7395
rect 32999 7361 33011 7395
rect 32953 7355 33011 7361
rect 33229 7395 33287 7401
rect 33229 7361 33241 7395
rect 33275 7361 33287 7395
rect 33229 7355 33287 7361
rect 33505 7395 33563 7401
rect 33505 7361 33517 7395
rect 33551 7361 33563 7395
rect 33505 7355 33563 7361
rect 32582 7284 32588 7336
rect 32640 7284 32646 7336
rect 32858 7284 32864 7336
rect 32916 7324 32922 7336
rect 33520 7324 33548 7355
rect 33686 7352 33692 7404
rect 33744 7392 33750 7404
rect 34057 7395 34115 7401
rect 34057 7392 34069 7395
rect 33744 7364 34069 7392
rect 33744 7352 33750 7364
rect 34057 7361 34069 7364
rect 34103 7361 34115 7395
rect 34057 7355 34115 7361
rect 34790 7352 34796 7404
rect 34848 7352 34854 7404
rect 35342 7352 35348 7404
rect 35400 7352 35406 7404
rect 35894 7352 35900 7404
rect 35952 7352 35958 7404
rect 37093 7395 37151 7401
rect 37093 7361 37105 7395
rect 37139 7361 37151 7395
rect 37093 7355 37151 7361
rect 37369 7395 37427 7401
rect 37369 7361 37381 7395
rect 37415 7392 37427 7395
rect 37550 7392 37556 7404
rect 37415 7364 37556 7392
rect 37415 7361 37427 7364
rect 37369 7355 37427 7361
rect 32916 7296 33548 7324
rect 32916 7284 32922 7296
rect 35710 7284 35716 7336
rect 35768 7324 35774 7336
rect 37108 7324 37136 7355
rect 37550 7352 37556 7364
rect 37608 7352 37614 7404
rect 37918 7352 37924 7404
rect 37976 7352 37982 7404
rect 38488 7401 38516 7432
rect 40497 7429 40509 7463
rect 40543 7429 40555 7463
rect 40497 7423 40555 7429
rect 38473 7395 38531 7401
rect 38473 7361 38485 7395
rect 38519 7361 38531 7395
rect 38473 7355 38531 7361
rect 39022 7352 39028 7404
rect 39080 7352 39086 7404
rect 39666 7352 39672 7404
rect 39724 7352 39730 7404
rect 39945 7395 40003 7401
rect 39945 7361 39957 7395
rect 39991 7361 40003 7395
rect 39945 7355 40003 7361
rect 41141 7395 41199 7401
rect 41141 7361 41153 7395
rect 41187 7361 41199 7395
rect 41141 7355 41199 7361
rect 35768 7296 37136 7324
rect 35768 7284 35774 7296
rect 37826 7284 37832 7336
rect 37884 7324 37890 7336
rect 39960 7324 39988 7355
rect 37884 7296 39988 7324
rect 41156 7324 41184 7355
rect 41414 7352 41420 7404
rect 41472 7352 41478 7404
rect 43346 7324 43352 7336
rect 41156 7296 43352 7324
rect 37884 7284 37890 7296
rect 43346 7284 43352 7296
rect 43404 7284 43410 7336
rect 31996 7228 32536 7256
rect 32600 7256 32628 7284
rect 33137 7259 33195 7265
rect 33137 7256 33149 7259
rect 32600 7228 33149 7256
rect 31996 7216 32002 7228
rect 33137 7225 33149 7228
rect 33183 7225 33195 7259
rect 33137 7219 33195 7225
rect 36538 7216 36544 7268
rect 36596 7256 36602 7268
rect 36596 7228 37504 7256
rect 36596 7216 36602 7228
rect 29144 7160 29316 7188
rect 29144 7148 29150 7160
rect 29546 7148 29552 7200
rect 29604 7148 29610 7200
rect 29822 7148 29828 7200
rect 29880 7148 29886 7200
rect 30098 7148 30104 7200
rect 30156 7148 30162 7200
rect 30374 7148 30380 7200
rect 30432 7148 30438 7200
rect 30650 7148 30656 7200
rect 30708 7188 30714 7200
rect 30837 7191 30895 7197
rect 30837 7188 30849 7191
rect 30708 7160 30849 7188
rect 30708 7148 30714 7160
rect 30837 7157 30849 7160
rect 30883 7157 30895 7191
rect 30837 7151 30895 7157
rect 30926 7148 30932 7200
rect 30984 7188 30990 7200
rect 31113 7191 31171 7197
rect 31113 7188 31125 7191
rect 30984 7160 31125 7188
rect 30984 7148 30990 7160
rect 31113 7157 31125 7160
rect 31159 7157 31171 7191
rect 31113 7151 31171 7157
rect 31202 7148 31208 7200
rect 31260 7188 31266 7200
rect 31665 7191 31723 7197
rect 31665 7188 31677 7191
rect 31260 7160 31677 7188
rect 31260 7148 31266 7160
rect 31665 7157 31677 7160
rect 31711 7157 31723 7191
rect 31665 7151 31723 7157
rect 32306 7148 32312 7200
rect 32364 7148 32370 7200
rect 32582 7148 32588 7200
rect 32640 7148 32646 7200
rect 32674 7148 32680 7200
rect 32732 7188 32738 7200
rect 32861 7191 32919 7197
rect 32861 7188 32873 7191
rect 32732 7160 32873 7188
rect 32732 7148 32738 7160
rect 32861 7157 32873 7160
rect 32907 7157 32919 7191
rect 32861 7151 32919 7157
rect 35158 7148 35164 7200
rect 35216 7188 35222 7200
rect 35989 7191 36047 7197
rect 35989 7188 36001 7191
rect 35216 7160 36001 7188
rect 35216 7148 35222 7160
rect 35989 7157 36001 7160
rect 36035 7157 36047 7191
rect 35989 7151 36047 7157
rect 36906 7148 36912 7200
rect 36964 7148 36970 7200
rect 37476 7197 37504 7228
rect 39574 7216 39580 7268
rect 39632 7256 39638 7268
rect 39632 7228 40632 7256
rect 39632 7216 39638 7228
rect 37461 7191 37519 7197
rect 37461 7157 37473 7191
rect 37507 7157 37519 7191
rect 37461 7151 37519 7157
rect 38746 7148 38752 7200
rect 38804 7148 38810 7200
rect 39114 7148 39120 7200
rect 39172 7148 39178 7200
rect 39482 7148 39488 7200
rect 39540 7148 39546 7200
rect 40604 7197 40632 7228
rect 40589 7191 40647 7197
rect 40589 7157 40601 7191
rect 40635 7157 40647 7191
rect 40589 7151 40647 7157
rect 40954 7148 40960 7200
rect 41012 7148 41018 7200
rect 1104 7098 43884 7120
rect 1104 7046 6297 7098
rect 6349 7046 6361 7098
rect 6413 7046 6425 7098
rect 6477 7046 6489 7098
rect 6541 7046 6553 7098
rect 6605 7046 16991 7098
rect 17043 7046 17055 7098
rect 17107 7046 17119 7098
rect 17171 7046 17183 7098
rect 17235 7046 17247 7098
rect 17299 7046 27685 7098
rect 27737 7046 27749 7098
rect 27801 7046 27813 7098
rect 27865 7046 27877 7098
rect 27929 7046 27941 7098
rect 27993 7046 38379 7098
rect 38431 7046 38443 7098
rect 38495 7046 38507 7098
rect 38559 7046 38571 7098
rect 38623 7046 38635 7098
rect 38687 7046 43884 7098
rect 1104 7024 43884 7046
rect 5166 6944 5172 6996
rect 5224 6944 5230 6996
rect 5718 6944 5724 6996
rect 5776 6944 5782 6996
rect 6822 6944 6828 6996
rect 6880 6944 6886 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 12250 6984 12256 6996
rect 7340 6956 12256 6984
rect 7340 6944 7346 6956
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 13078 6944 13084 6996
rect 13136 6944 13142 6996
rect 13630 6944 13636 6996
rect 13688 6944 13694 6996
rect 14182 6944 14188 6996
rect 14240 6944 14246 6996
rect 14550 6944 14556 6996
rect 14608 6944 14614 6996
rect 16298 6944 16304 6996
rect 16356 6984 16362 6996
rect 17954 6984 17960 6996
rect 16356 6956 17960 6984
rect 16356 6944 16362 6956
rect 17954 6944 17960 6956
rect 18012 6944 18018 6996
rect 18877 6987 18935 6993
rect 18877 6953 18889 6987
rect 18923 6984 18935 6987
rect 19978 6984 19984 6996
rect 18923 6956 19984 6984
rect 18923 6953 18935 6956
rect 18877 6947 18935 6953
rect 19978 6944 19984 6956
rect 20036 6944 20042 6996
rect 20438 6944 20444 6996
rect 20496 6984 20502 6996
rect 21450 6984 21456 6996
rect 20496 6956 21456 6984
rect 20496 6944 20502 6956
rect 21450 6944 21456 6956
rect 21508 6944 21514 6996
rect 26142 6984 26148 6996
rect 25148 6956 26148 6984
rect 9398 6916 9404 6928
rect 9232 6888 9404 6916
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 7561 6851 7619 6857
rect 7561 6848 7573 6851
rect 7156 6820 7573 6848
rect 7156 6808 7162 6820
rect 7561 6817 7573 6820
rect 7607 6817 7619 6851
rect 7561 6811 7619 6817
rect 7650 6808 7656 6860
rect 7708 6848 7714 6860
rect 8113 6851 8171 6857
rect 8113 6848 8125 6851
rect 7708 6820 8125 6848
rect 7708 6808 7714 6820
rect 8113 6817 8125 6820
rect 8159 6817 8171 6851
rect 8113 6811 8171 6817
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 8665 6851 8723 6857
rect 8665 6848 8677 6851
rect 8260 6820 8677 6848
rect 8260 6808 8266 6820
rect 8665 6817 8677 6820
rect 8711 6817 8723 6851
rect 8665 6811 8723 6817
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 6638 6780 6644 6792
rect 6227 6752 6644 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6780 6791 6783
rect 7742 6780 7748 6792
rect 6779 6752 7748 6780
rect 6779 6749 6791 6752
rect 6733 6743 6791 6749
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6780 7895 6783
rect 9232 6780 9260 6888
rect 9398 6876 9404 6888
rect 9456 6876 9462 6928
rect 14200 6916 14228 6944
rect 20254 6916 20260 6928
rect 14200 6888 20260 6916
rect 20254 6876 20260 6888
rect 20312 6876 20318 6928
rect 20346 6876 20352 6928
rect 20404 6916 20410 6928
rect 21729 6919 21787 6925
rect 21729 6916 21741 6919
rect 20404 6888 21741 6916
rect 20404 6876 20410 6888
rect 21729 6885 21741 6888
rect 21775 6885 21787 6919
rect 21729 6879 21787 6885
rect 9585 6851 9643 6857
rect 9585 6817 9597 6851
rect 9631 6848 9643 6851
rect 10134 6848 10140 6860
rect 9631 6820 10140 6848
rect 9631 6817 9643 6820
rect 9585 6811 9643 6817
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 10502 6808 10508 6860
rect 10560 6808 10566 6860
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 11020 6820 11069 6848
rect 11020 6808 11026 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 11606 6808 11612 6860
rect 11664 6808 11670 6860
rect 12342 6808 12348 6860
rect 12400 6848 12406 6860
rect 12713 6851 12771 6857
rect 12713 6848 12725 6851
rect 12400 6820 12725 6848
rect 12400 6808 12406 6820
rect 12713 6817 12725 6820
rect 12759 6817 12771 6851
rect 12713 6811 12771 6817
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 14884 6820 15301 6848
rect 14884 6808 14890 6820
rect 15289 6817 15301 6820
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 15841 6851 15899 6857
rect 15841 6848 15853 6851
rect 15436 6820 15853 6848
rect 15436 6808 15442 6820
rect 15841 6817 15853 6820
rect 15887 6817 15899 6851
rect 15841 6811 15899 6817
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 16393 6851 16451 6857
rect 16393 6848 16405 6851
rect 15988 6820 16405 6848
rect 15988 6808 15994 6820
rect 16393 6817 16405 6820
rect 16439 6817 16451 6851
rect 16393 6811 16451 6817
rect 16482 6808 16488 6860
rect 16540 6848 16546 6860
rect 16945 6851 17003 6857
rect 16945 6848 16957 6851
rect 16540 6820 16957 6848
rect 16540 6808 16546 6820
rect 16945 6817 16957 6820
rect 16991 6817 17003 6851
rect 16945 6811 17003 6817
rect 17034 6808 17040 6860
rect 17092 6848 17098 6860
rect 17497 6851 17555 6857
rect 17497 6848 17509 6851
rect 17092 6820 17509 6848
rect 17092 6808 17098 6820
rect 17497 6817 17509 6820
rect 17543 6817 17555 6851
rect 17497 6811 17555 6817
rect 17586 6808 17592 6860
rect 17644 6848 17650 6860
rect 18049 6851 18107 6857
rect 18049 6848 18061 6851
rect 17644 6820 18061 6848
rect 17644 6808 17650 6820
rect 18049 6817 18061 6820
rect 18095 6817 18107 6851
rect 18049 6811 18107 6817
rect 18138 6808 18144 6860
rect 18196 6848 18202 6860
rect 18601 6851 18659 6857
rect 18601 6848 18613 6851
rect 18196 6820 18613 6848
rect 18196 6808 18202 6820
rect 18601 6817 18613 6820
rect 18647 6817 18659 6851
rect 22094 6848 22100 6860
rect 18601 6811 18659 6817
rect 18708 6820 20392 6848
rect 7883 6752 9260 6780
rect 9291 6783 9349 6789
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 9291 6749 9303 6783
rect 9337 6780 9349 6783
rect 9398 6780 9404 6792
rect 9337 6752 9404 6780
rect 9337 6749 9349 6752
rect 9291 6743 9349 6749
rect 9398 6740 9404 6752
rect 9456 6740 9462 6792
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 11146 6780 11152 6792
rect 9548 6752 11152 6780
rect 9548 6740 9554 6752
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6780 12311 6783
rect 12618 6780 12624 6792
rect 12299 6752 12624 6780
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 14182 6780 14188 6792
rect 12912 6752 14188 6780
rect 5077 6715 5135 6721
rect 5077 6681 5089 6715
rect 5123 6681 5135 6715
rect 5077 6675 5135 6681
rect 5092 6644 5120 6675
rect 5626 6672 5632 6724
rect 5684 6672 5690 6724
rect 7285 6715 7343 6721
rect 7285 6681 7297 6715
rect 7331 6681 7343 6715
rect 7285 6675 7343 6681
rect 8389 6715 8447 6721
rect 8389 6681 8401 6715
rect 8435 6712 8447 6715
rect 10229 6715 10287 6721
rect 8435 6684 10180 6712
rect 8435 6681 8447 6684
rect 8389 6675 8447 6681
rect 6086 6644 6092 6656
rect 5092 6616 6092 6644
rect 6086 6604 6092 6616
rect 6144 6604 6150 6656
rect 6270 6604 6276 6656
rect 6328 6604 6334 6656
rect 7300 6644 7328 6675
rect 9858 6644 9864 6656
rect 7300 6616 9864 6644
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 10152 6644 10180 6684
rect 10229 6681 10241 6715
rect 10275 6712 10287 6715
rect 10686 6712 10692 6724
rect 10275 6684 10692 6712
rect 10275 6681 10287 6684
rect 10229 6675 10287 6681
rect 10686 6672 10692 6684
rect 10744 6672 10750 6724
rect 10778 6672 10784 6724
rect 10836 6672 10842 6724
rect 11330 6672 11336 6724
rect 11388 6672 11394 6724
rect 11885 6715 11943 6721
rect 11885 6681 11897 6715
rect 11931 6712 11943 6715
rect 12437 6715 12495 6721
rect 11931 6684 12204 6712
rect 11931 6681 11943 6684
rect 11885 6675 11943 6681
rect 12066 6644 12072 6656
rect 10152 6616 12072 6644
rect 12066 6604 12072 6616
rect 12124 6604 12130 6656
rect 12176 6644 12204 6684
rect 12437 6681 12449 6715
rect 12483 6712 12495 6715
rect 12912 6712 12940 6752
rect 14182 6740 14188 6752
rect 14240 6740 14246 6792
rect 14274 6740 14280 6792
rect 14332 6740 14338 6792
rect 15565 6783 15623 6789
rect 15565 6780 15577 6783
rect 14844 6752 15577 6780
rect 12483 6684 12940 6712
rect 12483 6681 12495 6684
rect 12437 6675 12495 6681
rect 12986 6672 12992 6724
rect 13044 6672 13050 6724
rect 13541 6715 13599 6721
rect 13541 6681 13553 6715
rect 13587 6712 13599 6715
rect 13906 6712 13912 6724
rect 13587 6684 13912 6712
rect 13587 6681 13599 6684
rect 13541 6675 13599 6681
rect 13906 6672 13912 6684
rect 13964 6672 13970 6724
rect 14461 6715 14519 6721
rect 14461 6681 14473 6715
rect 14507 6712 14519 6715
rect 14734 6712 14740 6724
rect 14507 6684 14740 6712
rect 14507 6681 14519 6684
rect 14461 6675 14519 6681
rect 14734 6672 14740 6684
rect 14792 6672 14798 6724
rect 13722 6644 13728 6656
rect 12176 6616 13728 6644
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 14093 6647 14151 6653
rect 14093 6613 14105 6647
rect 14139 6644 14151 6647
rect 14844 6644 14872 6752
rect 15565 6749 15577 6752
rect 15611 6749 15623 6783
rect 15565 6743 15623 6749
rect 16298 6740 16304 6792
rect 16356 6780 16362 6792
rect 18708 6780 18736 6820
rect 16356 6752 18736 6780
rect 16356 6740 16362 6752
rect 19058 6740 19064 6792
rect 19116 6740 19122 6792
rect 19334 6740 19340 6792
rect 19392 6740 19398 6792
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 19886 6740 19892 6792
rect 19944 6740 19950 6792
rect 20162 6740 20168 6792
rect 20220 6740 20226 6792
rect 15010 6672 15016 6724
rect 15068 6672 15074 6724
rect 15286 6672 15292 6724
rect 15344 6712 15350 6724
rect 16117 6715 16175 6721
rect 16117 6712 16129 6715
rect 15344 6684 16129 6712
rect 15344 6672 15350 6684
rect 16117 6681 16129 6684
rect 16163 6681 16175 6715
rect 16117 6675 16175 6681
rect 16666 6672 16672 6724
rect 16724 6672 16730 6724
rect 17218 6672 17224 6724
rect 17276 6672 17282 6724
rect 17402 6672 17408 6724
rect 17460 6712 17466 6724
rect 17773 6715 17831 6721
rect 17773 6712 17785 6715
rect 17460 6684 17785 6712
rect 17460 6672 17466 6684
rect 17773 6681 17785 6684
rect 17819 6681 17831 6715
rect 17773 6675 17831 6681
rect 18322 6672 18328 6724
rect 18380 6672 18386 6724
rect 18414 6672 18420 6724
rect 18472 6712 18478 6724
rect 18472 6684 20116 6712
rect 18472 6672 18478 6684
rect 14139 6616 14872 6644
rect 14139 6613 14151 6616
rect 14093 6607 14151 6613
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 19426 6644 19432 6656
rect 18564 6616 19432 6644
rect 18564 6604 18570 6616
rect 19426 6604 19432 6616
rect 19484 6604 19490 6656
rect 19518 6604 19524 6656
rect 19576 6604 19582 6656
rect 19794 6604 19800 6656
rect 19852 6604 19858 6656
rect 20088 6653 20116 6684
rect 20364 6653 20392 6820
rect 21008 6820 22100 6848
rect 20441 6783 20499 6789
rect 20441 6749 20453 6783
rect 20487 6780 20499 6783
rect 20530 6780 20536 6792
rect 20487 6752 20536 6780
rect 20487 6749 20499 6752
rect 20441 6743 20499 6749
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 20622 6740 20628 6792
rect 20680 6780 20686 6792
rect 21008 6789 21036 6820
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 20717 6783 20775 6789
rect 20717 6780 20729 6783
rect 20680 6752 20729 6780
rect 20680 6740 20686 6752
rect 20717 6749 20729 6752
rect 20763 6749 20775 6783
rect 20717 6743 20775 6749
rect 20993 6783 21051 6789
rect 20993 6749 21005 6783
rect 21039 6749 21051 6783
rect 20993 6743 21051 6749
rect 21269 6783 21327 6789
rect 21269 6749 21281 6783
rect 21315 6749 21327 6783
rect 21269 6743 21327 6749
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6780 21603 6783
rect 21818 6780 21824 6792
rect 21591 6752 21824 6780
rect 21591 6749 21603 6752
rect 21545 6743 21603 6749
rect 21284 6712 21312 6743
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 22002 6740 22008 6792
rect 22060 6780 22066 6792
rect 22060 6752 22692 6780
rect 22060 6740 22066 6752
rect 22664 6712 22692 6752
rect 22830 6740 22836 6792
rect 22888 6740 22894 6792
rect 23017 6783 23075 6789
rect 23017 6749 23029 6783
rect 23063 6780 23075 6783
rect 24026 6780 24032 6792
rect 23063 6752 24032 6780
rect 23063 6749 23075 6752
rect 23017 6743 23075 6749
rect 24026 6740 24032 6752
rect 24084 6740 24090 6792
rect 25148 6789 25176 6956
rect 26142 6944 26148 6956
rect 26200 6944 26206 6996
rect 26418 6944 26424 6996
rect 26476 6944 26482 6996
rect 26602 6944 26608 6996
rect 26660 6944 26666 6996
rect 27246 6944 27252 6996
rect 27304 6944 27310 6996
rect 28350 6944 28356 6996
rect 28408 6944 28414 6996
rect 28626 6944 28632 6996
rect 28684 6944 28690 6996
rect 36906 6944 36912 6996
rect 36964 6984 36970 6996
rect 36964 6956 39344 6984
rect 36964 6944 36970 6956
rect 26620 6916 26648 6944
rect 25424 6888 26648 6916
rect 25424 6789 25452 6888
rect 27264 6848 27292 6944
rect 28368 6916 28396 6944
rect 26252 6820 27292 6848
rect 27816 6888 28396 6916
rect 24857 6783 24915 6789
rect 24857 6749 24869 6783
rect 24903 6749 24915 6783
rect 24857 6743 24915 6749
rect 25133 6783 25191 6789
rect 25133 6749 25145 6783
rect 25179 6749 25191 6783
rect 25133 6743 25191 6749
rect 25409 6783 25467 6789
rect 25409 6749 25421 6783
rect 25455 6749 25467 6783
rect 25409 6743 25467 6749
rect 24872 6712 24900 6743
rect 26050 6740 26056 6792
rect 26108 6740 26114 6792
rect 26252 6789 26280 6820
rect 26237 6783 26295 6789
rect 26237 6749 26249 6783
rect 26283 6749 26295 6783
rect 26237 6743 26295 6749
rect 26513 6783 26571 6789
rect 26513 6749 26525 6783
rect 26559 6749 26571 6783
rect 26513 6743 26571 6749
rect 26789 6783 26847 6789
rect 26789 6749 26801 6783
rect 26835 6780 26847 6783
rect 27062 6780 27068 6792
rect 26835 6752 27068 6780
rect 26835 6749 26847 6752
rect 26789 6743 26847 6749
rect 26068 6712 26096 6740
rect 21284 6684 22094 6712
rect 22664 6684 23244 6712
rect 24872 6684 26096 6712
rect 20073 6647 20131 6653
rect 20073 6613 20085 6647
rect 20119 6613 20131 6647
rect 20073 6607 20131 6613
rect 20349 6647 20407 6653
rect 20349 6613 20361 6647
rect 20395 6613 20407 6647
rect 20349 6607 20407 6613
rect 20622 6604 20628 6656
rect 20680 6604 20686 6656
rect 20898 6604 20904 6656
rect 20956 6604 20962 6656
rect 21174 6604 21180 6656
rect 21232 6604 21238 6656
rect 21266 6604 21272 6656
rect 21324 6644 21330 6656
rect 21453 6647 21511 6653
rect 21453 6644 21465 6647
rect 21324 6616 21465 6644
rect 21324 6604 21330 6616
rect 21453 6613 21465 6616
rect 21499 6613 21511 6647
rect 22066 6644 22094 6684
rect 23216 6653 23244 6684
rect 26142 6672 26148 6724
rect 26200 6712 26206 6724
rect 26528 6712 26556 6743
rect 27062 6740 27068 6752
rect 27120 6740 27126 6792
rect 27157 6783 27215 6789
rect 27157 6749 27169 6783
rect 27203 6780 27215 6783
rect 27430 6780 27436 6792
rect 27203 6752 27436 6780
rect 27203 6749 27215 6752
rect 27157 6743 27215 6749
rect 27430 6740 27436 6752
rect 27488 6740 27494 6792
rect 27525 6783 27583 6789
rect 27525 6749 27537 6783
rect 27571 6780 27583 6783
rect 27816 6780 27844 6888
rect 28644 6848 28672 6944
rect 38102 6876 38108 6928
rect 38160 6916 38166 6928
rect 38160 6888 38424 6916
rect 38160 6876 38166 6888
rect 27908 6820 28672 6848
rect 27908 6789 27936 6820
rect 33594 6808 33600 6860
rect 33652 6848 33658 6860
rect 33652 6820 34284 6848
rect 33652 6808 33658 6820
rect 27571 6752 27844 6780
rect 27893 6783 27951 6789
rect 27571 6749 27583 6752
rect 27525 6743 27583 6749
rect 27893 6749 27905 6783
rect 27939 6749 27951 6783
rect 27893 6743 27951 6749
rect 28261 6783 28319 6789
rect 28261 6749 28273 6783
rect 28307 6749 28319 6783
rect 28261 6743 28319 6749
rect 28721 6783 28779 6789
rect 28721 6749 28733 6783
rect 28767 6780 28779 6783
rect 28810 6780 28816 6792
rect 28767 6752 28816 6780
rect 28767 6749 28779 6752
rect 28721 6743 28779 6749
rect 28276 6712 28304 6743
rect 28810 6740 28816 6752
rect 28868 6740 28874 6792
rect 28902 6740 28908 6792
rect 28960 6740 28966 6792
rect 29181 6783 29239 6789
rect 29181 6749 29193 6783
rect 29227 6780 29239 6783
rect 29546 6780 29552 6792
rect 29227 6752 29552 6780
rect 29227 6749 29239 6752
rect 29181 6743 29239 6749
rect 29546 6740 29552 6752
rect 29604 6740 29610 6792
rect 29641 6783 29699 6789
rect 29641 6749 29653 6783
rect 29687 6780 29699 6783
rect 29822 6780 29828 6792
rect 29687 6752 29828 6780
rect 29687 6749 29699 6752
rect 29641 6743 29699 6749
rect 29822 6740 29828 6752
rect 29880 6740 29886 6792
rect 30009 6783 30067 6789
rect 30009 6749 30021 6783
rect 30055 6780 30067 6783
rect 30098 6780 30104 6792
rect 30055 6752 30104 6780
rect 30055 6749 30067 6752
rect 30009 6743 30067 6749
rect 30098 6740 30104 6752
rect 30156 6740 30162 6792
rect 30285 6783 30343 6789
rect 30285 6749 30297 6783
rect 30331 6780 30343 6783
rect 30374 6780 30380 6792
rect 30331 6752 30380 6780
rect 30331 6749 30343 6752
rect 30285 6743 30343 6749
rect 30374 6740 30380 6752
rect 30432 6740 30438 6792
rect 31202 6740 31208 6792
rect 31260 6740 31266 6792
rect 31754 6740 31760 6792
rect 31812 6780 31818 6792
rect 32585 6783 32643 6789
rect 32585 6780 32597 6783
rect 31812 6752 32597 6780
rect 31812 6740 31818 6752
rect 32585 6749 32597 6752
rect 32631 6749 32643 6783
rect 32585 6743 32643 6749
rect 32950 6740 32956 6792
rect 33008 6780 33014 6792
rect 33137 6783 33195 6789
rect 33137 6780 33149 6783
rect 33008 6752 33149 6780
rect 33008 6740 33014 6752
rect 33137 6749 33149 6752
rect 33183 6749 33195 6783
rect 33137 6743 33195 6749
rect 33410 6740 33416 6792
rect 33468 6740 33474 6792
rect 33686 6740 33692 6792
rect 33744 6740 33750 6792
rect 33870 6740 33876 6792
rect 33928 6740 33934 6792
rect 34054 6740 34060 6792
rect 34112 6780 34118 6792
rect 34256 6789 34284 6820
rect 35250 6808 35256 6860
rect 35308 6848 35314 6860
rect 35713 6851 35771 6857
rect 35713 6848 35725 6851
rect 35308 6820 35725 6848
rect 35308 6808 35314 6820
rect 35713 6817 35725 6820
rect 35759 6817 35771 6851
rect 35713 6811 35771 6817
rect 35802 6808 35808 6860
rect 35860 6848 35866 6860
rect 36265 6851 36323 6857
rect 36265 6848 36277 6851
rect 35860 6820 36277 6848
rect 35860 6808 35866 6820
rect 36265 6817 36277 6820
rect 36311 6817 36323 6851
rect 36265 6811 36323 6817
rect 37182 6808 37188 6860
rect 37240 6848 37246 6860
rect 37921 6851 37979 6857
rect 37921 6848 37933 6851
rect 37240 6820 37933 6848
rect 37240 6808 37246 6820
rect 37921 6817 37933 6820
rect 37967 6817 37979 6851
rect 38396 6848 38424 6888
rect 38562 6876 38568 6928
rect 38620 6916 38626 6928
rect 38930 6916 38936 6928
rect 38620 6888 38936 6916
rect 38620 6876 38626 6888
rect 38930 6876 38936 6888
rect 38988 6876 38994 6928
rect 39114 6848 39120 6860
rect 38396 6820 39120 6848
rect 37921 6811 37979 6817
rect 39114 6808 39120 6820
rect 39172 6808 39178 6860
rect 34149 6783 34207 6789
rect 34149 6780 34161 6783
rect 34112 6752 34161 6780
rect 34112 6740 34118 6752
rect 34149 6749 34161 6752
rect 34195 6749 34207 6783
rect 34149 6743 34207 6749
rect 34241 6783 34299 6789
rect 34241 6749 34253 6783
rect 34287 6749 34299 6783
rect 34241 6743 34299 6749
rect 34885 6783 34943 6789
rect 34885 6749 34897 6783
rect 34931 6749 34943 6783
rect 34885 6743 34943 6749
rect 28920 6712 28948 6740
rect 33704 6712 33732 6740
rect 34900 6712 34928 6743
rect 35158 6740 35164 6792
rect 35216 6740 35222 6792
rect 37458 6740 37464 6792
rect 37516 6780 37522 6792
rect 38654 6780 38660 6792
rect 37516 6752 38660 6780
rect 37516 6740 37522 6752
rect 38654 6740 38660 6752
rect 38712 6740 38718 6792
rect 39316 6789 39344 6956
rect 39850 6808 39856 6860
rect 39908 6848 39914 6860
rect 40773 6851 40831 6857
rect 40773 6848 40785 6851
rect 39908 6820 40785 6848
rect 39908 6808 39914 6820
rect 40773 6817 40785 6820
rect 40819 6817 40831 6851
rect 40773 6811 40831 6817
rect 39301 6783 39359 6789
rect 39301 6749 39313 6783
rect 39347 6749 39359 6783
rect 39301 6743 39359 6749
rect 39482 6740 39488 6792
rect 39540 6780 39546 6792
rect 39945 6783 40003 6789
rect 39945 6780 39957 6783
rect 39540 6752 39957 6780
rect 39540 6740 39546 6752
rect 39945 6749 39957 6752
rect 39991 6749 40003 6783
rect 39945 6743 40003 6749
rect 40497 6783 40555 6789
rect 40497 6749 40509 6783
rect 40543 6780 40555 6783
rect 40954 6780 40960 6792
rect 40543 6752 40960 6780
rect 40543 6749 40555 6752
rect 40497 6743 40555 6749
rect 40954 6740 40960 6752
rect 41012 6740 41018 6792
rect 26200 6684 26464 6712
rect 26528 6684 27568 6712
rect 28276 6684 28948 6712
rect 32416 6684 33732 6712
rect 34164 6684 34928 6712
rect 26200 6672 26206 6684
rect 22649 6647 22707 6653
rect 22649 6644 22661 6647
rect 22066 6616 22661 6644
rect 21453 6607 21511 6613
rect 22649 6613 22661 6616
rect 22695 6613 22707 6647
rect 22649 6607 22707 6613
rect 23201 6647 23259 6653
rect 23201 6613 23213 6647
rect 23247 6613 23259 6647
rect 23201 6607 23259 6613
rect 23382 6604 23388 6656
rect 23440 6644 23446 6656
rect 25041 6647 25099 6653
rect 25041 6644 25053 6647
rect 23440 6616 25053 6644
rect 23440 6604 23446 6616
rect 25041 6613 25053 6616
rect 25087 6613 25099 6647
rect 25041 6607 25099 6613
rect 25314 6604 25320 6656
rect 25372 6604 25378 6656
rect 25590 6604 25596 6656
rect 25648 6604 25654 6656
rect 26436 6644 26464 6684
rect 27540 6656 27568 6684
rect 26697 6647 26755 6653
rect 26697 6644 26709 6647
rect 26436 6616 26709 6644
rect 26697 6613 26709 6616
rect 26743 6613 26755 6647
rect 26697 6607 26755 6613
rect 26970 6604 26976 6656
rect 27028 6604 27034 6656
rect 27338 6604 27344 6656
rect 27396 6604 27402 6656
rect 27522 6604 27528 6656
rect 27580 6604 27586 6656
rect 27614 6604 27620 6656
rect 27672 6644 27678 6656
rect 27709 6647 27767 6653
rect 27709 6644 27721 6647
rect 27672 6616 27721 6644
rect 27672 6604 27678 6616
rect 27709 6613 27721 6616
rect 27755 6613 27767 6647
rect 27709 6607 27767 6613
rect 28074 6604 28080 6656
rect 28132 6604 28138 6656
rect 28442 6604 28448 6656
rect 28500 6604 28506 6656
rect 28902 6604 28908 6656
rect 28960 6604 28966 6656
rect 29362 6604 29368 6656
rect 29420 6604 29426 6656
rect 29822 6604 29828 6656
rect 29880 6604 29886 6656
rect 30190 6604 30196 6656
rect 30248 6604 30254 6656
rect 30282 6604 30288 6656
rect 30340 6644 30346 6656
rect 30469 6647 30527 6653
rect 30469 6644 30481 6647
rect 30340 6616 30481 6644
rect 30340 6604 30346 6616
rect 30469 6613 30481 6616
rect 30515 6613 30527 6647
rect 30469 6607 30527 6613
rect 31386 6604 31392 6656
rect 31444 6604 31450 6656
rect 32416 6653 32444 6684
rect 34164 6656 34192 6684
rect 35434 6672 35440 6724
rect 35492 6672 35498 6724
rect 35986 6672 35992 6724
rect 36044 6672 36050 6724
rect 36538 6672 36544 6724
rect 36596 6672 36602 6724
rect 37090 6672 37096 6724
rect 37148 6672 37154 6724
rect 37642 6672 37648 6724
rect 37700 6672 37706 6724
rect 38194 6672 38200 6724
rect 38252 6672 38258 6724
rect 38378 6672 38384 6724
rect 38436 6712 38442 6724
rect 38749 6715 38807 6721
rect 38749 6712 38761 6715
rect 38436 6684 38761 6712
rect 38436 6672 38442 6684
rect 38749 6681 38761 6684
rect 38795 6681 38807 6715
rect 38749 6675 38807 6681
rect 39206 6672 39212 6724
rect 39264 6712 39270 6724
rect 39264 6684 40080 6712
rect 39264 6672 39270 6684
rect 32401 6647 32459 6653
rect 32401 6613 32413 6647
rect 32447 6613 32459 6647
rect 32401 6607 32459 6613
rect 33318 6604 33324 6656
rect 33376 6604 33382 6656
rect 33594 6604 33600 6656
rect 33652 6604 33658 6656
rect 33686 6604 33692 6656
rect 33744 6604 33750 6656
rect 33962 6604 33968 6656
rect 34020 6604 34026 6656
rect 34146 6604 34152 6656
rect 34204 6604 34210 6656
rect 34422 6604 34428 6656
rect 34480 6604 34486 6656
rect 34977 6647 35035 6653
rect 34977 6613 34989 6647
rect 35023 6644 35035 6647
rect 35894 6644 35900 6656
rect 35023 6616 35900 6644
rect 35023 6613 35035 6616
rect 34977 6607 35035 6613
rect 35894 6604 35900 6616
rect 35952 6604 35958 6656
rect 36078 6604 36084 6656
rect 36136 6644 36142 6656
rect 36633 6647 36691 6653
rect 36633 6644 36645 6647
rect 36136 6616 36645 6644
rect 36136 6604 36142 6616
rect 36633 6613 36645 6616
rect 36679 6613 36691 6647
rect 36633 6607 36691 6613
rect 36722 6604 36728 6656
rect 36780 6644 36786 6656
rect 37185 6647 37243 6653
rect 37185 6644 37197 6647
rect 36780 6616 37197 6644
rect 36780 6604 36786 6616
rect 37185 6613 37197 6616
rect 37231 6613 37243 6647
rect 37185 6607 37243 6613
rect 37734 6604 37740 6656
rect 37792 6644 37798 6656
rect 38289 6647 38347 6653
rect 38289 6644 38301 6647
rect 37792 6616 38301 6644
rect 37792 6604 37798 6616
rect 38289 6613 38301 6616
rect 38335 6613 38347 6647
rect 38289 6607 38347 6613
rect 38470 6604 38476 6656
rect 38528 6644 38534 6656
rect 38841 6647 38899 6653
rect 38841 6644 38853 6647
rect 38528 6616 38853 6644
rect 38528 6604 38534 6616
rect 38841 6613 38853 6616
rect 38887 6613 38899 6647
rect 38841 6607 38899 6613
rect 38930 6604 38936 6656
rect 38988 6644 38994 6656
rect 40052 6653 40080 6684
rect 39393 6647 39451 6653
rect 39393 6644 39405 6647
rect 38988 6616 39405 6644
rect 38988 6604 38994 6616
rect 39393 6613 39405 6616
rect 39439 6613 39451 6647
rect 39393 6607 39451 6613
rect 40037 6647 40095 6653
rect 40037 6613 40049 6647
rect 40083 6613 40095 6647
rect 40037 6607 40095 6613
rect 1104 6554 44040 6576
rect 1104 6502 11644 6554
rect 11696 6502 11708 6554
rect 11760 6502 11772 6554
rect 11824 6502 11836 6554
rect 11888 6502 11900 6554
rect 11952 6502 22338 6554
rect 22390 6502 22402 6554
rect 22454 6502 22466 6554
rect 22518 6502 22530 6554
rect 22582 6502 22594 6554
rect 22646 6502 33032 6554
rect 33084 6502 33096 6554
rect 33148 6502 33160 6554
rect 33212 6502 33224 6554
rect 33276 6502 33288 6554
rect 33340 6502 43726 6554
rect 43778 6502 43790 6554
rect 43842 6502 43854 6554
rect 43906 6502 43918 6554
rect 43970 6502 43982 6554
rect 44034 6502 44040 6554
rect 1104 6480 44040 6502
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5684 6412 6009 6440
rect 5684 6400 5690 6412
rect 5997 6409 6009 6412
rect 6043 6409 6055 6443
rect 5997 6403 6055 6409
rect 6086 6400 6092 6452
rect 6144 6440 6150 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 6144 6412 7849 6440
rect 6144 6400 6150 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 7837 6403 7895 6409
rect 8662 6400 8668 6452
rect 8720 6400 8726 6452
rect 9214 6400 9220 6452
rect 9272 6400 9278 6452
rect 9766 6400 9772 6452
rect 9824 6400 9830 6452
rect 10502 6440 10508 6452
rect 10152 6412 10508 6440
rect 5920 6344 9628 6372
rect 5920 6313 5948 6344
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 6178 6264 6184 6316
rect 6236 6264 6242 6316
rect 8018 6264 8024 6316
rect 8076 6264 8082 6316
rect 8570 6264 8576 6316
rect 8628 6264 8634 6316
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9600 6304 9628 6344
rect 9674 6332 9680 6384
rect 9732 6332 9738 6384
rect 10152 6304 10180 6412
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 10686 6400 10692 6452
rect 10744 6440 10750 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 10744 6412 11529 6440
rect 10744 6400 10750 6412
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 11517 6403 11575 6409
rect 11974 6400 11980 6452
rect 12032 6400 12038 6452
rect 13817 6443 13875 6449
rect 13817 6409 13829 6443
rect 13863 6409 13875 6443
rect 13817 6403 13875 6409
rect 10229 6375 10287 6381
rect 10229 6341 10241 6375
rect 10275 6372 10287 6375
rect 13630 6372 13636 6384
rect 10275 6344 13636 6372
rect 10275 6341 10287 6344
rect 10229 6335 10287 6341
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 13832 6372 13860 6403
rect 13998 6400 14004 6452
rect 14056 6440 14062 6452
rect 14277 6443 14335 6449
rect 14277 6440 14289 6443
rect 14056 6412 14289 6440
rect 14056 6400 14062 6412
rect 14277 6409 14289 6412
rect 14323 6409 14335 6443
rect 14277 6403 14335 6409
rect 14458 6400 14464 6452
rect 14516 6440 14522 6452
rect 14645 6443 14703 6449
rect 14645 6440 14657 6443
rect 14516 6412 14657 6440
rect 14516 6400 14522 6412
rect 14645 6409 14657 6412
rect 14691 6409 14703 6443
rect 14645 6403 14703 6409
rect 14734 6400 14740 6452
rect 14792 6440 14798 6452
rect 14792 6412 15240 6440
rect 14792 6400 14798 6412
rect 15010 6372 15016 6384
rect 13832 6344 15016 6372
rect 15010 6332 15016 6344
rect 15068 6332 15074 6384
rect 15212 6372 15240 6412
rect 15286 6400 15292 6452
rect 15344 6400 15350 6452
rect 15562 6400 15568 6452
rect 15620 6440 15626 6452
rect 15657 6443 15715 6449
rect 15657 6440 15669 6443
rect 15620 6412 15669 6440
rect 15620 6400 15626 6412
rect 15657 6409 15669 6412
rect 15703 6409 15715 6443
rect 15657 6403 15715 6409
rect 16117 6443 16175 6449
rect 16117 6409 16129 6443
rect 16163 6440 16175 6443
rect 16666 6440 16672 6452
rect 16163 6412 16672 6440
rect 16163 6409 16175 6412
rect 16117 6403 16175 6409
rect 16666 6400 16672 6412
rect 16724 6400 16730 6452
rect 17218 6400 17224 6452
rect 17276 6440 17282 6452
rect 17589 6443 17647 6449
rect 17589 6440 17601 6443
rect 17276 6412 17601 6440
rect 17276 6400 17282 6412
rect 17589 6409 17601 6412
rect 17635 6409 17647 6443
rect 17589 6403 17647 6409
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 18049 6443 18107 6449
rect 18049 6440 18061 6443
rect 17920 6412 18061 6440
rect 17920 6400 17926 6412
rect 18049 6409 18061 6412
rect 18095 6409 18107 6443
rect 18049 6403 18107 6409
rect 18322 6400 18328 6452
rect 18380 6400 18386 6452
rect 18598 6400 18604 6452
rect 18656 6400 18662 6452
rect 18966 6400 18972 6452
rect 19024 6400 19030 6452
rect 19058 6400 19064 6452
rect 19116 6400 19122 6452
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 22002 6440 22008 6452
rect 19392 6412 22008 6440
rect 19392 6400 19398 6412
rect 22002 6400 22008 6412
rect 22060 6400 22066 6452
rect 22186 6400 22192 6452
rect 22244 6440 22250 6452
rect 22465 6443 22523 6449
rect 22465 6440 22477 6443
rect 22244 6412 22477 6440
rect 22244 6400 22250 6412
rect 22465 6409 22477 6412
rect 22511 6409 22523 6443
rect 22922 6440 22928 6452
rect 22465 6403 22523 6409
rect 22572 6412 22928 6440
rect 18138 6372 18144 6384
rect 15212 6344 18144 6372
rect 18138 6332 18144 6344
rect 18196 6332 18202 6384
rect 9600 6276 10180 6304
rect 9125 6267 9183 6273
rect 5534 6196 5540 6248
rect 5592 6196 5598 6248
rect 9140 6236 9168 6267
rect 11054 6264 11060 6316
rect 11112 6264 11118 6316
rect 11698 6264 11704 6316
rect 11756 6264 11762 6316
rect 11882 6264 11888 6316
rect 11940 6264 11946 6316
rect 14001 6307 14059 6313
rect 13740 6276 13952 6304
rect 13740 6236 13768 6276
rect 9140 6208 13768 6236
rect 13924 6236 13952 6276
rect 14001 6273 14013 6307
rect 14047 6304 14059 6307
rect 14090 6304 14096 6316
rect 14047 6276 14096 6304
rect 14047 6273 14059 6276
rect 14001 6267 14059 6273
rect 14090 6264 14096 6276
rect 14148 6264 14154 6316
rect 14185 6307 14243 6313
rect 14185 6273 14197 6307
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 14200 6236 14228 6267
rect 14826 6264 14832 6316
rect 14884 6264 14890 6316
rect 15470 6264 15476 6316
rect 15528 6264 15534 6316
rect 15838 6264 15844 6316
rect 15896 6264 15902 6316
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 16390 6304 16396 6316
rect 16347 6276 16396 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6304 16911 6307
rect 17221 6307 17279 6313
rect 17221 6304 17233 6307
rect 16899 6276 17233 6304
rect 16899 6273 16911 6276
rect 16853 6267 16911 6273
rect 17221 6273 17233 6276
rect 17267 6304 17279 6307
rect 17402 6304 17408 6316
rect 17267 6276 17408 6304
rect 17267 6273 17279 6276
rect 17221 6267 17279 6273
rect 17402 6264 17408 6276
rect 17460 6264 17466 6316
rect 17494 6264 17500 6316
rect 17552 6264 17558 6316
rect 17770 6264 17776 6316
rect 17828 6264 17834 6316
rect 18230 6264 18236 6316
rect 18288 6264 18294 6316
rect 18506 6264 18512 6316
rect 18564 6264 18570 6316
rect 18782 6264 18788 6316
rect 18840 6264 18846 6316
rect 17862 6236 17868 6248
rect 13924 6208 14044 6236
rect 14200 6208 17868 6236
rect 5552 6168 5580 6196
rect 5721 6171 5779 6177
rect 5721 6168 5733 6171
rect 5552 6140 5733 6168
rect 5721 6137 5733 6140
rect 5767 6137 5779 6171
rect 5721 6131 5779 6137
rect 9398 6128 9404 6180
rect 9456 6168 9462 6180
rect 10873 6171 10931 6177
rect 10873 6168 10885 6171
rect 9456 6140 10885 6168
rect 9456 6128 9462 6140
rect 10873 6137 10885 6140
rect 10919 6137 10931 6171
rect 10873 6131 10931 6137
rect 9306 6060 9312 6112
rect 9364 6100 9370 6112
rect 10321 6103 10379 6109
rect 10321 6100 10333 6103
rect 9364 6072 10333 6100
rect 9364 6060 9370 6072
rect 10321 6069 10333 6072
rect 10367 6069 10379 6103
rect 10321 6063 10379 6069
rect 10410 6060 10416 6112
rect 10468 6100 10474 6112
rect 13630 6100 13636 6112
rect 10468 6072 13636 6100
rect 10468 6060 10474 6072
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 14016 6100 14044 6208
rect 17862 6196 17868 6208
rect 17920 6196 17926 6248
rect 19076 6236 19104 6400
rect 19168 6344 22232 6372
rect 19168 6313 19196 6344
rect 19153 6307 19211 6313
rect 19153 6273 19165 6307
rect 19199 6273 19211 6307
rect 19153 6267 19211 6273
rect 20438 6264 20444 6316
rect 20496 6264 20502 6316
rect 21821 6307 21879 6313
rect 21821 6273 21833 6307
rect 21867 6304 21879 6307
rect 21910 6304 21916 6316
rect 21867 6276 21916 6304
rect 21867 6273 21879 6276
rect 21821 6267 21879 6273
rect 21910 6264 21916 6276
rect 21968 6264 21974 6316
rect 22094 6236 22100 6248
rect 19076 6208 22100 6236
rect 22094 6196 22100 6208
rect 22152 6196 22158 6248
rect 22204 6236 22232 6344
rect 22281 6307 22339 6313
rect 22281 6273 22293 6307
rect 22327 6304 22339 6307
rect 22572 6304 22600 6412
rect 22922 6400 22928 6412
rect 22980 6400 22986 6452
rect 25958 6400 25964 6452
rect 26016 6440 26022 6452
rect 27338 6440 27344 6452
rect 26016 6412 27344 6440
rect 26016 6400 26022 6412
rect 27338 6400 27344 6412
rect 27396 6400 27402 6452
rect 33686 6400 33692 6452
rect 33744 6440 33750 6452
rect 34790 6440 34796 6452
rect 33744 6412 34796 6440
rect 33744 6400 33750 6412
rect 34790 6400 34796 6412
rect 34848 6400 34854 6452
rect 37277 6443 37335 6449
rect 37277 6409 37289 6443
rect 37323 6440 37335 6443
rect 38194 6440 38200 6452
rect 37323 6412 38200 6440
rect 37323 6409 37335 6412
rect 37277 6403 37335 6409
rect 38194 6400 38200 6412
rect 38252 6400 38258 6452
rect 38378 6400 38384 6452
rect 38436 6400 38442 6452
rect 30926 6372 30932 6384
rect 22327 6276 22600 6304
rect 22664 6344 30932 6372
rect 22327 6273 22339 6276
rect 22281 6267 22339 6273
rect 22664 6236 22692 6344
rect 30926 6332 30932 6344
rect 30984 6332 30990 6384
rect 33962 6332 33968 6384
rect 34020 6372 34026 6384
rect 38396 6372 38424 6400
rect 34020 6344 38424 6372
rect 34020 6332 34026 6344
rect 22741 6307 22799 6313
rect 22741 6273 22753 6307
rect 22787 6304 22799 6307
rect 22940 6304 23152 6308
rect 23474 6304 23480 6316
rect 22787 6280 23480 6304
rect 22787 6276 22968 6280
rect 23124 6276 23480 6280
rect 22787 6273 22799 6276
rect 22741 6267 22799 6273
rect 23474 6264 23480 6276
rect 23532 6264 23538 6316
rect 25777 6307 25835 6313
rect 25777 6273 25789 6307
rect 25823 6304 25835 6307
rect 25866 6304 25872 6316
rect 25823 6276 25872 6304
rect 25823 6273 25835 6276
rect 25777 6267 25835 6273
rect 25866 6264 25872 6276
rect 25924 6264 25930 6316
rect 34238 6264 34244 6316
rect 34296 6264 34302 6316
rect 37090 6304 37096 6316
rect 35866 6276 37096 6304
rect 22204 6208 22692 6236
rect 23106 6196 23112 6248
rect 23164 6236 23170 6248
rect 30282 6236 30288 6248
rect 23164 6208 30288 6236
rect 23164 6196 23170 6208
rect 30282 6196 30288 6208
rect 30340 6196 30346 6248
rect 30374 6196 30380 6248
rect 30432 6236 30438 6248
rect 35866 6236 35894 6276
rect 37090 6264 37096 6276
rect 37148 6264 37154 6316
rect 37274 6264 37280 6316
rect 37332 6304 37338 6316
rect 37461 6307 37519 6313
rect 37461 6304 37473 6307
rect 37332 6276 37473 6304
rect 37332 6264 37338 6276
rect 37461 6273 37473 6276
rect 37507 6273 37519 6307
rect 37461 6267 37519 6273
rect 37737 6307 37795 6313
rect 37737 6273 37749 6307
rect 37783 6273 37795 6307
rect 37737 6267 37795 6273
rect 30432 6208 35894 6236
rect 30432 6196 30438 6208
rect 36722 6196 36728 6248
rect 36780 6236 36786 6248
rect 37752 6236 37780 6267
rect 36780 6208 37780 6236
rect 36780 6196 36786 6208
rect 39022 6196 39028 6248
rect 39080 6196 39086 6248
rect 16574 6128 16580 6180
rect 16632 6168 16638 6180
rect 16669 6171 16727 6177
rect 16669 6168 16681 6171
rect 16632 6140 16681 6168
rect 16632 6128 16638 6140
rect 16669 6137 16681 6140
rect 16715 6137 16727 6171
rect 16669 6131 16727 6137
rect 17310 6128 17316 6180
rect 17368 6128 17374 6180
rect 17402 6128 17408 6180
rect 17460 6168 17466 6180
rect 20898 6168 20904 6180
rect 17460 6140 20904 6168
rect 17460 6128 17466 6140
rect 20898 6128 20904 6140
rect 20956 6128 20962 6180
rect 25314 6168 25320 6180
rect 21008 6140 25320 6168
rect 20625 6103 20683 6109
rect 20625 6100 20637 6103
rect 14016 6072 20637 6100
rect 20625 6069 20637 6072
rect 20671 6069 20683 6103
rect 20625 6063 20683 6069
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 21008 6100 21036 6140
rect 25314 6128 25320 6140
rect 25372 6128 25378 6180
rect 37553 6171 37611 6177
rect 37553 6137 37565 6171
rect 37599 6168 37611 6171
rect 39040 6168 39068 6196
rect 37599 6140 39068 6168
rect 37599 6137 37611 6140
rect 37553 6131 37611 6137
rect 20772 6072 21036 6100
rect 20772 6060 20778 6072
rect 22002 6060 22008 6112
rect 22060 6060 22066 6112
rect 22925 6103 22983 6109
rect 22925 6069 22937 6103
rect 22971 6100 22983 6103
rect 23014 6100 23020 6112
rect 22971 6072 23020 6100
rect 22971 6069 22983 6072
rect 22925 6063 22983 6069
rect 23014 6060 23020 6072
rect 23072 6060 23078 6112
rect 24026 6060 24032 6112
rect 24084 6100 24090 6112
rect 25961 6103 26019 6109
rect 25961 6100 25973 6103
rect 24084 6072 25973 6100
rect 24084 6060 24090 6072
rect 25961 6069 25973 6072
rect 26007 6069 26019 6103
rect 25961 6063 26019 6069
rect 34057 6103 34115 6109
rect 34057 6069 34069 6103
rect 34103 6100 34115 6103
rect 35342 6100 35348 6112
rect 34103 6072 35348 6100
rect 34103 6069 34115 6072
rect 34057 6063 34115 6069
rect 35342 6060 35348 6072
rect 35400 6060 35406 6112
rect 1104 6010 43884 6032
rect 1104 5958 6297 6010
rect 6349 5958 6361 6010
rect 6413 5958 6425 6010
rect 6477 5958 6489 6010
rect 6541 5958 6553 6010
rect 6605 5958 16991 6010
rect 17043 5958 17055 6010
rect 17107 5958 17119 6010
rect 17171 5958 17183 6010
rect 17235 5958 17247 6010
rect 17299 5958 27685 6010
rect 27737 5958 27749 6010
rect 27801 5958 27813 6010
rect 27865 5958 27877 6010
rect 27929 5958 27941 6010
rect 27993 5958 38379 6010
rect 38431 5958 38443 6010
rect 38495 5958 38507 6010
rect 38559 5958 38571 6010
rect 38623 5958 38635 6010
rect 38687 5958 43884 6010
rect 1104 5936 43884 5958
rect 6178 5856 6184 5908
rect 6236 5856 6242 5908
rect 8018 5856 8024 5908
rect 8076 5896 8082 5908
rect 10410 5896 10416 5908
rect 8076 5868 10416 5896
rect 8076 5856 8082 5868
rect 10410 5856 10416 5868
rect 10468 5856 10474 5908
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 12989 5899 13047 5905
rect 11756 5868 12434 5896
rect 11756 5856 11762 5868
rect 6196 5760 6224 5856
rect 12406 5828 12434 5868
rect 12989 5865 13001 5899
rect 13035 5896 13047 5899
rect 13354 5896 13360 5908
rect 13035 5868 13360 5896
rect 13035 5865 13047 5868
rect 12989 5859 13047 5865
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 13630 5856 13636 5908
rect 13688 5896 13694 5908
rect 16298 5896 16304 5908
rect 13688 5868 16304 5896
rect 13688 5856 13694 5868
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 17402 5856 17408 5908
rect 17460 5856 17466 5908
rect 18230 5856 18236 5908
rect 18288 5856 18294 5908
rect 20806 5856 20812 5908
rect 20864 5896 20870 5908
rect 29362 5896 29368 5908
rect 20864 5868 29368 5896
rect 20864 5856 20870 5868
rect 29362 5856 29368 5868
rect 29420 5856 29426 5908
rect 17420 5828 17448 5856
rect 12406 5800 17448 5828
rect 18248 5828 18276 5856
rect 18248 5800 22094 5828
rect 19794 5760 19800 5772
rect 6196 5732 19800 5760
rect 19794 5720 19800 5732
rect 19852 5720 19858 5772
rect 22066 5760 22094 5800
rect 22186 5788 22192 5840
rect 22244 5828 22250 5840
rect 23290 5828 23296 5840
rect 22244 5800 23296 5828
rect 22244 5788 22250 5800
rect 23290 5788 23296 5800
rect 23348 5788 23354 5840
rect 26970 5788 26976 5840
rect 27028 5788 27034 5840
rect 23198 5760 23204 5772
rect 22066 5732 23204 5760
rect 23198 5720 23204 5732
rect 23256 5720 23262 5772
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 11112 5664 12434 5692
rect 11112 5652 11118 5664
rect 12406 5624 12434 5664
rect 12802 5652 12808 5704
rect 12860 5652 12866 5704
rect 12986 5652 12992 5704
rect 13044 5692 13050 5704
rect 26988 5692 27016 5788
rect 13044 5664 27016 5692
rect 13044 5652 13050 5664
rect 16482 5624 16488 5636
rect 12406 5596 16488 5624
rect 16482 5584 16488 5596
rect 16540 5584 16546 5636
rect 17494 5584 17500 5636
rect 17552 5624 17558 5636
rect 32306 5624 32312 5636
rect 17552 5596 32312 5624
rect 17552 5584 17558 5596
rect 32306 5584 32312 5596
rect 32364 5584 32370 5636
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 12066 5556 12072 5568
rect 8628 5528 12072 5556
rect 8628 5516 8634 5528
rect 12066 5516 12072 5528
rect 12124 5516 12130 5568
rect 17678 5516 17684 5568
rect 17736 5556 17742 5568
rect 31386 5556 31392 5568
rect 17736 5528 31392 5556
rect 17736 5516 17742 5528
rect 31386 5516 31392 5528
rect 31444 5516 31450 5568
rect 1104 5466 44040 5488
rect 1104 5414 11644 5466
rect 11696 5414 11708 5466
rect 11760 5414 11772 5466
rect 11824 5414 11836 5466
rect 11888 5414 11900 5466
rect 11952 5414 22338 5466
rect 22390 5414 22402 5466
rect 22454 5414 22466 5466
rect 22518 5414 22530 5466
rect 22582 5414 22594 5466
rect 22646 5414 33032 5466
rect 33084 5414 33096 5466
rect 33148 5414 33160 5466
rect 33212 5414 33224 5466
rect 33276 5414 33288 5466
rect 33340 5414 43726 5466
rect 43778 5414 43790 5466
rect 43842 5414 43854 5466
rect 43906 5414 43918 5466
rect 43970 5414 43982 5466
rect 44034 5414 44040 5466
rect 1104 5392 44040 5414
rect 18138 5312 18144 5364
rect 18196 5352 18202 5364
rect 23382 5352 23388 5364
rect 18196 5324 23388 5352
rect 18196 5312 18202 5324
rect 23382 5312 23388 5324
rect 23440 5312 23446 5364
rect 13722 5244 13728 5296
rect 13780 5284 13786 5296
rect 25958 5284 25964 5296
rect 13780 5256 25964 5284
rect 13780 5244 13786 5256
rect 25958 5244 25964 5256
rect 26016 5244 26022 5296
rect 20438 5176 20444 5228
rect 20496 5216 20502 5228
rect 20809 5219 20867 5225
rect 20809 5216 20821 5219
rect 20496 5188 20821 5216
rect 20496 5176 20502 5188
rect 20809 5185 20821 5188
rect 20855 5185 20867 5219
rect 20809 5179 20867 5185
rect 11974 5108 11980 5160
rect 12032 5148 12038 5160
rect 28074 5148 28080 5160
rect 12032 5120 28080 5148
rect 12032 5108 12038 5120
rect 28074 5108 28080 5120
rect 28132 5108 28138 5160
rect 14182 5040 14188 5092
rect 14240 5080 14246 5092
rect 27614 5080 27620 5092
rect 14240 5052 27620 5080
rect 14240 5040 14246 5052
rect 27614 5040 27620 5052
rect 27672 5040 27678 5092
rect 6730 4972 6736 5024
rect 6788 5012 6794 5024
rect 19518 5012 19524 5024
rect 6788 4984 19524 5012
rect 6788 4972 6794 4984
rect 19518 4972 19524 4984
rect 19576 4972 19582 5024
rect 20993 5015 21051 5021
rect 20993 4981 21005 5015
rect 21039 5012 21051 5015
rect 30374 5012 30380 5024
rect 21039 4984 30380 5012
rect 21039 4981 21051 4984
rect 20993 4975 21051 4981
rect 30374 4972 30380 4984
rect 30432 4972 30438 5024
rect 1104 4922 43884 4944
rect 1104 4870 6297 4922
rect 6349 4870 6361 4922
rect 6413 4870 6425 4922
rect 6477 4870 6489 4922
rect 6541 4870 6553 4922
rect 6605 4870 16991 4922
rect 17043 4870 17055 4922
rect 17107 4870 17119 4922
rect 17171 4870 17183 4922
rect 17235 4870 17247 4922
rect 17299 4870 27685 4922
rect 27737 4870 27749 4922
rect 27801 4870 27813 4922
rect 27865 4870 27877 4922
rect 27929 4870 27941 4922
rect 27993 4870 38379 4922
rect 38431 4870 38443 4922
rect 38495 4870 38507 4922
rect 38559 4870 38571 4922
rect 38623 4870 38635 4922
rect 38687 4870 43884 4922
rect 1104 4848 43884 4870
rect 10594 4768 10600 4820
rect 10652 4808 10658 4820
rect 30190 4808 30196 4820
rect 10652 4780 30196 4808
rect 10652 4768 10658 4780
rect 30190 4768 30196 4780
rect 30248 4768 30254 4820
rect 10778 4700 10784 4752
rect 10836 4740 10842 4752
rect 29822 4740 29828 4752
rect 10836 4712 29828 4740
rect 10836 4700 10842 4712
rect 29822 4700 29828 4712
rect 29880 4700 29886 4752
rect 13906 4632 13912 4684
rect 13964 4672 13970 4684
rect 26418 4672 26424 4684
rect 13964 4644 26424 4672
rect 13964 4632 13970 4644
rect 26418 4632 26424 4644
rect 26476 4632 26482 4684
rect 11330 4564 11336 4616
rect 11388 4604 11394 4616
rect 28902 4604 28908 4616
rect 11388 4576 28908 4604
rect 11388 4564 11394 4576
rect 28902 4564 28908 4576
rect 28960 4564 28966 4616
rect 33410 4564 33416 4616
rect 33468 4604 33474 4616
rect 36538 4604 36544 4616
rect 33468 4576 36544 4604
rect 33468 4564 33474 4576
rect 36538 4564 36544 4576
rect 36596 4564 36602 4616
rect 1104 4378 44040 4400
rect 1104 4326 11644 4378
rect 11696 4326 11708 4378
rect 11760 4326 11772 4378
rect 11824 4326 11836 4378
rect 11888 4326 11900 4378
rect 11952 4326 22338 4378
rect 22390 4326 22402 4378
rect 22454 4326 22466 4378
rect 22518 4326 22530 4378
rect 22582 4326 22594 4378
rect 22646 4326 33032 4378
rect 33084 4326 33096 4378
rect 33148 4326 33160 4378
rect 33212 4326 33224 4378
rect 33276 4326 33288 4378
rect 33340 4326 43726 4378
rect 43778 4326 43790 4378
rect 43842 4326 43854 4378
rect 43906 4326 43918 4378
rect 43970 4326 43982 4378
rect 44034 4326 44040 4378
rect 1104 4304 44040 4326
rect 1104 3834 43884 3856
rect 1104 3782 6297 3834
rect 6349 3782 6361 3834
rect 6413 3782 6425 3834
rect 6477 3782 6489 3834
rect 6541 3782 6553 3834
rect 6605 3782 16991 3834
rect 17043 3782 17055 3834
rect 17107 3782 17119 3834
rect 17171 3782 17183 3834
rect 17235 3782 17247 3834
rect 17299 3782 27685 3834
rect 27737 3782 27749 3834
rect 27801 3782 27813 3834
rect 27865 3782 27877 3834
rect 27929 3782 27941 3834
rect 27993 3782 38379 3834
rect 38431 3782 38443 3834
rect 38495 3782 38507 3834
rect 38559 3782 38571 3834
rect 38623 3782 38635 3834
rect 38687 3782 43884 3834
rect 1104 3760 43884 3782
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 35158 3516 35164 3528
rect 11020 3488 35164 3516
rect 11020 3476 11026 3488
rect 35158 3476 35164 3488
rect 35216 3476 35222 3528
rect 6638 3408 6644 3460
rect 6696 3448 6702 3460
rect 34238 3448 34244 3460
rect 6696 3420 34244 3448
rect 6696 3408 6702 3420
rect 34238 3408 34244 3420
rect 34296 3408 34302 3460
rect 1104 3290 44040 3312
rect 1104 3238 11644 3290
rect 11696 3238 11708 3290
rect 11760 3238 11772 3290
rect 11824 3238 11836 3290
rect 11888 3238 11900 3290
rect 11952 3238 22338 3290
rect 22390 3238 22402 3290
rect 22454 3238 22466 3290
rect 22518 3238 22530 3290
rect 22582 3238 22594 3290
rect 22646 3238 33032 3290
rect 33084 3238 33096 3290
rect 33148 3238 33160 3290
rect 33212 3238 33224 3290
rect 33276 3238 33288 3290
rect 33340 3238 43726 3290
rect 43778 3238 43790 3290
rect 43842 3238 43854 3290
rect 43906 3238 43918 3290
rect 43970 3238 43982 3290
rect 44034 3238 44040 3290
rect 1104 3216 44040 3238
rect 18877 3179 18935 3185
rect 18877 3145 18889 3179
rect 18923 3176 18935 3179
rect 18923 3148 31754 3176
rect 18923 3145 18935 3148
rect 18877 3139 18935 3145
rect 31726 3108 31754 3148
rect 37550 3108 37556 3120
rect 31726 3080 37556 3108
rect 37550 3068 37556 3080
rect 37608 3068 37614 3120
rect 18690 3000 18696 3052
rect 18748 3000 18754 3052
rect 22922 3000 22928 3052
rect 22980 3000 22986 3052
rect 25038 3000 25044 3052
rect 25096 3000 25102 3052
rect 28966 2944 31800 2972
rect 23109 2907 23167 2913
rect 23109 2873 23121 2907
rect 23155 2904 23167 2907
rect 28966 2904 28994 2944
rect 23155 2876 28994 2904
rect 31772 2904 31800 2944
rect 33134 2932 33140 2984
rect 33192 2972 33198 2984
rect 35986 2972 35992 2984
rect 33192 2944 35992 2972
rect 33192 2932 33198 2944
rect 35986 2932 35992 2944
rect 36044 2932 36050 2984
rect 37918 2904 37924 2916
rect 31772 2876 37924 2904
rect 23155 2873 23167 2876
rect 23109 2867 23167 2873
rect 37918 2864 37924 2876
rect 37976 2864 37982 2916
rect 25225 2839 25283 2845
rect 25225 2805 25237 2839
rect 25271 2836 25283 2839
rect 37642 2836 37648 2848
rect 25271 2808 37648 2836
rect 25271 2805 25283 2808
rect 25225 2799 25283 2805
rect 37642 2796 37648 2808
rect 37700 2796 37706 2848
rect 1104 2746 43884 2768
rect 1104 2694 6297 2746
rect 6349 2694 6361 2746
rect 6413 2694 6425 2746
rect 6477 2694 6489 2746
rect 6541 2694 6553 2746
rect 6605 2694 16991 2746
rect 17043 2694 17055 2746
rect 17107 2694 17119 2746
rect 17171 2694 17183 2746
rect 17235 2694 17247 2746
rect 17299 2694 27685 2746
rect 27737 2694 27749 2746
rect 27801 2694 27813 2746
rect 27865 2694 27877 2746
rect 27929 2694 27941 2746
rect 27993 2694 38379 2746
rect 38431 2694 38443 2746
rect 38495 2694 38507 2746
rect 38559 2694 38571 2746
rect 38623 2694 38635 2746
rect 38687 2694 43884 2746
rect 1104 2672 43884 2694
rect 3973 2635 4031 2641
rect 3973 2601 3985 2635
rect 4019 2632 4031 2635
rect 6914 2632 6920 2644
rect 4019 2604 6920 2632
rect 4019 2601 4031 2604
rect 3973 2595 4031 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 11977 2635 12035 2641
rect 11977 2601 11989 2635
rect 12023 2632 12035 2635
rect 12802 2632 12808 2644
rect 12023 2604 12808 2632
rect 12023 2601 12035 2604
rect 11977 2595 12035 2601
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 18325 2635 18383 2641
rect 18325 2601 18337 2635
rect 18371 2632 18383 2635
rect 18690 2632 18696 2644
rect 18371 2604 18696 2632
rect 18371 2601 18383 2604
rect 18325 2595 18383 2601
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 20438 2592 20444 2644
rect 20496 2592 20502 2644
rect 22557 2635 22615 2641
rect 22557 2601 22569 2635
rect 22603 2632 22615 2635
rect 22922 2632 22928 2644
rect 22603 2604 22928 2632
rect 22603 2601 22615 2604
rect 22557 2595 22615 2601
rect 22922 2592 22928 2604
rect 22980 2592 22986 2644
rect 24673 2635 24731 2641
rect 24673 2601 24685 2635
rect 24719 2632 24731 2635
rect 25038 2632 25044 2644
rect 24719 2604 25044 2632
rect 24719 2601 24731 2604
rect 24673 2595 24731 2601
rect 25038 2592 25044 2604
rect 25096 2592 25102 2644
rect 33137 2635 33195 2641
rect 26206 2604 29224 2632
rect 16209 2567 16267 2573
rect 16209 2533 16221 2567
rect 16255 2533 16267 2567
rect 16209 2527 16267 2533
rect 16853 2567 16911 2573
rect 16853 2533 16865 2567
rect 16899 2564 16911 2567
rect 26206 2564 26234 2604
rect 16899 2536 26234 2564
rect 29089 2567 29147 2573
rect 16899 2533 16911 2536
rect 16853 2527 16911 2533
rect 29089 2533 29101 2567
rect 29135 2533 29147 2567
rect 29196 2564 29224 2604
rect 33137 2601 33149 2635
rect 33183 2632 33195 2635
rect 34054 2632 34060 2644
rect 33183 2604 34060 2632
rect 33183 2601 33195 2604
rect 33137 2595 33195 2601
rect 34054 2592 34060 2604
rect 34112 2592 34118 2644
rect 34701 2635 34759 2641
rect 34701 2601 34713 2635
rect 34747 2632 34759 2635
rect 35434 2632 35440 2644
rect 34747 2604 35440 2632
rect 34747 2601 34759 2604
rect 34701 2595 34759 2601
rect 35434 2592 35440 2604
rect 35492 2592 35498 2644
rect 35710 2592 35716 2644
rect 35768 2592 35774 2644
rect 36814 2592 36820 2644
rect 36872 2592 36878 2644
rect 37826 2592 37832 2644
rect 37884 2592 37890 2644
rect 39485 2635 39543 2641
rect 39485 2601 39497 2635
rect 39531 2632 39543 2635
rect 39666 2632 39672 2644
rect 39531 2604 39672 2632
rect 39531 2601 39543 2604
rect 39485 2595 39543 2601
rect 39666 2592 39672 2604
rect 39724 2592 39730 2644
rect 41414 2592 41420 2644
rect 41472 2632 41478 2644
rect 41601 2635 41659 2641
rect 41601 2632 41613 2635
rect 41472 2604 41613 2632
rect 41472 2592 41478 2604
rect 41601 2601 41613 2604
rect 41647 2601 41659 2635
rect 41601 2595 41659 2601
rect 43346 2592 43352 2644
rect 43404 2592 43410 2644
rect 33410 2564 33416 2576
rect 29196 2536 33416 2564
rect 29089 2527 29147 2533
rect 6638 2456 6644 2508
rect 6696 2456 6702 2508
rect 8021 2499 8079 2505
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 10962 2496 10968 2508
rect 8067 2468 10968 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 16224 2496 16252 2527
rect 29104 2496 29132 2527
rect 33410 2524 33416 2536
rect 33468 2524 33474 2576
rect 35253 2567 35311 2573
rect 35253 2533 35265 2567
rect 35299 2564 35311 2567
rect 35728 2564 35756 2592
rect 37274 2564 37280 2576
rect 35299 2536 35756 2564
rect 35866 2536 37280 2564
rect 35299 2533 35311 2536
rect 35253 2527 35311 2533
rect 35866 2496 35894 2536
rect 37274 2524 37280 2536
rect 37332 2524 37338 2576
rect 37369 2567 37427 2573
rect 37369 2533 37381 2567
rect 37415 2533 37427 2567
rect 37369 2527 37427 2533
rect 16224 2468 16574 2496
rect 29104 2468 35894 2496
rect 37384 2496 37412 2527
rect 37384 2468 38056 2496
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1360 2400 1409 2428
rect 1360 2388 1366 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5592 2400 6377 2428
rect 5592 2388 5598 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 7742 2388 7748 2440
rect 7800 2388 7806 2440
rect 9858 2388 9864 2440
rect 9916 2388 9922 2440
rect 12158 2388 12164 2440
rect 12216 2388 12222 2440
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14056 2400 14289 2428
rect 14056 2388 14062 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 16390 2388 16396 2440
rect 16448 2388 16454 2440
rect 16546 2428 16574 2468
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16546 2400 16681 2428
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 18230 2388 18236 2440
rect 18288 2428 18294 2440
rect 18509 2431 18567 2437
rect 18509 2428 18521 2431
rect 18288 2400 18521 2428
rect 18288 2388 18294 2400
rect 18509 2397 18521 2400
rect 18555 2397 18567 2431
rect 18509 2391 18567 2397
rect 20622 2388 20628 2440
rect 20680 2388 20686 2440
rect 22738 2388 22744 2440
rect 22796 2388 22802 2440
rect 24854 2388 24860 2440
rect 24912 2388 24918 2440
rect 26694 2388 26700 2440
rect 26752 2428 26758 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 26752 2400 27169 2428
rect 26752 2388 26758 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 28902 2388 28908 2440
rect 28960 2388 28966 2440
rect 31018 2388 31024 2440
rect 31076 2388 31082 2440
rect 32858 2428 32864 2440
rect 31128 2400 32864 2428
rect 3418 2320 3424 2372
rect 3476 2360 3482 2372
rect 3881 2363 3939 2369
rect 3881 2360 3893 2363
rect 3476 2332 3893 2360
rect 3476 2320 3482 2332
rect 3881 2329 3893 2332
rect 3927 2329 3939 2363
rect 3881 2323 3939 2329
rect 14645 2363 14703 2369
rect 14645 2329 14657 2363
rect 14691 2329 14703 2363
rect 14645 2323 14703 2329
rect 14829 2363 14887 2369
rect 14829 2329 14841 2363
rect 14875 2360 14887 2363
rect 31128 2360 31156 2400
rect 32858 2388 32864 2400
rect 32916 2388 32922 2440
rect 32950 2388 32956 2440
rect 33008 2428 33014 2440
rect 33321 2431 33379 2437
rect 33321 2428 33333 2431
rect 33008 2400 33333 2428
rect 33008 2388 33014 2400
rect 33321 2397 33333 2400
rect 33367 2397 33379 2431
rect 33321 2391 33379 2397
rect 34882 2388 34888 2440
rect 34940 2388 34946 2440
rect 35158 2388 35164 2440
rect 35216 2428 35222 2440
rect 35437 2431 35495 2437
rect 35437 2428 35449 2431
rect 35216 2400 35449 2428
rect 35216 2388 35222 2400
rect 35437 2397 35449 2400
rect 35483 2397 35495 2431
rect 35437 2391 35495 2397
rect 36998 2388 37004 2440
rect 37056 2388 37062 2440
rect 37550 2388 37556 2440
rect 37608 2388 37614 2440
rect 38028 2437 38056 2468
rect 38013 2431 38071 2437
rect 38013 2397 38025 2431
rect 38059 2397 38071 2431
rect 38013 2391 38071 2397
rect 39666 2388 39672 2440
rect 39724 2388 39730 2440
rect 41782 2388 41788 2440
rect 41840 2388 41846 2440
rect 43530 2388 43536 2440
rect 43588 2388 43594 2440
rect 36722 2360 36728 2372
rect 14875 2332 31156 2360
rect 31220 2332 36728 2360
rect 14875 2329 14887 2332
rect 14829 2323 14887 2329
rect 10042 2252 10048 2304
rect 10100 2252 10106 2304
rect 14093 2295 14151 2301
rect 14093 2261 14105 2295
rect 14139 2292 14151 2295
rect 14660 2292 14688 2323
rect 14139 2264 14688 2292
rect 14139 2261 14151 2264
rect 14093 2255 14151 2261
rect 26970 2252 26976 2304
rect 27028 2252 27034 2304
rect 31220 2301 31248 2332
rect 36722 2320 36728 2332
rect 36780 2320 36786 2372
rect 31205 2295 31263 2301
rect 31205 2261 31217 2295
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 1104 2202 44040 2224
rect 1104 2150 11644 2202
rect 11696 2150 11708 2202
rect 11760 2150 11772 2202
rect 11824 2150 11836 2202
rect 11888 2150 11900 2202
rect 11952 2150 22338 2202
rect 22390 2150 22402 2202
rect 22454 2150 22466 2202
rect 22518 2150 22530 2202
rect 22582 2150 22594 2202
rect 22646 2150 33032 2202
rect 33084 2150 33096 2202
rect 33148 2150 33160 2202
rect 33212 2150 33224 2202
rect 33276 2150 33288 2202
rect 33340 2150 43726 2202
rect 43778 2150 43790 2202
rect 43842 2150 43854 2202
rect 43906 2150 43918 2202
rect 43970 2150 43982 2202
rect 44034 2150 44040 2202
rect 1104 2128 44040 2150
rect 1670 2048 1676 2100
rect 1728 2088 1734 2100
rect 1728 2060 9674 2088
rect 1728 2048 1734 2060
rect 9646 1952 9674 2060
rect 10042 2048 10048 2100
rect 10100 2088 10106 2100
rect 10100 2060 16574 2088
rect 10100 2048 10106 2060
rect 16546 2020 16574 2060
rect 26970 2048 26976 2100
rect 27028 2088 27034 2100
rect 36998 2088 37004 2100
rect 27028 2060 37004 2088
rect 27028 2048 27034 2060
rect 36998 2048 37004 2060
rect 37056 2048 37062 2100
rect 34882 2020 34888 2032
rect 16546 1992 34888 2020
rect 34882 1980 34888 1992
rect 34940 1980 34946 2032
rect 31754 1952 31760 1964
rect 9646 1924 31760 1952
rect 31754 1912 31760 1924
rect 31812 1912 31818 1964
<< via1 >>
rect 16396 8508 16448 8560
rect 32588 8508 32640 8560
rect 15844 8440 15896 8492
rect 33508 8440 33560 8492
rect 15476 8372 15528 8424
rect 33692 8372 33744 8424
rect 13360 8304 13412 8356
rect 36176 8304 36228 8356
rect 13820 8236 13872 8288
rect 14280 8236 14332 8288
rect 25320 8236 25372 8288
rect 25964 8236 26016 8288
rect 28816 8236 28868 8288
rect 29736 8236 29788 8288
rect 29920 8236 29972 8288
rect 30748 8236 30800 8288
rect 7748 8032 7800 8084
rect 23204 8168 23256 8220
rect 12440 8100 12492 8152
rect 16120 8100 16172 8152
rect 16304 8100 16356 8152
rect 19432 8100 19484 8152
rect 13636 8032 13688 8084
rect 22100 8032 22152 8084
rect 29184 8100 29236 8152
rect 30288 8100 30340 8152
rect 31208 8032 31260 8084
rect 11060 7964 11112 8016
rect 11796 7964 11848 8016
rect 12164 7964 12216 8016
rect 20720 7964 20772 8016
rect 23296 7964 23348 8016
rect 30656 7964 30708 8016
rect 14096 7896 14148 7948
rect 25320 7896 25372 7948
rect 26792 7896 26844 7948
rect 31392 7896 31444 7948
rect 31484 7896 31536 7948
rect 8392 7760 8444 7812
rect 20352 7828 20404 7880
rect 26884 7828 26936 7880
rect 32680 7828 32732 7880
rect 16304 7760 16356 7812
rect 22928 7760 22980 7812
rect 27436 7760 27488 7812
rect 28540 7760 28592 7812
rect 6736 7692 6788 7744
rect 21088 7692 21140 7744
rect 27252 7692 27304 7744
rect 28448 7692 28500 7744
rect 11644 7590 11696 7642
rect 11708 7590 11760 7642
rect 11772 7590 11824 7642
rect 11836 7590 11888 7642
rect 11900 7590 11952 7642
rect 22338 7590 22390 7642
rect 22402 7590 22454 7642
rect 22466 7590 22518 7642
rect 22530 7590 22582 7642
rect 22594 7590 22646 7642
rect 33032 7590 33084 7642
rect 33096 7590 33148 7642
rect 33160 7590 33212 7642
rect 33224 7590 33276 7642
rect 33288 7590 33340 7642
rect 43726 7590 43778 7642
rect 43790 7590 43842 7642
rect 43854 7590 43906 7642
rect 43918 7590 43970 7642
rect 43982 7590 44034 7642
rect 5448 7488 5500 7540
rect 6000 7488 6052 7540
rect 7380 7488 7432 7540
rect 7932 7488 7984 7540
rect 8484 7488 8536 7540
rect 9036 7488 9088 7540
rect 10692 7488 10744 7540
rect 11060 7488 11112 7540
rect 6736 7463 6788 7472
rect 6736 7429 6745 7463
rect 6745 7429 6779 7463
rect 6779 7429 6788 7463
rect 6736 7420 6788 7429
rect 5540 7352 5592 7404
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 8392 7463 8444 7472
rect 8392 7429 8401 7463
rect 8401 7429 8435 7463
rect 8435 7429 8444 7463
rect 8392 7420 8444 7429
rect 10048 7420 10100 7472
rect 6736 7284 6788 7336
rect 10600 7352 10652 7404
rect 12072 7488 12124 7540
rect 12164 7531 12216 7540
rect 12164 7497 12173 7531
rect 12173 7497 12207 7531
rect 12207 7497 12216 7531
rect 12164 7488 12216 7497
rect 13176 7488 13228 7540
rect 13728 7488 13780 7540
rect 13820 7531 13872 7540
rect 13820 7497 13829 7531
rect 13829 7497 13863 7531
rect 13863 7497 13872 7531
rect 13820 7488 13872 7497
rect 15108 7488 15160 7540
rect 15660 7488 15712 7540
rect 16212 7488 16264 7540
rect 16764 7488 16816 7540
rect 17316 7531 17368 7540
rect 17316 7497 17325 7531
rect 17325 7497 17359 7531
rect 17359 7497 17368 7531
rect 17316 7488 17368 7497
rect 17868 7531 17920 7540
rect 17868 7497 17877 7531
rect 17877 7497 17911 7531
rect 17911 7497 17920 7531
rect 17868 7488 17920 7497
rect 18420 7531 18472 7540
rect 18420 7497 18429 7531
rect 18429 7497 18463 7531
rect 18463 7497 18472 7531
rect 18420 7488 18472 7497
rect 14648 7420 14700 7472
rect 19156 7420 19208 7472
rect 21088 7488 21140 7540
rect 22928 7488 22980 7540
rect 20996 7420 21048 7472
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 13268 7352 13320 7404
rect 14188 7352 14240 7404
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 16580 7352 16632 7404
rect 17316 7352 17368 7404
rect 17868 7352 17920 7404
rect 18604 7352 18656 7404
rect 18972 7352 19024 7404
rect 6552 7216 6604 7268
rect 9680 7216 9732 7268
rect 11244 7216 11296 7268
rect 12072 7216 12124 7268
rect 12256 7216 12308 7268
rect 13636 7216 13688 7268
rect 14648 7216 14700 7268
rect 17684 7284 17736 7336
rect 19984 7395 20036 7404
rect 19984 7361 19993 7395
rect 19993 7361 20027 7395
rect 20027 7361 20036 7395
rect 19984 7352 20036 7361
rect 20812 7352 20864 7404
rect 21180 7352 21232 7404
rect 21364 7395 21416 7404
rect 21364 7361 21373 7395
rect 21373 7361 21407 7395
rect 21407 7361 21416 7395
rect 21364 7352 21416 7361
rect 21640 7395 21692 7404
rect 21640 7361 21649 7395
rect 21649 7361 21683 7395
rect 21683 7361 21692 7395
rect 21640 7352 21692 7361
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 22284 7395 22336 7404
rect 22284 7361 22293 7395
rect 22293 7361 22327 7395
rect 22327 7361 22336 7395
rect 22284 7352 22336 7361
rect 22836 7395 22888 7404
rect 22836 7361 22845 7395
rect 22845 7361 22879 7395
rect 22879 7361 22888 7395
rect 22836 7352 22888 7361
rect 23112 7395 23164 7404
rect 23112 7361 23121 7395
rect 23121 7361 23155 7395
rect 23155 7361 23164 7395
rect 23112 7352 23164 7361
rect 23388 7352 23440 7404
rect 23940 7395 23992 7404
rect 23940 7361 23949 7395
rect 23949 7361 23983 7395
rect 23983 7361 23992 7395
rect 23940 7352 23992 7361
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 25320 7488 25372 7540
rect 26148 7488 26200 7540
rect 24676 7420 24728 7472
rect 24492 7352 24544 7404
rect 25504 7420 25556 7472
rect 25872 7420 25924 7472
rect 16304 7148 16356 7200
rect 17408 7148 17460 7200
rect 18788 7191 18840 7200
rect 18788 7157 18797 7191
rect 18797 7157 18831 7191
rect 18831 7157 18840 7191
rect 18788 7148 18840 7157
rect 19248 7148 19300 7200
rect 20536 7216 20588 7268
rect 21916 7216 21968 7268
rect 23112 7216 23164 7268
rect 24584 7259 24636 7268
rect 24584 7225 24593 7259
rect 24593 7225 24627 7259
rect 24627 7225 24636 7259
rect 24584 7216 24636 7225
rect 24768 7216 24820 7268
rect 21456 7191 21508 7200
rect 21456 7157 21465 7191
rect 21465 7157 21499 7191
rect 21499 7157 21508 7191
rect 21456 7148 21508 7157
rect 21824 7191 21876 7200
rect 21824 7157 21833 7191
rect 21833 7157 21867 7191
rect 21867 7157 21876 7191
rect 21824 7148 21876 7157
rect 22100 7191 22152 7200
rect 22100 7157 22109 7191
rect 22109 7157 22143 7191
rect 22143 7157 22152 7191
rect 22100 7148 22152 7157
rect 22928 7191 22980 7200
rect 22928 7157 22937 7191
rect 22937 7157 22971 7191
rect 22971 7157 22980 7191
rect 22928 7148 22980 7157
rect 23480 7191 23532 7200
rect 23480 7157 23489 7191
rect 23489 7157 23523 7191
rect 23523 7157 23532 7191
rect 23480 7148 23532 7157
rect 24032 7191 24084 7200
rect 24032 7157 24041 7191
rect 24041 7157 24075 7191
rect 24075 7157 24084 7191
rect 24032 7148 24084 7157
rect 25136 7191 25188 7200
rect 25136 7157 25145 7191
rect 25145 7157 25179 7191
rect 25179 7157 25188 7191
rect 25136 7148 25188 7157
rect 25964 7352 26016 7404
rect 27068 7488 27120 7540
rect 28356 7488 28408 7540
rect 26976 7420 27028 7472
rect 27896 7420 27948 7472
rect 25872 7284 25924 7336
rect 26700 7284 26752 7336
rect 27528 7284 27580 7336
rect 28448 7352 28500 7404
rect 28540 7395 28592 7404
rect 28540 7361 28549 7395
rect 28549 7361 28583 7395
rect 28583 7361 28592 7395
rect 28540 7352 28592 7361
rect 29460 7488 29512 7540
rect 28356 7284 28408 7336
rect 29736 7395 29788 7404
rect 29736 7361 29745 7395
rect 29745 7361 29779 7395
rect 29779 7361 29788 7395
rect 29736 7352 29788 7361
rect 27436 7216 27488 7268
rect 28816 7216 28868 7268
rect 30288 7395 30340 7404
rect 30288 7361 30297 7395
rect 30297 7361 30331 7395
rect 30331 7361 30340 7395
rect 30288 7352 30340 7361
rect 30472 7488 30524 7540
rect 30748 7352 30800 7404
rect 31392 7531 31444 7540
rect 31392 7497 31401 7531
rect 31401 7497 31435 7531
rect 31435 7497 31444 7531
rect 31392 7488 31444 7497
rect 31484 7488 31536 7540
rect 32496 7488 32548 7540
rect 31300 7420 31352 7472
rect 30196 7284 30248 7336
rect 31484 7395 31536 7404
rect 31484 7361 31493 7395
rect 31493 7361 31527 7395
rect 31527 7361 31536 7395
rect 31484 7352 31536 7361
rect 32220 7420 32272 7472
rect 33508 7488 33560 7540
rect 33692 7531 33744 7540
rect 33692 7497 33701 7531
rect 33701 7497 33735 7531
rect 33735 7497 33744 7531
rect 33692 7488 33744 7497
rect 33876 7488 33928 7540
rect 34612 7488 34664 7540
rect 34704 7420 34756 7472
rect 35716 7488 35768 7540
rect 37096 7488 37148 7540
rect 39120 7488 39172 7540
rect 36176 7420 36228 7472
rect 36820 7420 36872 7472
rect 31024 7284 31076 7336
rect 31852 7284 31904 7336
rect 25872 7148 25924 7200
rect 26056 7191 26108 7200
rect 26056 7157 26065 7191
rect 26065 7157 26099 7191
rect 26099 7157 26108 7191
rect 26056 7148 26108 7157
rect 26148 7148 26200 7200
rect 26608 7191 26660 7200
rect 26608 7157 26617 7191
rect 26617 7157 26651 7191
rect 26651 7157 26660 7191
rect 26608 7148 26660 7157
rect 27252 7191 27304 7200
rect 27252 7157 27261 7191
rect 27261 7157 27295 7191
rect 27295 7157 27304 7191
rect 27252 7148 27304 7157
rect 27528 7191 27580 7200
rect 27528 7157 27537 7191
rect 27537 7157 27571 7191
rect 27571 7157 27580 7191
rect 27528 7148 27580 7157
rect 28356 7191 28408 7200
rect 28356 7157 28365 7191
rect 28365 7157 28399 7191
rect 28399 7157 28408 7191
rect 28356 7148 28408 7157
rect 28632 7191 28684 7200
rect 28632 7157 28641 7191
rect 28641 7157 28675 7191
rect 28675 7157 28684 7191
rect 28632 7148 28684 7157
rect 28908 7191 28960 7200
rect 28908 7157 28917 7191
rect 28917 7157 28951 7191
rect 28951 7157 28960 7191
rect 28908 7148 28960 7157
rect 29092 7148 29144 7200
rect 30564 7216 30616 7268
rect 31484 7216 31536 7268
rect 31944 7216 31996 7268
rect 32588 7284 32640 7336
rect 32864 7284 32916 7336
rect 33692 7352 33744 7404
rect 34796 7395 34848 7404
rect 34796 7361 34805 7395
rect 34805 7361 34839 7395
rect 34839 7361 34848 7395
rect 34796 7352 34848 7361
rect 35348 7395 35400 7404
rect 35348 7361 35357 7395
rect 35357 7361 35391 7395
rect 35391 7361 35400 7395
rect 35348 7352 35400 7361
rect 35900 7395 35952 7404
rect 35900 7361 35909 7395
rect 35909 7361 35943 7395
rect 35943 7361 35952 7395
rect 35900 7352 35952 7361
rect 35716 7284 35768 7336
rect 37556 7352 37608 7404
rect 37924 7395 37976 7404
rect 37924 7361 37933 7395
rect 37933 7361 37967 7395
rect 37967 7361 37976 7395
rect 37924 7352 37976 7361
rect 39028 7395 39080 7404
rect 39028 7361 39037 7395
rect 39037 7361 39071 7395
rect 39071 7361 39080 7395
rect 39028 7352 39080 7361
rect 39672 7395 39724 7404
rect 39672 7361 39681 7395
rect 39681 7361 39715 7395
rect 39715 7361 39724 7395
rect 39672 7352 39724 7361
rect 37832 7284 37884 7336
rect 41420 7395 41472 7404
rect 41420 7361 41429 7395
rect 41429 7361 41463 7395
rect 41463 7361 41472 7395
rect 41420 7352 41472 7361
rect 43352 7284 43404 7336
rect 36544 7216 36596 7268
rect 29552 7191 29604 7200
rect 29552 7157 29561 7191
rect 29561 7157 29595 7191
rect 29595 7157 29604 7191
rect 29552 7148 29604 7157
rect 29828 7191 29880 7200
rect 29828 7157 29837 7191
rect 29837 7157 29871 7191
rect 29871 7157 29880 7191
rect 29828 7148 29880 7157
rect 30104 7191 30156 7200
rect 30104 7157 30113 7191
rect 30113 7157 30147 7191
rect 30147 7157 30156 7191
rect 30104 7148 30156 7157
rect 30380 7191 30432 7200
rect 30380 7157 30389 7191
rect 30389 7157 30423 7191
rect 30423 7157 30432 7191
rect 30380 7148 30432 7157
rect 30656 7148 30708 7200
rect 30932 7148 30984 7200
rect 31208 7148 31260 7200
rect 32312 7191 32364 7200
rect 32312 7157 32321 7191
rect 32321 7157 32355 7191
rect 32355 7157 32364 7191
rect 32312 7148 32364 7157
rect 32588 7191 32640 7200
rect 32588 7157 32597 7191
rect 32597 7157 32631 7191
rect 32631 7157 32640 7191
rect 32588 7148 32640 7157
rect 32680 7148 32732 7200
rect 35164 7148 35216 7200
rect 36912 7191 36964 7200
rect 36912 7157 36921 7191
rect 36921 7157 36955 7191
rect 36955 7157 36964 7191
rect 36912 7148 36964 7157
rect 39580 7216 39632 7268
rect 38752 7191 38804 7200
rect 38752 7157 38761 7191
rect 38761 7157 38795 7191
rect 38795 7157 38804 7191
rect 38752 7148 38804 7157
rect 39120 7191 39172 7200
rect 39120 7157 39129 7191
rect 39129 7157 39163 7191
rect 39163 7157 39172 7191
rect 39120 7148 39172 7157
rect 39488 7191 39540 7200
rect 39488 7157 39497 7191
rect 39497 7157 39531 7191
rect 39531 7157 39540 7191
rect 39488 7148 39540 7157
rect 40960 7191 41012 7200
rect 40960 7157 40969 7191
rect 40969 7157 41003 7191
rect 41003 7157 41012 7191
rect 40960 7148 41012 7157
rect 6297 7046 6349 7098
rect 6361 7046 6413 7098
rect 6425 7046 6477 7098
rect 6489 7046 6541 7098
rect 6553 7046 6605 7098
rect 16991 7046 17043 7098
rect 17055 7046 17107 7098
rect 17119 7046 17171 7098
rect 17183 7046 17235 7098
rect 17247 7046 17299 7098
rect 27685 7046 27737 7098
rect 27749 7046 27801 7098
rect 27813 7046 27865 7098
rect 27877 7046 27929 7098
rect 27941 7046 27993 7098
rect 38379 7046 38431 7098
rect 38443 7046 38495 7098
rect 38507 7046 38559 7098
rect 38571 7046 38623 7098
rect 38635 7046 38687 7098
rect 5172 6987 5224 6996
rect 5172 6953 5181 6987
rect 5181 6953 5215 6987
rect 5215 6953 5224 6987
rect 5172 6944 5224 6953
rect 5724 6987 5776 6996
rect 5724 6953 5733 6987
rect 5733 6953 5767 6987
rect 5767 6953 5776 6987
rect 5724 6944 5776 6953
rect 6828 6987 6880 6996
rect 6828 6953 6837 6987
rect 6837 6953 6871 6987
rect 6871 6953 6880 6987
rect 6828 6944 6880 6953
rect 7288 6944 7340 6996
rect 12256 6944 12308 6996
rect 13084 6987 13136 6996
rect 13084 6953 13093 6987
rect 13093 6953 13127 6987
rect 13127 6953 13136 6987
rect 13084 6944 13136 6953
rect 13636 6987 13688 6996
rect 13636 6953 13645 6987
rect 13645 6953 13679 6987
rect 13679 6953 13688 6987
rect 13636 6944 13688 6953
rect 14188 6944 14240 6996
rect 14556 6987 14608 6996
rect 14556 6953 14565 6987
rect 14565 6953 14599 6987
rect 14599 6953 14608 6987
rect 14556 6944 14608 6953
rect 16304 6944 16356 6996
rect 17960 6944 18012 6996
rect 19984 6944 20036 6996
rect 20444 6944 20496 6996
rect 21456 6944 21508 6996
rect 7104 6808 7156 6860
rect 7656 6808 7708 6860
rect 8208 6808 8260 6860
rect 6644 6740 6696 6792
rect 7748 6740 7800 6792
rect 9404 6876 9456 6928
rect 20260 6876 20312 6928
rect 20352 6876 20404 6928
rect 10140 6808 10192 6860
rect 10508 6851 10560 6860
rect 10508 6817 10517 6851
rect 10517 6817 10551 6851
rect 10551 6817 10560 6851
rect 10508 6808 10560 6817
rect 10968 6808 11020 6860
rect 11612 6851 11664 6860
rect 11612 6817 11621 6851
rect 11621 6817 11655 6851
rect 11655 6817 11664 6851
rect 11612 6808 11664 6817
rect 12348 6808 12400 6860
rect 14832 6808 14884 6860
rect 15384 6808 15436 6860
rect 15936 6808 15988 6860
rect 16488 6808 16540 6860
rect 17040 6808 17092 6860
rect 17592 6808 17644 6860
rect 18144 6808 18196 6860
rect 9404 6740 9456 6792
rect 9496 6740 9548 6792
rect 11152 6740 11204 6792
rect 12624 6740 12676 6792
rect 5632 6715 5684 6724
rect 5632 6681 5641 6715
rect 5641 6681 5675 6715
rect 5675 6681 5684 6715
rect 5632 6672 5684 6681
rect 6092 6604 6144 6656
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 9864 6604 9916 6656
rect 10692 6672 10744 6724
rect 10784 6715 10836 6724
rect 10784 6681 10793 6715
rect 10793 6681 10827 6715
rect 10827 6681 10836 6715
rect 10784 6672 10836 6681
rect 11336 6715 11388 6724
rect 11336 6681 11345 6715
rect 11345 6681 11379 6715
rect 11379 6681 11388 6715
rect 11336 6672 11388 6681
rect 12072 6604 12124 6656
rect 14188 6740 14240 6792
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 12992 6715 13044 6724
rect 12992 6681 13001 6715
rect 13001 6681 13035 6715
rect 13035 6681 13044 6715
rect 12992 6672 13044 6681
rect 13912 6672 13964 6724
rect 14740 6672 14792 6724
rect 13728 6604 13780 6656
rect 16304 6740 16356 6792
rect 19064 6783 19116 6792
rect 19064 6749 19073 6783
rect 19073 6749 19107 6783
rect 19107 6749 19116 6783
rect 19064 6740 19116 6749
rect 19340 6783 19392 6792
rect 19340 6749 19349 6783
rect 19349 6749 19383 6783
rect 19383 6749 19392 6783
rect 19340 6740 19392 6749
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 19892 6783 19944 6792
rect 19892 6749 19901 6783
rect 19901 6749 19935 6783
rect 19935 6749 19944 6783
rect 19892 6740 19944 6749
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 15016 6715 15068 6724
rect 15016 6681 15025 6715
rect 15025 6681 15059 6715
rect 15059 6681 15068 6715
rect 15016 6672 15068 6681
rect 15292 6672 15344 6724
rect 16672 6715 16724 6724
rect 16672 6681 16681 6715
rect 16681 6681 16715 6715
rect 16715 6681 16724 6715
rect 16672 6672 16724 6681
rect 17224 6715 17276 6724
rect 17224 6681 17233 6715
rect 17233 6681 17267 6715
rect 17267 6681 17276 6715
rect 17224 6672 17276 6681
rect 17408 6672 17460 6724
rect 18328 6715 18380 6724
rect 18328 6681 18337 6715
rect 18337 6681 18371 6715
rect 18371 6681 18380 6715
rect 18328 6672 18380 6681
rect 18420 6672 18472 6724
rect 18512 6604 18564 6656
rect 19432 6604 19484 6656
rect 19524 6647 19576 6656
rect 19524 6613 19533 6647
rect 19533 6613 19567 6647
rect 19567 6613 19576 6647
rect 19524 6604 19576 6613
rect 19800 6647 19852 6656
rect 19800 6613 19809 6647
rect 19809 6613 19843 6647
rect 19843 6613 19852 6647
rect 19800 6604 19852 6613
rect 20536 6740 20588 6792
rect 20628 6740 20680 6792
rect 22100 6808 22152 6860
rect 21824 6740 21876 6792
rect 22008 6740 22060 6792
rect 22836 6783 22888 6792
rect 22836 6749 22845 6783
rect 22845 6749 22879 6783
rect 22879 6749 22888 6783
rect 22836 6740 22888 6749
rect 24032 6740 24084 6792
rect 26148 6944 26200 6996
rect 26424 6987 26476 6996
rect 26424 6953 26433 6987
rect 26433 6953 26467 6987
rect 26467 6953 26476 6987
rect 26424 6944 26476 6953
rect 26608 6944 26660 6996
rect 27252 6944 27304 6996
rect 28356 6944 28408 6996
rect 28632 6944 28684 6996
rect 36912 6944 36964 6996
rect 26056 6740 26108 6792
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 20904 6647 20956 6656
rect 20904 6613 20913 6647
rect 20913 6613 20947 6647
rect 20947 6613 20956 6647
rect 20904 6604 20956 6613
rect 21180 6647 21232 6656
rect 21180 6613 21189 6647
rect 21189 6613 21223 6647
rect 21223 6613 21232 6647
rect 21180 6604 21232 6613
rect 21272 6604 21324 6656
rect 26148 6672 26200 6724
rect 27068 6740 27120 6792
rect 27436 6740 27488 6792
rect 38108 6876 38160 6928
rect 33600 6808 33652 6860
rect 28816 6740 28868 6792
rect 28908 6740 28960 6792
rect 29552 6740 29604 6792
rect 29828 6740 29880 6792
rect 30104 6740 30156 6792
rect 30380 6740 30432 6792
rect 31208 6783 31260 6792
rect 31208 6749 31217 6783
rect 31217 6749 31251 6783
rect 31251 6749 31260 6783
rect 31208 6740 31260 6749
rect 31760 6740 31812 6792
rect 32956 6740 33008 6792
rect 33416 6783 33468 6792
rect 33416 6749 33425 6783
rect 33425 6749 33459 6783
rect 33459 6749 33468 6783
rect 33416 6740 33468 6749
rect 33692 6740 33744 6792
rect 33876 6783 33928 6792
rect 33876 6749 33885 6783
rect 33885 6749 33919 6783
rect 33919 6749 33928 6783
rect 33876 6740 33928 6749
rect 34060 6740 34112 6792
rect 35256 6808 35308 6860
rect 35808 6808 35860 6860
rect 37188 6808 37240 6860
rect 38568 6876 38620 6928
rect 38936 6876 38988 6928
rect 39120 6808 39172 6860
rect 35164 6783 35216 6792
rect 35164 6749 35173 6783
rect 35173 6749 35207 6783
rect 35207 6749 35216 6783
rect 35164 6740 35216 6749
rect 37464 6740 37516 6792
rect 38660 6740 38712 6792
rect 39856 6808 39908 6860
rect 39488 6740 39540 6792
rect 40960 6740 41012 6792
rect 23388 6604 23440 6656
rect 25320 6647 25372 6656
rect 25320 6613 25329 6647
rect 25329 6613 25363 6647
rect 25363 6613 25372 6647
rect 25320 6604 25372 6613
rect 25596 6647 25648 6656
rect 25596 6613 25605 6647
rect 25605 6613 25639 6647
rect 25639 6613 25648 6647
rect 25596 6604 25648 6613
rect 26976 6647 27028 6656
rect 26976 6613 26985 6647
rect 26985 6613 27019 6647
rect 27019 6613 27028 6647
rect 26976 6604 27028 6613
rect 27344 6647 27396 6656
rect 27344 6613 27353 6647
rect 27353 6613 27387 6647
rect 27387 6613 27396 6647
rect 27344 6604 27396 6613
rect 27528 6604 27580 6656
rect 27620 6604 27672 6656
rect 28080 6647 28132 6656
rect 28080 6613 28089 6647
rect 28089 6613 28123 6647
rect 28123 6613 28132 6647
rect 28080 6604 28132 6613
rect 28448 6647 28500 6656
rect 28448 6613 28457 6647
rect 28457 6613 28491 6647
rect 28491 6613 28500 6647
rect 28448 6604 28500 6613
rect 28908 6647 28960 6656
rect 28908 6613 28917 6647
rect 28917 6613 28951 6647
rect 28951 6613 28960 6647
rect 28908 6604 28960 6613
rect 29368 6647 29420 6656
rect 29368 6613 29377 6647
rect 29377 6613 29411 6647
rect 29411 6613 29420 6647
rect 29368 6604 29420 6613
rect 29828 6647 29880 6656
rect 29828 6613 29837 6647
rect 29837 6613 29871 6647
rect 29871 6613 29880 6647
rect 29828 6604 29880 6613
rect 30196 6647 30248 6656
rect 30196 6613 30205 6647
rect 30205 6613 30239 6647
rect 30239 6613 30248 6647
rect 30196 6604 30248 6613
rect 30288 6604 30340 6656
rect 31392 6647 31444 6656
rect 31392 6613 31401 6647
rect 31401 6613 31435 6647
rect 31435 6613 31444 6647
rect 31392 6604 31444 6613
rect 35440 6715 35492 6724
rect 35440 6681 35449 6715
rect 35449 6681 35483 6715
rect 35483 6681 35492 6715
rect 35440 6672 35492 6681
rect 35992 6715 36044 6724
rect 35992 6681 36001 6715
rect 36001 6681 36035 6715
rect 36035 6681 36044 6715
rect 35992 6672 36044 6681
rect 36544 6715 36596 6724
rect 36544 6681 36553 6715
rect 36553 6681 36587 6715
rect 36587 6681 36596 6715
rect 36544 6672 36596 6681
rect 37096 6715 37148 6724
rect 37096 6681 37105 6715
rect 37105 6681 37139 6715
rect 37139 6681 37148 6715
rect 37096 6672 37148 6681
rect 37648 6715 37700 6724
rect 37648 6681 37657 6715
rect 37657 6681 37691 6715
rect 37691 6681 37700 6715
rect 37648 6672 37700 6681
rect 38200 6715 38252 6724
rect 38200 6681 38209 6715
rect 38209 6681 38243 6715
rect 38243 6681 38252 6715
rect 38200 6672 38252 6681
rect 38384 6672 38436 6724
rect 39212 6672 39264 6724
rect 33324 6647 33376 6656
rect 33324 6613 33333 6647
rect 33333 6613 33367 6647
rect 33367 6613 33376 6647
rect 33324 6604 33376 6613
rect 33600 6647 33652 6656
rect 33600 6613 33609 6647
rect 33609 6613 33643 6647
rect 33643 6613 33652 6647
rect 33600 6604 33652 6613
rect 33692 6647 33744 6656
rect 33692 6613 33701 6647
rect 33701 6613 33735 6647
rect 33735 6613 33744 6647
rect 33692 6604 33744 6613
rect 33968 6647 34020 6656
rect 33968 6613 33977 6647
rect 33977 6613 34011 6647
rect 34011 6613 34020 6647
rect 33968 6604 34020 6613
rect 34152 6604 34204 6656
rect 34428 6647 34480 6656
rect 34428 6613 34437 6647
rect 34437 6613 34471 6647
rect 34471 6613 34480 6647
rect 34428 6604 34480 6613
rect 35900 6604 35952 6656
rect 36084 6604 36136 6656
rect 36728 6604 36780 6656
rect 37740 6604 37792 6656
rect 38476 6604 38528 6656
rect 38936 6604 38988 6656
rect 11644 6502 11696 6554
rect 11708 6502 11760 6554
rect 11772 6502 11824 6554
rect 11836 6502 11888 6554
rect 11900 6502 11952 6554
rect 22338 6502 22390 6554
rect 22402 6502 22454 6554
rect 22466 6502 22518 6554
rect 22530 6502 22582 6554
rect 22594 6502 22646 6554
rect 33032 6502 33084 6554
rect 33096 6502 33148 6554
rect 33160 6502 33212 6554
rect 33224 6502 33276 6554
rect 33288 6502 33340 6554
rect 43726 6502 43778 6554
rect 43790 6502 43842 6554
rect 43854 6502 43906 6554
rect 43918 6502 43970 6554
rect 43982 6502 44034 6554
rect 5632 6400 5684 6452
rect 6092 6400 6144 6452
rect 8668 6443 8720 6452
rect 8668 6409 8677 6443
rect 8677 6409 8711 6443
rect 8711 6409 8720 6443
rect 8668 6400 8720 6409
rect 9220 6443 9272 6452
rect 9220 6409 9229 6443
rect 9229 6409 9263 6443
rect 9263 6409 9272 6443
rect 9220 6400 9272 6409
rect 9772 6443 9824 6452
rect 9772 6409 9781 6443
rect 9781 6409 9815 6443
rect 9815 6409 9824 6443
rect 9772 6400 9824 6409
rect 6184 6307 6236 6316
rect 6184 6273 6193 6307
rect 6193 6273 6227 6307
rect 6227 6273 6236 6307
rect 6184 6264 6236 6273
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 9680 6375 9732 6384
rect 9680 6341 9689 6375
rect 9689 6341 9723 6375
rect 9723 6341 9732 6375
rect 9680 6332 9732 6341
rect 10508 6400 10560 6452
rect 10692 6400 10744 6452
rect 11980 6443 12032 6452
rect 11980 6409 11989 6443
rect 11989 6409 12023 6443
rect 12023 6409 12032 6443
rect 11980 6400 12032 6409
rect 13636 6332 13688 6384
rect 14004 6400 14056 6452
rect 14464 6400 14516 6452
rect 14740 6400 14792 6452
rect 15016 6332 15068 6384
rect 15292 6443 15344 6452
rect 15292 6409 15301 6443
rect 15301 6409 15335 6443
rect 15335 6409 15344 6443
rect 15292 6400 15344 6409
rect 15568 6400 15620 6452
rect 16672 6400 16724 6452
rect 17224 6400 17276 6452
rect 17868 6400 17920 6452
rect 18328 6443 18380 6452
rect 18328 6409 18337 6443
rect 18337 6409 18371 6443
rect 18371 6409 18380 6443
rect 18328 6400 18380 6409
rect 18604 6443 18656 6452
rect 18604 6409 18613 6443
rect 18613 6409 18647 6443
rect 18647 6409 18656 6443
rect 18604 6400 18656 6409
rect 18972 6443 19024 6452
rect 18972 6409 18981 6443
rect 18981 6409 19015 6443
rect 19015 6409 19024 6443
rect 18972 6400 19024 6409
rect 19064 6400 19116 6452
rect 19340 6400 19392 6452
rect 22008 6400 22060 6452
rect 22192 6400 22244 6452
rect 18144 6332 18196 6384
rect 5540 6196 5592 6248
rect 11060 6307 11112 6316
rect 11060 6273 11069 6307
rect 11069 6273 11103 6307
rect 11103 6273 11112 6307
rect 11060 6264 11112 6273
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 14096 6264 14148 6316
rect 14832 6307 14884 6316
rect 14832 6273 14841 6307
rect 14841 6273 14875 6307
rect 14875 6273 14884 6307
rect 14832 6264 14884 6273
rect 15476 6307 15528 6316
rect 15476 6273 15485 6307
rect 15485 6273 15519 6307
rect 15519 6273 15528 6307
rect 15476 6264 15528 6273
rect 15844 6307 15896 6316
rect 15844 6273 15853 6307
rect 15853 6273 15887 6307
rect 15887 6273 15896 6307
rect 15844 6264 15896 6273
rect 16396 6264 16448 6316
rect 17408 6264 17460 6316
rect 17500 6307 17552 6316
rect 17500 6273 17509 6307
rect 17509 6273 17543 6307
rect 17543 6273 17552 6307
rect 17500 6264 17552 6273
rect 17776 6307 17828 6316
rect 17776 6273 17785 6307
rect 17785 6273 17819 6307
rect 17819 6273 17828 6307
rect 17776 6264 17828 6273
rect 18236 6307 18288 6316
rect 18236 6273 18245 6307
rect 18245 6273 18279 6307
rect 18279 6273 18288 6307
rect 18236 6264 18288 6273
rect 18512 6307 18564 6316
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 18788 6307 18840 6316
rect 18788 6273 18797 6307
rect 18797 6273 18831 6307
rect 18831 6273 18840 6307
rect 18788 6264 18840 6273
rect 9404 6128 9456 6180
rect 9312 6060 9364 6112
rect 10416 6060 10468 6112
rect 13636 6060 13688 6112
rect 17868 6196 17920 6248
rect 20444 6307 20496 6316
rect 20444 6273 20453 6307
rect 20453 6273 20487 6307
rect 20487 6273 20496 6307
rect 20444 6264 20496 6273
rect 21916 6264 21968 6316
rect 22100 6196 22152 6248
rect 22928 6400 22980 6452
rect 25964 6400 26016 6452
rect 27344 6400 27396 6452
rect 33692 6400 33744 6452
rect 34796 6400 34848 6452
rect 38200 6400 38252 6452
rect 38384 6400 38436 6452
rect 30932 6332 30984 6384
rect 33968 6332 34020 6384
rect 23480 6264 23532 6316
rect 25872 6264 25924 6316
rect 34244 6307 34296 6316
rect 34244 6273 34253 6307
rect 34253 6273 34287 6307
rect 34287 6273 34296 6307
rect 34244 6264 34296 6273
rect 23112 6196 23164 6248
rect 30288 6196 30340 6248
rect 30380 6196 30432 6248
rect 37096 6264 37148 6316
rect 37280 6264 37332 6316
rect 36728 6196 36780 6248
rect 39028 6196 39080 6248
rect 16580 6128 16632 6180
rect 17316 6171 17368 6180
rect 17316 6137 17325 6171
rect 17325 6137 17359 6171
rect 17359 6137 17368 6171
rect 17316 6128 17368 6137
rect 17408 6128 17460 6180
rect 20904 6128 20956 6180
rect 20720 6060 20772 6112
rect 25320 6128 25372 6180
rect 22008 6103 22060 6112
rect 22008 6069 22017 6103
rect 22017 6069 22051 6103
rect 22051 6069 22060 6103
rect 22008 6060 22060 6069
rect 23020 6060 23072 6112
rect 24032 6060 24084 6112
rect 35348 6060 35400 6112
rect 6297 5958 6349 6010
rect 6361 5958 6413 6010
rect 6425 5958 6477 6010
rect 6489 5958 6541 6010
rect 6553 5958 6605 6010
rect 16991 5958 17043 6010
rect 17055 5958 17107 6010
rect 17119 5958 17171 6010
rect 17183 5958 17235 6010
rect 17247 5958 17299 6010
rect 27685 5958 27737 6010
rect 27749 5958 27801 6010
rect 27813 5958 27865 6010
rect 27877 5958 27929 6010
rect 27941 5958 27993 6010
rect 38379 5958 38431 6010
rect 38443 5958 38495 6010
rect 38507 5958 38559 6010
rect 38571 5958 38623 6010
rect 38635 5958 38687 6010
rect 6184 5856 6236 5908
rect 8024 5856 8076 5908
rect 10416 5856 10468 5908
rect 11704 5856 11756 5908
rect 13360 5856 13412 5908
rect 13636 5856 13688 5908
rect 16304 5856 16356 5908
rect 17408 5856 17460 5908
rect 18236 5856 18288 5908
rect 20812 5856 20864 5908
rect 29368 5856 29420 5908
rect 19800 5720 19852 5772
rect 22192 5788 22244 5840
rect 23296 5788 23348 5840
rect 26976 5788 27028 5840
rect 23204 5720 23256 5772
rect 11060 5652 11112 5704
rect 12808 5695 12860 5704
rect 12808 5661 12817 5695
rect 12817 5661 12851 5695
rect 12851 5661 12860 5695
rect 12808 5652 12860 5661
rect 12992 5652 13044 5704
rect 16488 5584 16540 5636
rect 17500 5584 17552 5636
rect 32312 5584 32364 5636
rect 8576 5516 8628 5568
rect 12072 5516 12124 5568
rect 17684 5516 17736 5568
rect 31392 5516 31444 5568
rect 11644 5414 11696 5466
rect 11708 5414 11760 5466
rect 11772 5414 11824 5466
rect 11836 5414 11888 5466
rect 11900 5414 11952 5466
rect 22338 5414 22390 5466
rect 22402 5414 22454 5466
rect 22466 5414 22518 5466
rect 22530 5414 22582 5466
rect 22594 5414 22646 5466
rect 33032 5414 33084 5466
rect 33096 5414 33148 5466
rect 33160 5414 33212 5466
rect 33224 5414 33276 5466
rect 33288 5414 33340 5466
rect 43726 5414 43778 5466
rect 43790 5414 43842 5466
rect 43854 5414 43906 5466
rect 43918 5414 43970 5466
rect 43982 5414 44034 5466
rect 18144 5312 18196 5364
rect 23388 5312 23440 5364
rect 13728 5244 13780 5296
rect 25964 5244 26016 5296
rect 20444 5176 20496 5228
rect 11980 5108 12032 5160
rect 28080 5108 28132 5160
rect 14188 5040 14240 5092
rect 27620 5040 27672 5092
rect 6736 4972 6788 5024
rect 19524 4972 19576 5024
rect 30380 4972 30432 5024
rect 6297 4870 6349 4922
rect 6361 4870 6413 4922
rect 6425 4870 6477 4922
rect 6489 4870 6541 4922
rect 6553 4870 6605 4922
rect 16991 4870 17043 4922
rect 17055 4870 17107 4922
rect 17119 4870 17171 4922
rect 17183 4870 17235 4922
rect 17247 4870 17299 4922
rect 27685 4870 27737 4922
rect 27749 4870 27801 4922
rect 27813 4870 27865 4922
rect 27877 4870 27929 4922
rect 27941 4870 27993 4922
rect 38379 4870 38431 4922
rect 38443 4870 38495 4922
rect 38507 4870 38559 4922
rect 38571 4870 38623 4922
rect 38635 4870 38687 4922
rect 10600 4768 10652 4820
rect 30196 4768 30248 4820
rect 10784 4700 10836 4752
rect 29828 4700 29880 4752
rect 13912 4632 13964 4684
rect 26424 4632 26476 4684
rect 11336 4564 11388 4616
rect 28908 4564 28960 4616
rect 33416 4564 33468 4616
rect 36544 4564 36596 4616
rect 11644 4326 11696 4378
rect 11708 4326 11760 4378
rect 11772 4326 11824 4378
rect 11836 4326 11888 4378
rect 11900 4326 11952 4378
rect 22338 4326 22390 4378
rect 22402 4326 22454 4378
rect 22466 4326 22518 4378
rect 22530 4326 22582 4378
rect 22594 4326 22646 4378
rect 33032 4326 33084 4378
rect 33096 4326 33148 4378
rect 33160 4326 33212 4378
rect 33224 4326 33276 4378
rect 33288 4326 33340 4378
rect 43726 4326 43778 4378
rect 43790 4326 43842 4378
rect 43854 4326 43906 4378
rect 43918 4326 43970 4378
rect 43982 4326 44034 4378
rect 6297 3782 6349 3834
rect 6361 3782 6413 3834
rect 6425 3782 6477 3834
rect 6489 3782 6541 3834
rect 6553 3782 6605 3834
rect 16991 3782 17043 3834
rect 17055 3782 17107 3834
rect 17119 3782 17171 3834
rect 17183 3782 17235 3834
rect 17247 3782 17299 3834
rect 27685 3782 27737 3834
rect 27749 3782 27801 3834
rect 27813 3782 27865 3834
rect 27877 3782 27929 3834
rect 27941 3782 27993 3834
rect 38379 3782 38431 3834
rect 38443 3782 38495 3834
rect 38507 3782 38559 3834
rect 38571 3782 38623 3834
rect 38635 3782 38687 3834
rect 10968 3476 11020 3528
rect 35164 3476 35216 3528
rect 6644 3408 6696 3460
rect 34244 3408 34296 3460
rect 11644 3238 11696 3290
rect 11708 3238 11760 3290
rect 11772 3238 11824 3290
rect 11836 3238 11888 3290
rect 11900 3238 11952 3290
rect 22338 3238 22390 3290
rect 22402 3238 22454 3290
rect 22466 3238 22518 3290
rect 22530 3238 22582 3290
rect 22594 3238 22646 3290
rect 33032 3238 33084 3290
rect 33096 3238 33148 3290
rect 33160 3238 33212 3290
rect 33224 3238 33276 3290
rect 33288 3238 33340 3290
rect 43726 3238 43778 3290
rect 43790 3238 43842 3290
rect 43854 3238 43906 3290
rect 43918 3238 43970 3290
rect 43982 3238 44034 3290
rect 37556 3068 37608 3120
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 18696 3000 18748 3009
rect 22928 3043 22980 3052
rect 22928 3009 22937 3043
rect 22937 3009 22971 3043
rect 22971 3009 22980 3043
rect 22928 3000 22980 3009
rect 25044 3043 25096 3052
rect 25044 3009 25053 3043
rect 25053 3009 25087 3043
rect 25087 3009 25096 3043
rect 25044 3000 25096 3009
rect 33140 2932 33192 2984
rect 35992 2932 36044 2984
rect 37924 2864 37976 2916
rect 37648 2796 37700 2848
rect 6297 2694 6349 2746
rect 6361 2694 6413 2746
rect 6425 2694 6477 2746
rect 6489 2694 6541 2746
rect 6553 2694 6605 2746
rect 16991 2694 17043 2746
rect 17055 2694 17107 2746
rect 17119 2694 17171 2746
rect 17183 2694 17235 2746
rect 17247 2694 17299 2746
rect 27685 2694 27737 2746
rect 27749 2694 27801 2746
rect 27813 2694 27865 2746
rect 27877 2694 27929 2746
rect 27941 2694 27993 2746
rect 38379 2694 38431 2746
rect 38443 2694 38495 2746
rect 38507 2694 38559 2746
rect 38571 2694 38623 2746
rect 38635 2694 38687 2746
rect 6920 2592 6972 2644
rect 12808 2592 12860 2644
rect 18696 2592 18748 2644
rect 20444 2635 20496 2644
rect 20444 2601 20453 2635
rect 20453 2601 20487 2635
rect 20487 2601 20496 2635
rect 20444 2592 20496 2601
rect 22928 2592 22980 2644
rect 25044 2592 25096 2644
rect 34060 2592 34112 2644
rect 35440 2592 35492 2644
rect 35716 2592 35768 2644
rect 36820 2635 36872 2644
rect 36820 2601 36829 2635
rect 36829 2601 36863 2635
rect 36863 2601 36872 2635
rect 36820 2592 36872 2601
rect 37832 2635 37884 2644
rect 37832 2601 37841 2635
rect 37841 2601 37875 2635
rect 37875 2601 37884 2635
rect 37832 2592 37884 2601
rect 39672 2592 39724 2644
rect 41420 2592 41472 2644
rect 43352 2635 43404 2644
rect 43352 2601 43361 2635
rect 43361 2601 43395 2635
rect 43395 2601 43404 2635
rect 43352 2592 43404 2601
rect 6644 2499 6696 2508
rect 6644 2465 6653 2499
rect 6653 2465 6687 2499
rect 6687 2465 6696 2499
rect 6644 2456 6696 2465
rect 10968 2456 11020 2508
rect 33416 2524 33468 2576
rect 37280 2524 37332 2576
rect 1308 2388 1360 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 5540 2388 5592 2440
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 12164 2431 12216 2440
rect 12164 2397 12173 2431
rect 12173 2397 12207 2431
rect 12207 2397 12216 2431
rect 12164 2388 12216 2397
rect 14004 2388 14056 2440
rect 16396 2431 16448 2440
rect 16396 2397 16405 2431
rect 16405 2397 16439 2431
rect 16439 2397 16448 2431
rect 16396 2388 16448 2397
rect 18236 2388 18288 2440
rect 20628 2431 20680 2440
rect 20628 2397 20637 2431
rect 20637 2397 20671 2431
rect 20671 2397 20680 2431
rect 20628 2388 20680 2397
rect 22744 2431 22796 2440
rect 22744 2397 22753 2431
rect 22753 2397 22787 2431
rect 22787 2397 22796 2431
rect 22744 2388 22796 2397
rect 24860 2431 24912 2440
rect 24860 2397 24869 2431
rect 24869 2397 24903 2431
rect 24903 2397 24912 2431
rect 24860 2388 24912 2397
rect 26700 2388 26752 2440
rect 28908 2431 28960 2440
rect 28908 2397 28917 2431
rect 28917 2397 28951 2431
rect 28951 2397 28960 2431
rect 28908 2388 28960 2397
rect 31024 2431 31076 2440
rect 31024 2397 31033 2431
rect 31033 2397 31067 2431
rect 31067 2397 31076 2431
rect 31024 2388 31076 2397
rect 3424 2320 3476 2372
rect 32864 2388 32916 2440
rect 32956 2388 33008 2440
rect 34888 2431 34940 2440
rect 34888 2397 34897 2431
rect 34897 2397 34931 2431
rect 34931 2397 34940 2431
rect 34888 2388 34940 2397
rect 35164 2388 35216 2440
rect 37004 2431 37056 2440
rect 37004 2397 37013 2431
rect 37013 2397 37047 2431
rect 37047 2397 37056 2431
rect 37004 2388 37056 2397
rect 37556 2431 37608 2440
rect 37556 2397 37565 2431
rect 37565 2397 37599 2431
rect 37599 2397 37608 2431
rect 37556 2388 37608 2397
rect 39672 2431 39724 2440
rect 39672 2397 39681 2431
rect 39681 2397 39715 2431
rect 39715 2397 39724 2431
rect 39672 2388 39724 2397
rect 41788 2431 41840 2440
rect 41788 2397 41797 2431
rect 41797 2397 41831 2431
rect 41831 2397 41840 2431
rect 41788 2388 41840 2397
rect 43536 2431 43588 2440
rect 43536 2397 43545 2431
rect 43545 2397 43579 2431
rect 43579 2397 43588 2431
rect 43536 2388 43588 2397
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 26976 2295 27028 2304
rect 26976 2261 26985 2295
rect 26985 2261 27019 2295
rect 27019 2261 27028 2295
rect 26976 2252 27028 2261
rect 36728 2320 36780 2372
rect 11644 2150 11696 2202
rect 11708 2150 11760 2202
rect 11772 2150 11824 2202
rect 11836 2150 11888 2202
rect 11900 2150 11952 2202
rect 22338 2150 22390 2202
rect 22402 2150 22454 2202
rect 22466 2150 22518 2202
rect 22530 2150 22582 2202
rect 22594 2150 22646 2202
rect 33032 2150 33084 2202
rect 33096 2150 33148 2202
rect 33160 2150 33212 2202
rect 33224 2150 33276 2202
rect 33288 2150 33340 2202
rect 43726 2150 43778 2202
rect 43790 2150 43842 2202
rect 43854 2150 43906 2202
rect 43918 2150 43970 2202
rect 43982 2150 44034 2202
rect 1676 2048 1728 2100
rect 10048 2048 10100 2100
rect 26976 2048 27028 2100
rect 37004 2048 37056 2100
rect 34888 1980 34940 2032
rect 31760 1912 31812 1964
<< metal2 >>
rect 5170 9840 5226 10000
rect 5446 9840 5502 10000
rect 5722 9840 5778 10000
rect 5998 9840 6054 10000
rect 6274 9840 6330 10000
rect 6550 9840 6606 10000
rect 6826 9840 6882 10000
rect 7102 9840 7158 10000
rect 7378 9840 7434 10000
rect 7654 9840 7710 10000
rect 7930 9840 7986 10000
rect 8206 9840 8262 10000
rect 8482 9840 8538 10000
rect 8758 9840 8814 10000
rect 9034 9840 9090 10000
rect 9310 9840 9366 10000
rect 9586 9840 9642 10000
rect 9862 9840 9918 10000
rect 10138 9840 10194 10000
rect 10414 9840 10470 10000
rect 10690 9840 10746 10000
rect 10966 9840 11022 10000
rect 11242 9840 11298 10000
rect 11518 9840 11574 10000
rect 11794 9840 11850 10000
rect 12070 9840 12126 10000
rect 12346 9840 12402 10000
rect 12622 9840 12678 10000
rect 12898 9840 12954 10000
rect 13174 9840 13230 10000
rect 13450 9840 13506 10000
rect 13726 9840 13782 10000
rect 14002 9840 14058 10000
rect 14278 9840 14334 10000
rect 14554 9840 14610 10000
rect 14830 9840 14886 10000
rect 15106 9840 15162 10000
rect 15382 9840 15438 10000
rect 15658 9840 15714 10000
rect 15934 9840 15990 10000
rect 16210 9840 16266 10000
rect 16486 9840 16542 10000
rect 16762 9840 16818 10000
rect 17038 9840 17094 10000
rect 17314 9840 17370 10000
rect 17590 9840 17646 10000
rect 17866 9840 17922 10000
rect 18142 9840 18198 10000
rect 18418 9840 18474 10000
rect 18694 9840 18750 10000
rect 18970 9840 19026 10000
rect 19246 9840 19302 10000
rect 19522 9840 19578 10000
rect 19798 9840 19854 10000
rect 20074 9840 20130 10000
rect 20350 9840 20406 10000
rect 20626 9840 20682 10000
rect 20902 9840 20958 10000
rect 21178 9840 21234 10000
rect 21454 9840 21510 10000
rect 21730 9840 21786 10000
rect 22006 9840 22062 10000
rect 22282 9840 22338 10000
rect 22558 9840 22614 10000
rect 22834 9840 22890 10000
rect 23110 9840 23166 10000
rect 23386 9840 23442 10000
rect 23662 9840 23718 10000
rect 23938 9840 23994 10000
rect 24214 9840 24270 10000
rect 24490 9840 24546 10000
rect 24766 9840 24822 10000
rect 25042 9840 25098 10000
rect 25318 9840 25374 10000
rect 25594 9840 25650 10000
rect 25870 9840 25926 10000
rect 26146 9840 26202 10000
rect 26422 9840 26478 10000
rect 26698 9840 26754 10000
rect 26974 9840 27030 10000
rect 27250 9840 27306 10000
rect 27526 9840 27582 10000
rect 27802 9840 27858 10000
rect 28078 9840 28134 10000
rect 28354 9840 28410 10000
rect 28630 9840 28686 10000
rect 28906 9840 28962 10000
rect 29182 9840 29238 10000
rect 29458 9840 29514 10000
rect 29734 9840 29790 10000
rect 30010 9840 30066 10000
rect 30286 9840 30342 10000
rect 30562 9840 30618 10000
rect 30838 9840 30894 10000
rect 31114 9840 31170 10000
rect 31390 9840 31446 10000
rect 31666 9840 31722 10000
rect 31942 9840 31998 10000
rect 32218 9840 32274 10000
rect 32494 9840 32550 10000
rect 32770 9840 32826 10000
rect 33046 9840 33102 10000
rect 33322 9840 33378 10000
rect 33598 9840 33654 10000
rect 33874 9840 33930 10000
rect 34150 9840 34206 10000
rect 34426 9840 34482 10000
rect 34702 9840 34758 10000
rect 34978 9840 35034 10000
rect 35254 9840 35310 10000
rect 35530 9840 35586 10000
rect 35806 9840 35862 10000
rect 36082 9840 36138 10000
rect 36358 9840 36414 10000
rect 36634 9840 36690 10000
rect 36910 9840 36966 10000
rect 37186 9840 37242 10000
rect 37462 9840 37518 10000
rect 37738 9840 37794 10000
rect 38014 9840 38070 10000
rect 38290 9840 38346 10000
rect 38566 9840 38622 10000
rect 38842 9840 38898 10000
rect 39118 9840 39174 10000
rect 39394 9840 39450 10000
rect 39670 9840 39726 10000
rect 5184 7002 5212 9840
rect 5460 7546 5488 9840
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5552 6254 5580 7346
rect 5736 7002 5764 9840
rect 6012 7546 6040 9840
rect 6288 8242 6316 9840
rect 6196 8214 6316 8242
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5828 7313 5856 7346
rect 5814 7304 5870 7313
rect 5814 7239 5870 7248
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 6196 6780 6224 8214
rect 6564 7274 6592 9840
rect 6642 8120 6698 8129
rect 6642 8055 6698 8064
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 6297 7100 6605 7109
rect 6297 7098 6303 7100
rect 6359 7098 6383 7100
rect 6439 7098 6463 7100
rect 6519 7098 6543 7100
rect 6599 7098 6605 7100
rect 6359 7046 6361 7098
rect 6541 7046 6543 7098
rect 6297 7044 6303 7046
rect 6359 7044 6383 7046
rect 6439 7044 6463 7046
rect 6519 7044 6543 7046
rect 6599 7044 6605 7046
rect 6297 7035 6605 7044
rect 6656 6798 6684 8055
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6748 7478 6776 7686
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6644 6792 6696 6798
rect 6196 6752 6316 6780
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5644 6458 5672 6666
rect 6288 6662 6316 6752
rect 6644 6734 6696 6740
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6104 6458 6132 6598
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 6196 5914 6224 6258
rect 6297 6012 6605 6021
rect 6297 6010 6303 6012
rect 6359 6010 6383 6012
rect 6439 6010 6463 6012
rect 6519 6010 6543 6012
rect 6599 6010 6605 6012
rect 6359 5958 6361 6010
rect 6541 5958 6543 6010
rect 6297 5956 6303 5958
rect 6359 5956 6383 5958
rect 6439 5956 6463 5958
rect 6519 5956 6543 5958
rect 6599 5956 6605 5958
rect 6297 5947 6605 5956
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6748 5030 6776 7278
rect 6840 7002 6868 9840
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 7116 6866 7144 9840
rect 7392 7546 7420 9840
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7300 7002 7328 7346
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7668 6866 7696 9840
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7760 6798 7788 8026
rect 7944 7546 7972 9840
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 8220 6866 8248 9840
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8404 7478 8432 7754
rect 8496 7546 8524 9840
rect 8772 7970 8800 9840
rect 8680 7942 8800 7970
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 8680 6458 8708 7942
rect 9048 7546 9076 9840
rect 9324 7970 9352 9840
rect 9232 7942 9352 7970
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9232 6458 9260 7942
rect 9600 7834 9628 9840
rect 9876 7970 9904 9840
rect 9324 7806 9628 7834
rect 9784 7942 9904 7970
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8036 5914 8064 6258
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8588 5574 8616 6258
rect 9324 6118 9352 7806
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9404 6928 9456 6934
rect 9456 6876 9536 6882
rect 9404 6870 9536 6876
rect 9416 6854 9536 6870
rect 9508 6798 9536 6854
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9416 6186 9444 6734
rect 9692 6390 9720 7210
rect 9784 6458 9812 7942
rect 10046 7848 10102 7857
rect 10046 7783 10102 7792
rect 10060 7478 10088 7783
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10152 6866 10180 9840
rect 10428 8242 10456 9840
rect 10428 8214 10548 8242
rect 10520 6866 10548 8214
rect 10704 7546 10732 9840
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10506 6760 10562 6769
rect 10506 6695 10562 6704
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9876 6225 9904 6598
rect 10520 6458 10548 6695
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 9862 6216 9918 6225
rect 9404 6180 9456 6186
rect 9862 6151 9918 6160
rect 9404 6122 9456 6128
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10428 5914 10456 6054
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 6918 5128 6974 5137
rect 6918 5063 6974 5072
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6297 4924 6605 4933
rect 6297 4922 6303 4924
rect 6359 4922 6383 4924
rect 6439 4922 6463 4924
rect 6519 4922 6543 4924
rect 6599 4922 6605 4924
rect 6359 4870 6361 4922
rect 6541 4870 6543 4922
rect 6297 4868 6303 4870
rect 6359 4868 6383 4870
rect 6439 4868 6463 4870
rect 6519 4868 6543 4870
rect 6599 4868 6605 4870
rect 6297 4859 6605 4868
rect 6297 3836 6605 3845
rect 6297 3834 6303 3836
rect 6359 3834 6383 3836
rect 6439 3834 6463 3836
rect 6519 3834 6543 3836
rect 6599 3834 6605 3836
rect 6359 3782 6361 3834
rect 6541 3782 6543 3834
rect 6297 3780 6303 3782
rect 6359 3780 6383 3782
rect 6439 3780 6463 3782
rect 6519 3780 6543 3782
rect 6599 3780 6605 3782
rect 6297 3771 6605 3780
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6297 2748 6605 2757
rect 6297 2746 6303 2748
rect 6359 2746 6383 2748
rect 6439 2746 6463 2748
rect 6519 2746 6543 2748
rect 6599 2746 6605 2748
rect 6359 2694 6361 2746
rect 6541 2694 6543 2746
rect 6297 2692 6303 2694
rect 6359 2692 6383 2694
rect 6439 2692 6463 2694
rect 6519 2692 6543 2694
rect 6599 2692 6605 2694
rect 6297 2683 6605 2692
rect 6656 2514 6684 3402
rect 6932 2650 6960 5063
rect 10612 4826 10640 7346
rect 10980 6866 11008 9840
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11150 7984 11206 7993
rect 11072 7546 11100 7958
rect 11150 7919 11206 7928
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11164 6798 11192 7919
rect 11256 7274 11284 9840
rect 11532 7426 11560 9840
rect 11808 8022 11836 9840
rect 11796 8016 11848 8022
rect 12084 7970 12112 9840
rect 11796 7958 11848 7964
rect 11992 7942 12112 7970
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 11644 7644 11952 7653
rect 11644 7642 11650 7644
rect 11706 7642 11730 7644
rect 11786 7642 11810 7644
rect 11866 7642 11890 7644
rect 11946 7642 11952 7644
rect 11706 7590 11708 7642
rect 11888 7590 11890 7642
rect 11644 7588 11650 7590
rect 11706 7588 11730 7590
rect 11786 7588 11810 7590
rect 11866 7588 11890 7590
rect 11946 7588 11952 7590
rect 11644 7579 11952 7588
rect 11532 7398 11652 7426
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11624 6866 11652 7398
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 10704 6458 10732 6666
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10796 4758 10824 6666
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11072 5710 11100 6258
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 11348 4622 11376 6666
rect 11644 6556 11952 6565
rect 11644 6554 11650 6556
rect 11706 6554 11730 6556
rect 11786 6554 11810 6556
rect 11866 6554 11890 6556
rect 11946 6554 11952 6556
rect 11706 6502 11708 6554
rect 11888 6502 11890 6554
rect 11644 6500 11650 6502
rect 11706 6500 11730 6502
rect 11786 6500 11810 6502
rect 11866 6500 11890 6502
rect 11946 6500 11952 6502
rect 11644 6491 11952 6500
rect 11992 6458 12020 7942
rect 12176 7546 12204 7958
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12084 7274 12112 7482
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 12268 7002 12296 7210
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12360 6866 12388 9840
rect 12440 8152 12492 8158
rect 12440 8094 12492 8100
rect 12452 7410 12480 8094
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12636 6798 12664 9840
rect 12912 6984 12940 9840
rect 13188 7546 13216 9840
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13084 6996 13136 7002
rect 12912 6956 13084 6984
rect 13084 6938 13136 6944
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11716 5914 11744 6258
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11900 5692 11928 6258
rect 11900 5664 12020 5692
rect 11644 5468 11952 5477
rect 11644 5466 11650 5468
rect 11706 5466 11730 5468
rect 11786 5466 11810 5468
rect 11866 5466 11890 5468
rect 11946 5466 11952 5468
rect 11706 5414 11708 5466
rect 11888 5414 11890 5466
rect 11644 5412 11650 5414
rect 11706 5412 11730 5414
rect 11786 5412 11810 5414
rect 11866 5412 11890 5414
rect 11946 5412 11952 5414
rect 11644 5403 11952 5412
rect 11992 5166 12020 5664
rect 12084 5658 12112 6598
rect 13004 5710 13032 6666
rect 12808 5704 12860 5710
rect 12084 5630 12204 5658
rect 12808 5646 12860 5652
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12072 5568 12124 5574
rect 12070 5536 12072 5545
rect 12124 5536 12126 5545
rect 12070 5471 12126 5480
rect 12176 5409 12204 5630
rect 12162 5400 12218 5409
rect 12162 5335 12218 5344
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11644 4380 11952 4389
rect 11644 4378 11650 4380
rect 11706 4378 11730 4380
rect 11786 4378 11810 4380
rect 11866 4378 11890 4380
rect 11946 4378 11952 4380
rect 11706 4326 11708 4378
rect 11888 4326 11890 4378
rect 11644 4324 11650 4326
rect 11706 4324 11730 4326
rect 11786 4324 11810 4326
rect 11866 4324 11890 4326
rect 11946 4324 11952 4326
rect 11644 4315 11952 4324
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 10980 2514 11008 3470
rect 11644 3292 11952 3301
rect 11644 3290 11650 3292
rect 11706 3290 11730 3292
rect 11786 3290 11810 3292
rect 11866 3290 11890 3292
rect 11946 3290 11952 3292
rect 11706 3238 11708 3290
rect 11888 3238 11890 3290
rect 11644 3236 11650 3238
rect 11706 3236 11730 3238
rect 11786 3236 11810 3238
rect 11866 3236 11890 3238
rect 11946 3236 11952 3238
rect 11644 3227 11952 3236
rect 12820 2650 12848 5646
rect 13280 4593 13308 7346
rect 13372 5914 13400 8298
rect 13464 6984 13492 9840
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13648 7274 13676 8026
rect 13740 7546 13768 9840
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 7546 13860 8230
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 13636 6996 13688 7002
rect 13464 6956 13636 6984
rect 13636 6938 13688 6944
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13634 6488 13690 6497
rect 13634 6423 13690 6432
rect 13648 6390 13676 6423
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13648 5914 13676 6054
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13740 5302 13768 6598
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 13924 4690 13952 6666
rect 14016 6458 14044 9840
rect 14292 8294 14320 9840
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14108 6322 14136 7890
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14200 7002 14228 7346
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14292 6905 14320 7346
rect 14278 6896 14334 6905
rect 14278 6831 14334 6840
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14200 5098 14228 6734
rect 14292 5273 14320 6734
rect 14476 6458 14504 7346
rect 14568 7002 14596 9840
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14660 7274 14688 7414
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14844 6866 14872 9840
rect 15120 7546 15148 9840
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15396 6866 15424 9840
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 14740 6724 14792 6730
rect 14740 6666 14792 6672
rect 15016 6724 15068 6730
rect 15016 6666 15068 6672
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 14752 6458 14780 6666
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 15028 6390 15056 6666
rect 15304 6458 15332 6666
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 15488 6322 15516 8366
rect 15672 7546 15700 9840
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15580 6458 15608 7346
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15856 6322 15884 8434
rect 15948 6866 15976 9840
rect 16120 8152 16172 8158
rect 16120 8094 16172 8100
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 14278 5264 14334 5273
rect 14278 5199 14334 5208
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 14844 4729 14872 6258
rect 14830 4720 14886 4729
rect 13912 4684 13964 4690
rect 14830 4655 14886 4664
rect 13912 4626 13964 4632
rect 13266 4584 13322 4593
rect 13266 4519 13322 4528
rect 16132 4185 16160 8094
rect 16224 7546 16252 9840
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16304 8152 16356 8158
rect 16304 8094 16356 8100
rect 16316 7818 16344 8094
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16316 7002 16344 7142
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16316 5914 16344 6734
rect 16408 6322 16436 8502
rect 16500 6866 16528 9840
rect 16776 7546 16804 9840
rect 17052 8242 17080 9840
rect 16868 8214 17080 8242
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16486 6624 16542 6633
rect 16486 6559 16542 6568
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16500 5642 16528 6559
rect 16592 6186 16620 7346
rect 16868 6848 16896 8214
rect 17328 7546 17356 9840
rect 17498 8256 17554 8265
rect 17498 8191 17554 8200
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 16991 7100 17299 7109
rect 16991 7098 16997 7100
rect 17053 7098 17077 7100
rect 17133 7098 17157 7100
rect 17213 7098 17237 7100
rect 17293 7098 17299 7100
rect 17053 7046 17055 7098
rect 17235 7046 17237 7098
rect 16991 7044 16997 7046
rect 17053 7044 17077 7046
rect 17133 7044 17157 7046
rect 17213 7044 17237 7046
rect 17293 7044 17299 7046
rect 16991 7035 17299 7044
rect 17040 6860 17092 6866
rect 16868 6820 17040 6848
rect 17040 6802 17092 6808
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 16684 6458 16712 6666
rect 17236 6458 17264 6666
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17328 6186 17356 7346
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17420 6730 17448 7142
rect 17408 6724 17460 6730
rect 17408 6666 17460 6672
rect 17512 6474 17540 8191
rect 17604 6866 17632 9840
rect 17880 7546 17908 9840
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17420 6446 17540 6474
rect 17420 6322 17448 6446
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 16580 6180 16632 6186
rect 16580 6122 16632 6128
rect 17316 6180 17368 6186
rect 17316 6122 17368 6128
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 16991 6012 17299 6021
rect 16991 6010 16997 6012
rect 17053 6010 17077 6012
rect 17133 6010 17157 6012
rect 17213 6010 17237 6012
rect 17293 6010 17299 6012
rect 17053 5958 17055 6010
rect 17235 5958 17237 6010
rect 16991 5956 16997 5958
rect 17053 5956 17077 5958
rect 17133 5956 17157 5958
rect 17213 5956 17237 5958
rect 17293 5956 17299 5958
rect 16991 5947 17299 5956
rect 17420 5914 17448 6122
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17512 5642 17540 6258
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 17500 5636 17552 5642
rect 17500 5578 17552 5584
rect 17696 5574 17724 7278
rect 17880 6458 17908 7346
rect 17958 7168 18014 7177
rect 17958 7103 18014 7112
rect 17972 7002 18000 7103
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 18156 6866 18184 9840
rect 18432 7546 18460 9840
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18418 6760 18474 6769
rect 18328 6724 18380 6730
rect 18418 6695 18420 6704
rect 18328 6666 18380 6672
rect 18472 6695 18474 6704
rect 18420 6666 18472 6672
rect 18340 6458 18368 6666
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18144 6384 18196 6390
rect 17774 6352 17830 6361
rect 18144 6326 18196 6332
rect 17774 6287 17776 6296
rect 17828 6287 17830 6296
rect 17776 6258 17828 6264
rect 17868 6248 17920 6254
rect 17866 6216 17868 6225
rect 17920 6216 17922 6225
rect 17866 6151 17922 6160
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 18156 5370 18184 6326
rect 18524 6322 18552 6598
rect 18616 6458 18644 7346
rect 18708 7188 18736 9840
rect 18984 8514 19012 9840
rect 18984 8486 19196 8514
rect 19168 7478 19196 8486
rect 19156 7472 19208 7478
rect 19156 7414 19208 7420
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18788 7200 18840 7206
rect 18708 7160 18788 7188
rect 18788 7142 18840 7148
rect 18786 7032 18842 7041
rect 18786 6967 18842 6976
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18800 6322 18828 6967
rect 18984 6458 19012 7346
rect 19260 7206 19288 9840
rect 19536 8378 19564 9840
rect 19812 8378 19840 9840
rect 20088 8378 20116 9840
rect 20364 8378 20392 9840
rect 19352 8350 19564 8378
rect 19628 8350 19840 8378
rect 19904 8350 20116 8378
rect 20180 8350 20392 8378
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 19352 6798 19380 8350
rect 19432 8152 19484 8158
rect 19432 8094 19484 8100
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19076 6458 19104 6734
rect 19444 6662 19472 8094
rect 19628 6798 19656 8350
rect 19904 6798 19932 8350
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 19996 7002 20024 7346
rect 19984 6996 20036 7002
rect 19984 6938 20036 6944
rect 20180 6798 20208 8350
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20364 6934 20392 7822
rect 20536 7268 20588 7274
rect 20536 7210 20588 7216
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20260 6928 20312 6934
rect 20260 6870 20312 6876
rect 20352 6928 20404 6934
rect 20352 6870 20404 6876
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18248 5914 18276 6258
rect 19352 6089 19380 6394
rect 19338 6080 19394 6089
rect 19338 6015 19394 6024
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 19536 5030 19564 6598
rect 19812 5778 19840 6598
rect 20272 6202 20300 6870
rect 20456 6322 20484 6938
rect 20548 6798 20576 7210
rect 20640 6798 20668 9840
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 20732 7449 20760 7958
rect 20718 7440 20774 7449
rect 20718 7375 20774 7384
rect 20812 7404 20864 7410
rect 20916 7392 20944 9840
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21100 7546 21128 7686
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20996 7472 21048 7478
rect 20996 7414 21048 7420
rect 20864 7364 20944 7392
rect 20812 7346 20864 7352
rect 20810 7168 20866 7177
rect 20810 7103 20866 7112
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20640 6497 20668 6598
rect 20626 6488 20682 6497
rect 20626 6423 20682 6432
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20272 6174 20760 6202
rect 20732 6118 20760 6174
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20824 5914 20852 7103
rect 20904 6656 20956 6662
rect 21008 6633 21036 7414
rect 21192 7410 21220 9840
rect 21270 7848 21326 7857
rect 21270 7783 21326 7792
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21284 6662 21312 7783
rect 21364 7404 21416 7410
rect 21468 7392 21496 9840
rect 21416 7364 21496 7392
rect 21640 7404 21692 7410
rect 21364 7346 21416 7352
rect 21744 7392 21772 9840
rect 22020 7410 22048 9840
rect 22296 8650 22324 9840
rect 22204 8622 22324 8650
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 21692 7364 21772 7392
rect 22008 7404 22060 7410
rect 21640 7346 21692 7352
rect 22008 7346 22060 7352
rect 22112 7290 22140 8026
rect 22204 7392 22232 8622
rect 22572 8378 22600 9840
rect 22572 8350 22784 8378
rect 22338 7644 22646 7653
rect 22338 7642 22344 7644
rect 22400 7642 22424 7644
rect 22480 7642 22504 7644
rect 22560 7642 22584 7644
rect 22640 7642 22646 7644
rect 22400 7590 22402 7642
rect 22582 7590 22584 7642
rect 22338 7588 22344 7590
rect 22400 7588 22424 7590
rect 22480 7588 22504 7590
rect 22560 7588 22584 7590
rect 22640 7588 22646 7590
rect 22338 7579 22646 7588
rect 22284 7404 22336 7410
rect 22204 7364 22284 7392
rect 22284 7346 22336 7352
rect 21916 7268 21968 7274
rect 22112 7262 22232 7290
rect 21916 7210 21968 7216
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21824 7200 21876 7206
rect 21824 7142 21876 7148
rect 21468 7002 21496 7142
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21836 6798 21864 7142
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21180 6656 21232 6662
rect 20904 6598 20956 6604
rect 20994 6624 21050 6633
rect 20916 6186 20944 6598
rect 21180 6598 21232 6604
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 20994 6559 21050 6568
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 21192 5545 21220 6598
rect 21928 6322 21956 7210
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22112 6866 22140 7142
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22008 6792 22060 6798
rect 22008 6734 22060 6740
rect 22020 6458 22048 6734
rect 22204 6458 22232 7262
rect 22756 6780 22784 8350
rect 22848 7410 22876 9840
rect 22926 7984 22982 7993
rect 22982 7942 23060 7970
rect 22926 7919 22982 7928
rect 22928 7812 22980 7818
rect 22928 7754 22980 7760
rect 22940 7546 22968 7754
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 22928 7200 22980 7206
rect 22928 7142 22980 7148
rect 22836 6792 22888 6798
rect 22756 6752 22836 6780
rect 22836 6734 22888 6740
rect 22338 6556 22646 6565
rect 22338 6554 22344 6556
rect 22400 6554 22424 6556
rect 22480 6554 22504 6556
rect 22560 6554 22584 6556
rect 22640 6554 22646 6556
rect 22400 6502 22402 6554
rect 22582 6502 22584 6554
rect 22338 6500 22344 6502
rect 22400 6500 22424 6502
rect 22480 6500 22504 6502
rect 22560 6500 22584 6502
rect 22640 6500 22646 6502
rect 22338 6491 22646 6500
rect 22940 6458 22968 7142
rect 22008 6452 22060 6458
rect 22008 6394 22060 6400
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22928 6452 22980 6458
rect 22928 6394 22980 6400
rect 21916 6316 21968 6322
rect 21916 6258 21968 6264
rect 22100 6248 22152 6254
rect 22152 6196 22232 6202
rect 22100 6190 22232 6196
rect 22112 6174 22232 6190
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 21178 5536 21234 5545
rect 21178 5471 21234 5480
rect 22020 5409 22048 6054
rect 22204 5846 22232 6174
rect 23032 6118 23060 7942
rect 23124 7410 23152 9840
rect 23204 8220 23256 8226
rect 23204 8162 23256 8168
rect 23112 7404 23164 7410
rect 23112 7346 23164 7352
rect 23112 7268 23164 7274
rect 23112 7210 23164 7216
rect 23124 6254 23152 7210
rect 23112 6248 23164 6254
rect 23112 6190 23164 6196
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 22192 5840 22244 5846
rect 22192 5782 22244 5788
rect 23216 5778 23244 8162
rect 23296 8016 23348 8022
rect 23296 7958 23348 7964
rect 23308 5846 23336 7958
rect 23400 7410 23428 9840
rect 23388 7404 23440 7410
rect 23676 7392 23704 9840
rect 23952 8650 23980 9840
rect 24228 8650 24256 9840
rect 24504 8650 24532 9840
rect 23952 8622 24072 8650
rect 24228 8622 24348 8650
rect 24504 8622 24716 8650
rect 23940 7404 23992 7410
rect 23676 7364 23940 7392
rect 23388 7346 23440 7352
rect 24044 7392 24072 8622
rect 24216 7404 24268 7410
rect 24044 7364 24216 7392
rect 23940 7346 23992 7352
rect 24320 7392 24348 8622
rect 24688 7478 24716 8622
rect 24676 7472 24728 7478
rect 24676 7414 24728 7420
rect 24492 7404 24544 7410
rect 24320 7364 24492 7392
rect 24216 7346 24268 7352
rect 24492 7346 24544 7352
rect 24582 7304 24638 7313
rect 24780 7274 24808 9840
rect 25056 8650 25084 9840
rect 25056 8622 25268 8650
rect 25134 8120 25190 8129
rect 25240 8106 25268 8622
rect 25332 8294 25360 9840
rect 25320 8288 25372 8294
rect 25320 8230 25372 8236
rect 25240 8078 25544 8106
rect 25134 8055 25190 8064
rect 24582 7239 24584 7248
rect 24636 7239 24638 7248
rect 24768 7268 24820 7274
rect 24584 7210 24636 7216
rect 24768 7210 24820 7216
rect 25148 7206 25176 8055
rect 25320 7948 25372 7954
rect 25320 7890 25372 7896
rect 25332 7546 25360 7890
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25516 7478 25544 8078
rect 25504 7472 25556 7478
rect 25504 7414 25556 7420
rect 25608 7324 25636 9840
rect 25884 7478 25912 9840
rect 25964 8288 26016 8294
rect 25964 8230 26016 8236
rect 25872 7472 25924 7478
rect 25872 7414 25924 7420
rect 25976 7410 26004 8230
rect 26160 7546 26188 9840
rect 26148 7540 26200 7546
rect 26148 7482 26200 7488
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 25872 7336 25924 7342
rect 25608 7296 25872 7324
rect 26436 7324 26464 9840
rect 26712 8650 26740 9840
rect 26988 8786 27016 9840
rect 26988 8758 27200 8786
rect 26712 8622 27016 8650
rect 26882 8256 26938 8265
rect 26882 8191 26938 8200
rect 26792 7948 26844 7954
rect 26792 7890 26844 7896
rect 26700 7336 26752 7342
rect 26436 7296 26700 7324
rect 25872 7278 25924 7284
rect 26700 7278 26752 7284
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 24032 7200 24084 7206
rect 24032 7142 24084 7148
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 25872 7200 25924 7206
rect 25872 7142 25924 7148
rect 26056 7200 26108 7206
rect 26056 7142 26108 7148
rect 26148 7200 26200 7206
rect 26148 7142 26200 7148
rect 26608 7200 26660 7206
rect 26608 7142 26660 7148
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 23296 5840 23348 5846
rect 23296 5782 23348 5788
rect 23204 5772 23256 5778
rect 23204 5714 23256 5720
rect 22338 5468 22646 5477
rect 22338 5466 22344 5468
rect 22400 5466 22424 5468
rect 22480 5466 22504 5468
rect 22560 5466 22584 5468
rect 22640 5466 22646 5468
rect 22400 5414 22402 5466
rect 22582 5414 22584 5466
rect 22338 5412 22344 5414
rect 22400 5412 22424 5414
rect 22480 5412 22504 5414
rect 22560 5412 22584 5414
rect 22640 5412 22646 5414
rect 22006 5400 22062 5409
rect 22338 5403 22646 5412
rect 23400 5370 23428 6598
rect 23492 6322 23520 7142
rect 24044 6798 24072 7142
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 25320 6656 25372 6662
rect 25320 6598 25372 6604
rect 25596 6656 25648 6662
rect 25596 6598 25648 6604
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 25332 6186 25360 6598
rect 25608 6225 25636 6598
rect 25884 6322 25912 7142
rect 26068 6798 26096 7142
rect 26160 7002 26188 7142
rect 26620 7002 26648 7142
rect 26804 7041 26832 7890
rect 26896 7886 26924 8191
rect 26884 7880 26936 7886
rect 26884 7822 26936 7828
rect 26988 7478 27016 8622
rect 27172 7562 27200 8758
rect 27264 7750 27292 9840
rect 27540 8922 27568 9840
rect 27448 8894 27568 8922
rect 27448 7818 27476 8894
rect 27816 8650 27844 9840
rect 27816 8622 27936 8650
rect 27436 7812 27488 7818
rect 27436 7754 27488 7760
rect 27252 7744 27304 7750
rect 27252 7686 27304 7692
rect 27068 7540 27120 7546
rect 27172 7534 27568 7562
rect 27068 7482 27120 7488
rect 26976 7472 27028 7478
rect 26976 7414 27028 7420
rect 26790 7032 26846 7041
rect 26148 6996 26200 7002
rect 26148 6938 26200 6944
rect 26424 6996 26476 7002
rect 26424 6938 26476 6944
rect 26608 6996 26660 7002
rect 26790 6967 26846 6976
rect 26608 6938 26660 6944
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26148 6724 26200 6730
rect 26148 6666 26200 6672
rect 25964 6452 26016 6458
rect 25964 6394 26016 6400
rect 25872 6316 25924 6322
rect 25872 6258 25924 6264
rect 25594 6216 25650 6225
rect 25320 6180 25372 6186
rect 25594 6151 25650 6160
rect 25320 6122 25372 6128
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 22006 5335 22062 5344
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 16991 4924 17299 4933
rect 16991 4922 16997 4924
rect 17053 4922 17077 4924
rect 17133 4922 17157 4924
rect 17213 4922 17237 4924
rect 17293 4922 17299 4924
rect 17053 4870 17055 4922
rect 17235 4870 17237 4922
rect 16991 4868 16997 4870
rect 17053 4868 17077 4870
rect 17133 4868 17157 4870
rect 17213 4868 17237 4870
rect 17293 4868 17299 4870
rect 16991 4859 17299 4868
rect 16118 4176 16174 4185
rect 16118 4111 16174 4120
rect 16991 3836 17299 3845
rect 16991 3834 16997 3836
rect 17053 3834 17077 3836
rect 17133 3834 17157 3836
rect 17213 3834 17237 3836
rect 17293 3834 17299 3836
rect 17053 3782 17055 3834
rect 17235 3782 17237 3834
rect 16991 3780 16997 3782
rect 17053 3780 17077 3782
rect 17133 3780 17157 3782
rect 17213 3780 17237 3782
rect 17293 3780 17299 3782
rect 16991 3771 17299 3780
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 16991 2748 17299 2757
rect 16991 2746 16997 2748
rect 17053 2746 17077 2748
rect 17133 2746 17157 2748
rect 17213 2746 17237 2748
rect 17293 2746 17299 2748
rect 17053 2694 17055 2746
rect 17235 2694 17237 2746
rect 16991 2692 16997 2694
rect 17053 2692 17077 2694
rect 17133 2692 17157 2694
rect 17213 2692 17237 2694
rect 17293 2692 17299 2694
rect 16991 2683 17299 2692
rect 18708 2650 18736 2994
rect 20456 2650 20484 5170
rect 24044 4593 24072 6054
rect 25976 5302 26004 6394
rect 25964 5296 26016 5302
rect 25964 5238 26016 5244
rect 24030 4584 24086 4593
rect 24030 4519 24086 4528
rect 22338 4380 22646 4389
rect 22338 4378 22344 4380
rect 22400 4378 22424 4380
rect 22480 4378 22504 4380
rect 22560 4378 22584 4380
rect 22640 4378 22646 4380
rect 22400 4326 22402 4378
rect 22582 4326 22584 4378
rect 22338 4324 22344 4326
rect 22400 4324 22424 4326
rect 22480 4324 22504 4326
rect 22560 4324 22584 4326
rect 22640 4324 22646 4326
rect 22338 4315 22646 4324
rect 26160 4185 26188 6666
rect 26436 4690 26464 6938
rect 27080 6798 27108 7482
rect 27540 7342 27568 7534
rect 27908 7478 27936 8622
rect 27896 7472 27948 7478
rect 27896 7414 27948 7420
rect 27528 7336 27580 7342
rect 28092 7324 28120 9840
rect 28368 7546 28396 9840
rect 28644 8650 28672 9840
rect 28644 8622 28856 8650
rect 28828 8294 28856 8622
rect 28816 8288 28868 8294
rect 28816 8230 28868 8236
rect 28540 7812 28592 7818
rect 28540 7754 28592 7760
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 28356 7540 28408 7546
rect 28356 7482 28408 7488
rect 28460 7410 28488 7686
rect 28552 7410 28580 7754
rect 28448 7404 28500 7410
rect 28448 7346 28500 7352
rect 28540 7404 28592 7410
rect 28540 7346 28592 7352
rect 28356 7336 28408 7342
rect 28092 7296 28356 7324
rect 27528 7278 27580 7284
rect 28356 7278 28408 7284
rect 28446 7304 28502 7313
rect 27436 7268 27488 7274
rect 28920 7290 28948 9840
rect 29196 8158 29224 9840
rect 29184 8152 29236 8158
rect 29184 8094 29236 8100
rect 29472 7546 29500 9840
rect 29748 8650 29776 9840
rect 29748 8622 29960 8650
rect 29932 8294 29960 8622
rect 29736 8288 29788 8294
rect 29736 8230 29788 8236
rect 29920 8288 29972 8294
rect 29920 8230 29972 8236
rect 29460 7540 29512 7546
rect 29460 7482 29512 7488
rect 29748 7410 29776 8230
rect 29736 7404 29788 7410
rect 29736 7346 29788 7352
rect 30024 7324 30052 9840
rect 30300 8242 30328 9840
rect 30300 8214 30512 8242
rect 30288 8152 30340 8158
rect 30288 8094 30340 8100
rect 30300 7410 30328 8094
rect 30484 7546 30512 8214
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 30288 7404 30340 7410
rect 30288 7346 30340 7352
rect 30196 7336 30248 7342
rect 30024 7296 30196 7324
rect 28446 7239 28502 7248
rect 28816 7268 28868 7274
rect 27436 7210 27488 7216
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 27264 7002 27292 7142
rect 27252 6996 27304 7002
rect 27252 6938 27304 6944
rect 27448 6798 27476 7210
rect 27528 7200 27580 7206
rect 27528 7142 27580 7148
rect 28356 7200 28408 7206
rect 28356 7142 28408 7148
rect 27068 6792 27120 6798
rect 27068 6734 27120 6740
rect 27436 6792 27488 6798
rect 27436 6734 27488 6740
rect 27540 6662 27568 7142
rect 27685 7100 27993 7109
rect 27685 7098 27691 7100
rect 27747 7098 27771 7100
rect 27827 7098 27851 7100
rect 27907 7098 27931 7100
rect 27987 7098 27993 7100
rect 27747 7046 27749 7098
rect 27929 7046 27931 7098
rect 27685 7044 27691 7046
rect 27747 7044 27771 7046
rect 27827 7044 27851 7046
rect 27907 7044 27931 7046
rect 27987 7044 27993 7046
rect 27685 7035 27993 7044
rect 28368 7002 28396 7142
rect 28356 6996 28408 7002
rect 28356 6938 28408 6944
rect 28460 6662 28488 7239
rect 28920 7262 29040 7290
rect 30196 7278 30248 7284
rect 30576 7274 30604 9840
rect 30748 8288 30800 8294
rect 30748 8230 30800 8236
rect 30656 8016 30708 8022
rect 30656 7958 30708 7964
rect 28816 7210 28868 7216
rect 28632 7200 28684 7206
rect 28632 7142 28684 7148
rect 28644 7002 28672 7142
rect 28632 6996 28684 7002
rect 28632 6938 28684 6944
rect 28828 6798 28856 7210
rect 28908 7200 28960 7206
rect 29012 7188 29040 7262
rect 30564 7268 30616 7274
rect 30564 7210 30616 7216
rect 30668 7206 30696 7958
rect 30760 7410 30788 8230
rect 30748 7404 30800 7410
rect 30748 7346 30800 7352
rect 30852 7324 30880 9840
rect 31024 7336 31076 7342
rect 30852 7296 31024 7324
rect 31024 7278 31076 7284
rect 29092 7200 29144 7206
rect 29012 7160 29092 7188
rect 28908 7142 28960 7148
rect 29092 7142 29144 7148
rect 29552 7200 29604 7206
rect 29552 7142 29604 7148
rect 29828 7200 29880 7206
rect 29828 7142 29880 7148
rect 30104 7200 30156 7206
rect 30104 7142 30156 7148
rect 30380 7200 30432 7206
rect 30380 7142 30432 7148
rect 30656 7200 30708 7206
rect 30656 7142 30708 7148
rect 30932 7200 30984 7206
rect 30932 7142 30984 7148
rect 28920 6798 28948 7142
rect 29564 6798 29592 7142
rect 29840 6798 29868 7142
rect 30116 6798 30144 7142
rect 30392 6798 30420 7142
rect 28816 6792 28868 6798
rect 28816 6734 28868 6740
rect 28908 6792 28960 6798
rect 28908 6734 28960 6740
rect 29552 6792 29604 6798
rect 29552 6734 29604 6740
rect 29828 6792 29880 6798
rect 29828 6734 29880 6740
rect 30104 6792 30156 6798
rect 30104 6734 30156 6740
rect 30380 6792 30432 6798
rect 30380 6734 30432 6740
rect 26976 6656 27028 6662
rect 26976 6598 27028 6604
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 27528 6656 27580 6662
rect 27528 6598 27580 6604
rect 27620 6656 27672 6662
rect 27620 6598 27672 6604
rect 28080 6656 28132 6662
rect 28080 6598 28132 6604
rect 28448 6656 28500 6662
rect 28448 6598 28500 6604
rect 28908 6656 28960 6662
rect 28908 6598 28960 6604
rect 29368 6656 29420 6662
rect 29368 6598 29420 6604
rect 29828 6656 29880 6662
rect 29828 6598 29880 6604
rect 30196 6656 30248 6662
rect 30196 6598 30248 6604
rect 30288 6656 30340 6662
rect 30288 6598 30340 6604
rect 26988 5846 27016 6598
rect 27356 6458 27384 6598
rect 27344 6452 27396 6458
rect 27344 6394 27396 6400
rect 27632 6066 27660 6598
rect 27540 6038 27660 6066
rect 27540 5930 27568 6038
rect 27685 6012 27993 6021
rect 27685 6010 27691 6012
rect 27747 6010 27771 6012
rect 27827 6010 27851 6012
rect 27907 6010 27931 6012
rect 27987 6010 27993 6012
rect 27747 5958 27749 6010
rect 27929 5958 27931 6010
rect 27685 5956 27691 5958
rect 27747 5956 27771 5958
rect 27827 5956 27851 5958
rect 27907 5956 27931 5958
rect 27987 5956 27993 5958
rect 27685 5947 27993 5956
rect 27540 5902 27660 5930
rect 26976 5840 27028 5846
rect 26976 5782 27028 5788
rect 27632 5098 27660 5902
rect 28092 5166 28120 6598
rect 28080 5160 28132 5166
rect 28080 5102 28132 5108
rect 27620 5092 27672 5098
rect 27620 5034 27672 5040
rect 27685 4924 27993 4933
rect 27685 4922 27691 4924
rect 27747 4922 27771 4924
rect 27827 4922 27851 4924
rect 27907 4922 27931 4924
rect 27987 4922 27993 4924
rect 27747 4870 27749 4922
rect 27929 4870 27931 4922
rect 27685 4868 27691 4870
rect 27747 4868 27771 4870
rect 27827 4868 27851 4870
rect 27907 4868 27931 4870
rect 27987 4868 27993 4870
rect 27685 4859 27993 4868
rect 26424 4684 26476 4690
rect 26424 4626 26476 4632
rect 28920 4622 28948 6598
rect 29380 5914 29408 6598
rect 29368 5908 29420 5914
rect 29368 5850 29420 5856
rect 29840 4758 29868 6598
rect 30208 4826 30236 6598
rect 30300 6254 30328 6598
rect 30944 6390 30972 7142
rect 31128 6780 31156 9840
rect 31404 8650 31432 9840
rect 31680 8786 31708 9840
rect 31312 8622 31432 8650
rect 31588 8758 31708 8786
rect 31208 8084 31260 8090
rect 31208 8026 31260 8032
rect 31220 7206 31248 8026
rect 31312 7478 31340 8622
rect 31392 7948 31444 7954
rect 31392 7890 31444 7896
rect 31484 7948 31536 7954
rect 31484 7890 31536 7896
rect 31404 7546 31432 7890
rect 31496 7546 31524 7890
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 31484 7540 31536 7546
rect 31484 7482 31536 7488
rect 31300 7472 31352 7478
rect 31300 7414 31352 7420
rect 31484 7404 31536 7410
rect 31484 7346 31536 7352
rect 31496 7274 31524 7346
rect 31588 7324 31616 8758
rect 31852 7336 31904 7342
rect 31588 7296 31852 7324
rect 31852 7278 31904 7284
rect 31956 7274 31984 9840
rect 32232 7478 32260 9840
rect 32508 7546 32536 9840
rect 32588 8560 32640 8566
rect 32588 8502 32640 8508
rect 32496 7540 32548 7546
rect 32496 7482 32548 7488
rect 32220 7472 32272 7478
rect 32220 7414 32272 7420
rect 32600 7342 32628 8502
rect 32680 7880 32732 7886
rect 32680 7822 32732 7828
rect 32588 7336 32640 7342
rect 32588 7278 32640 7284
rect 31484 7268 31536 7274
rect 31484 7210 31536 7216
rect 31944 7268 31996 7274
rect 31944 7210 31996 7216
rect 32692 7206 32720 7822
rect 32784 7324 32812 9840
rect 33060 8922 33088 9840
rect 32968 8894 33088 8922
rect 33336 8922 33364 9840
rect 33336 8894 33456 8922
rect 32864 7336 32916 7342
rect 32784 7296 32864 7324
rect 32864 7278 32916 7284
rect 31208 7200 31260 7206
rect 31208 7142 31260 7148
rect 32312 7200 32364 7206
rect 32312 7142 32364 7148
rect 32588 7200 32640 7206
rect 32588 7142 32640 7148
rect 32680 7200 32732 7206
rect 32680 7142 32732 7148
rect 31208 6792 31260 6798
rect 31128 6752 31208 6780
rect 31208 6734 31260 6740
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 31392 6656 31444 6662
rect 31392 6598 31444 6604
rect 30932 6384 30984 6390
rect 30932 6326 30984 6332
rect 30288 6248 30340 6254
rect 30288 6190 30340 6196
rect 30380 6248 30432 6254
rect 30380 6190 30432 6196
rect 30392 5030 30420 6190
rect 31404 5574 31432 6598
rect 31392 5568 31444 5574
rect 31392 5510 31444 5516
rect 30380 5024 30432 5030
rect 30380 4966 30432 4972
rect 30196 4820 30248 4826
rect 30196 4762 30248 4768
rect 29828 4752 29880 4758
rect 29828 4694 29880 4700
rect 28908 4616 28960 4622
rect 28908 4558 28960 4564
rect 26146 4176 26202 4185
rect 26146 4111 26202 4120
rect 27685 3836 27993 3845
rect 27685 3834 27691 3836
rect 27747 3834 27771 3836
rect 27827 3834 27851 3836
rect 27907 3834 27931 3836
rect 27987 3834 27993 3836
rect 27747 3782 27749 3834
rect 27929 3782 27931 3834
rect 27685 3780 27691 3782
rect 27747 3780 27771 3782
rect 27827 3780 27851 3782
rect 27907 3780 27931 3782
rect 27987 3780 27993 3782
rect 27685 3771 27993 3780
rect 22338 3292 22646 3301
rect 22338 3290 22344 3292
rect 22400 3290 22424 3292
rect 22480 3290 22504 3292
rect 22560 3290 22584 3292
rect 22640 3290 22646 3292
rect 22400 3238 22402 3290
rect 22582 3238 22584 3290
rect 22338 3236 22344 3238
rect 22400 3236 22424 3238
rect 22480 3236 22504 3238
rect 22560 3236 22584 3238
rect 22640 3236 22646 3238
rect 22338 3227 22646 3236
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 25044 3052 25096 3058
rect 25044 2994 25096 3000
rect 22940 2650 22968 2994
rect 25056 2650 25084 2994
rect 27685 2748 27993 2757
rect 27685 2746 27691 2748
rect 27747 2746 27771 2748
rect 27827 2746 27851 2748
rect 27907 2746 27931 2748
rect 27987 2746 27993 2748
rect 27747 2694 27749 2746
rect 27929 2694 27931 2746
rect 27685 2692 27691 2694
rect 27747 2692 27771 2694
rect 27827 2692 27851 2694
rect 27907 2692 27931 2694
rect 27987 2692 27993 2694
rect 27685 2683 27993 2692
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 25044 2644 25096 2650
rect 25044 2586 25096 2592
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 22744 2440 22796 2446
rect 24860 2440 24912 2446
rect 22744 2382 22796 2388
rect 24780 2400 24860 2428
rect 1320 160 1348 2382
rect 1688 2106 1716 2382
rect 3424 2372 3476 2378
rect 3424 2314 3476 2320
rect 1676 2100 1728 2106
rect 1676 2042 1728 2048
rect 3436 160 3464 2314
rect 5552 160 5580 2382
rect 1306 0 1362 160
rect 3422 0 3478 160
rect 5538 0 5594 160
rect 7654 82 7710 160
rect 7760 82 7788 2382
rect 7654 54 7788 82
rect 9770 82 9826 160
rect 9876 82 9904 2382
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 10060 2106 10088 2246
rect 11644 2204 11952 2213
rect 11644 2202 11650 2204
rect 11706 2202 11730 2204
rect 11786 2202 11810 2204
rect 11866 2202 11890 2204
rect 11946 2202 11952 2204
rect 11706 2150 11708 2202
rect 11888 2150 11890 2202
rect 11644 2148 11650 2150
rect 11706 2148 11730 2150
rect 11786 2148 11810 2150
rect 11866 2148 11890 2150
rect 11946 2148 11952 2150
rect 11644 2139 11952 2148
rect 10048 2100 10100 2106
rect 10048 2042 10100 2048
rect 9770 54 9904 82
rect 11886 82 11942 160
rect 12176 82 12204 2382
rect 14016 160 14044 2382
rect 11886 54 12204 82
rect 7654 0 7710 54
rect 9770 0 9826 54
rect 11886 0 11942 54
rect 14002 0 14058 160
rect 16118 82 16174 160
rect 16408 82 16436 2382
rect 18248 160 18276 2382
rect 16118 54 16436 82
rect 16118 0 16174 54
rect 18234 0 18290 160
rect 20350 82 20406 160
rect 20640 82 20668 2382
rect 22338 2204 22646 2213
rect 22338 2202 22344 2204
rect 22400 2202 22424 2204
rect 22480 2202 22504 2204
rect 22560 2202 22584 2204
rect 22640 2202 22646 2204
rect 22400 2150 22402 2202
rect 22582 2150 22584 2202
rect 22338 2148 22344 2150
rect 22400 2148 22424 2150
rect 22480 2148 22504 2150
rect 22560 2148 22584 2150
rect 22640 2148 22646 2150
rect 22338 2139 22646 2148
rect 20350 54 20668 82
rect 22466 82 22522 160
rect 22756 82 22784 2382
rect 22466 54 22784 82
rect 24582 82 24638 160
rect 24780 82 24808 2400
rect 24860 2382 24912 2388
rect 26700 2440 26752 2446
rect 26700 2382 26752 2388
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 26712 160 26740 2382
rect 26976 2304 27028 2310
rect 26976 2246 27028 2252
rect 26988 2106 27016 2246
rect 26976 2100 27028 2106
rect 26976 2042 27028 2048
rect 24582 54 24808 82
rect 20350 0 20406 54
rect 22466 0 22522 54
rect 24582 0 24638 54
rect 26698 0 26754 160
rect 28814 82 28870 160
rect 28920 82 28948 2382
rect 28814 54 28948 82
rect 30930 82 30986 160
rect 31036 82 31064 2382
rect 31772 1970 31800 6734
rect 32324 5642 32352 7142
rect 32600 6361 32628 7142
rect 32968 6798 32996 8894
rect 33032 7644 33340 7653
rect 33032 7642 33038 7644
rect 33094 7642 33118 7644
rect 33174 7642 33198 7644
rect 33254 7642 33278 7644
rect 33334 7642 33340 7644
rect 33094 7590 33096 7642
rect 33276 7590 33278 7642
rect 33032 7588 33038 7590
rect 33094 7588 33118 7590
rect 33174 7588 33198 7590
rect 33254 7588 33278 7590
rect 33334 7588 33340 7590
rect 33032 7579 33340 7588
rect 33428 6798 33456 8894
rect 33508 8492 33560 8498
rect 33508 8434 33560 8440
rect 33520 7546 33548 8434
rect 33508 7540 33560 7546
rect 33508 7482 33560 7488
rect 33612 6866 33640 9840
rect 33692 8424 33744 8430
rect 33692 8366 33744 8372
rect 33704 7546 33732 8366
rect 33888 7546 33916 9840
rect 33692 7540 33744 7546
rect 33692 7482 33744 7488
rect 33876 7540 33928 7546
rect 33876 7482 33928 7488
rect 33692 7404 33744 7410
rect 33692 7346 33744 7352
rect 33600 6860 33652 6866
rect 33600 6802 33652 6808
rect 33704 6798 33732 7346
rect 32956 6792 33008 6798
rect 33416 6792 33468 6798
rect 32956 6734 33008 6740
rect 33322 6760 33378 6769
rect 33416 6734 33468 6740
rect 33692 6792 33744 6798
rect 33692 6734 33744 6740
rect 33876 6792 33928 6798
rect 33876 6734 33928 6740
rect 34060 6792 34112 6798
rect 34060 6734 34112 6740
rect 33322 6695 33378 6704
rect 33336 6662 33364 6695
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 33600 6656 33652 6662
rect 33600 6598 33652 6604
rect 33692 6656 33744 6662
rect 33692 6598 33744 6604
rect 33032 6556 33340 6565
rect 33032 6554 33038 6556
rect 33094 6554 33118 6556
rect 33174 6554 33198 6556
rect 33254 6554 33278 6556
rect 33334 6554 33340 6556
rect 33094 6502 33096 6554
rect 33276 6502 33278 6554
rect 33032 6500 33038 6502
rect 33094 6500 33118 6502
rect 33174 6500 33198 6502
rect 33254 6500 33278 6502
rect 33334 6500 33340 6502
rect 33032 6491 33340 6500
rect 32586 6352 32642 6361
rect 32586 6287 32642 6296
rect 32312 5636 32364 5642
rect 32312 5578 32364 5584
rect 33032 5468 33340 5477
rect 33032 5466 33038 5468
rect 33094 5466 33118 5468
rect 33174 5466 33198 5468
rect 33254 5466 33278 5468
rect 33334 5466 33340 5468
rect 33094 5414 33096 5466
rect 33276 5414 33278 5466
rect 33032 5412 33038 5414
rect 33094 5412 33118 5414
rect 33174 5412 33198 5414
rect 33254 5412 33278 5414
rect 33334 5412 33340 5414
rect 33032 5403 33340 5412
rect 33612 5273 33640 6598
rect 33704 6458 33732 6598
rect 33692 6452 33744 6458
rect 33692 6394 33744 6400
rect 33598 5264 33654 5273
rect 33598 5199 33654 5208
rect 33888 5137 33916 6734
rect 33968 6656 34020 6662
rect 33968 6598 34020 6604
rect 33980 6390 34008 6598
rect 33968 6384 34020 6390
rect 33968 6326 34020 6332
rect 33874 5128 33930 5137
rect 33874 5063 33930 5072
rect 33416 4616 33468 4622
rect 33416 4558 33468 4564
rect 33032 4380 33340 4389
rect 33032 4378 33038 4380
rect 33094 4378 33118 4380
rect 33174 4378 33198 4380
rect 33254 4378 33278 4380
rect 33334 4378 33340 4380
rect 33094 4326 33096 4378
rect 33276 4326 33278 4378
rect 33032 4324 33038 4326
rect 33094 4324 33118 4326
rect 33174 4324 33198 4326
rect 33254 4324 33278 4326
rect 33334 4324 33340 4326
rect 33032 4315 33340 4324
rect 33032 3292 33340 3301
rect 33032 3290 33038 3292
rect 33094 3290 33118 3292
rect 33174 3290 33198 3292
rect 33254 3290 33278 3292
rect 33334 3290 33340 3292
rect 33094 3238 33096 3290
rect 33276 3238 33278 3290
rect 33032 3236 33038 3238
rect 33094 3236 33118 3238
rect 33174 3236 33198 3238
rect 33254 3236 33278 3238
rect 33334 3236 33340 3238
rect 33032 3227 33340 3236
rect 33140 2984 33192 2990
rect 33140 2926 33192 2932
rect 33152 2530 33180 2926
rect 33428 2582 33456 4558
rect 34072 2650 34100 6734
rect 34164 6662 34192 9840
rect 34440 7528 34468 9840
rect 34612 7540 34664 7546
rect 34440 7500 34612 7528
rect 34612 7482 34664 7488
rect 34716 7478 34744 9840
rect 34704 7472 34756 7478
rect 34704 7414 34756 7420
rect 34796 7404 34848 7410
rect 34796 7346 34848 7352
rect 34152 6656 34204 6662
rect 34152 6598 34204 6604
rect 34428 6656 34480 6662
rect 34428 6598 34480 6604
rect 34244 6316 34296 6322
rect 34244 6258 34296 6264
rect 34256 3466 34284 6258
rect 34440 4729 34468 6598
rect 34808 6458 34836 7346
rect 34992 7188 35020 9840
rect 35164 7200 35216 7206
rect 34992 7160 35164 7188
rect 35164 7142 35216 7148
rect 35268 6866 35296 9840
rect 35544 7528 35572 9840
rect 35716 7540 35768 7546
rect 35544 7500 35716 7528
rect 35716 7482 35768 7488
rect 35348 7404 35400 7410
rect 35348 7346 35400 7352
rect 35256 6860 35308 6866
rect 35256 6802 35308 6808
rect 35164 6792 35216 6798
rect 35164 6734 35216 6740
rect 34796 6452 34848 6458
rect 34796 6394 34848 6400
rect 34426 4720 34482 4729
rect 34426 4655 34482 4664
rect 35176 3534 35204 6734
rect 35360 6118 35388 7346
rect 35716 7336 35768 7342
rect 35716 7278 35768 7284
rect 35440 6724 35492 6730
rect 35440 6666 35492 6672
rect 35348 6112 35400 6118
rect 35348 6054 35400 6060
rect 35164 3528 35216 3534
rect 35164 3470 35216 3476
rect 34244 3460 34296 3466
rect 34244 3402 34296 3408
rect 35452 2650 35480 6666
rect 35728 2650 35756 7278
rect 35820 6866 35848 9840
rect 35900 7404 35952 7410
rect 35900 7346 35952 7352
rect 35808 6860 35860 6866
rect 35808 6802 35860 6808
rect 35912 6662 35940 7346
rect 35992 6724 36044 6730
rect 35992 6666 36044 6672
rect 35900 6656 35952 6662
rect 35900 6598 35952 6604
rect 36004 2990 36032 6666
rect 36096 6662 36124 9840
rect 36372 8514 36400 9840
rect 36372 8486 36584 8514
rect 36176 8356 36228 8362
rect 36176 8298 36228 8304
rect 36188 7478 36216 8298
rect 36176 7472 36228 7478
rect 36176 7414 36228 7420
rect 36556 7274 36584 8486
rect 36544 7268 36596 7274
rect 36544 7210 36596 7216
rect 36648 6914 36676 9840
rect 36924 7528 36952 9840
rect 37096 7540 37148 7546
rect 36924 7500 37096 7528
rect 37096 7482 37148 7488
rect 36820 7472 36872 7478
rect 36820 7414 36872 7420
rect 36648 6886 36768 6914
rect 36544 6724 36596 6730
rect 36544 6666 36596 6672
rect 36084 6656 36136 6662
rect 36084 6598 36136 6604
rect 36556 4622 36584 6666
rect 36740 6662 36768 6886
rect 36728 6656 36780 6662
rect 36728 6598 36780 6604
rect 36728 6248 36780 6254
rect 36728 6190 36780 6196
rect 36544 4616 36596 4622
rect 36544 4558 36596 4564
rect 35992 2984 36044 2990
rect 35992 2926 36044 2932
rect 34060 2644 34112 2650
rect 34060 2586 34112 2592
rect 35440 2644 35492 2650
rect 35440 2586 35492 2592
rect 35716 2644 35768 2650
rect 35716 2586 35768 2592
rect 32876 2502 33180 2530
rect 33416 2576 33468 2582
rect 33416 2518 33468 2524
rect 32876 2446 32904 2502
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 32956 2440 33008 2446
rect 32956 2382 33008 2388
rect 34888 2440 34940 2446
rect 34888 2382 34940 2388
rect 35164 2440 35216 2446
rect 35164 2382 35216 2388
rect 31760 1964 31812 1970
rect 31760 1906 31812 1912
rect 30930 54 31064 82
rect 32968 82 32996 2382
rect 33032 2204 33340 2213
rect 33032 2202 33038 2204
rect 33094 2202 33118 2204
rect 33174 2202 33198 2204
rect 33254 2202 33278 2204
rect 33334 2202 33340 2204
rect 33094 2150 33096 2202
rect 33276 2150 33278 2202
rect 33032 2148 33038 2150
rect 33094 2148 33118 2150
rect 33174 2148 33198 2150
rect 33254 2148 33278 2150
rect 33334 2148 33340 2150
rect 33032 2139 33340 2148
rect 34900 2038 34928 2382
rect 34888 2032 34940 2038
rect 34888 1974 34940 1980
rect 35176 160 35204 2382
rect 36740 2378 36768 6190
rect 36832 2650 36860 7414
rect 36912 7200 36964 7206
rect 36912 7142 36964 7148
rect 36924 7002 36952 7142
rect 36912 6996 36964 7002
rect 36912 6938 36964 6944
rect 37200 6866 37228 9840
rect 37188 6860 37240 6866
rect 37188 6802 37240 6808
rect 37476 6798 37504 9840
rect 37556 7404 37608 7410
rect 37556 7346 37608 7352
rect 37464 6792 37516 6798
rect 37464 6734 37516 6740
rect 37096 6724 37148 6730
rect 37096 6666 37148 6672
rect 37108 6322 37136 6666
rect 37096 6316 37148 6322
rect 37096 6258 37148 6264
rect 37280 6316 37332 6322
rect 37280 6258 37332 6264
rect 36820 2644 36872 2650
rect 36820 2586 36872 2592
rect 37292 2582 37320 6258
rect 37568 3126 37596 7346
rect 37648 6724 37700 6730
rect 37648 6666 37700 6672
rect 37556 3120 37608 3126
rect 37556 3062 37608 3068
rect 37660 2854 37688 6666
rect 37752 6662 37780 9840
rect 38028 8922 38056 9840
rect 38028 8894 38148 8922
rect 37924 7404 37976 7410
rect 37924 7346 37976 7352
rect 37832 7336 37884 7342
rect 37832 7278 37884 7284
rect 37740 6656 37792 6662
rect 37740 6598 37792 6604
rect 37648 2848 37700 2854
rect 37648 2790 37700 2796
rect 37844 2650 37872 7278
rect 37936 2922 37964 7346
rect 38120 6934 38148 8894
rect 38108 6928 38160 6934
rect 38304 6914 38332 9840
rect 38580 7290 38608 9840
rect 38856 7528 38884 9840
rect 39132 9330 39160 9840
rect 39132 9302 39252 9330
rect 39120 7540 39172 7546
rect 38856 7500 39120 7528
rect 39120 7482 39172 7488
rect 39028 7404 39080 7410
rect 39028 7346 39080 7352
rect 38580 7262 38976 7290
rect 38752 7200 38804 7206
rect 38752 7142 38804 7148
rect 38379 7100 38687 7109
rect 38379 7098 38385 7100
rect 38441 7098 38465 7100
rect 38521 7098 38545 7100
rect 38601 7098 38625 7100
rect 38681 7098 38687 7100
rect 38441 7046 38443 7098
rect 38623 7046 38625 7098
rect 38379 7044 38385 7046
rect 38441 7044 38465 7046
rect 38521 7044 38545 7046
rect 38601 7044 38625 7046
rect 38681 7044 38687 7046
rect 38379 7035 38687 7044
rect 38108 6870 38160 6876
rect 38212 6886 38332 6914
rect 38568 6928 38620 6934
rect 38212 6848 38240 6886
rect 38764 6914 38792 7142
rect 38948 6934 38976 7262
rect 38568 6870 38620 6876
rect 38672 6886 38792 6914
rect 38936 6928 38988 6934
rect 38212 6820 38516 6848
rect 38200 6724 38252 6730
rect 38200 6666 38252 6672
rect 38384 6724 38436 6730
rect 38384 6666 38436 6672
rect 38212 6458 38240 6666
rect 38396 6458 38424 6666
rect 38488 6662 38516 6820
rect 38476 6656 38528 6662
rect 38476 6598 38528 6604
rect 38580 6610 38608 6870
rect 38672 6798 38700 6886
rect 38936 6870 38988 6876
rect 38660 6792 38712 6798
rect 38660 6734 38712 6740
rect 38936 6656 38988 6662
rect 38580 6604 38936 6610
rect 38580 6598 38988 6604
rect 38580 6582 38976 6598
rect 38200 6452 38252 6458
rect 38200 6394 38252 6400
rect 38384 6452 38436 6458
rect 38384 6394 38436 6400
rect 39040 6254 39068 7346
rect 39120 7200 39172 7206
rect 39120 7142 39172 7148
rect 39132 6866 39160 7142
rect 39120 6860 39172 6866
rect 39120 6802 39172 6808
rect 39224 6730 39252 9302
rect 39408 8514 39436 9840
rect 39408 8486 39620 8514
rect 39592 7274 39620 8486
rect 39684 8378 39712 9840
rect 39684 8350 39896 8378
rect 39672 7404 39724 7410
rect 39672 7346 39724 7352
rect 39580 7268 39632 7274
rect 39580 7210 39632 7216
rect 39488 7200 39540 7206
rect 39488 7142 39540 7148
rect 39500 6798 39528 7142
rect 39488 6792 39540 6798
rect 39488 6734 39540 6740
rect 39212 6724 39264 6730
rect 39212 6666 39264 6672
rect 39028 6248 39080 6254
rect 39028 6190 39080 6196
rect 38379 6012 38687 6021
rect 38379 6010 38385 6012
rect 38441 6010 38465 6012
rect 38521 6010 38545 6012
rect 38601 6010 38625 6012
rect 38681 6010 38687 6012
rect 38441 5958 38443 6010
rect 38623 5958 38625 6010
rect 38379 5956 38385 5958
rect 38441 5956 38465 5958
rect 38521 5956 38545 5958
rect 38601 5956 38625 5958
rect 38681 5956 38687 5958
rect 38379 5947 38687 5956
rect 38379 4924 38687 4933
rect 38379 4922 38385 4924
rect 38441 4922 38465 4924
rect 38521 4922 38545 4924
rect 38601 4922 38625 4924
rect 38681 4922 38687 4924
rect 38441 4870 38443 4922
rect 38623 4870 38625 4922
rect 38379 4868 38385 4870
rect 38441 4868 38465 4870
rect 38521 4868 38545 4870
rect 38601 4868 38625 4870
rect 38681 4868 38687 4870
rect 38379 4859 38687 4868
rect 38379 3836 38687 3845
rect 38379 3834 38385 3836
rect 38441 3834 38465 3836
rect 38521 3834 38545 3836
rect 38601 3834 38625 3836
rect 38681 3834 38687 3836
rect 38441 3782 38443 3834
rect 38623 3782 38625 3834
rect 38379 3780 38385 3782
rect 38441 3780 38465 3782
rect 38521 3780 38545 3782
rect 38601 3780 38625 3782
rect 38681 3780 38687 3782
rect 38379 3771 38687 3780
rect 37924 2916 37976 2922
rect 37924 2858 37976 2864
rect 38379 2748 38687 2757
rect 38379 2746 38385 2748
rect 38441 2746 38465 2748
rect 38521 2746 38545 2748
rect 38601 2746 38625 2748
rect 38681 2746 38687 2748
rect 38441 2694 38443 2746
rect 38623 2694 38625 2746
rect 38379 2692 38385 2694
rect 38441 2692 38465 2694
rect 38521 2692 38545 2694
rect 38601 2692 38625 2694
rect 38681 2692 38687 2694
rect 38379 2683 38687 2692
rect 39684 2650 39712 7346
rect 39868 6866 39896 8350
rect 43726 7644 44034 7653
rect 43726 7642 43732 7644
rect 43788 7642 43812 7644
rect 43868 7642 43892 7644
rect 43948 7642 43972 7644
rect 44028 7642 44034 7644
rect 43788 7590 43790 7642
rect 43970 7590 43972 7642
rect 43726 7588 43732 7590
rect 43788 7588 43812 7590
rect 43868 7588 43892 7590
rect 43948 7588 43972 7590
rect 44028 7588 44034 7590
rect 43726 7579 44034 7588
rect 41420 7404 41472 7410
rect 41420 7346 41472 7352
rect 40960 7200 41012 7206
rect 40960 7142 41012 7148
rect 39856 6860 39908 6866
rect 39856 6802 39908 6808
rect 40972 6798 41000 7142
rect 40960 6792 41012 6798
rect 40960 6734 41012 6740
rect 41432 2650 41460 7346
rect 43352 7336 43404 7342
rect 43352 7278 43404 7284
rect 43364 2650 43392 7278
rect 43726 6556 44034 6565
rect 43726 6554 43732 6556
rect 43788 6554 43812 6556
rect 43868 6554 43892 6556
rect 43948 6554 43972 6556
rect 44028 6554 44034 6556
rect 43788 6502 43790 6554
rect 43970 6502 43972 6554
rect 43726 6500 43732 6502
rect 43788 6500 43812 6502
rect 43868 6500 43892 6502
rect 43948 6500 43972 6502
rect 44028 6500 44034 6502
rect 43726 6491 44034 6500
rect 43726 5468 44034 5477
rect 43726 5466 43732 5468
rect 43788 5466 43812 5468
rect 43868 5466 43892 5468
rect 43948 5466 43972 5468
rect 44028 5466 44034 5468
rect 43788 5414 43790 5466
rect 43970 5414 43972 5466
rect 43726 5412 43732 5414
rect 43788 5412 43812 5414
rect 43868 5412 43892 5414
rect 43948 5412 43972 5414
rect 44028 5412 44034 5414
rect 43726 5403 44034 5412
rect 43726 4380 44034 4389
rect 43726 4378 43732 4380
rect 43788 4378 43812 4380
rect 43868 4378 43892 4380
rect 43948 4378 43972 4380
rect 44028 4378 44034 4380
rect 43788 4326 43790 4378
rect 43970 4326 43972 4378
rect 43726 4324 43732 4326
rect 43788 4324 43812 4326
rect 43868 4324 43892 4326
rect 43948 4324 43972 4326
rect 44028 4324 44034 4326
rect 43726 4315 44034 4324
rect 43726 3292 44034 3301
rect 43726 3290 43732 3292
rect 43788 3290 43812 3292
rect 43868 3290 43892 3292
rect 43948 3290 43972 3292
rect 44028 3290 44034 3292
rect 43788 3238 43790 3290
rect 43970 3238 43972 3290
rect 43726 3236 43732 3238
rect 43788 3236 43812 3238
rect 43868 3236 43892 3238
rect 43948 3236 43972 3238
rect 44028 3236 44034 3238
rect 43726 3227 44034 3236
rect 37832 2644 37884 2650
rect 37832 2586 37884 2592
rect 39672 2644 39724 2650
rect 39672 2586 39724 2592
rect 41420 2644 41472 2650
rect 41420 2586 41472 2592
rect 43352 2644 43404 2650
rect 43352 2586 43404 2592
rect 37280 2576 37332 2582
rect 37280 2518 37332 2524
rect 37004 2440 37056 2446
rect 37004 2382 37056 2388
rect 37556 2440 37608 2446
rect 37556 2382 37608 2388
rect 39672 2440 39724 2446
rect 39672 2382 39724 2388
rect 41788 2440 41840 2446
rect 41788 2382 41840 2388
rect 43536 2440 43588 2446
rect 43536 2382 43588 2388
rect 36728 2372 36780 2378
rect 36728 2314 36780 2320
rect 37016 2106 37044 2382
rect 37004 2100 37056 2106
rect 37004 2042 37056 2048
rect 33046 82 33102 160
rect 32968 54 33102 82
rect 28814 0 28870 54
rect 30930 0 30986 54
rect 33046 0 33102 54
rect 35162 0 35218 160
rect 37278 82 37334 160
rect 37568 82 37596 2382
rect 37278 54 37596 82
rect 39394 82 39450 160
rect 39684 82 39712 2382
rect 39394 54 39712 82
rect 41510 82 41566 160
rect 41800 82 41828 2382
rect 41510 54 41828 82
rect 43548 82 43576 2382
rect 43726 2204 44034 2213
rect 43726 2202 43732 2204
rect 43788 2202 43812 2204
rect 43868 2202 43892 2204
rect 43948 2202 43972 2204
rect 44028 2202 44034 2204
rect 43788 2150 43790 2202
rect 43970 2150 43972 2202
rect 43726 2148 43732 2150
rect 43788 2148 43812 2150
rect 43868 2148 43892 2150
rect 43948 2148 43972 2150
rect 44028 2148 44034 2150
rect 43726 2139 44034 2148
rect 43626 82 43682 160
rect 43548 54 43682 82
rect 37278 0 37334 54
rect 39394 0 39450 54
rect 41510 0 41566 54
rect 43626 0 43682 54
<< via2 >>
rect 5814 7248 5870 7304
rect 6642 8064 6698 8120
rect 6303 7098 6359 7100
rect 6383 7098 6439 7100
rect 6463 7098 6519 7100
rect 6543 7098 6599 7100
rect 6303 7046 6349 7098
rect 6349 7046 6359 7098
rect 6383 7046 6413 7098
rect 6413 7046 6425 7098
rect 6425 7046 6439 7098
rect 6463 7046 6477 7098
rect 6477 7046 6489 7098
rect 6489 7046 6519 7098
rect 6543 7046 6553 7098
rect 6553 7046 6599 7098
rect 6303 7044 6359 7046
rect 6383 7044 6439 7046
rect 6463 7044 6519 7046
rect 6543 7044 6599 7046
rect 6303 6010 6359 6012
rect 6383 6010 6439 6012
rect 6463 6010 6519 6012
rect 6543 6010 6599 6012
rect 6303 5958 6349 6010
rect 6349 5958 6359 6010
rect 6383 5958 6413 6010
rect 6413 5958 6425 6010
rect 6425 5958 6439 6010
rect 6463 5958 6477 6010
rect 6477 5958 6489 6010
rect 6489 5958 6519 6010
rect 6543 5958 6553 6010
rect 6553 5958 6599 6010
rect 6303 5956 6359 5958
rect 6383 5956 6439 5958
rect 6463 5956 6519 5958
rect 6543 5956 6599 5958
rect 10046 7792 10102 7848
rect 10506 6704 10562 6760
rect 9862 6160 9918 6216
rect 6918 5072 6974 5128
rect 6303 4922 6359 4924
rect 6383 4922 6439 4924
rect 6463 4922 6519 4924
rect 6543 4922 6599 4924
rect 6303 4870 6349 4922
rect 6349 4870 6359 4922
rect 6383 4870 6413 4922
rect 6413 4870 6425 4922
rect 6425 4870 6439 4922
rect 6463 4870 6477 4922
rect 6477 4870 6489 4922
rect 6489 4870 6519 4922
rect 6543 4870 6553 4922
rect 6553 4870 6599 4922
rect 6303 4868 6359 4870
rect 6383 4868 6439 4870
rect 6463 4868 6519 4870
rect 6543 4868 6599 4870
rect 6303 3834 6359 3836
rect 6383 3834 6439 3836
rect 6463 3834 6519 3836
rect 6543 3834 6599 3836
rect 6303 3782 6349 3834
rect 6349 3782 6359 3834
rect 6383 3782 6413 3834
rect 6413 3782 6425 3834
rect 6425 3782 6439 3834
rect 6463 3782 6477 3834
rect 6477 3782 6489 3834
rect 6489 3782 6519 3834
rect 6543 3782 6553 3834
rect 6553 3782 6599 3834
rect 6303 3780 6359 3782
rect 6383 3780 6439 3782
rect 6463 3780 6519 3782
rect 6543 3780 6599 3782
rect 6303 2746 6359 2748
rect 6383 2746 6439 2748
rect 6463 2746 6519 2748
rect 6543 2746 6599 2748
rect 6303 2694 6349 2746
rect 6349 2694 6359 2746
rect 6383 2694 6413 2746
rect 6413 2694 6425 2746
rect 6425 2694 6439 2746
rect 6463 2694 6477 2746
rect 6477 2694 6489 2746
rect 6489 2694 6519 2746
rect 6543 2694 6553 2746
rect 6553 2694 6599 2746
rect 6303 2692 6359 2694
rect 6383 2692 6439 2694
rect 6463 2692 6519 2694
rect 6543 2692 6599 2694
rect 11150 7928 11206 7984
rect 11650 7642 11706 7644
rect 11730 7642 11786 7644
rect 11810 7642 11866 7644
rect 11890 7642 11946 7644
rect 11650 7590 11696 7642
rect 11696 7590 11706 7642
rect 11730 7590 11760 7642
rect 11760 7590 11772 7642
rect 11772 7590 11786 7642
rect 11810 7590 11824 7642
rect 11824 7590 11836 7642
rect 11836 7590 11866 7642
rect 11890 7590 11900 7642
rect 11900 7590 11946 7642
rect 11650 7588 11706 7590
rect 11730 7588 11786 7590
rect 11810 7588 11866 7590
rect 11890 7588 11946 7590
rect 11650 6554 11706 6556
rect 11730 6554 11786 6556
rect 11810 6554 11866 6556
rect 11890 6554 11946 6556
rect 11650 6502 11696 6554
rect 11696 6502 11706 6554
rect 11730 6502 11760 6554
rect 11760 6502 11772 6554
rect 11772 6502 11786 6554
rect 11810 6502 11824 6554
rect 11824 6502 11836 6554
rect 11836 6502 11866 6554
rect 11890 6502 11900 6554
rect 11900 6502 11946 6554
rect 11650 6500 11706 6502
rect 11730 6500 11786 6502
rect 11810 6500 11866 6502
rect 11890 6500 11946 6502
rect 11650 5466 11706 5468
rect 11730 5466 11786 5468
rect 11810 5466 11866 5468
rect 11890 5466 11946 5468
rect 11650 5414 11696 5466
rect 11696 5414 11706 5466
rect 11730 5414 11760 5466
rect 11760 5414 11772 5466
rect 11772 5414 11786 5466
rect 11810 5414 11824 5466
rect 11824 5414 11836 5466
rect 11836 5414 11866 5466
rect 11890 5414 11900 5466
rect 11900 5414 11946 5466
rect 11650 5412 11706 5414
rect 11730 5412 11786 5414
rect 11810 5412 11866 5414
rect 11890 5412 11946 5414
rect 12070 5516 12072 5536
rect 12072 5516 12124 5536
rect 12124 5516 12126 5536
rect 12070 5480 12126 5516
rect 12162 5344 12218 5400
rect 11650 4378 11706 4380
rect 11730 4378 11786 4380
rect 11810 4378 11866 4380
rect 11890 4378 11946 4380
rect 11650 4326 11696 4378
rect 11696 4326 11706 4378
rect 11730 4326 11760 4378
rect 11760 4326 11772 4378
rect 11772 4326 11786 4378
rect 11810 4326 11824 4378
rect 11824 4326 11836 4378
rect 11836 4326 11866 4378
rect 11890 4326 11900 4378
rect 11900 4326 11946 4378
rect 11650 4324 11706 4326
rect 11730 4324 11786 4326
rect 11810 4324 11866 4326
rect 11890 4324 11946 4326
rect 11650 3290 11706 3292
rect 11730 3290 11786 3292
rect 11810 3290 11866 3292
rect 11890 3290 11946 3292
rect 11650 3238 11696 3290
rect 11696 3238 11706 3290
rect 11730 3238 11760 3290
rect 11760 3238 11772 3290
rect 11772 3238 11786 3290
rect 11810 3238 11824 3290
rect 11824 3238 11836 3290
rect 11836 3238 11866 3290
rect 11890 3238 11900 3290
rect 11900 3238 11946 3290
rect 11650 3236 11706 3238
rect 11730 3236 11786 3238
rect 11810 3236 11866 3238
rect 11890 3236 11946 3238
rect 13634 6432 13690 6488
rect 14278 6840 14334 6896
rect 14278 5208 14334 5264
rect 14830 4664 14886 4720
rect 13266 4528 13322 4584
rect 16486 6568 16542 6624
rect 17498 8200 17554 8256
rect 16997 7098 17053 7100
rect 17077 7098 17133 7100
rect 17157 7098 17213 7100
rect 17237 7098 17293 7100
rect 16997 7046 17043 7098
rect 17043 7046 17053 7098
rect 17077 7046 17107 7098
rect 17107 7046 17119 7098
rect 17119 7046 17133 7098
rect 17157 7046 17171 7098
rect 17171 7046 17183 7098
rect 17183 7046 17213 7098
rect 17237 7046 17247 7098
rect 17247 7046 17293 7098
rect 16997 7044 17053 7046
rect 17077 7044 17133 7046
rect 17157 7044 17213 7046
rect 17237 7044 17293 7046
rect 16997 6010 17053 6012
rect 17077 6010 17133 6012
rect 17157 6010 17213 6012
rect 17237 6010 17293 6012
rect 16997 5958 17043 6010
rect 17043 5958 17053 6010
rect 17077 5958 17107 6010
rect 17107 5958 17119 6010
rect 17119 5958 17133 6010
rect 17157 5958 17171 6010
rect 17171 5958 17183 6010
rect 17183 5958 17213 6010
rect 17237 5958 17247 6010
rect 17247 5958 17293 6010
rect 16997 5956 17053 5958
rect 17077 5956 17133 5958
rect 17157 5956 17213 5958
rect 17237 5956 17293 5958
rect 17958 7112 18014 7168
rect 18418 6724 18474 6760
rect 18418 6704 18420 6724
rect 18420 6704 18472 6724
rect 18472 6704 18474 6724
rect 17774 6316 17830 6352
rect 17774 6296 17776 6316
rect 17776 6296 17828 6316
rect 17828 6296 17830 6316
rect 17866 6196 17868 6216
rect 17868 6196 17920 6216
rect 17920 6196 17922 6216
rect 17866 6160 17922 6196
rect 18786 6976 18842 7032
rect 19338 6024 19394 6080
rect 20718 7384 20774 7440
rect 20810 7112 20866 7168
rect 20626 6432 20682 6488
rect 21270 7792 21326 7848
rect 22344 7642 22400 7644
rect 22424 7642 22480 7644
rect 22504 7642 22560 7644
rect 22584 7642 22640 7644
rect 22344 7590 22390 7642
rect 22390 7590 22400 7642
rect 22424 7590 22454 7642
rect 22454 7590 22466 7642
rect 22466 7590 22480 7642
rect 22504 7590 22518 7642
rect 22518 7590 22530 7642
rect 22530 7590 22560 7642
rect 22584 7590 22594 7642
rect 22594 7590 22640 7642
rect 22344 7588 22400 7590
rect 22424 7588 22480 7590
rect 22504 7588 22560 7590
rect 22584 7588 22640 7590
rect 20994 6568 21050 6624
rect 22926 7928 22982 7984
rect 22344 6554 22400 6556
rect 22424 6554 22480 6556
rect 22504 6554 22560 6556
rect 22584 6554 22640 6556
rect 22344 6502 22390 6554
rect 22390 6502 22400 6554
rect 22424 6502 22454 6554
rect 22454 6502 22466 6554
rect 22466 6502 22480 6554
rect 22504 6502 22518 6554
rect 22518 6502 22530 6554
rect 22530 6502 22560 6554
rect 22584 6502 22594 6554
rect 22594 6502 22640 6554
rect 22344 6500 22400 6502
rect 22424 6500 22480 6502
rect 22504 6500 22560 6502
rect 22584 6500 22640 6502
rect 21178 5480 21234 5536
rect 24582 7268 24638 7304
rect 25134 8064 25190 8120
rect 24582 7248 24584 7268
rect 24584 7248 24636 7268
rect 24636 7248 24638 7268
rect 26882 8200 26938 8256
rect 22344 5466 22400 5468
rect 22424 5466 22480 5468
rect 22504 5466 22560 5468
rect 22584 5466 22640 5468
rect 22344 5414 22390 5466
rect 22390 5414 22400 5466
rect 22424 5414 22454 5466
rect 22454 5414 22466 5466
rect 22466 5414 22480 5466
rect 22504 5414 22518 5466
rect 22518 5414 22530 5466
rect 22530 5414 22560 5466
rect 22584 5414 22594 5466
rect 22594 5414 22640 5466
rect 22344 5412 22400 5414
rect 22424 5412 22480 5414
rect 22504 5412 22560 5414
rect 22584 5412 22640 5414
rect 22006 5344 22062 5400
rect 26790 6976 26846 7032
rect 25594 6160 25650 6216
rect 16997 4922 17053 4924
rect 17077 4922 17133 4924
rect 17157 4922 17213 4924
rect 17237 4922 17293 4924
rect 16997 4870 17043 4922
rect 17043 4870 17053 4922
rect 17077 4870 17107 4922
rect 17107 4870 17119 4922
rect 17119 4870 17133 4922
rect 17157 4870 17171 4922
rect 17171 4870 17183 4922
rect 17183 4870 17213 4922
rect 17237 4870 17247 4922
rect 17247 4870 17293 4922
rect 16997 4868 17053 4870
rect 17077 4868 17133 4870
rect 17157 4868 17213 4870
rect 17237 4868 17293 4870
rect 16118 4120 16174 4176
rect 16997 3834 17053 3836
rect 17077 3834 17133 3836
rect 17157 3834 17213 3836
rect 17237 3834 17293 3836
rect 16997 3782 17043 3834
rect 17043 3782 17053 3834
rect 17077 3782 17107 3834
rect 17107 3782 17119 3834
rect 17119 3782 17133 3834
rect 17157 3782 17171 3834
rect 17171 3782 17183 3834
rect 17183 3782 17213 3834
rect 17237 3782 17247 3834
rect 17247 3782 17293 3834
rect 16997 3780 17053 3782
rect 17077 3780 17133 3782
rect 17157 3780 17213 3782
rect 17237 3780 17293 3782
rect 16997 2746 17053 2748
rect 17077 2746 17133 2748
rect 17157 2746 17213 2748
rect 17237 2746 17293 2748
rect 16997 2694 17043 2746
rect 17043 2694 17053 2746
rect 17077 2694 17107 2746
rect 17107 2694 17119 2746
rect 17119 2694 17133 2746
rect 17157 2694 17171 2746
rect 17171 2694 17183 2746
rect 17183 2694 17213 2746
rect 17237 2694 17247 2746
rect 17247 2694 17293 2746
rect 16997 2692 17053 2694
rect 17077 2692 17133 2694
rect 17157 2692 17213 2694
rect 17237 2692 17293 2694
rect 24030 4528 24086 4584
rect 22344 4378 22400 4380
rect 22424 4378 22480 4380
rect 22504 4378 22560 4380
rect 22584 4378 22640 4380
rect 22344 4326 22390 4378
rect 22390 4326 22400 4378
rect 22424 4326 22454 4378
rect 22454 4326 22466 4378
rect 22466 4326 22480 4378
rect 22504 4326 22518 4378
rect 22518 4326 22530 4378
rect 22530 4326 22560 4378
rect 22584 4326 22594 4378
rect 22594 4326 22640 4378
rect 22344 4324 22400 4326
rect 22424 4324 22480 4326
rect 22504 4324 22560 4326
rect 22584 4324 22640 4326
rect 28446 7248 28502 7304
rect 27691 7098 27747 7100
rect 27771 7098 27827 7100
rect 27851 7098 27907 7100
rect 27931 7098 27987 7100
rect 27691 7046 27737 7098
rect 27737 7046 27747 7098
rect 27771 7046 27801 7098
rect 27801 7046 27813 7098
rect 27813 7046 27827 7098
rect 27851 7046 27865 7098
rect 27865 7046 27877 7098
rect 27877 7046 27907 7098
rect 27931 7046 27941 7098
rect 27941 7046 27987 7098
rect 27691 7044 27747 7046
rect 27771 7044 27827 7046
rect 27851 7044 27907 7046
rect 27931 7044 27987 7046
rect 27691 6010 27747 6012
rect 27771 6010 27827 6012
rect 27851 6010 27907 6012
rect 27931 6010 27987 6012
rect 27691 5958 27737 6010
rect 27737 5958 27747 6010
rect 27771 5958 27801 6010
rect 27801 5958 27813 6010
rect 27813 5958 27827 6010
rect 27851 5958 27865 6010
rect 27865 5958 27877 6010
rect 27877 5958 27907 6010
rect 27931 5958 27941 6010
rect 27941 5958 27987 6010
rect 27691 5956 27747 5958
rect 27771 5956 27827 5958
rect 27851 5956 27907 5958
rect 27931 5956 27987 5958
rect 27691 4922 27747 4924
rect 27771 4922 27827 4924
rect 27851 4922 27907 4924
rect 27931 4922 27987 4924
rect 27691 4870 27737 4922
rect 27737 4870 27747 4922
rect 27771 4870 27801 4922
rect 27801 4870 27813 4922
rect 27813 4870 27827 4922
rect 27851 4870 27865 4922
rect 27865 4870 27877 4922
rect 27877 4870 27907 4922
rect 27931 4870 27941 4922
rect 27941 4870 27987 4922
rect 27691 4868 27747 4870
rect 27771 4868 27827 4870
rect 27851 4868 27907 4870
rect 27931 4868 27987 4870
rect 26146 4120 26202 4176
rect 27691 3834 27747 3836
rect 27771 3834 27827 3836
rect 27851 3834 27907 3836
rect 27931 3834 27987 3836
rect 27691 3782 27737 3834
rect 27737 3782 27747 3834
rect 27771 3782 27801 3834
rect 27801 3782 27813 3834
rect 27813 3782 27827 3834
rect 27851 3782 27865 3834
rect 27865 3782 27877 3834
rect 27877 3782 27907 3834
rect 27931 3782 27941 3834
rect 27941 3782 27987 3834
rect 27691 3780 27747 3782
rect 27771 3780 27827 3782
rect 27851 3780 27907 3782
rect 27931 3780 27987 3782
rect 22344 3290 22400 3292
rect 22424 3290 22480 3292
rect 22504 3290 22560 3292
rect 22584 3290 22640 3292
rect 22344 3238 22390 3290
rect 22390 3238 22400 3290
rect 22424 3238 22454 3290
rect 22454 3238 22466 3290
rect 22466 3238 22480 3290
rect 22504 3238 22518 3290
rect 22518 3238 22530 3290
rect 22530 3238 22560 3290
rect 22584 3238 22594 3290
rect 22594 3238 22640 3290
rect 22344 3236 22400 3238
rect 22424 3236 22480 3238
rect 22504 3236 22560 3238
rect 22584 3236 22640 3238
rect 27691 2746 27747 2748
rect 27771 2746 27827 2748
rect 27851 2746 27907 2748
rect 27931 2746 27987 2748
rect 27691 2694 27737 2746
rect 27737 2694 27747 2746
rect 27771 2694 27801 2746
rect 27801 2694 27813 2746
rect 27813 2694 27827 2746
rect 27851 2694 27865 2746
rect 27865 2694 27877 2746
rect 27877 2694 27907 2746
rect 27931 2694 27941 2746
rect 27941 2694 27987 2746
rect 27691 2692 27747 2694
rect 27771 2692 27827 2694
rect 27851 2692 27907 2694
rect 27931 2692 27987 2694
rect 11650 2202 11706 2204
rect 11730 2202 11786 2204
rect 11810 2202 11866 2204
rect 11890 2202 11946 2204
rect 11650 2150 11696 2202
rect 11696 2150 11706 2202
rect 11730 2150 11760 2202
rect 11760 2150 11772 2202
rect 11772 2150 11786 2202
rect 11810 2150 11824 2202
rect 11824 2150 11836 2202
rect 11836 2150 11866 2202
rect 11890 2150 11900 2202
rect 11900 2150 11946 2202
rect 11650 2148 11706 2150
rect 11730 2148 11786 2150
rect 11810 2148 11866 2150
rect 11890 2148 11946 2150
rect 22344 2202 22400 2204
rect 22424 2202 22480 2204
rect 22504 2202 22560 2204
rect 22584 2202 22640 2204
rect 22344 2150 22390 2202
rect 22390 2150 22400 2202
rect 22424 2150 22454 2202
rect 22454 2150 22466 2202
rect 22466 2150 22480 2202
rect 22504 2150 22518 2202
rect 22518 2150 22530 2202
rect 22530 2150 22560 2202
rect 22584 2150 22594 2202
rect 22594 2150 22640 2202
rect 22344 2148 22400 2150
rect 22424 2148 22480 2150
rect 22504 2148 22560 2150
rect 22584 2148 22640 2150
rect 33038 7642 33094 7644
rect 33118 7642 33174 7644
rect 33198 7642 33254 7644
rect 33278 7642 33334 7644
rect 33038 7590 33084 7642
rect 33084 7590 33094 7642
rect 33118 7590 33148 7642
rect 33148 7590 33160 7642
rect 33160 7590 33174 7642
rect 33198 7590 33212 7642
rect 33212 7590 33224 7642
rect 33224 7590 33254 7642
rect 33278 7590 33288 7642
rect 33288 7590 33334 7642
rect 33038 7588 33094 7590
rect 33118 7588 33174 7590
rect 33198 7588 33254 7590
rect 33278 7588 33334 7590
rect 33322 6704 33378 6760
rect 33038 6554 33094 6556
rect 33118 6554 33174 6556
rect 33198 6554 33254 6556
rect 33278 6554 33334 6556
rect 33038 6502 33084 6554
rect 33084 6502 33094 6554
rect 33118 6502 33148 6554
rect 33148 6502 33160 6554
rect 33160 6502 33174 6554
rect 33198 6502 33212 6554
rect 33212 6502 33224 6554
rect 33224 6502 33254 6554
rect 33278 6502 33288 6554
rect 33288 6502 33334 6554
rect 33038 6500 33094 6502
rect 33118 6500 33174 6502
rect 33198 6500 33254 6502
rect 33278 6500 33334 6502
rect 32586 6296 32642 6352
rect 33038 5466 33094 5468
rect 33118 5466 33174 5468
rect 33198 5466 33254 5468
rect 33278 5466 33334 5468
rect 33038 5414 33084 5466
rect 33084 5414 33094 5466
rect 33118 5414 33148 5466
rect 33148 5414 33160 5466
rect 33160 5414 33174 5466
rect 33198 5414 33212 5466
rect 33212 5414 33224 5466
rect 33224 5414 33254 5466
rect 33278 5414 33288 5466
rect 33288 5414 33334 5466
rect 33038 5412 33094 5414
rect 33118 5412 33174 5414
rect 33198 5412 33254 5414
rect 33278 5412 33334 5414
rect 33598 5208 33654 5264
rect 33874 5072 33930 5128
rect 33038 4378 33094 4380
rect 33118 4378 33174 4380
rect 33198 4378 33254 4380
rect 33278 4378 33334 4380
rect 33038 4326 33084 4378
rect 33084 4326 33094 4378
rect 33118 4326 33148 4378
rect 33148 4326 33160 4378
rect 33160 4326 33174 4378
rect 33198 4326 33212 4378
rect 33212 4326 33224 4378
rect 33224 4326 33254 4378
rect 33278 4326 33288 4378
rect 33288 4326 33334 4378
rect 33038 4324 33094 4326
rect 33118 4324 33174 4326
rect 33198 4324 33254 4326
rect 33278 4324 33334 4326
rect 33038 3290 33094 3292
rect 33118 3290 33174 3292
rect 33198 3290 33254 3292
rect 33278 3290 33334 3292
rect 33038 3238 33084 3290
rect 33084 3238 33094 3290
rect 33118 3238 33148 3290
rect 33148 3238 33160 3290
rect 33160 3238 33174 3290
rect 33198 3238 33212 3290
rect 33212 3238 33224 3290
rect 33224 3238 33254 3290
rect 33278 3238 33288 3290
rect 33288 3238 33334 3290
rect 33038 3236 33094 3238
rect 33118 3236 33174 3238
rect 33198 3236 33254 3238
rect 33278 3236 33334 3238
rect 34426 4664 34482 4720
rect 33038 2202 33094 2204
rect 33118 2202 33174 2204
rect 33198 2202 33254 2204
rect 33278 2202 33334 2204
rect 33038 2150 33084 2202
rect 33084 2150 33094 2202
rect 33118 2150 33148 2202
rect 33148 2150 33160 2202
rect 33160 2150 33174 2202
rect 33198 2150 33212 2202
rect 33212 2150 33224 2202
rect 33224 2150 33254 2202
rect 33278 2150 33288 2202
rect 33288 2150 33334 2202
rect 33038 2148 33094 2150
rect 33118 2148 33174 2150
rect 33198 2148 33254 2150
rect 33278 2148 33334 2150
rect 38385 7098 38441 7100
rect 38465 7098 38521 7100
rect 38545 7098 38601 7100
rect 38625 7098 38681 7100
rect 38385 7046 38431 7098
rect 38431 7046 38441 7098
rect 38465 7046 38495 7098
rect 38495 7046 38507 7098
rect 38507 7046 38521 7098
rect 38545 7046 38559 7098
rect 38559 7046 38571 7098
rect 38571 7046 38601 7098
rect 38625 7046 38635 7098
rect 38635 7046 38681 7098
rect 38385 7044 38441 7046
rect 38465 7044 38521 7046
rect 38545 7044 38601 7046
rect 38625 7044 38681 7046
rect 38385 6010 38441 6012
rect 38465 6010 38521 6012
rect 38545 6010 38601 6012
rect 38625 6010 38681 6012
rect 38385 5958 38431 6010
rect 38431 5958 38441 6010
rect 38465 5958 38495 6010
rect 38495 5958 38507 6010
rect 38507 5958 38521 6010
rect 38545 5958 38559 6010
rect 38559 5958 38571 6010
rect 38571 5958 38601 6010
rect 38625 5958 38635 6010
rect 38635 5958 38681 6010
rect 38385 5956 38441 5958
rect 38465 5956 38521 5958
rect 38545 5956 38601 5958
rect 38625 5956 38681 5958
rect 38385 4922 38441 4924
rect 38465 4922 38521 4924
rect 38545 4922 38601 4924
rect 38625 4922 38681 4924
rect 38385 4870 38431 4922
rect 38431 4870 38441 4922
rect 38465 4870 38495 4922
rect 38495 4870 38507 4922
rect 38507 4870 38521 4922
rect 38545 4870 38559 4922
rect 38559 4870 38571 4922
rect 38571 4870 38601 4922
rect 38625 4870 38635 4922
rect 38635 4870 38681 4922
rect 38385 4868 38441 4870
rect 38465 4868 38521 4870
rect 38545 4868 38601 4870
rect 38625 4868 38681 4870
rect 38385 3834 38441 3836
rect 38465 3834 38521 3836
rect 38545 3834 38601 3836
rect 38625 3834 38681 3836
rect 38385 3782 38431 3834
rect 38431 3782 38441 3834
rect 38465 3782 38495 3834
rect 38495 3782 38507 3834
rect 38507 3782 38521 3834
rect 38545 3782 38559 3834
rect 38559 3782 38571 3834
rect 38571 3782 38601 3834
rect 38625 3782 38635 3834
rect 38635 3782 38681 3834
rect 38385 3780 38441 3782
rect 38465 3780 38521 3782
rect 38545 3780 38601 3782
rect 38625 3780 38681 3782
rect 38385 2746 38441 2748
rect 38465 2746 38521 2748
rect 38545 2746 38601 2748
rect 38625 2746 38681 2748
rect 38385 2694 38431 2746
rect 38431 2694 38441 2746
rect 38465 2694 38495 2746
rect 38495 2694 38507 2746
rect 38507 2694 38521 2746
rect 38545 2694 38559 2746
rect 38559 2694 38571 2746
rect 38571 2694 38601 2746
rect 38625 2694 38635 2746
rect 38635 2694 38681 2746
rect 38385 2692 38441 2694
rect 38465 2692 38521 2694
rect 38545 2692 38601 2694
rect 38625 2692 38681 2694
rect 43732 7642 43788 7644
rect 43812 7642 43868 7644
rect 43892 7642 43948 7644
rect 43972 7642 44028 7644
rect 43732 7590 43778 7642
rect 43778 7590 43788 7642
rect 43812 7590 43842 7642
rect 43842 7590 43854 7642
rect 43854 7590 43868 7642
rect 43892 7590 43906 7642
rect 43906 7590 43918 7642
rect 43918 7590 43948 7642
rect 43972 7590 43982 7642
rect 43982 7590 44028 7642
rect 43732 7588 43788 7590
rect 43812 7588 43868 7590
rect 43892 7588 43948 7590
rect 43972 7588 44028 7590
rect 43732 6554 43788 6556
rect 43812 6554 43868 6556
rect 43892 6554 43948 6556
rect 43972 6554 44028 6556
rect 43732 6502 43778 6554
rect 43778 6502 43788 6554
rect 43812 6502 43842 6554
rect 43842 6502 43854 6554
rect 43854 6502 43868 6554
rect 43892 6502 43906 6554
rect 43906 6502 43918 6554
rect 43918 6502 43948 6554
rect 43972 6502 43982 6554
rect 43982 6502 44028 6554
rect 43732 6500 43788 6502
rect 43812 6500 43868 6502
rect 43892 6500 43948 6502
rect 43972 6500 44028 6502
rect 43732 5466 43788 5468
rect 43812 5466 43868 5468
rect 43892 5466 43948 5468
rect 43972 5466 44028 5468
rect 43732 5414 43778 5466
rect 43778 5414 43788 5466
rect 43812 5414 43842 5466
rect 43842 5414 43854 5466
rect 43854 5414 43868 5466
rect 43892 5414 43906 5466
rect 43906 5414 43918 5466
rect 43918 5414 43948 5466
rect 43972 5414 43982 5466
rect 43982 5414 44028 5466
rect 43732 5412 43788 5414
rect 43812 5412 43868 5414
rect 43892 5412 43948 5414
rect 43972 5412 44028 5414
rect 43732 4378 43788 4380
rect 43812 4378 43868 4380
rect 43892 4378 43948 4380
rect 43972 4378 44028 4380
rect 43732 4326 43778 4378
rect 43778 4326 43788 4378
rect 43812 4326 43842 4378
rect 43842 4326 43854 4378
rect 43854 4326 43868 4378
rect 43892 4326 43906 4378
rect 43906 4326 43918 4378
rect 43918 4326 43948 4378
rect 43972 4326 43982 4378
rect 43982 4326 44028 4378
rect 43732 4324 43788 4326
rect 43812 4324 43868 4326
rect 43892 4324 43948 4326
rect 43972 4324 44028 4326
rect 43732 3290 43788 3292
rect 43812 3290 43868 3292
rect 43892 3290 43948 3292
rect 43972 3290 44028 3292
rect 43732 3238 43778 3290
rect 43778 3238 43788 3290
rect 43812 3238 43842 3290
rect 43842 3238 43854 3290
rect 43854 3238 43868 3290
rect 43892 3238 43906 3290
rect 43906 3238 43918 3290
rect 43918 3238 43948 3290
rect 43972 3238 43982 3290
rect 43982 3238 44028 3290
rect 43732 3236 43788 3238
rect 43812 3236 43868 3238
rect 43892 3236 43948 3238
rect 43972 3236 44028 3238
rect 43732 2202 43788 2204
rect 43812 2202 43868 2204
rect 43892 2202 43948 2204
rect 43972 2202 44028 2204
rect 43732 2150 43778 2202
rect 43778 2150 43788 2202
rect 43812 2150 43842 2202
rect 43842 2150 43854 2202
rect 43854 2150 43868 2202
rect 43892 2150 43906 2202
rect 43906 2150 43918 2202
rect 43918 2150 43948 2202
rect 43972 2150 43982 2202
rect 43982 2150 44028 2202
rect 43732 2148 43788 2150
rect 43812 2148 43868 2150
rect 43892 2148 43948 2150
rect 43972 2148 44028 2150
<< metal3 >>
rect 17493 8258 17559 8261
rect 26877 8258 26943 8261
rect 17493 8256 26943 8258
rect 17493 8200 17498 8256
rect 17554 8200 26882 8256
rect 26938 8200 26943 8256
rect 17493 8198 26943 8200
rect 17493 8195 17559 8198
rect 26877 8195 26943 8198
rect 6637 8122 6703 8125
rect 25129 8122 25195 8125
rect 6637 8120 25195 8122
rect 6637 8064 6642 8120
rect 6698 8064 25134 8120
rect 25190 8064 25195 8120
rect 6637 8062 25195 8064
rect 6637 8059 6703 8062
rect 25129 8059 25195 8062
rect 11145 7986 11211 7989
rect 22921 7986 22987 7989
rect 11145 7984 22987 7986
rect 11145 7928 11150 7984
rect 11206 7928 22926 7984
rect 22982 7928 22987 7984
rect 11145 7926 22987 7928
rect 11145 7923 11211 7926
rect 22921 7923 22987 7926
rect 10041 7850 10107 7853
rect 21265 7850 21331 7853
rect 10041 7848 21331 7850
rect 10041 7792 10046 7848
rect 10102 7792 21270 7848
rect 21326 7792 21331 7848
rect 10041 7790 21331 7792
rect 10041 7787 10107 7790
rect 21265 7787 21331 7790
rect 11640 7648 11956 7649
rect 11640 7584 11646 7648
rect 11710 7584 11726 7648
rect 11790 7584 11806 7648
rect 11870 7584 11886 7648
rect 11950 7584 11956 7648
rect 11640 7583 11956 7584
rect 22334 7648 22650 7649
rect 22334 7584 22340 7648
rect 22404 7584 22420 7648
rect 22484 7584 22500 7648
rect 22564 7584 22580 7648
rect 22644 7584 22650 7648
rect 22334 7583 22650 7584
rect 33028 7648 33344 7649
rect 33028 7584 33034 7648
rect 33098 7584 33114 7648
rect 33178 7584 33194 7648
rect 33258 7584 33274 7648
rect 33338 7584 33344 7648
rect 33028 7583 33344 7584
rect 43722 7648 44038 7649
rect 43722 7584 43728 7648
rect 43792 7584 43808 7648
rect 43872 7584 43888 7648
rect 43952 7584 43968 7648
rect 44032 7584 44038 7648
rect 43722 7583 44038 7584
rect 20713 7442 20779 7445
rect 20713 7440 28458 7442
rect 20713 7384 20718 7440
rect 20774 7384 28458 7440
rect 20713 7382 28458 7384
rect 20713 7379 20779 7382
rect 28398 7309 28458 7382
rect 5809 7306 5875 7309
rect 24577 7306 24643 7309
rect 5809 7304 24643 7306
rect 5809 7248 5814 7304
rect 5870 7248 24582 7304
rect 24638 7248 24643 7304
rect 5809 7246 24643 7248
rect 28398 7304 28507 7309
rect 28398 7248 28446 7304
rect 28502 7248 28507 7304
rect 28398 7246 28507 7248
rect 5809 7243 5875 7246
rect 24577 7243 24643 7246
rect 28441 7243 28507 7246
rect 17953 7170 18019 7173
rect 20805 7170 20871 7173
rect 17953 7168 20871 7170
rect 17953 7112 17958 7168
rect 18014 7112 20810 7168
rect 20866 7112 20871 7168
rect 17953 7110 20871 7112
rect 17953 7107 18019 7110
rect 20805 7107 20871 7110
rect 6293 7104 6609 7105
rect 6293 7040 6299 7104
rect 6363 7040 6379 7104
rect 6443 7040 6459 7104
rect 6523 7040 6539 7104
rect 6603 7040 6609 7104
rect 6293 7039 6609 7040
rect 16987 7104 17303 7105
rect 16987 7040 16993 7104
rect 17057 7040 17073 7104
rect 17137 7040 17153 7104
rect 17217 7040 17233 7104
rect 17297 7040 17303 7104
rect 16987 7039 17303 7040
rect 27681 7104 27997 7105
rect 27681 7040 27687 7104
rect 27751 7040 27767 7104
rect 27831 7040 27847 7104
rect 27911 7040 27927 7104
rect 27991 7040 27997 7104
rect 27681 7039 27997 7040
rect 38375 7104 38691 7105
rect 38375 7040 38381 7104
rect 38445 7040 38461 7104
rect 38525 7040 38541 7104
rect 38605 7040 38621 7104
rect 38685 7040 38691 7104
rect 38375 7039 38691 7040
rect 18781 7034 18847 7037
rect 26785 7034 26851 7037
rect 18781 7032 26851 7034
rect 18781 6976 18786 7032
rect 18842 6976 26790 7032
rect 26846 6976 26851 7032
rect 18781 6974 26851 6976
rect 18781 6971 18847 6974
rect 26785 6971 26851 6974
rect 14273 6898 14339 6901
rect 14273 6896 22110 6898
rect 14273 6840 14278 6896
rect 14334 6840 22110 6896
rect 14273 6838 22110 6840
rect 14273 6835 14339 6838
rect 10501 6762 10567 6765
rect 18413 6762 18479 6765
rect 10501 6760 18479 6762
rect 10501 6704 10506 6760
rect 10562 6704 18418 6760
rect 18474 6704 18479 6760
rect 10501 6702 18479 6704
rect 22050 6762 22110 6838
rect 33317 6762 33383 6765
rect 22050 6760 33383 6762
rect 22050 6704 33322 6760
rect 33378 6704 33383 6760
rect 22050 6702 33383 6704
rect 10501 6699 10567 6702
rect 18413 6699 18479 6702
rect 33317 6699 33383 6702
rect 16481 6626 16547 6629
rect 20989 6626 21055 6629
rect 16481 6624 21055 6626
rect 16481 6568 16486 6624
rect 16542 6568 20994 6624
rect 21050 6568 21055 6624
rect 16481 6566 21055 6568
rect 16481 6563 16547 6566
rect 20989 6563 21055 6566
rect 11640 6560 11956 6561
rect 11640 6496 11646 6560
rect 11710 6496 11726 6560
rect 11790 6496 11806 6560
rect 11870 6496 11886 6560
rect 11950 6496 11956 6560
rect 11640 6495 11956 6496
rect 22334 6560 22650 6561
rect 22334 6496 22340 6560
rect 22404 6496 22420 6560
rect 22484 6496 22500 6560
rect 22564 6496 22580 6560
rect 22644 6496 22650 6560
rect 22334 6495 22650 6496
rect 33028 6560 33344 6561
rect 33028 6496 33034 6560
rect 33098 6496 33114 6560
rect 33178 6496 33194 6560
rect 33258 6496 33274 6560
rect 33338 6496 33344 6560
rect 33028 6495 33344 6496
rect 43722 6560 44038 6561
rect 43722 6496 43728 6560
rect 43792 6496 43808 6560
rect 43872 6496 43888 6560
rect 43952 6496 43968 6560
rect 44032 6496 44038 6560
rect 43722 6495 44038 6496
rect 13629 6490 13695 6493
rect 20621 6490 20687 6493
rect 13629 6488 20687 6490
rect 13629 6432 13634 6488
rect 13690 6432 20626 6488
rect 20682 6432 20687 6488
rect 13629 6430 20687 6432
rect 13629 6427 13695 6430
rect 20621 6427 20687 6430
rect 17769 6354 17835 6357
rect 32581 6354 32647 6357
rect 17769 6352 32647 6354
rect 17769 6296 17774 6352
rect 17830 6296 32586 6352
rect 32642 6296 32647 6352
rect 17769 6294 32647 6296
rect 17769 6291 17835 6294
rect 32581 6291 32647 6294
rect 9857 6218 9923 6221
rect 17861 6218 17927 6221
rect 25589 6218 25655 6221
rect 9857 6216 17602 6218
rect 9857 6160 9862 6216
rect 9918 6160 17602 6216
rect 9857 6158 17602 6160
rect 9857 6155 9923 6158
rect 17542 6082 17602 6158
rect 17861 6216 25655 6218
rect 17861 6160 17866 6216
rect 17922 6160 25594 6216
rect 25650 6160 25655 6216
rect 17861 6158 25655 6160
rect 17861 6155 17927 6158
rect 25589 6155 25655 6158
rect 19333 6082 19399 6085
rect 17542 6080 19399 6082
rect 17542 6024 19338 6080
rect 19394 6024 19399 6080
rect 17542 6022 19399 6024
rect 19333 6019 19399 6022
rect 6293 6016 6609 6017
rect 6293 5952 6299 6016
rect 6363 5952 6379 6016
rect 6443 5952 6459 6016
rect 6523 5952 6539 6016
rect 6603 5952 6609 6016
rect 6293 5951 6609 5952
rect 16987 6016 17303 6017
rect 16987 5952 16993 6016
rect 17057 5952 17073 6016
rect 17137 5952 17153 6016
rect 17217 5952 17233 6016
rect 17297 5952 17303 6016
rect 16987 5951 17303 5952
rect 27681 6016 27997 6017
rect 27681 5952 27687 6016
rect 27751 5952 27767 6016
rect 27831 5952 27847 6016
rect 27911 5952 27927 6016
rect 27991 5952 27997 6016
rect 27681 5951 27997 5952
rect 38375 6016 38691 6017
rect 38375 5952 38381 6016
rect 38445 5952 38461 6016
rect 38525 5952 38541 6016
rect 38605 5952 38621 6016
rect 38685 5952 38691 6016
rect 38375 5951 38691 5952
rect 12065 5538 12131 5541
rect 21173 5538 21239 5541
rect 12065 5536 21239 5538
rect 12065 5480 12070 5536
rect 12126 5480 21178 5536
rect 21234 5480 21239 5536
rect 12065 5478 21239 5480
rect 12065 5475 12131 5478
rect 21173 5475 21239 5478
rect 11640 5472 11956 5473
rect 11640 5408 11646 5472
rect 11710 5408 11726 5472
rect 11790 5408 11806 5472
rect 11870 5408 11886 5472
rect 11950 5408 11956 5472
rect 11640 5407 11956 5408
rect 22334 5472 22650 5473
rect 22334 5408 22340 5472
rect 22404 5408 22420 5472
rect 22484 5408 22500 5472
rect 22564 5408 22580 5472
rect 22644 5408 22650 5472
rect 22334 5407 22650 5408
rect 33028 5472 33344 5473
rect 33028 5408 33034 5472
rect 33098 5408 33114 5472
rect 33178 5408 33194 5472
rect 33258 5408 33274 5472
rect 33338 5408 33344 5472
rect 33028 5407 33344 5408
rect 43722 5472 44038 5473
rect 43722 5408 43728 5472
rect 43792 5408 43808 5472
rect 43872 5408 43888 5472
rect 43952 5408 43968 5472
rect 44032 5408 44038 5472
rect 43722 5407 44038 5408
rect 12157 5402 12223 5405
rect 22001 5402 22067 5405
rect 12157 5400 22067 5402
rect 12157 5344 12162 5400
rect 12218 5344 22006 5400
rect 22062 5344 22067 5400
rect 12157 5342 22067 5344
rect 12157 5339 12223 5342
rect 22001 5339 22067 5342
rect 14273 5266 14339 5269
rect 33593 5266 33659 5269
rect 14273 5264 33659 5266
rect 14273 5208 14278 5264
rect 14334 5208 33598 5264
rect 33654 5208 33659 5264
rect 14273 5206 33659 5208
rect 14273 5203 14339 5206
rect 33593 5203 33659 5206
rect 6913 5130 6979 5133
rect 33869 5130 33935 5133
rect 6913 5128 33935 5130
rect 6913 5072 6918 5128
rect 6974 5072 33874 5128
rect 33930 5072 33935 5128
rect 6913 5070 33935 5072
rect 6913 5067 6979 5070
rect 33869 5067 33935 5070
rect 6293 4928 6609 4929
rect 6293 4864 6299 4928
rect 6363 4864 6379 4928
rect 6443 4864 6459 4928
rect 6523 4864 6539 4928
rect 6603 4864 6609 4928
rect 6293 4863 6609 4864
rect 16987 4928 17303 4929
rect 16987 4864 16993 4928
rect 17057 4864 17073 4928
rect 17137 4864 17153 4928
rect 17217 4864 17233 4928
rect 17297 4864 17303 4928
rect 16987 4863 17303 4864
rect 27681 4928 27997 4929
rect 27681 4864 27687 4928
rect 27751 4864 27767 4928
rect 27831 4864 27847 4928
rect 27911 4864 27927 4928
rect 27991 4864 27997 4928
rect 27681 4863 27997 4864
rect 38375 4928 38691 4929
rect 38375 4864 38381 4928
rect 38445 4864 38461 4928
rect 38525 4864 38541 4928
rect 38605 4864 38621 4928
rect 38685 4864 38691 4928
rect 38375 4863 38691 4864
rect 14825 4722 14891 4725
rect 34421 4722 34487 4725
rect 14825 4720 34487 4722
rect 14825 4664 14830 4720
rect 14886 4664 34426 4720
rect 34482 4664 34487 4720
rect 14825 4662 34487 4664
rect 14825 4659 14891 4662
rect 34421 4659 34487 4662
rect 13261 4586 13327 4589
rect 24025 4586 24091 4589
rect 13261 4584 24091 4586
rect 13261 4528 13266 4584
rect 13322 4528 24030 4584
rect 24086 4528 24091 4584
rect 13261 4526 24091 4528
rect 13261 4523 13327 4526
rect 24025 4523 24091 4526
rect 11640 4384 11956 4385
rect 11640 4320 11646 4384
rect 11710 4320 11726 4384
rect 11790 4320 11806 4384
rect 11870 4320 11886 4384
rect 11950 4320 11956 4384
rect 11640 4319 11956 4320
rect 22334 4384 22650 4385
rect 22334 4320 22340 4384
rect 22404 4320 22420 4384
rect 22484 4320 22500 4384
rect 22564 4320 22580 4384
rect 22644 4320 22650 4384
rect 22334 4319 22650 4320
rect 33028 4384 33344 4385
rect 33028 4320 33034 4384
rect 33098 4320 33114 4384
rect 33178 4320 33194 4384
rect 33258 4320 33274 4384
rect 33338 4320 33344 4384
rect 33028 4319 33344 4320
rect 43722 4384 44038 4385
rect 43722 4320 43728 4384
rect 43792 4320 43808 4384
rect 43872 4320 43888 4384
rect 43952 4320 43968 4384
rect 44032 4320 44038 4384
rect 43722 4319 44038 4320
rect 16113 4178 16179 4181
rect 26141 4178 26207 4181
rect 16113 4176 26207 4178
rect 16113 4120 16118 4176
rect 16174 4120 26146 4176
rect 26202 4120 26207 4176
rect 16113 4118 26207 4120
rect 16113 4115 16179 4118
rect 26141 4115 26207 4118
rect 6293 3840 6609 3841
rect 6293 3776 6299 3840
rect 6363 3776 6379 3840
rect 6443 3776 6459 3840
rect 6523 3776 6539 3840
rect 6603 3776 6609 3840
rect 6293 3775 6609 3776
rect 16987 3840 17303 3841
rect 16987 3776 16993 3840
rect 17057 3776 17073 3840
rect 17137 3776 17153 3840
rect 17217 3776 17233 3840
rect 17297 3776 17303 3840
rect 16987 3775 17303 3776
rect 27681 3840 27997 3841
rect 27681 3776 27687 3840
rect 27751 3776 27767 3840
rect 27831 3776 27847 3840
rect 27911 3776 27927 3840
rect 27991 3776 27997 3840
rect 27681 3775 27997 3776
rect 38375 3840 38691 3841
rect 38375 3776 38381 3840
rect 38445 3776 38461 3840
rect 38525 3776 38541 3840
rect 38605 3776 38621 3840
rect 38685 3776 38691 3840
rect 38375 3775 38691 3776
rect 11640 3296 11956 3297
rect 11640 3232 11646 3296
rect 11710 3232 11726 3296
rect 11790 3232 11806 3296
rect 11870 3232 11886 3296
rect 11950 3232 11956 3296
rect 11640 3231 11956 3232
rect 22334 3296 22650 3297
rect 22334 3232 22340 3296
rect 22404 3232 22420 3296
rect 22484 3232 22500 3296
rect 22564 3232 22580 3296
rect 22644 3232 22650 3296
rect 22334 3231 22650 3232
rect 33028 3296 33344 3297
rect 33028 3232 33034 3296
rect 33098 3232 33114 3296
rect 33178 3232 33194 3296
rect 33258 3232 33274 3296
rect 33338 3232 33344 3296
rect 33028 3231 33344 3232
rect 43722 3296 44038 3297
rect 43722 3232 43728 3296
rect 43792 3232 43808 3296
rect 43872 3232 43888 3296
rect 43952 3232 43968 3296
rect 44032 3232 44038 3296
rect 43722 3231 44038 3232
rect 6293 2752 6609 2753
rect 6293 2688 6299 2752
rect 6363 2688 6379 2752
rect 6443 2688 6459 2752
rect 6523 2688 6539 2752
rect 6603 2688 6609 2752
rect 6293 2687 6609 2688
rect 16987 2752 17303 2753
rect 16987 2688 16993 2752
rect 17057 2688 17073 2752
rect 17137 2688 17153 2752
rect 17217 2688 17233 2752
rect 17297 2688 17303 2752
rect 16987 2687 17303 2688
rect 27681 2752 27997 2753
rect 27681 2688 27687 2752
rect 27751 2688 27767 2752
rect 27831 2688 27847 2752
rect 27911 2688 27927 2752
rect 27991 2688 27997 2752
rect 27681 2687 27997 2688
rect 38375 2752 38691 2753
rect 38375 2688 38381 2752
rect 38445 2688 38461 2752
rect 38525 2688 38541 2752
rect 38605 2688 38621 2752
rect 38685 2688 38691 2752
rect 38375 2687 38691 2688
rect 11640 2208 11956 2209
rect 11640 2144 11646 2208
rect 11710 2144 11726 2208
rect 11790 2144 11806 2208
rect 11870 2144 11886 2208
rect 11950 2144 11956 2208
rect 11640 2143 11956 2144
rect 22334 2208 22650 2209
rect 22334 2144 22340 2208
rect 22404 2144 22420 2208
rect 22484 2144 22500 2208
rect 22564 2144 22580 2208
rect 22644 2144 22650 2208
rect 22334 2143 22650 2144
rect 33028 2208 33344 2209
rect 33028 2144 33034 2208
rect 33098 2144 33114 2208
rect 33178 2144 33194 2208
rect 33258 2144 33274 2208
rect 33338 2144 33344 2208
rect 33028 2143 33344 2144
rect 43722 2208 44038 2209
rect 43722 2144 43728 2208
rect 43792 2144 43808 2208
rect 43872 2144 43888 2208
rect 43952 2144 43968 2208
rect 44032 2144 44038 2208
rect 43722 2143 44038 2144
<< via3 >>
rect 11646 7644 11710 7648
rect 11646 7588 11650 7644
rect 11650 7588 11706 7644
rect 11706 7588 11710 7644
rect 11646 7584 11710 7588
rect 11726 7644 11790 7648
rect 11726 7588 11730 7644
rect 11730 7588 11786 7644
rect 11786 7588 11790 7644
rect 11726 7584 11790 7588
rect 11806 7644 11870 7648
rect 11806 7588 11810 7644
rect 11810 7588 11866 7644
rect 11866 7588 11870 7644
rect 11806 7584 11870 7588
rect 11886 7644 11950 7648
rect 11886 7588 11890 7644
rect 11890 7588 11946 7644
rect 11946 7588 11950 7644
rect 11886 7584 11950 7588
rect 22340 7644 22404 7648
rect 22340 7588 22344 7644
rect 22344 7588 22400 7644
rect 22400 7588 22404 7644
rect 22340 7584 22404 7588
rect 22420 7644 22484 7648
rect 22420 7588 22424 7644
rect 22424 7588 22480 7644
rect 22480 7588 22484 7644
rect 22420 7584 22484 7588
rect 22500 7644 22564 7648
rect 22500 7588 22504 7644
rect 22504 7588 22560 7644
rect 22560 7588 22564 7644
rect 22500 7584 22564 7588
rect 22580 7644 22644 7648
rect 22580 7588 22584 7644
rect 22584 7588 22640 7644
rect 22640 7588 22644 7644
rect 22580 7584 22644 7588
rect 33034 7644 33098 7648
rect 33034 7588 33038 7644
rect 33038 7588 33094 7644
rect 33094 7588 33098 7644
rect 33034 7584 33098 7588
rect 33114 7644 33178 7648
rect 33114 7588 33118 7644
rect 33118 7588 33174 7644
rect 33174 7588 33178 7644
rect 33114 7584 33178 7588
rect 33194 7644 33258 7648
rect 33194 7588 33198 7644
rect 33198 7588 33254 7644
rect 33254 7588 33258 7644
rect 33194 7584 33258 7588
rect 33274 7644 33338 7648
rect 33274 7588 33278 7644
rect 33278 7588 33334 7644
rect 33334 7588 33338 7644
rect 33274 7584 33338 7588
rect 43728 7644 43792 7648
rect 43728 7588 43732 7644
rect 43732 7588 43788 7644
rect 43788 7588 43792 7644
rect 43728 7584 43792 7588
rect 43808 7644 43872 7648
rect 43808 7588 43812 7644
rect 43812 7588 43868 7644
rect 43868 7588 43872 7644
rect 43808 7584 43872 7588
rect 43888 7644 43952 7648
rect 43888 7588 43892 7644
rect 43892 7588 43948 7644
rect 43948 7588 43952 7644
rect 43888 7584 43952 7588
rect 43968 7644 44032 7648
rect 43968 7588 43972 7644
rect 43972 7588 44028 7644
rect 44028 7588 44032 7644
rect 43968 7584 44032 7588
rect 6299 7100 6363 7104
rect 6299 7044 6303 7100
rect 6303 7044 6359 7100
rect 6359 7044 6363 7100
rect 6299 7040 6363 7044
rect 6379 7100 6443 7104
rect 6379 7044 6383 7100
rect 6383 7044 6439 7100
rect 6439 7044 6443 7100
rect 6379 7040 6443 7044
rect 6459 7100 6523 7104
rect 6459 7044 6463 7100
rect 6463 7044 6519 7100
rect 6519 7044 6523 7100
rect 6459 7040 6523 7044
rect 6539 7100 6603 7104
rect 6539 7044 6543 7100
rect 6543 7044 6599 7100
rect 6599 7044 6603 7100
rect 6539 7040 6603 7044
rect 16993 7100 17057 7104
rect 16993 7044 16997 7100
rect 16997 7044 17053 7100
rect 17053 7044 17057 7100
rect 16993 7040 17057 7044
rect 17073 7100 17137 7104
rect 17073 7044 17077 7100
rect 17077 7044 17133 7100
rect 17133 7044 17137 7100
rect 17073 7040 17137 7044
rect 17153 7100 17217 7104
rect 17153 7044 17157 7100
rect 17157 7044 17213 7100
rect 17213 7044 17217 7100
rect 17153 7040 17217 7044
rect 17233 7100 17297 7104
rect 17233 7044 17237 7100
rect 17237 7044 17293 7100
rect 17293 7044 17297 7100
rect 17233 7040 17297 7044
rect 27687 7100 27751 7104
rect 27687 7044 27691 7100
rect 27691 7044 27747 7100
rect 27747 7044 27751 7100
rect 27687 7040 27751 7044
rect 27767 7100 27831 7104
rect 27767 7044 27771 7100
rect 27771 7044 27827 7100
rect 27827 7044 27831 7100
rect 27767 7040 27831 7044
rect 27847 7100 27911 7104
rect 27847 7044 27851 7100
rect 27851 7044 27907 7100
rect 27907 7044 27911 7100
rect 27847 7040 27911 7044
rect 27927 7100 27991 7104
rect 27927 7044 27931 7100
rect 27931 7044 27987 7100
rect 27987 7044 27991 7100
rect 27927 7040 27991 7044
rect 38381 7100 38445 7104
rect 38381 7044 38385 7100
rect 38385 7044 38441 7100
rect 38441 7044 38445 7100
rect 38381 7040 38445 7044
rect 38461 7100 38525 7104
rect 38461 7044 38465 7100
rect 38465 7044 38521 7100
rect 38521 7044 38525 7100
rect 38461 7040 38525 7044
rect 38541 7100 38605 7104
rect 38541 7044 38545 7100
rect 38545 7044 38601 7100
rect 38601 7044 38605 7100
rect 38541 7040 38605 7044
rect 38621 7100 38685 7104
rect 38621 7044 38625 7100
rect 38625 7044 38681 7100
rect 38681 7044 38685 7100
rect 38621 7040 38685 7044
rect 11646 6556 11710 6560
rect 11646 6500 11650 6556
rect 11650 6500 11706 6556
rect 11706 6500 11710 6556
rect 11646 6496 11710 6500
rect 11726 6556 11790 6560
rect 11726 6500 11730 6556
rect 11730 6500 11786 6556
rect 11786 6500 11790 6556
rect 11726 6496 11790 6500
rect 11806 6556 11870 6560
rect 11806 6500 11810 6556
rect 11810 6500 11866 6556
rect 11866 6500 11870 6556
rect 11806 6496 11870 6500
rect 11886 6556 11950 6560
rect 11886 6500 11890 6556
rect 11890 6500 11946 6556
rect 11946 6500 11950 6556
rect 11886 6496 11950 6500
rect 22340 6556 22404 6560
rect 22340 6500 22344 6556
rect 22344 6500 22400 6556
rect 22400 6500 22404 6556
rect 22340 6496 22404 6500
rect 22420 6556 22484 6560
rect 22420 6500 22424 6556
rect 22424 6500 22480 6556
rect 22480 6500 22484 6556
rect 22420 6496 22484 6500
rect 22500 6556 22564 6560
rect 22500 6500 22504 6556
rect 22504 6500 22560 6556
rect 22560 6500 22564 6556
rect 22500 6496 22564 6500
rect 22580 6556 22644 6560
rect 22580 6500 22584 6556
rect 22584 6500 22640 6556
rect 22640 6500 22644 6556
rect 22580 6496 22644 6500
rect 33034 6556 33098 6560
rect 33034 6500 33038 6556
rect 33038 6500 33094 6556
rect 33094 6500 33098 6556
rect 33034 6496 33098 6500
rect 33114 6556 33178 6560
rect 33114 6500 33118 6556
rect 33118 6500 33174 6556
rect 33174 6500 33178 6556
rect 33114 6496 33178 6500
rect 33194 6556 33258 6560
rect 33194 6500 33198 6556
rect 33198 6500 33254 6556
rect 33254 6500 33258 6556
rect 33194 6496 33258 6500
rect 33274 6556 33338 6560
rect 33274 6500 33278 6556
rect 33278 6500 33334 6556
rect 33334 6500 33338 6556
rect 33274 6496 33338 6500
rect 43728 6556 43792 6560
rect 43728 6500 43732 6556
rect 43732 6500 43788 6556
rect 43788 6500 43792 6556
rect 43728 6496 43792 6500
rect 43808 6556 43872 6560
rect 43808 6500 43812 6556
rect 43812 6500 43868 6556
rect 43868 6500 43872 6556
rect 43808 6496 43872 6500
rect 43888 6556 43952 6560
rect 43888 6500 43892 6556
rect 43892 6500 43948 6556
rect 43948 6500 43952 6556
rect 43888 6496 43952 6500
rect 43968 6556 44032 6560
rect 43968 6500 43972 6556
rect 43972 6500 44028 6556
rect 44028 6500 44032 6556
rect 43968 6496 44032 6500
rect 6299 6012 6363 6016
rect 6299 5956 6303 6012
rect 6303 5956 6359 6012
rect 6359 5956 6363 6012
rect 6299 5952 6363 5956
rect 6379 6012 6443 6016
rect 6379 5956 6383 6012
rect 6383 5956 6439 6012
rect 6439 5956 6443 6012
rect 6379 5952 6443 5956
rect 6459 6012 6523 6016
rect 6459 5956 6463 6012
rect 6463 5956 6519 6012
rect 6519 5956 6523 6012
rect 6459 5952 6523 5956
rect 6539 6012 6603 6016
rect 6539 5956 6543 6012
rect 6543 5956 6599 6012
rect 6599 5956 6603 6012
rect 6539 5952 6603 5956
rect 16993 6012 17057 6016
rect 16993 5956 16997 6012
rect 16997 5956 17053 6012
rect 17053 5956 17057 6012
rect 16993 5952 17057 5956
rect 17073 6012 17137 6016
rect 17073 5956 17077 6012
rect 17077 5956 17133 6012
rect 17133 5956 17137 6012
rect 17073 5952 17137 5956
rect 17153 6012 17217 6016
rect 17153 5956 17157 6012
rect 17157 5956 17213 6012
rect 17213 5956 17217 6012
rect 17153 5952 17217 5956
rect 17233 6012 17297 6016
rect 17233 5956 17237 6012
rect 17237 5956 17293 6012
rect 17293 5956 17297 6012
rect 17233 5952 17297 5956
rect 27687 6012 27751 6016
rect 27687 5956 27691 6012
rect 27691 5956 27747 6012
rect 27747 5956 27751 6012
rect 27687 5952 27751 5956
rect 27767 6012 27831 6016
rect 27767 5956 27771 6012
rect 27771 5956 27827 6012
rect 27827 5956 27831 6012
rect 27767 5952 27831 5956
rect 27847 6012 27911 6016
rect 27847 5956 27851 6012
rect 27851 5956 27907 6012
rect 27907 5956 27911 6012
rect 27847 5952 27911 5956
rect 27927 6012 27991 6016
rect 27927 5956 27931 6012
rect 27931 5956 27987 6012
rect 27987 5956 27991 6012
rect 27927 5952 27991 5956
rect 38381 6012 38445 6016
rect 38381 5956 38385 6012
rect 38385 5956 38441 6012
rect 38441 5956 38445 6012
rect 38381 5952 38445 5956
rect 38461 6012 38525 6016
rect 38461 5956 38465 6012
rect 38465 5956 38521 6012
rect 38521 5956 38525 6012
rect 38461 5952 38525 5956
rect 38541 6012 38605 6016
rect 38541 5956 38545 6012
rect 38545 5956 38601 6012
rect 38601 5956 38605 6012
rect 38541 5952 38605 5956
rect 38621 6012 38685 6016
rect 38621 5956 38625 6012
rect 38625 5956 38681 6012
rect 38681 5956 38685 6012
rect 38621 5952 38685 5956
rect 11646 5468 11710 5472
rect 11646 5412 11650 5468
rect 11650 5412 11706 5468
rect 11706 5412 11710 5468
rect 11646 5408 11710 5412
rect 11726 5468 11790 5472
rect 11726 5412 11730 5468
rect 11730 5412 11786 5468
rect 11786 5412 11790 5468
rect 11726 5408 11790 5412
rect 11806 5468 11870 5472
rect 11806 5412 11810 5468
rect 11810 5412 11866 5468
rect 11866 5412 11870 5468
rect 11806 5408 11870 5412
rect 11886 5468 11950 5472
rect 11886 5412 11890 5468
rect 11890 5412 11946 5468
rect 11946 5412 11950 5468
rect 11886 5408 11950 5412
rect 22340 5468 22404 5472
rect 22340 5412 22344 5468
rect 22344 5412 22400 5468
rect 22400 5412 22404 5468
rect 22340 5408 22404 5412
rect 22420 5468 22484 5472
rect 22420 5412 22424 5468
rect 22424 5412 22480 5468
rect 22480 5412 22484 5468
rect 22420 5408 22484 5412
rect 22500 5468 22564 5472
rect 22500 5412 22504 5468
rect 22504 5412 22560 5468
rect 22560 5412 22564 5468
rect 22500 5408 22564 5412
rect 22580 5468 22644 5472
rect 22580 5412 22584 5468
rect 22584 5412 22640 5468
rect 22640 5412 22644 5468
rect 22580 5408 22644 5412
rect 33034 5468 33098 5472
rect 33034 5412 33038 5468
rect 33038 5412 33094 5468
rect 33094 5412 33098 5468
rect 33034 5408 33098 5412
rect 33114 5468 33178 5472
rect 33114 5412 33118 5468
rect 33118 5412 33174 5468
rect 33174 5412 33178 5468
rect 33114 5408 33178 5412
rect 33194 5468 33258 5472
rect 33194 5412 33198 5468
rect 33198 5412 33254 5468
rect 33254 5412 33258 5468
rect 33194 5408 33258 5412
rect 33274 5468 33338 5472
rect 33274 5412 33278 5468
rect 33278 5412 33334 5468
rect 33334 5412 33338 5468
rect 33274 5408 33338 5412
rect 43728 5468 43792 5472
rect 43728 5412 43732 5468
rect 43732 5412 43788 5468
rect 43788 5412 43792 5468
rect 43728 5408 43792 5412
rect 43808 5468 43872 5472
rect 43808 5412 43812 5468
rect 43812 5412 43868 5468
rect 43868 5412 43872 5468
rect 43808 5408 43872 5412
rect 43888 5468 43952 5472
rect 43888 5412 43892 5468
rect 43892 5412 43948 5468
rect 43948 5412 43952 5468
rect 43888 5408 43952 5412
rect 43968 5468 44032 5472
rect 43968 5412 43972 5468
rect 43972 5412 44028 5468
rect 44028 5412 44032 5468
rect 43968 5408 44032 5412
rect 6299 4924 6363 4928
rect 6299 4868 6303 4924
rect 6303 4868 6359 4924
rect 6359 4868 6363 4924
rect 6299 4864 6363 4868
rect 6379 4924 6443 4928
rect 6379 4868 6383 4924
rect 6383 4868 6439 4924
rect 6439 4868 6443 4924
rect 6379 4864 6443 4868
rect 6459 4924 6523 4928
rect 6459 4868 6463 4924
rect 6463 4868 6519 4924
rect 6519 4868 6523 4924
rect 6459 4864 6523 4868
rect 6539 4924 6603 4928
rect 6539 4868 6543 4924
rect 6543 4868 6599 4924
rect 6599 4868 6603 4924
rect 6539 4864 6603 4868
rect 16993 4924 17057 4928
rect 16993 4868 16997 4924
rect 16997 4868 17053 4924
rect 17053 4868 17057 4924
rect 16993 4864 17057 4868
rect 17073 4924 17137 4928
rect 17073 4868 17077 4924
rect 17077 4868 17133 4924
rect 17133 4868 17137 4924
rect 17073 4864 17137 4868
rect 17153 4924 17217 4928
rect 17153 4868 17157 4924
rect 17157 4868 17213 4924
rect 17213 4868 17217 4924
rect 17153 4864 17217 4868
rect 17233 4924 17297 4928
rect 17233 4868 17237 4924
rect 17237 4868 17293 4924
rect 17293 4868 17297 4924
rect 17233 4864 17297 4868
rect 27687 4924 27751 4928
rect 27687 4868 27691 4924
rect 27691 4868 27747 4924
rect 27747 4868 27751 4924
rect 27687 4864 27751 4868
rect 27767 4924 27831 4928
rect 27767 4868 27771 4924
rect 27771 4868 27827 4924
rect 27827 4868 27831 4924
rect 27767 4864 27831 4868
rect 27847 4924 27911 4928
rect 27847 4868 27851 4924
rect 27851 4868 27907 4924
rect 27907 4868 27911 4924
rect 27847 4864 27911 4868
rect 27927 4924 27991 4928
rect 27927 4868 27931 4924
rect 27931 4868 27987 4924
rect 27987 4868 27991 4924
rect 27927 4864 27991 4868
rect 38381 4924 38445 4928
rect 38381 4868 38385 4924
rect 38385 4868 38441 4924
rect 38441 4868 38445 4924
rect 38381 4864 38445 4868
rect 38461 4924 38525 4928
rect 38461 4868 38465 4924
rect 38465 4868 38521 4924
rect 38521 4868 38525 4924
rect 38461 4864 38525 4868
rect 38541 4924 38605 4928
rect 38541 4868 38545 4924
rect 38545 4868 38601 4924
rect 38601 4868 38605 4924
rect 38541 4864 38605 4868
rect 38621 4924 38685 4928
rect 38621 4868 38625 4924
rect 38625 4868 38681 4924
rect 38681 4868 38685 4924
rect 38621 4864 38685 4868
rect 11646 4380 11710 4384
rect 11646 4324 11650 4380
rect 11650 4324 11706 4380
rect 11706 4324 11710 4380
rect 11646 4320 11710 4324
rect 11726 4380 11790 4384
rect 11726 4324 11730 4380
rect 11730 4324 11786 4380
rect 11786 4324 11790 4380
rect 11726 4320 11790 4324
rect 11806 4380 11870 4384
rect 11806 4324 11810 4380
rect 11810 4324 11866 4380
rect 11866 4324 11870 4380
rect 11806 4320 11870 4324
rect 11886 4380 11950 4384
rect 11886 4324 11890 4380
rect 11890 4324 11946 4380
rect 11946 4324 11950 4380
rect 11886 4320 11950 4324
rect 22340 4380 22404 4384
rect 22340 4324 22344 4380
rect 22344 4324 22400 4380
rect 22400 4324 22404 4380
rect 22340 4320 22404 4324
rect 22420 4380 22484 4384
rect 22420 4324 22424 4380
rect 22424 4324 22480 4380
rect 22480 4324 22484 4380
rect 22420 4320 22484 4324
rect 22500 4380 22564 4384
rect 22500 4324 22504 4380
rect 22504 4324 22560 4380
rect 22560 4324 22564 4380
rect 22500 4320 22564 4324
rect 22580 4380 22644 4384
rect 22580 4324 22584 4380
rect 22584 4324 22640 4380
rect 22640 4324 22644 4380
rect 22580 4320 22644 4324
rect 33034 4380 33098 4384
rect 33034 4324 33038 4380
rect 33038 4324 33094 4380
rect 33094 4324 33098 4380
rect 33034 4320 33098 4324
rect 33114 4380 33178 4384
rect 33114 4324 33118 4380
rect 33118 4324 33174 4380
rect 33174 4324 33178 4380
rect 33114 4320 33178 4324
rect 33194 4380 33258 4384
rect 33194 4324 33198 4380
rect 33198 4324 33254 4380
rect 33254 4324 33258 4380
rect 33194 4320 33258 4324
rect 33274 4380 33338 4384
rect 33274 4324 33278 4380
rect 33278 4324 33334 4380
rect 33334 4324 33338 4380
rect 33274 4320 33338 4324
rect 43728 4380 43792 4384
rect 43728 4324 43732 4380
rect 43732 4324 43788 4380
rect 43788 4324 43792 4380
rect 43728 4320 43792 4324
rect 43808 4380 43872 4384
rect 43808 4324 43812 4380
rect 43812 4324 43868 4380
rect 43868 4324 43872 4380
rect 43808 4320 43872 4324
rect 43888 4380 43952 4384
rect 43888 4324 43892 4380
rect 43892 4324 43948 4380
rect 43948 4324 43952 4380
rect 43888 4320 43952 4324
rect 43968 4380 44032 4384
rect 43968 4324 43972 4380
rect 43972 4324 44028 4380
rect 44028 4324 44032 4380
rect 43968 4320 44032 4324
rect 6299 3836 6363 3840
rect 6299 3780 6303 3836
rect 6303 3780 6359 3836
rect 6359 3780 6363 3836
rect 6299 3776 6363 3780
rect 6379 3836 6443 3840
rect 6379 3780 6383 3836
rect 6383 3780 6439 3836
rect 6439 3780 6443 3836
rect 6379 3776 6443 3780
rect 6459 3836 6523 3840
rect 6459 3780 6463 3836
rect 6463 3780 6519 3836
rect 6519 3780 6523 3836
rect 6459 3776 6523 3780
rect 6539 3836 6603 3840
rect 6539 3780 6543 3836
rect 6543 3780 6599 3836
rect 6599 3780 6603 3836
rect 6539 3776 6603 3780
rect 16993 3836 17057 3840
rect 16993 3780 16997 3836
rect 16997 3780 17053 3836
rect 17053 3780 17057 3836
rect 16993 3776 17057 3780
rect 17073 3836 17137 3840
rect 17073 3780 17077 3836
rect 17077 3780 17133 3836
rect 17133 3780 17137 3836
rect 17073 3776 17137 3780
rect 17153 3836 17217 3840
rect 17153 3780 17157 3836
rect 17157 3780 17213 3836
rect 17213 3780 17217 3836
rect 17153 3776 17217 3780
rect 17233 3836 17297 3840
rect 17233 3780 17237 3836
rect 17237 3780 17293 3836
rect 17293 3780 17297 3836
rect 17233 3776 17297 3780
rect 27687 3836 27751 3840
rect 27687 3780 27691 3836
rect 27691 3780 27747 3836
rect 27747 3780 27751 3836
rect 27687 3776 27751 3780
rect 27767 3836 27831 3840
rect 27767 3780 27771 3836
rect 27771 3780 27827 3836
rect 27827 3780 27831 3836
rect 27767 3776 27831 3780
rect 27847 3836 27911 3840
rect 27847 3780 27851 3836
rect 27851 3780 27907 3836
rect 27907 3780 27911 3836
rect 27847 3776 27911 3780
rect 27927 3836 27991 3840
rect 27927 3780 27931 3836
rect 27931 3780 27987 3836
rect 27987 3780 27991 3836
rect 27927 3776 27991 3780
rect 38381 3836 38445 3840
rect 38381 3780 38385 3836
rect 38385 3780 38441 3836
rect 38441 3780 38445 3836
rect 38381 3776 38445 3780
rect 38461 3836 38525 3840
rect 38461 3780 38465 3836
rect 38465 3780 38521 3836
rect 38521 3780 38525 3836
rect 38461 3776 38525 3780
rect 38541 3836 38605 3840
rect 38541 3780 38545 3836
rect 38545 3780 38601 3836
rect 38601 3780 38605 3836
rect 38541 3776 38605 3780
rect 38621 3836 38685 3840
rect 38621 3780 38625 3836
rect 38625 3780 38681 3836
rect 38681 3780 38685 3836
rect 38621 3776 38685 3780
rect 11646 3292 11710 3296
rect 11646 3236 11650 3292
rect 11650 3236 11706 3292
rect 11706 3236 11710 3292
rect 11646 3232 11710 3236
rect 11726 3292 11790 3296
rect 11726 3236 11730 3292
rect 11730 3236 11786 3292
rect 11786 3236 11790 3292
rect 11726 3232 11790 3236
rect 11806 3292 11870 3296
rect 11806 3236 11810 3292
rect 11810 3236 11866 3292
rect 11866 3236 11870 3292
rect 11806 3232 11870 3236
rect 11886 3292 11950 3296
rect 11886 3236 11890 3292
rect 11890 3236 11946 3292
rect 11946 3236 11950 3292
rect 11886 3232 11950 3236
rect 22340 3292 22404 3296
rect 22340 3236 22344 3292
rect 22344 3236 22400 3292
rect 22400 3236 22404 3292
rect 22340 3232 22404 3236
rect 22420 3292 22484 3296
rect 22420 3236 22424 3292
rect 22424 3236 22480 3292
rect 22480 3236 22484 3292
rect 22420 3232 22484 3236
rect 22500 3292 22564 3296
rect 22500 3236 22504 3292
rect 22504 3236 22560 3292
rect 22560 3236 22564 3292
rect 22500 3232 22564 3236
rect 22580 3292 22644 3296
rect 22580 3236 22584 3292
rect 22584 3236 22640 3292
rect 22640 3236 22644 3292
rect 22580 3232 22644 3236
rect 33034 3292 33098 3296
rect 33034 3236 33038 3292
rect 33038 3236 33094 3292
rect 33094 3236 33098 3292
rect 33034 3232 33098 3236
rect 33114 3292 33178 3296
rect 33114 3236 33118 3292
rect 33118 3236 33174 3292
rect 33174 3236 33178 3292
rect 33114 3232 33178 3236
rect 33194 3292 33258 3296
rect 33194 3236 33198 3292
rect 33198 3236 33254 3292
rect 33254 3236 33258 3292
rect 33194 3232 33258 3236
rect 33274 3292 33338 3296
rect 33274 3236 33278 3292
rect 33278 3236 33334 3292
rect 33334 3236 33338 3292
rect 33274 3232 33338 3236
rect 43728 3292 43792 3296
rect 43728 3236 43732 3292
rect 43732 3236 43788 3292
rect 43788 3236 43792 3292
rect 43728 3232 43792 3236
rect 43808 3292 43872 3296
rect 43808 3236 43812 3292
rect 43812 3236 43868 3292
rect 43868 3236 43872 3292
rect 43808 3232 43872 3236
rect 43888 3292 43952 3296
rect 43888 3236 43892 3292
rect 43892 3236 43948 3292
rect 43948 3236 43952 3292
rect 43888 3232 43952 3236
rect 43968 3292 44032 3296
rect 43968 3236 43972 3292
rect 43972 3236 44028 3292
rect 44028 3236 44032 3292
rect 43968 3232 44032 3236
rect 6299 2748 6363 2752
rect 6299 2692 6303 2748
rect 6303 2692 6359 2748
rect 6359 2692 6363 2748
rect 6299 2688 6363 2692
rect 6379 2748 6443 2752
rect 6379 2692 6383 2748
rect 6383 2692 6439 2748
rect 6439 2692 6443 2748
rect 6379 2688 6443 2692
rect 6459 2748 6523 2752
rect 6459 2692 6463 2748
rect 6463 2692 6519 2748
rect 6519 2692 6523 2748
rect 6459 2688 6523 2692
rect 6539 2748 6603 2752
rect 6539 2692 6543 2748
rect 6543 2692 6599 2748
rect 6599 2692 6603 2748
rect 6539 2688 6603 2692
rect 16993 2748 17057 2752
rect 16993 2692 16997 2748
rect 16997 2692 17053 2748
rect 17053 2692 17057 2748
rect 16993 2688 17057 2692
rect 17073 2748 17137 2752
rect 17073 2692 17077 2748
rect 17077 2692 17133 2748
rect 17133 2692 17137 2748
rect 17073 2688 17137 2692
rect 17153 2748 17217 2752
rect 17153 2692 17157 2748
rect 17157 2692 17213 2748
rect 17213 2692 17217 2748
rect 17153 2688 17217 2692
rect 17233 2748 17297 2752
rect 17233 2692 17237 2748
rect 17237 2692 17293 2748
rect 17293 2692 17297 2748
rect 17233 2688 17297 2692
rect 27687 2748 27751 2752
rect 27687 2692 27691 2748
rect 27691 2692 27747 2748
rect 27747 2692 27751 2748
rect 27687 2688 27751 2692
rect 27767 2748 27831 2752
rect 27767 2692 27771 2748
rect 27771 2692 27827 2748
rect 27827 2692 27831 2748
rect 27767 2688 27831 2692
rect 27847 2748 27911 2752
rect 27847 2692 27851 2748
rect 27851 2692 27907 2748
rect 27907 2692 27911 2748
rect 27847 2688 27911 2692
rect 27927 2748 27991 2752
rect 27927 2692 27931 2748
rect 27931 2692 27987 2748
rect 27987 2692 27991 2748
rect 27927 2688 27991 2692
rect 38381 2748 38445 2752
rect 38381 2692 38385 2748
rect 38385 2692 38441 2748
rect 38441 2692 38445 2748
rect 38381 2688 38445 2692
rect 38461 2748 38525 2752
rect 38461 2692 38465 2748
rect 38465 2692 38521 2748
rect 38521 2692 38525 2748
rect 38461 2688 38525 2692
rect 38541 2748 38605 2752
rect 38541 2692 38545 2748
rect 38545 2692 38601 2748
rect 38601 2692 38605 2748
rect 38541 2688 38605 2692
rect 38621 2748 38685 2752
rect 38621 2692 38625 2748
rect 38625 2692 38681 2748
rect 38681 2692 38685 2748
rect 38621 2688 38685 2692
rect 11646 2204 11710 2208
rect 11646 2148 11650 2204
rect 11650 2148 11706 2204
rect 11706 2148 11710 2204
rect 11646 2144 11710 2148
rect 11726 2204 11790 2208
rect 11726 2148 11730 2204
rect 11730 2148 11786 2204
rect 11786 2148 11790 2204
rect 11726 2144 11790 2148
rect 11806 2204 11870 2208
rect 11806 2148 11810 2204
rect 11810 2148 11866 2204
rect 11866 2148 11870 2204
rect 11806 2144 11870 2148
rect 11886 2204 11950 2208
rect 11886 2148 11890 2204
rect 11890 2148 11946 2204
rect 11946 2148 11950 2204
rect 11886 2144 11950 2148
rect 22340 2204 22404 2208
rect 22340 2148 22344 2204
rect 22344 2148 22400 2204
rect 22400 2148 22404 2204
rect 22340 2144 22404 2148
rect 22420 2204 22484 2208
rect 22420 2148 22424 2204
rect 22424 2148 22480 2204
rect 22480 2148 22484 2204
rect 22420 2144 22484 2148
rect 22500 2204 22564 2208
rect 22500 2148 22504 2204
rect 22504 2148 22560 2204
rect 22560 2148 22564 2204
rect 22500 2144 22564 2148
rect 22580 2204 22644 2208
rect 22580 2148 22584 2204
rect 22584 2148 22640 2204
rect 22640 2148 22644 2204
rect 22580 2144 22644 2148
rect 33034 2204 33098 2208
rect 33034 2148 33038 2204
rect 33038 2148 33094 2204
rect 33094 2148 33098 2204
rect 33034 2144 33098 2148
rect 33114 2204 33178 2208
rect 33114 2148 33118 2204
rect 33118 2148 33174 2204
rect 33174 2148 33178 2204
rect 33114 2144 33178 2148
rect 33194 2204 33258 2208
rect 33194 2148 33198 2204
rect 33198 2148 33254 2204
rect 33254 2148 33258 2204
rect 33194 2144 33258 2148
rect 33274 2204 33338 2208
rect 33274 2148 33278 2204
rect 33278 2148 33334 2204
rect 33334 2148 33338 2204
rect 33274 2144 33338 2148
rect 43728 2204 43792 2208
rect 43728 2148 43732 2204
rect 43732 2148 43788 2204
rect 43788 2148 43792 2204
rect 43728 2144 43792 2148
rect 43808 2204 43872 2208
rect 43808 2148 43812 2204
rect 43812 2148 43868 2204
rect 43868 2148 43872 2204
rect 43808 2144 43872 2148
rect 43888 2204 43952 2208
rect 43888 2148 43892 2204
rect 43892 2148 43948 2204
rect 43948 2148 43952 2204
rect 43888 2144 43952 2148
rect 43968 2204 44032 2208
rect 43968 2148 43972 2204
rect 43972 2148 44028 2204
rect 44028 2148 44032 2204
rect 43968 2144 44032 2148
<< metal4 >>
rect 6291 7104 6611 7664
rect 6291 7040 6299 7104
rect 6363 7040 6379 7104
rect 6443 7040 6459 7104
rect 6523 7040 6539 7104
rect 6603 7040 6611 7104
rect 6291 6016 6611 7040
rect 6291 5952 6299 6016
rect 6363 5952 6379 6016
rect 6443 5952 6459 6016
rect 6523 5952 6539 6016
rect 6603 5952 6611 6016
rect 6291 4928 6611 5952
rect 6291 4864 6299 4928
rect 6363 4864 6379 4928
rect 6443 4864 6459 4928
rect 6523 4864 6539 4928
rect 6603 4864 6611 4928
rect 6291 3840 6611 4864
rect 6291 3776 6299 3840
rect 6363 3776 6379 3840
rect 6443 3776 6459 3840
rect 6523 3776 6539 3840
rect 6603 3776 6611 3840
rect 6291 2752 6611 3776
rect 6291 2688 6299 2752
rect 6363 2688 6379 2752
rect 6443 2688 6459 2752
rect 6523 2688 6539 2752
rect 6603 2688 6611 2752
rect 6291 2128 6611 2688
rect 11638 7648 11958 7664
rect 11638 7584 11646 7648
rect 11710 7584 11726 7648
rect 11790 7584 11806 7648
rect 11870 7584 11886 7648
rect 11950 7584 11958 7648
rect 11638 6560 11958 7584
rect 11638 6496 11646 6560
rect 11710 6496 11726 6560
rect 11790 6496 11806 6560
rect 11870 6496 11886 6560
rect 11950 6496 11958 6560
rect 11638 5472 11958 6496
rect 11638 5408 11646 5472
rect 11710 5408 11726 5472
rect 11790 5408 11806 5472
rect 11870 5408 11886 5472
rect 11950 5408 11958 5472
rect 11638 4384 11958 5408
rect 11638 4320 11646 4384
rect 11710 4320 11726 4384
rect 11790 4320 11806 4384
rect 11870 4320 11886 4384
rect 11950 4320 11958 4384
rect 11638 3296 11958 4320
rect 11638 3232 11646 3296
rect 11710 3232 11726 3296
rect 11790 3232 11806 3296
rect 11870 3232 11886 3296
rect 11950 3232 11958 3296
rect 11638 2208 11958 3232
rect 11638 2144 11646 2208
rect 11710 2144 11726 2208
rect 11790 2144 11806 2208
rect 11870 2144 11886 2208
rect 11950 2144 11958 2208
rect 11638 2128 11958 2144
rect 16985 7104 17305 7664
rect 16985 7040 16993 7104
rect 17057 7040 17073 7104
rect 17137 7040 17153 7104
rect 17217 7040 17233 7104
rect 17297 7040 17305 7104
rect 16985 6016 17305 7040
rect 16985 5952 16993 6016
rect 17057 5952 17073 6016
rect 17137 5952 17153 6016
rect 17217 5952 17233 6016
rect 17297 5952 17305 6016
rect 16985 4928 17305 5952
rect 16985 4864 16993 4928
rect 17057 4864 17073 4928
rect 17137 4864 17153 4928
rect 17217 4864 17233 4928
rect 17297 4864 17305 4928
rect 16985 3840 17305 4864
rect 16985 3776 16993 3840
rect 17057 3776 17073 3840
rect 17137 3776 17153 3840
rect 17217 3776 17233 3840
rect 17297 3776 17305 3840
rect 16985 2752 17305 3776
rect 16985 2688 16993 2752
rect 17057 2688 17073 2752
rect 17137 2688 17153 2752
rect 17217 2688 17233 2752
rect 17297 2688 17305 2752
rect 16985 2128 17305 2688
rect 22332 7648 22652 7664
rect 22332 7584 22340 7648
rect 22404 7584 22420 7648
rect 22484 7584 22500 7648
rect 22564 7584 22580 7648
rect 22644 7584 22652 7648
rect 22332 6560 22652 7584
rect 22332 6496 22340 6560
rect 22404 6496 22420 6560
rect 22484 6496 22500 6560
rect 22564 6496 22580 6560
rect 22644 6496 22652 6560
rect 22332 5472 22652 6496
rect 22332 5408 22340 5472
rect 22404 5408 22420 5472
rect 22484 5408 22500 5472
rect 22564 5408 22580 5472
rect 22644 5408 22652 5472
rect 22332 4384 22652 5408
rect 22332 4320 22340 4384
rect 22404 4320 22420 4384
rect 22484 4320 22500 4384
rect 22564 4320 22580 4384
rect 22644 4320 22652 4384
rect 22332 3296 22652 4320
rect 22332 3232 22340 3296
rect 22404 3232 22420 3296
rect 22484 3232 22500 3296
rect 22564 3232 22580 3296
rect 22644 3232 22652 3296
rect 22332 2208 22652 3232
rect 22332 2144 22340 2208
rect 22404 2144 22420 2208
rect 22484 2144 22500 2208
rect 22564 2144 22580 2208
rect 22644 2144 22652 2208
rect 22332 2128 22652 2144
rect 27679 7104 27999 7664
rect 27679 7040 27687 7104
rect 27751 7040 27767 7104
rect 27831 7040 27847 7104
rect 27911 7040 27927 7104
rect 27991 7040 27999 7104
rect 27679 6016 27999 7040
rect 27679 5952 27687 6016
rect 27751 5952 27767 6016
rect 27831 5952 27847 6016
rect 27911 5952 27927 6016
rect 27991 5952 27999 6016
rect 27679 4928 27999 5952
rect 27679 4864 27687 4928
rect 27751 4864 27767 4928
rect 27831 4864 27847 4928
rect 27911 4864 27927 4928
rect 27991 4864 27999 4928
rect 27679 3840 27999 4864
rect 27679 3776 27687 3840
rect 27751 3776 27767 3840
rect 27831 3776 27847 3840
rect 27911 3776 27927 3840
rect 27991 3776 27999 3840
rect 27679 2752 27999 3776
rect 27679 2688 27687 2752
rect 27751 2688 27767 2752
rect 27831 2688 27847 2752
rect 27911 2688 27927 2752
rect 27991 2688 27999 2752
rect 27679 2128 27999 2688
rect 33026 7648 33346 7664
rect 33026 7584 33034 7648
rect 33098 7584 33114 7648
rect 33178 7584 33194 7648
rect 33258 7584 33274 7648
rect 33338 7584 33346 7648
rect 33026 6560 33346 7584
rect 33026 6496 33034 6560
rect 33098 6496 33114 6560
rect 33178 6496 33194 6560
rect 33258 6496 33274 6560
rect 33338 6496 33346 6560
rect 33026 5472 33346 6496
rect 33026 5408 33034 5472
rect 33098 5408 33114 5472
rect 33178 5408 33194 5472
rect 33258 5408 33274 5472
rect 33338 5408 33346 5472
rect 33026 4384 33346 5408
rect 33026 4320 33034 4384
rect 33098 4320 33114 4384
rect 33178 4320 33194 4384
rect 33258 4320 33274 4384
rect 33338 4320 33346 4384
rect 33026 3296 33346 4320
rect 33026 3232 33034 3296
rect 33098 3232 33114 3296
rect 33178 3232 33194 3296
rect 33258 3232 33274 3296
rect 33338 3232 33346 3296
rect 33026 2208 33346 3232
rect 33026 2144 33034 2208
rect 33098 2144 33114 2208
rect 33178 2144 33194 2208
rect 33258 2144 33274 2208
rect 33338 2144 33346 2208
rect 33026 2128 33346 2144
rect 38373 7104 38693 7664
rect 38373 7040 38381 7104
rect 38445 7040 38461 7104
rect 38525 7040 38541 7104
rect 38605 7040 38621 7104
rect 38685 7040 38693 7104
rect 38373 6016 38693 7040
rect 38373 5952 38381 6016
rect 38445 5952 38461 6016
rect 38525 5952 38541 6016
rect 38605 5952 38621 6016
rect 38685 5952 38693 6016
rect 38373 4928 38693 5952
rect 38373 4864 38381 4928
rect 38445 4864 38461 4928
rect 38525 4864 38541 4928
rect 38605 4864 38621 4928
rect 38685 4864 38693 4928
rect 38373 3840 38693 4864
rect 38373 3776 38381 3840
rect 38445 3776 38461 3840
rect 38525 3776 38541 3840
rect 38605 3776 38621 3840
rect 38685 3776 38693 3840
rect 38373 2752 38693 3776
rect 38373 2688 38381 2752
rect 38445 2688 38461 2752
rect 38525 2688 38541 2752
rect 38605 2688 38621 2752
rect 38685 2688 38693 2752
rect 38373 2128 38693 2688
rect 43720 7648 44040 7664
rect 43720 7584 43728 7648
rect 43792 7584 43808 7648
rect 43872 7584 43888 7648
rect 43952 7584 43968 7648
rect 44032 7584 44040 7648
rect 43720 6560 44040 7584
rect 43720 6496 43728 6560
rect 43792 6496 43808 6560
rect 43872 6496 43888 6560
rect 43952 6496 43968 6560
rect 44032 6496 44040 6560
rect 43720 5472 44040 6496
rect 43720 5408 43728 5472
rect 43792 5408 43808 5472
rect 43872 5408 43888 5472
rect 43952 5408 43968 5472
rect 44032 5408 44040 5472
rect 43720 4384 44040 5408
rect 43720 4320 43728 4384
rect 43792 4320 43808 4384
rect 43872 4320 43888 4384
rect 43952 4320 43968 4384
rect 44032 4320 44040 4384
rect 43720 3296 44040 4320
rect 43720 3232 43728 3296
rect 43792 3232 43808 3296
rect 43872 3232 43888 3296
rect 43952 3232 43968 3296
rect 44032 3232 44040 3296
rect 43720 2208 44040 3232
rect 43720 2144 43728 2208
rect 43792 2144 43808 2208
rect 43872 2144 43888 2208
rect 43952 2144 43968 2208
rect 44032 2144 44040 2208
rect 43720 2128 44040 2144
use sky130_fd_sc_hd__clkbuf_2  _01_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _02_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _03_
timestamp 1688980957
transform 1 0 18676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _04_
timestamp 1688980957
transform 1 0 20792 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _05_
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _06_
timestamp 1688980957
transform 1 0 25024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1688980957
transform 1 0 37536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _11_
timestamp 1688980957
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1688980957
transform 1 0 41216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1688980957
transform 1 0 40940 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1688980957
transform 1 0 7820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1688980957
transform 1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1688980957
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _20_
timestamp 1688980957
transform 1 0 24932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _21_
timestamp 1688980957
transform 1 0 24380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _22_
timestamp 1688980957
transform 1 0 23184 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _23_
timestamp 1688980957
transform 1 0 23000 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _24_
timestamp 1688980957
transform 1 0 22356 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _25_
timestamp 1688980957
transform 1 0 22724 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _26_
timestamp 1688980957
transform 1 0 22264 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _27_
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _28_
timestamp 1688980957
transform 1 0 21252 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _29_
timestamp 1688980957
transform 1 0 20976 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _30_
timestamp 1688980957
transform 1 0 21528 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _31_
timestamp 1688980957
transform 1 0 20424 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _32_
timestamp 1688980957
transform 1 0 20424 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1688980957
transform 1 0 8924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1688980957
transform 1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _36_
timestamp 1688980957
transform 1 0 29992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _37_
timestamp 1688980957
transform 1 0 29624 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _38_
timestamp 1688980957
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _39_
timestamp 1688980957
transform 1 0 28704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _40_
timestamp 1688980957
transform 1 0 28244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _41_
timestamp 1688980957
transform 1 0 27876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _42_
timestamp 1688980957
transform 1 0 27508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _43_
timestamp 1688980957
transform 1 0 27140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _44_
timestamp 1688980957
transform 1 0 26772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _45_
timestamp 1688980957
transform 1 0 26496 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _46_
timestamp 1688980957
transform 1 0 26220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _47_
timestamp 1688980957
transform 1 0 25760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _48_
timestamp 1688980957
transform 1 0 25392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _49_
timestamp 1688980957
transform 1 0 25116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _50_
timestamp 1688980957
transform 1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1688980957
transform 1 0 13800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1688980957
transform 1 0 14628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1688980957
transform 1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1688980957
transform 1 0 15272 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1688980957
transform 1 0 15640 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1688980957
transform 1 0 16100 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1688980957
transform 1 0 17572 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1688980957
transform 1 0 17296 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1688980957
transform 1 0 18032 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1688980957
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1688980957
transform 1 0 18584 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1688980957
transform 1 0 18952 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _67_
timestamp 1688980957
transform 1 0 30268 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1688980957
transform 1 0 32384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1688980957
transform 1 0 33672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1688980957
transform 1 0 34040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1688980957
transform 1 0 34960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _73_
timestamp 1688980957
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform -1 0 9568 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform -1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform -1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_13 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_33
timestamp 1688980957
transform 1 0 4140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_45 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_67 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_71 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_93
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_98
timestamp 1688980957
transform 1 0 10120 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 1688980957
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_117
timestamp 1688980957
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_133 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_144
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_150
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_162
timestamp 1688980957
transform 1 0 16008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_172
timestamp 1688980957
transform 1 0 16928 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_184
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_190
timestamp 1688980957
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_213
timestamp 1688980957
transform 1 0 20700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_236
timestamp 1688980957
transform 1 0 22816 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_248
timestamp 1688980957
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_259
timestamp 1688980957
transform 1 0 24932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_271
timestamp 1688980957
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_284
timestamp 1688980957
transform 1 0 27232 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_296
timestamp 1688980957
transform 1 0 28336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_328
timestamp 1688980957
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_345
timestamp 1688980957
transform 1 0 32844 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_351
timestamp 1688980957
transform 1 0 33396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_368
timestamp 1688980957
transform 1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_374
timestamp 1688980957
transform 1 0 35512 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_386
timestamp 1688980957
transform 1 0 36616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_391
timestamp 1688980957
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_397
timestamp 1688980957
transform 1 0 37628 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_402
timestamp 1688980957
transform 1 0 38088 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_414
timestamp 1688980957
transform 1 0 39192 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_439
timestamp 1688980957
transform 1 0 41492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_443
timestamp 1688980957
transform 1 0 41860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_447
timestamp 1688980957
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_457
timestamp 1688980957
transform 1 0 43148 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_189
timestamp 1688980957
transform 1 0 18492 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_194
timestamp 1688980957
transform 1 0 18952 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_206
timestamp 1688980957
transform 1 0 20056 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_218
timestamp 1688980957
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_240
timestamp 1688980957
transform 1 0 23184 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_252
timestamp 1688980957
transform 1 0 24288 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_263
timestamp 1688980957
transform 1 0 25300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_275
timestamp 1688980957
transform 1 0 26404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_461
timestamp 1688980957
transform 1 0 43516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_461
timestamp 1688980957
transform 1 0 43516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_213
timestamp 1688980957
transform 1 0 20700 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_130
timestamp 1688980957
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1688980957
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_461
timestamp 1688980957
transform 1 0 43516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_47
timestamp 1688980957
transform 1 0 5428 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_76
timestamp 1688980957
transform 1 0 8096 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_104
timestamp 1688980957
transform 1 0 10672 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 1688980957
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_122
timestamp 1688980957
transform 1 0 12328 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_134
timestamp 1688980957
transform 1 0 13432 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_150
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_157
timestamp 1688980957
transform 1 0 15548 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1688980957
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_172
timestamp 1688980957
transform 1 0 16928 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_182
timestamp 1688980957
transform 1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_197
timestamp 1688980957
transform 1 0 19228 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_209
timestamp 1688980957
transform 1 0 20332 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_213
timestamp 1688980957
transform 1 0 20700 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_221
timestamp 1688980957
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_228
timestamp 1688980957
transform 1 0 22080 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_233
timestamp 1688980957
transform 1 0 22540 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_238
timestamp 1688980957
transform 1 0 23000 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_250
timestamp 1688980957
transform 1 0 24104 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_262
timestamp 1688980957
transform 1 0 25208 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_271
timestamp 1688980957
transform 1 0 26036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_357
timestamp 1688980957
transform 1 0 33948 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_399
timestamp 1688980957
transform 1 0 37812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_411
timestamp 1688980957
transform 1 0 38916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_423
timestamp 1688980957
transform 1 0 40020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_435
timestamp 1688980957
transform 1 0 41124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_94
timestamp 1688980957
transform 1 0 9752 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_192
timestamp 1688980957
transform 1 0 18768 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_225
timestamp 1688980957
transform 1 0 21804 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_237
timestamp 1688980957
transform 1 0 22908 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_241
timestamp 1688980957
transform 1 0 23276 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_249
timestamp 1688980957
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_257
timestamp 1688980957
transform 1 0 24748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_267
timestamp 1688980957
transform 1 0 25668 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_282
timestamp 1688980957
transform 1 0 27048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_286
timestamp 1688980957
transform 1 0 27416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_290
timestamp 1688980957
transform 1 0 27784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_294
timestamp 1688980957
transform 1 0 28152 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_298
timestamp 1688980957
transform 1 0 28520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_303
timestamp 1688980957
transform 1 0 28980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_313
timestamp 1688980957
transform 1 0 29900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_320
timestamp 1688980957
transform 1 0 30544 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_326
timestamp 1688980957
transform 1 0 31096 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_330
timestamp 1688980957
transform 1 0 31464 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_338
timestamp 1688980957
transform 1 0 32200 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_343
timestamp 1688980957
transform 1 0 32660 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_347
timestamp 1688980957
transform 1 0 33028 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_371
timestamp 1688980957
transform 1 0 35236 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_461
timestamp 1688980957
transform 1 0 43516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_29
timestamp 1688980957
transform 1 0 3772 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_37
timestamp 1688980957
transform 1 0 4508 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_88
timestamp 1688980957
transform 1 0 9200 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_92
timestamp 1688980957
transform 1 0 9568 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_117
timestamp 1688980957
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_121
timestamp 1688980957
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_197
timestamp 1688980957
transform 1 0 19228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_210
timestamp 1688980957
transform 1 0 20424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_355
timestamp 1688980957
transform 1 0 33764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_363
timestamp 1688980957
transform 1 0 34500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_439
timestamp 1688980957
transform 1 0 41492 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 24656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 31004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 33120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 35236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 37352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 41584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 16192 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 19320 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 19596 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 19872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 20148 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 20700 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 22080 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 22632 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 23736 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 24656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 25208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 25484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 25760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 28612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 29532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 29808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 30084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 26036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform 1 0 26312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 27784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 28336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 30360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1688980957
transform 1 0 32936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1688980957
transform 1 0 33488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform 1 0 33120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1688980957
transform 1 0 33396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1688980957
transform 1 0 34224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1688980957
transform 1 0 30636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1688980957
transform 1 0 30912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1688980957
transform 1 0 31188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1688980957
transform 1 0 31464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1688980957
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1688980957
transform 1 0 31188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1688980957
transform 1 0 32384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1688980957
transform 1 0 32660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 37536 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 38088 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 38916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 38640 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 39192 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 39836 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 40388 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 40388 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 35236 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 35788 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 35328 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 36340 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 35880 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 36432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 36984 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 37812 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 4968 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 4600 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output96
timestamp 1688980957
transform 1 0 5520 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 5152 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 6072 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 6624 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output101
timestamp 1688980957
transform 1 0 7176 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 6624 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 7728 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 7176 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 8464 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 8280 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 9016 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 9568 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 9200 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 10120 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform -1 0 10304 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 12880 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 14076 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 13432 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform 1 0 14352 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform 1 0 14904 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 10672 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform -1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 11224 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform -1 0 11408 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 11776 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 12328 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform 1 0 11776 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 12880 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 12328 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 14352 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 17480 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 18216 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output133
timestamp 1688980957
transform 1 0 18032 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output134
timestamp 1688980957
transform 1 0 18584 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 19872 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 19320 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 15456 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform 1 0 14904 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform 1 0 16008 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 15456 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 16560 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 17112 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 16928 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 17664 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform 1 0 33948 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 43884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 43884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 43884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 43884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 43884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 43884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 43884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  S_term_single_147 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
<< labels >>
flabel metal2 s 34150 9840 34206 10000 0 FreeSans 224 90 0 0 Co
port 0 nsew signal tristate
flabel metal2 s 3422 0 3478 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 1 nsew signal input
flabel metal2 s 24582 0 24638 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 2 nsew signal input
flabel metal2 s 26698 0 26754 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 3 nsew signal input
flabel metal2 s 28814 0 28870 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 4 nsew signal input
flabel metal2 s 30930 0 30986 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 5 nsew signal input
flabel metal2 s 33046 0 33102 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 6 nsew signal input
flabel metal2 s 35162 0 35218 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 7 nsew signal input
flabel metal2 s 37278 0 37334 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 8 nsew signal input
flabel metal2 s 39394 0 39450 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 9 nsew signal input
flabel metal2 s 41510 0 41566 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 10 nsew signal input
flabel metal2 s 43626 0 43682 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 11 nsew signal input
flabel metal2 s 5538 0 5594 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 12 nsew signal input
flabel metal2 s 7654 0 7710 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 13 nsew signal input
flabel metal2 s 9770 0 9826 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 14 nsew signal input
flabel metal2 s 11886 0 11942 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 15 nsew signal input
flabel metal2 s 14002 0 14058 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 16 nsew signal input
flabel metal2 s 16118 0 16174 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 17 nsew signal input
flabel metal2 s 18234 0 18290 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 18 nsew signal input
flabel metal2 s 20350 0 20406 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 19 nsew signal input
flabel metal2 s 22466 0 22522 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 20 nsew signal input
flabel metal2 s 34426 9840 34482 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 21 nsew signal tristate
flabel metal2 s 37186 9840 37242 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 22 nsew signal tristate
flabel metal2 s 37462 9840 37518 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 23 nsew signal tristate
flabel metal2 s 37738 9840 37794 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 24 nsew signal tristate
flabel metal2 s 38014 9840 38070 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 25 nsew signal tristate
flabel metal2 s 38290 9840 38346 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 26 nsew signal tristate
flabel metal2 s 38566 9840 38622 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 27 nsew signal tristate
flabel metal2 s 38842 9840 38898 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 28 nsew signal tristate
flabel metal2 s 39118 9840 39174 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 29 nsew signal tristate
flabel metal2 s 39394 9840 39450 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 30 nsew signal tristate
flabel metal2 s 39670 9840 39726 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 31 nsew signal tristate
flabel metal2 s 34702 9840 34758 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 32 nsew signal tristate
flabel metal2 s 34978 9840 35034 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 33 nsew signal tristate
flabel metal2 s 35254 9840 35310 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 34 nsew signal tristate
flabel metal2 s 35530 9840 35586 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 35 nsew signal tristate
flabel metal2 s 35806 9840 35862 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 36 nsew signal tristate
flabel metal2 s 36082 9840 36138 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 37 nsew signal tristate
flabel metal2 s 36358 9840 36414 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 38 nsew signal tristate
flabel metal2 s 36634 9840 36690 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 39 nsew signal tristate
flabel metal2 s 36910 9840 36966 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 40 nsew signal tristate
flabel metal2 s 5170 9840 5226 10000 0 FreeSans 224 90 0 0 N1BEG[0]
port 41 nsew signal tristate
flabel metal2 s 5446 9840 5502 10000 0 FreeSans 224 90 0 0 N1BEG[1]
port 42 nsew signal tristate
flabel metal2 s 5722 9840 5778 10000 0 FreeSans 224 90 0 0 N1BEG[2]
port 43 nsew signal tristate
flabel metal2 s 5998 9840 6054 10000 0 FreeSans 224 90 0 0 N1BEG[3]
port 44 nsew signal tristate
flabel metal2 s 6274 9840 6330 10000 0 FreeSans 224 90 0 0 N2BEG[0]
port 45 nsew signal tristate
flabel metal2 s 6550 9840 6606 10000 0 FreeSans 224 90 0 0 N2BEG[1]
port 46 nsew signal tristate
flabel metal2 s 6826 9840 6882 10000 0 FreeSans 224 90 0 0 N2BEG[2]
port 47 nsew signal tristate
flabel metal2 s 7102 9840 7158 10000 0 FreeSans 224 90 0 0 N2BEG[3]
port 48 nsew signal tristate
flabel metal2 s 7378 9840 7434 10000 0 FreeSans 224 90 0 0 N2BEG[4]
port 49 nsew signal tristate
flabel metal2 s 7654 9840 7710 10000 0 FreeSans 224 90 0 0 N2BEG[5]
port 50 nsew signal tristate
flabel metal2 s 7930 9840 7986 10000 0 FreeSans 224 90 0 0 N2BEG[6]
port 51 nsew signal tristate
flabel metal2 s 8206 9840 8262 10000 0 FreeSans 224 90 0 0 N2BEG[7]
port 52 nsew signal tristate
flabel metal2 s 8482 9840 8538 10000 0 FreeSans 224 90 0 0 N2BEGb[0]
port 53 nsew signal tristate
flabel metal2 s 8758 9840 8814 10000 0 FreeSans 224 90 0 0 N2BEGb[1]
port 54 nsew signal tristate
flabel metal2 s 9034 9840 9090 10000 0 FreeSans 224 90 0 0 N2BEGb[2]
port 55 nsew signal tristate
flabel metal2 s 9310 9840 9366 10000 0 FreeSans 224 90 0 0 N2BEGb[3]
port 56 nsew signal tristate
flabel metal2 s 9586 9840 9642 10000 0 FreeSans 224 90 0 0 N2BEGb[4]
port 57 nsew signal tristate
flabel metal2 s 9862 9840 9918 10000 0 FreeSans 224 90 0 0 N2BEGb[5]
port 58 nsew signal tristate
flabel metal2 s 10138 9840 10194 10000 0 FreeSans 224 90 0 0 N2BEGb[6]
port 59 nsew signal tristate
flabel metal2 s 10414 9840 10470 10000 0 FreeSans 224 90 0 0 N2BEGb[7]
port 60 nsew signal tristate
flabel metal2 s 10690 9840 10746 10000 0 FreeSans 224 90 0 0 N4BEG[0]
port 61 nsew signal tristate
flabel metal2 s 13450 9840 13506 10000 0 FreeSans 224 90 0 0 N4BEG[10]
port 62 nsew signal tristate
flabel metal2 s 13726 9840 13782 10000 0 FreeSans 224 90 0 0 N4BEG[11]
port 63 nsew signal tristate
flabel metal2 s 14002 9840 14058 10000 0 FreeSans 224 90 0 0 N4BEG[12]
port 64 nsew signal tristate
flabel metal2 s 14278 9840 14334 10000 0 FreeSans 224 90 0 0 N4BEG[13]
port 65 nsew signal tristate
flabel metal2 s 14554 9840 14610 10000 0 FreeSans 224 90 0 0 N4BEG[14]
port 66 nsew signal tristate
flabel metal2 s 14830 9840 14886 10000 0 FreeSans 224 90 0 0 N4BEG[15]
port 67 nsew signal tristate
flabel metal2 s 10966 9840 11022 10000 0 FreeSans 224 90 0 0 N4BEG[1]
port 68 nsew signal tristate
flabel metal2 s 11242 9840 11298 10000 0 FreeSans 224 90 0 0 N4BEG[2]
port 69 nsew signal tristate
flabel metal2 s 11518 9840 11574 10000 0 FreeSans 224 90 0 0 N4BEG[3]
port 70 nsew signal tristate
flabel metal2 s 11794 9840 11850 10000 0 FreeSans 224 90 0 0 N4BEG[4]
port 71 nsew signal tristate
flabel metal2 s 12070 9840 12126 10000 0 FreeSans 224 90 0 0 N4BEG[5]
port 72 nsew signal tristate
flabel metal2 s 12346 9840 12402 10000 0 FreeSans 224 90 0 0 N4BEG[6]
port 73 nsew signal tristate
flabel metal2 s 12622 9840 12678 10000 0 FreeSans 224 90 0 0 N4BEG[7]
port 74 nsew signal tristate
flabel metal2 s 12898 9840 12954 10000 0 FreeSans 224 90 0 0 N4BEG[8]
port 75 nsew signal tristate
flabel metal2 s 13174 9840 13230 10000 0 FreeSans 224 90 0 0 N4BEG[9]
port 76 nsew signal tristate
flabel metal2 s 15106 9840 15162 10000 0 FreeSans 224 90 0 0 NN4BEG[0]
port 77 nsew signal tristate
flabel metal2 s 17866 9840 17922 10000 0 FreeSans 224 90 0 0 NN4BEG[10]
port 78 nsew signal tristate
flabel metal2 s 18142 9840 18198 10000 0 FreeSans 224 90 0 0 NN4BEG[11]
port 79 nsew signal tristate
flabel metal2 s 18418 9840 18474 10000 0 FreeSans 224 90 0 0 NN4BEG[12]
port 80 nsew signal tristate
flabel metal2 s 18694 9840 18750 10000 0 FreeSans 224 90 0 0 NN4BEG[13]
port 81 nsew signal tristate
flabel metal2 s 18970 9840 19026 10000 0 FreeSans 224 90 0 0 NN4BEG[14]
port 82 nsew signal tristate
flabel metal2 s 19246 9840 19302 10000 0 FreeSans 224 90 0 0 NN4BEG[15]
port 83 nsew signal tristate
flabel metal2 s 15382 9840 15438 10000 0 FreeSans 224 90 0 0 NN4BEG[1]
port 84 nsew signal tristate
flabel metal2 s 15658 9840 15714 10000 0 FreeSans 224 90 0 0 NN4BEG[2]
port 85 nsew signal tristate
flabel metal2 s 15934 9840 15990 10000 0 FreeSans 224 90 0 0 NN4BEG[3]
port 86 nsew signal tristate
flabel metal2 s 16210 9840 16266 10000 0 FreeSans 224 90 0 0 NN4BEG[4]
port 87 nsew signal tristate
flabel metal2 s 16486 9840 16542 10000 0 FreeSans 224 90 0 0 NN4BEG[5]
port 88 nsew signal tristate
flabel metal2 s 16762 9840 16818 10000 0 FreeSans 224 90 0 0 NN4BEG[6]
port 89 nsew signal tristate
flabel metal2 s 17038 9840 17094 10000 0 FreeSans 224 90 0 0 NN4BEG[7]
port 90 nsew signal tristate
flabel metal2 s 17314 9840 17370 10000 0 FreeSans 224 90 0 0 NN4BEG[8]
port 91 nsew signal tristate
flabel metal2 s 17590 9840 17646 10000 0 FreeSans 224 90 0 0 NN4BEG[9]
port 92 nsew signal tristate
flabel metal2 s 19522 9840 19578 10000 0 FreeSans 224 90 0 0 S1END[0]
port 93 nsew signal input
flabel metal2 s 19798 9840 19854 10000 0 FreeSans 224 90 0 0 S1END[1]
port 94 nsew signal input
flabel metal2 s 20074 9840 20130 10000 0 FreeSans 224 90 0 0 S1END[2]
port 95 nsew signal input
flabel metal2 s 20350 9840 20406 10000 0 FreeSans 224 90 0 0 S1END[3]
port 96 nsew signal input
flabel metal2 s 20626 9840 20682 10000 0 FreeSans 224 90 0 0 S2END[0]
port 97 nsew signal input
flabel metal2 s 20902 9840 20958 10000 0 FreeSans 224 90 0 0 S2END[1]
port 98 nsew signal input
flabel metal2 s 21178 9840 21234 10000 0 FreeSans 224 90 0 0 S2END[2]
port 99 nsew signal input
flabel metal2 s 21454 9840 21510 10000 0 FreeSans 224 90 0 0 S2END[3]
port 100 nsew signal input
flabel metal2 s 21730 9840 21786 10000 0 FreeSans 224 90 0 0 S2END[4]
port 101 nsew signal input
flabel metal2 s 22006 9840 22062 10000 0 FreeSans 224 90 0 0 S2END[5]
port 102 nsew signal input
flabel metal2 s 22282 9840 22338 10000 0 FreeSans 224 90 0 0 S2END[6]
port 103 nsew signal input
flabel metal2 s 22558 9840 22614 10000 0 FreeSans 224 90 0 0 S2END[7]
port 104 nsew signal input
flabel metal2 s 22834 9840 22890 10000 0 FreeSans 224 90 0 0 S2MID[0]
port 105 nsew signal input
flabel metal2 s 23110 9840 23166 10000 0 FreeSans 224 90 0 0 S2MID[1]
port 106 nsew signal input
flabel metal2 s 23386 9840 23442 10000 0 FreeSans 224 90 0 0 S2MID[2]
port 107 nsew signal input
flabel metal2 s 23662 9840 23718 10000 0 FreeSans 224 90 0 0 S2MID[3]
port 108 nsew signal input
flabel metal2 s 23938 9840 23994 10000 0 FreeSans 224 90 0 0 S2MID[4]
port 109 nsew signal input
flabel metal2 s 24214 9840 24270 10000 0 FreeSans 224 90 0 0 S2MID[5]
port 110 nsew signal input
flabel metal2 s 24490 9840 24546 10000 0 FreeSans 224 90 0 0 S2MID[6]
port 111 nsew signal input
flabel metal2 s 24766 9840 24822 10000 0 FreeSans 224 90 0 0 S2MID[7]
port 112 nsew signal input
flabel metal2 s 25042 9840 25098 10000 0 FreeSans 224 90 0 0 S4END[0]
port 113 nsew signal input
flabel metal2 s 27802 9840 27858 10000 0 FreeSans 224 90 0 0 S4END[10]
port 114 nsew signal input
flabel metal2 s 28078 9840 28134 10000 0 FreeSans 224 90 0 0 S4END[11]
port 115 nsew signal input
flabel metal2 s 28354 9840 28410 10000 0 FreeSans 224 90 0 0 S4END[12]
port 116 nsew signal input
flabel metal2 s 28630 9840 28686 10000 0 FreeSans 224 90 0 0 S4END[13]
port 117 nsew signal input
flabel metal2 s 28906 9840 28962 10000 0 FreeSans 224 90 0 0 S4END[14]
port 118 nsew signal input
flabel metal2 s 29182 9840 29238 10000 0 FreeSans 224 90 0 0 S4END[15]
port 119 nsew signal input
flabel metal2 s 25318 9840 25374 10000 0 FreeSans 224 90 0 0 S4END[1]
port 120 nsew signal input
flabel metal2 s 25594 9840 25650 10000 0 FreeSans 224 90 0 0 S4END[2]
port 121 nsew signal input
flabel metal2 s 25870 9840 25926 10000 0 FreeSans 224 90 0 0 S4END[3]
port 122 nsew signal input
flabel metal2 s 26146 9840 26202 10000 0 FreeSans 224 90 0 0 S4END[4]
port 123 nsew signal input
flabel metal2 s 26422 9840 26478 10000 0 FreeSans 224 90 0 0 S4END[5]
port 124 nsew signal input
flabel metal2 s 26698 9840 26754 10000 0 FreeSans 224 90 0 0 S4END[6]
port 125 nsew signal input
flabel metal2 s 26974 9840 27030 10000 0 FreeSans 224 90 0 0 S4END[7]
port 126 nsew signal input
flabel metal2 s 27250 9840 27306 10000 0 FreeSans 224 90 0 0 S4END[8]
port 127 nsew signal input
flabel metal2 s 27526 9840 27582 10000 0 FreeSans 224 90 0 0 S4END[9]
port 128 nsew signal input
flabel metal2 s 29458 9840 29514 10000 0 FreeSans 224 90 0 0 SS4END[0]
port 129 nsew signal input
flabel metal2 s 32218 9840 32274 10000 0 FreeSans 224 90 0 0 SS4END[10]
port 130 nsew signal input
flabel metal2 s 32494 9840 32550 10000 0 FreeSans 224 90 0 0 SS4END[11]
port 131 nsew signal input
flabel metal2 s 32770 9840 32826 10000 0 FreeSans 224 90 0 0 SS4END[12]
port 132 nsew signal input
flabel metal2 s 33046 9840 33102 10000 0 FreeSans 224 90 0 0 SS4END[13]
port 133 nsew signal input
flabel metal2 s 33322 9840 33378 10000 0 FreeSans 224 90 0 0 SS4END[14]
port 134 nsew signal input
flabel metal2 s 33598 9840 33654 10000 0 FreeSans 224 90 0 0 SS4END[15]
port 135 nsew signal input
flabel metal2 s 29734 9840 29790 10000 0 FreeSans 224 90 0 0 SS4END[1]
port 136 nsew signal input
flabel metal2 s 30010 9840 30066 10000 0 FreeSans 224 90 0 0 SS4END[2]
port 137 nsew signal input
flabel metal2 s 30286 9840 30342 10000 0 FreeSans 224 90 0 0 SS4END[3]
port 138 nsew signal input
flabel metal2 s 30562 9840 30618 10000 0 FreeSans 224 90 0 0 SS4END[4]
port 139 nsew signal input
flabel metal2 s 30838 9840 30894 10000 0 FreeSans 224 90 0 0 SS4END[5]
port 140 nsew signal input
flabel metal2 s 31114 9840 31170 10000 0 FreeSans 224 90 0 0 SS4END[6]
port 141 nsew signal input
flabel metal2 s 31390 9840 31446 10000 0 FreeSans 224 90 0 0 SS4END[7]
port 142 nsew signal input
flabel metal2 s 31666 9840 31722 10000 0 FreeSans 224 90 0 0 SS4END[8]
port 143 nsew signal input
flabel metal2 s 31942 9840 31998 10000 0 FreeSans 224 90 0 0 SS4END[9]
port 144 nsew signal input
flabel metal2 s 1306 0 1362 160 0 FreeSans 224 90 0 0 UserCLK
port 145 nsew signal input
flabel metal2 s 33874 9840 33930 10000 0 FreeSans 224 90 0 0 UserCLKo
port 146 nsew signal tristate
flabel metal4 s 6291 2128 6611 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 16985 2128 17305 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 27679 2128 27999 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 38373 2128 38693 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 11638 2128 11958 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
flabel metal4 s 22332 2128 22652 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
flabel metal4 s 33026 2128 33346 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
flabel metal4 s 43720 2128 44040 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
rlabel metal1 22494 7072 22494 7072 0 vccd1
rlabel via1 22572 7616 22572 7616 0 vssd1
rlabel metal2 3450 1214 3450 1214 0 FrameStrobe[0]
rlabel metal2 24709 68 24709 68 0 FrameStrobe[10]
rlabel metal2 26726 1248 26726 1248 0 FrameStrobe[11]
rlabel metal2 28895 68 28895 68 0 FrameStrobe[12]
rlabel metal2 31011 68 31011 68 0 FrameStrobe[13]
rlabel metal2 33021 68 33021 68 0 FrameStrobe[14]
rlabel metal2 35190 1248 35190 1248 0 FrameStrobe[15]
rlabel metal2 37451 68 37451 68 0 FrameStrobe[16]
rlabel metal2 39567 68 39567 68 0 FrameStrobe[17]
rlabel metal2 41683 68 41683 68 0 FrameStrobe[18]
rlabel metal2 43601 68 43601 68 0 FrameStrobe[19]
rlabel metal2 5566 1248 5566 1248 0 FrameStrobe[1]
rlabel metal2 7735 68 7735 68 0 FrameStrobe[2]
rlabel metal2 9851 68 9851 68 0 FrameStrobe[3]
rlabel metal2 12059 68 12059 68 0 FrameStrobe[4]
rlabel metal2 14030 1248 14030 1248 0 FrameStrobe[5]
rlabel metal2 16291 68 16291 68 0 FrameStrobe[6]
rlabel metal2 18262 1248 18262 1248 0 FrameStrobe[7]
rlabel metal2 20523 68 20523 68 0 FrameStrobe[8]
rlabel metal2 22639 68 22639 68 0 FrameStrobe[9]
rlabel metal2 34454 8680 34454 8680 0 FrameStrobe_O[0]
rlabel metal1 37582 6834 37582 6834 0 FrameStrobe_O[10]
rlabel metal1 38088 6766 38088 6766 0 FrameStrobe_O[11]
rlabel metal1 38042 6630 38042 6630 0 FrameStrobe_O[12]
rlabel metal1 38778 6834 38778 6834 0 FrameStrobe_O[13]
rlabel metal2 38364 6834 38364 6834 0 FrameStrobe_O[14]
rlabel metal2 38778 6596 38778 6596 0 FrameStrobe_O[15]
rlabel metal2 38870 8680 38870 8680 0 FrameStrobe_O[16]
rlabel metal1 39652 6698 39652 6698 0 FrameStrobe_O[17]
rlabel metal2 39422 9173 39422 9173 0 FrameStrobe_O[18]
rlabel metal1 40342 6834 40342 6834 0 FrameStrobe_O[19]
rlabel metal2 34730 8646 34730 8646 0 FrameStrobe_O[1]
rlabel metal2 35006 8510 35006 8510 0 FrameStrobe_O[2]
rlabel metal1 35512 6834 35512 6834 0 FrameStrobe_O[3]
rlabel metal2 35558 8680 35558 8680 0 FrameStrobe_O[4]
rlabel metal1 36064 6834 36064 6834 0 FrameStrobe_O[5]
rlabel metal1 36386 6630 36386 6630 0 FrameStrobe_O[6]
rlabel metal2 36386 9173 36386 9173 0 FrameStrobe_O[7]
rlabel metal1 36984 6630 36984 6630 0 FrameStrobe_O[8]
rlabel metal2 36938 8680 36938 8680 0 FrameStrobe_O[9]
rlabel metal2 5198 8408 5198 8408 0 N1BEG[0]
rlabel metal1 5244 7514 5244 7514 0 N1BEG[1]
rlabel metal2 5750 8408 5750 8408 0 N1BEG[2]
rlabel metal1 5796 7514 5796 7514 0 N1BEG[3]
rlabel metal2 6302 9037 6302 9037 0 N2BEG[0]
rlabel metal1 6348 7242 6348 7242 0 N2BEG[1]
rlabel metal2 6854 8408 6854 8408 0 N2BEG[2]
rlabel metal2 7130 8340 7130 8340 0 N2BEG[3]
rlabel metal1 7222 7514 7222 7514 0 N2BEG[4]
rlabel metal2 7682 8340 7682 8340 0 N2BEG[5]
rlabel metal1 7774 7514 7774 7514 0 N2BEG[6]
rlabel metal2 8234 8340 8234 8340 0 N2BEG[7]
rlabel metal1 8326 7514 8326 7514 0 N2BEGb[0]
rlabel metal2 8786 8901 8786 8901 0 N2BEGb[1]
rlabel metal1 8878 7514 8878 7514 0 N2BEGb[2]
rlabel metal2 9338 8901 9338 8901 0 N2BEGb[3]
rlabel metal2 9614 8833 9614 8833 0 N2BEGb[4]
rlabel metal2 9890 8901 9890 8901 0 N2BEGb[5]
rlabel metal2 10166 8340 10166 8340 0 N2BEGb[6]
rlabel metal2 10442 9037 10442 9037 0 N2BEGb[7]
rlabel metal1 10304 7514 10304 7514 0 N4BEG[0]
rlabel metal2 13478 8408 13478 8408 0 N4BEG[10]
rlabel metal1 13524 7514 13524 7514 0 N4BEG[11]
rlabel metal2 14030 8136 14030 8136 0 N4BEG[12]
rlabel metal2 13846 7888 13846 7888 0 N4BEG[13]
rlabel metal2 14582 8408 14582 8408 0 N4BEG[14]
rlabel metal2 14858 8340 14858 8340 0 N4BEG[15]
rlabel metal2 10994 8340 10994 8340 0 N4BEG[1]
rlabel metal1 10902 7242 10902 7242 0 N4BEG[2]
rlabel metal2 11546 8629 11546 8629 0 N4BEG[3]
rlabel metal1 11040 7514 11040 7514 0 N4BEG[4]
rlabel metal2 12098 8901 12098 8901 0 N4BEG[5]
rlabel metal2 12374 8340 12374 8340 0 N4BEG[6]
rlabel metal2 12650 8306 12650 8306 0 N4BEG[7]
rlabel metal2 12926 8408 12926 8408 0 N4BEG[8]
rlabel metal1 12972 7514 12972 7514 0 N4BEG[9]
rlabel metal1 14950 7514 14950 7514 0 NN4BEG[0]
rlabel metal2 17894 8680 17894 8680 0 NN4BEG[10]
rlabel metal2 18170 8340 18170 8340 0 NN4BEG[11]
rlabel metal2 18446 8680 18446 8680 0 NN4BEG[12]
rlabel metal2 18722 8510 18722 8510 0 NN4BEG[13]
rlabel metal2 18998 9173 18998 9173 0 NN4BEG[14]
rlabel metal2 19274 8510 19274 8510 0 NN4BEG[15]
rlabel metal2 15410 8340 15410 8340 0 NN4BEG[1]
rlabel metal1 15502 7514 15502 7514 0 NN4BEG[2]
rlabel metal2 15962 8340 15962 8340 0 NN4BEG[3]
rlabel metal1 16054 7514 16054 7514 0 NN4BEG[4]
rlabel metal2 16514 8340 16514 8340 0 NN4BEG[5]
rlabel metal1 16606 7514 16606 7514 0 NN4BEG[6]
rlabel metal2 17066 9037 17066 9037 0 NN4BEG[7]
rlabel metal2 17342 8680 17342 8680 0 NN4BEG[8]
rlabel metal2 17618 8340 17618 8340 0 NN4BEG[9]
rlabel metal2 19550 9105 19550 9105 0 S1END[0]
rlabel metal2 19826 9105 19826 9105 0 S1END[1]
rlabel metal2 20102 9105 20102 9105 0 S1END[2]
rlabel metal2 20378 9105 20378 9105 0 S1END[3]
rlabel metal2 20654 8306 20654 8306 0 S2END[0]
rlabel metal2 20930 8612 20930 8612 0 S2END[1]
rlabel metal2 21206 8612 21206 8612 0 S2END[2]
rlabel metal2 21482 8612 21482 8612 0 S2END[3]
rlabel metal2 21758 8612 21758 8612 0 S2END[4]
rlabel metal2 22034 8612 22034 8612 0 S2END[5]
rlabel metal2 22310 9241 22310 9241 0 S2END[6]
rlabel metal2 22586 9105 22586 9105 0 S2END[7]
rlabel metal2 22862 8612 22862 8612 0 S2MID[0]
rlabel metal2 23138 8612 23138 8612 0 S2MID[1]
rlabel metal2 23414 8612 23414 8612 0 S2MID[2]
rlabel metal2 23690 8612 23690 8612 0 S2MID[3]
rlabel metal2 23966 9241 23966 9241 0 S2MID[4]
rlabel metal2 24242 9241 24242 9241 0 S2MID[5]
rlabel metal2 24518 9241 24518 9241 0 S2MID[6]
rlabel metal2 24794 8544 24794 8544 0 S2MID[7]
rlabel metal2 25070 9241 25070 9241 0 S4END[0]
rlabel metal2 27830 9241 27830 9241 0 S4END[10]
rlabel metal2 28106 8578 28106 8578 0 S4END[11]
rlabel metal2 28382 8680 28382 8680 0 S4END[12]
rlabel metal2 28658 9241 28658 9241 0 S4END[13]
rlabel metal2 28934 8561 28934 8561 0 S4END[14]
rlabel metal2 29210 8986 29210 8986 0 S4END[15]
rlabel metal2 25346 9054 25346 9054 0 S4END[1]
rlabel metal2 25622 8578 25622 8578 0 S4END[2]
rlabel metal2 25898 8646 25898 8646 0 S4END[3]
rlabel metal2 26174 8680 26174 8680 0 S4END[4]
rlabel metal2 26450 8578 26450 8578 0 S4END[5]
rlabel metal2 26726 9241 26726 9241 0 S4END[6]
rlabel metal2 27002 9309 27002 9309 0 S4END[7]
rlabel metal2 27278 8782 27278 8782 0 S4END[8]
rlabel metal2 27554 9377 27554 9377 0 S4END[9]
rlabel metal2 29486 8680 29486 8680 0 SS4END[0]
rlabel metal2 32246 8646 32246 8646 0 SS4END[10]
rlabel metal2 32522 8680 32522 8680 0 SS4END[11]
rlabel metal2 32798 8578 32798 8578 0 SS4END[12]
rlabel metal1 33074 6766 33074 6766 0 SS4END[13]
rlabel metal2 33350 9377 33350 9377 0 SS4END[14]
rlabel metal1 33948 6834 33948 6834 0 SS4END[15]
rlabel metal2 29762 9241 29762 9241 0 SS4END[1]
rlabel metal2 30038 8578 30038 8578 0 SS4END[2]
rlabel metal2 30314 9037 30314 9037 0 SS4END[3]
rlabel metal2 30590 8544 30590 8544 0 SS4END[4]
rlabel metal1 31786 7344 31786 7344 0 SS4END[5]
rlabel metal2 31142 8306 31142 8306 0 SS4END[6]
rlabel metal1 32154 7412 32154 7412 0 SS4END[7]
rlabel metal1 32154 7310 32154 7310 0 SS4END[8]
rlabel metal2 31970 8544 31970 8544 0 SS4END[9]
rlabel metal2 1334 1248 1334 1248 0 UserCLK
rlabel metal2 33902 8680 33902 8680 0 UserCLKo
rlabel metal1 5474 2618 5474 2618 0 net1
rlabel metal1 41538 2618 41538 2618 0 net10
rlabel metal2 7774 7412 7774 7412 0 net100
rlabel metal3 17572 6120 17572 6120 0 net101
rlabel metal2 21114 7616 21114 7616 0 net102
rlabel metal2 11178 7361 11178 7361 0 net103
rlabel metal2 13662 7650 13662 7650 0 net104
rlabel metal2 22034 5729 22034 5729 0 net105
rlabel metal1 21390 6630 21390 6630 0 net106
rlabel metal2 21206 6069 21206 6069 0 net107
rlabel metal1 21068 6902 21068 6902 0 net108
rlabel metal1 9154 6256 9154 6256 0 net109
rlabel metal1 42274 7310 42274 7310 0 net11
rlabel metal2 20654 6545 20654 6545 0 net110
rlabel metal2 9706 6800 9706 6800 0 net111
rlabel metal2 9430 6460 9430 6460 0 net112
rlabel metal1 11132 6426 11132 6426 0 net113
rlabel metal1 10396 7378 10396 7378 0 net114
rlabel metal2 13938 5678 13938 5678 0 net115
rlabel metal2 24058 5321 24058 5321 0 net116
rlabel via2 17894 6205 17894 6205 0 net117
rlabel metal1 21022 6120 21022 6120 0 net118
rlabel metal2 18170 5848 18170 5848 0 net119
rlabel metal2 34270 4862 34270 4862 0 net12
rlabel metal1 13846 6392 13846 6392 0 net120
rlabel metal2 10810 5712 10810 5712 0 net121
rlabel metal2 16330 7072 16330 7072 0 net122
rlabel metal2 11362 5644 11362 5644 0 net123
rlabel metal2 20746 7701 20746 7701 0 net124
rlabel metal2 12006 5406 12006 5406 0 net125
rlabel metal2 14214 5916 14214 5916 0 net126
rlabel metal2 13754 5950 13754 5950 0 net127
rlabel metal2 13018 6188 13018 6188 0 net128
rlabel metal2 16146 6137 16146 6137 0 net129
rlabel metal1 9522 2482 9522 2482 0 net13
rlabel metal1 14582 6426 14582 6426 0 net130
rlabel metal1 17986 6426 17986 6426 0 net131
rlabel metal2 18354 6562 18354 6562 0 net132
rlabel metal2 18630 6902 18630 6902 0 net133
rlabel metal2 18998 6902 18998 6902 0 net134
rlabel metal1 19458 6970 19458 6970 0 net135
rlabel metal1 19458 7344 19458 7344 0 net136
rlabel metal1 15226 6766 15226 6766 0 net137
rlabel metal1 14858 7446 14858 7446 0 net138
rlabel metal2 15318 6562 15318 6562 0 net139
rlabel metal2 10074 2176 10074 2176 0 net14
rlabel metal1 15640 6426 15640 6426 0 net140
rlabel metal1 16422 6426 16422 6426 0 net141
rlabel metal1 16652 6154 16652 6154 0 net142
rlabel metal1 17434 6426 17434 6426 0 net143
rlabel metal2 17342 6766 17342 6766 0 net144
rlabel metal1 17618 6698 17618 6698 0 net145
rlabel metal1 32430 6664 32430 6664 0 net146
rlabel metal1 34914 6732 34914 6732 0 net147
rlabel metal1 12420 2618 12420 2618 0 net15
rlabel metal1 14674 2312 14674 2312 0 net16
rlabel metal1 16238 2516 16238 2516 0 net17
rlabel metal1 18538 2618 18538 2618 0 net18
rlabel metal1 20654 5202 20654 5202 0 net19
rlabel metal1 24886 2618 24886 2618 0 net2
rlabel metal1 22770 2618 22770 2618 0 net20
rlabel metal2 19550 5814 19550 5814 0 net21
rlabel metal2 19826 6188 19826 6188 0 net22
rlabel metal1 20102 6664 20102 6664 0 net23
rlabel metal2 13662 5984 13662 5984 0 net24
rlabel metal1 17434 5848 17434 5848 0 net25
rlabel metal2 16514 6103 16514 6103 0 net26
rlabel metal1 16790 7276 16790 7276 0 net27
rlabel metal1 20516 6766 20516 6766 0 net28
rlabel metal2 20470 6630 20470 6630 0 net29
rlabel metal2 37030 2244 37030 2244 0 net3
rlabel metal1 21712 6766 21712 6766 0 net30
rlabel metal1 21022 6800 21022 6800 0 net31
rlabel metal1 21298 6732 21298 6732 0 net32
rlabel metal2 21942 6766 21942 6766 0 net33
rlabel metal1 22448 6290 22448 6290 0 net34
rlabel metal1 22862 6290 22862 6290 0 net35
rlabel metal1 22402 7412 22402 7412 0 net36
rlabel metal1 23552 6766 23552 6766 0 net37
rlabel metal1 23230 7344 23230 7344 0 net38
rlabel metal1 24426 7446 24426 7446 0 net39
rlabel metal2 37306 4420 37306 4420 0 net4
rlabel metal1 24978 7344 24978 7344 0 net40
rlabel metal2 14122 7106 14122 7106 0 net41
rlabel metal1 27922 6800 27922 6800 0 net42
rlabel metal1 28290 6732 28290 6732 0 net43
rlabel metal1 28796 6766 28796 6766 0 net44
rlabel metal1 29394 6766 29394 6766 0 net45
rlabel metal1 29762 6766 29762 6766 0 net46
rlabel metal1 30084 6766 30084 6766 0 net47
rlabel metal1 24886 6732 24886 6732 0 net48
rlabel metal1 25162 6868 25162 6868 0 net49
rlabel metal2 36754 4284 36754 4284 0 net5
rlabel metal1 25438 6834 25438 6834 0 net50
rlabel metal1 25852 6290 25852 6290 0 net51
rlabel metal1 26266 6800 26266 6800 0 net52
rlabel metal1 26542 6732 26542 6732 0 net53
rlabel metal1 26956 6766 26956 6766 0 net54
rlabel metal1 27324 6766 27324 6766 0 net55
rlabel metal1 27692 6766 27692 6766 0 net56
rlabel metal1 30360 6766 30360 6766 0 net57
rlabel metal1 32890 7242 32890 7242 0 net58
rlabel metal1 33488 7514 33488 7514 0 net59
rlabel metal1 33626 2618 33626 2618 0 net6
rlabel metal2 33718 7956 33718 7956 0 net60
rlabel metal2 33350 6681 33350 6681 0 net61
rlabel metal2 33626 5933 33626 5933 0 net62
rlabel metal2 34454 5661 34454 5661 0 net63
rlabel metal1 19090 6324 19090 6324 0 net64
rlabel metal1 19182 6324 19182 6324 0 net65
rlabel metal2 18814 6647 18814 6647 0 net66
rlabel metal2 19458 7378 19458 7378 0 net67
rlabel metal1 18262 5848 18262 5848 0 net68
rlabel metal2 17710 6426 17710 6426 0 net69
rlabel metal1 37122 7344 37122 7344 0 net7
rlabel metal2 32338 6392 32338 6392 0 net70
rlabel metal2 32614 6749 32614 6749 0 net71
rlabel metal1 32798 7174 32798 7174 0 net72
rlabel metal1 9660 2006 9660 2006 0 net73
rlabel metal2 33718 6528 33718 6528 0 net74
rlabel metal2 37674 4760 37674 4760 0 net75
rlabel metal1 37674 7446 37674 7446 0 net76
rlabel metal1 37766 6426 37766 6426 0 net77
rlabel metal1 38318 6154 38318 6154 0 net78
rlabel metal1 38410 6392 38410 6392 0 net79
rlabel metal1 38042 2448 38042 2448 0 net8
rlabel metal1 38134 6970 38134 6970 0 net80
rlabel metal1 38916 7310 38916 7310 0 net81
rlabel metal1 39744 6766 39744 6766 0 net82
rlabel metal1 40526 7480 40526 7480 0 net83
rlabel metal1 40756 6766 40756 6766 0 net84
rlabel metal1 34730 6086 34730 6086 0 net85
rlabel metal2 35926 7004 35926 7004 0 net86
rlabel metal1 35098 2618 35098 2618 0 net87
rlabel metal1 36340 7446 36340 7446 0 net88
rlabel metal2 36018 4828 36018 4828 0 net89
rlabel metal1 39606 2618 39606 2618 0 net9
rlabel metal2 36570 5644 36570 5644 0 net90
rlabel metal1 37490 7378 37490 7378 0 net91
rlabel metal2 37122 6494 37122 6494 0 net92
rlabel metal1 26059 2890 26059 2890 0 net93
rlabel metal1 6992 6426 6992 6426 0 net94
rlabel metal1 5658 6154 5658 6154 0 net95
rlabel metal1 5842 6426 5842 6426 0 net96
rlabel metal1 5842 7446 5842 7446 0 net97
rlabel metal2 6670 7429 6670 7429 0 net98
rlabel metal2 5842 7327 5842 7327 0 net99
<< properties >>
string FIXED_BBOX 0 0 45000 10000
<< end >>
