magic
tech sky130A
magscale 1 2
timestamp 1733416662
<< obsli1 >>
rect 1104 1071 43884 89233
<< obsm1 >>
rect 14 76 44882 90024
<< metal2 >>
rect 5354 90640 5410 90800
rect 5630 90640 5686 90800
rect 5906 90640 5962 90800
rect 6182 90640 6238 90800
rect 6458 90640 6514 90800
rect 6734 90640 6790 90800
rect 7010 90640 7066 90800
rect 7286 90640 7342 90800
rect 7562 90640 7618 90800
rect 7838 90640 7894 90800
rect 8114 90640 8170 90800
rect 8390 90640 8446 90800
rect 8666 90640 8722 90800
rect 8942 90640 8998 90800
rect 9218 90640 9274 90800
rect 9494 90640 9550 90800
rect 9770 90640 9826 90800
rect 10046 90640 10102 90800
rect 10322 90640 10378 90800
rect 10598 90640 10654 90800
rect 10874 90640 10930 90800
rect 11150 90640 11206 90800
rect 11426 90640 11482 90800
rect 11702 90640 11758 90800
rect 11978 90640 12034 90800
rect 12254 90640 12310 90800
rect 12530 90640 12586 90800
rect 12806 90640 12862 90800
rect 13082 90640 13138 90800
rect 13358 90640 13414 90800
rect 13634 90640 13690 90800
rect 13910 90640 13966 90800
rect 14186 90640 14242 90800
rect 14462 90640 14518 90800
rect 14738 90640 14794 90800
rect 15014 90640 15070 90800
rect 15290 90640 15346 90800
rect 15566 90640 15622 90800
rect 15842 90640 15898 90800
rect 16118 90640 16174 90800
rect 16394 90640 16450 90800
rect 16670 90640 16726 90800
rect 16946 90640 17002 90800
rect 17222 90640 17278 90800
rect 17498 90640 17554 90800
rect 17774 90640 17830 90800
rect 18050 90640 18106 90800
rect 18326 90640 18382 90800
rect 18602 90640 18658 90800
rect 18878 90640 18934 90800
rect 19154 90640 19210 90800
rect 19430 90640 19486 90800
rect 19706 90640 19762 90800
rect 19982 90640 20038 90800
rect 20258 90640 20314 90800
rect 20534 90640 20590 90800
rect 20810 90640 20866 90800
rect 21086 90640 21142 90800
rect 21362 90640 21418 90800
rect 21638 90640 21694 90800
rect 21914 90640 21970 90800
rect 22190 90640 22246 90800
rect 22466 90640 22522 90800
rect 22742 90640 22798 90800
rect 23018 90640 23074 90800
rect 23294 90640 23350 90800
rect 23570 90640 23626 90800
rect 23846 90640 23902 90800
rect 24122 90640 24178 90800
rect 24398 90640 24454 90800
rect 24674 90640 24730 90800
rect 24950 90640 25006 90800
rect 25226 90640 25282 90800
rect 25502 90640 25558 90800
rect 25778 90640 25834 90800
rect 26054 90640 26110 90800
rect 26330 90640 26386 90800
rect 26606 90640 26662 90800
rect 26882 90640 26938 90800
rect 27158 90640 27214 90800
rect 27434 90640 27490 90800
rect 27710 90640 27766 90800
rect 27986 90640 28042 90800
rect 28262 90640 28318 90800
rect 28538 90640 28594 90800
rect 28814 90640 28870 90800
rect 29090 90640 29146 90800
rect 29366 90640 29422 90800
rect 29642 90640 29698 90800
rect 29918 90640 29974 90800
rect 30194 90640 30250 90800
rect 30470 90640 30526 90800
rect 30746 90640 30802 90800
rect 31022 90640 31078 90800
rect 31298 90640 31354 90800
rect 31574 90640 31630 90800
rect 31850 90640 31906 90800
rect 32126 90640 32182 90800
rect 32402 90640 32458 90800
rect 32678 90640 32734 90800
rect 32954 90640 33010 90800
rect 33230 90640 33286 90800
rect 33506 90640 33562 90800
rect 33782 90640 33838 90800
rect 34058 90640 34114 90800
rect 34334 90640 34390 90800
rect 34610 90640 34666 90800
rect 34886 90640 34942 90800
rect 35162 90640 35218 90800
rect 35438 90640 35494 90800
rect 35714 90640 35770 90800
rect 35990 90640 36046 90800
rect 36266 90640 36322 90800
rect 36542 90640 36598 90800
rect 36818 90640 36874 90800
rect 37094 90640 37150 90800
rect 37370 90640 37426 90800
rect 37646 90640 37702 90800
rect 37922 90640 37978 90800
rect 38198 90640 38254 90800
rect 38474 90640 38530 90800
rect 38750 90640 38806 90800
rect 39026 90640 39082 90800
rect 39302 90640 39358 90800
rect 39578 90640 39634 90800
rect 5354 0 5410 160
rect 5630 0 5686 160
rect 5906 0 5962 160
rect 6182 0 6238 160
rect 6458 0 6514 160
rect 6734 0 6790 160
rect 7010 0 7066 160
rect 7286 0 7342 160
rect 7562 0 7618 160
rect 7838 0 7894 160
rect 8114 0 8170 160
rect 8390 0 8446 160
rect 8666 0 8722 160
rect 8942 0 8998 160
rect 9218 0 9274 160
rect 9494 0 9550 160
rect 9770 0 9826 160
rect 10046 0 10102 160
rect 10322 0 10378 160
rect 10598 0 10654 160
rect 10874 0 10930 160
rect 11150 0 11206 160
rect 11426 0 11482 160
rect 11702 0 11758 160
rect 11978 0 12034 160
rect 12254 0 12310 160
rect 12530 0 12586 160
rect 12806 0 12862 160
rect 13082 0 13138 160
rect 13358 0 13414 160
rect 13634 0 13690 160
rect 13910 0 13966 160
rect 14186 0 14242 160
rect 14462 0 14518 160
rect 14738 0 14794 160
rect 15014 0 15070 160
rect 15290 0 15346 160
rect 15566 0 15622 160
rect 15842 0 15898 160
rect 16118 0 16174 160
rect 16394 0 16450 160
rect 16670 0 16726 160
rect 16946 0 17002 160
rect 17222 0 17278 160
rect 17498 0 17554 160
rect 17774 0 17830 160
rect 18050 0 18106 160
rect 18326 0 18382 160
rect 18602 0 18658 160
rect 18878 0 18934 160
rect 19154 0 19210 160
rect 19430 0 19486 160
rect 19706 0 19762 160
rect 19982 0 20038 160
rect 20258 0 20314 160
rect 20534 0 20590 160
rect 20810 0 20866 160
rect 21086 0 21142 160
rect 21362 0 21418 160
rect 21638 0 21694 160
rect 21914 0 21970 160
rect 22190 0 22246 160
rect 22466 0 22522 160
rect 22742 0 22798 160
rect 23018 0 23074 160
rect 23294 0 23350 160
rect 23570 0 23626 160
rect 23846 0 23902 160
rect 24122 0 24178 160
rect 24398 0 24454 160
rect 24674 0 24730 160
rect 24950 0 25006 160
rect 25226 0 25282 160
rect 25502 0 25558 160
rect 25778 0 25834 160
rect 26054 0 26110 160
rect 26330 0 26386 160
rect 26606 0 26662 160
rect 26882 0 26938 160
rect 27158 0 27214 160
rect 27434 0 27490 160
rect 27710 0 27766 160
rect 27986 0 28042 160
rect 28262 0 28318 160
rect 28538 0 28594 160
rect 28814 0 28870 160
rect 29090 0 29146 160
rect 29366 0 29422 160
rect 29642 0 29698 160
rect 29918 0 29974 160
rect 30194 0 30250 160
rect 30470 0 30526 160
rect 30746 0 30802 160
rect 31022 0 31078 160
rect 31298 0 31354 160
rect 31574 0 31630 160
rect 31850 0 31906 160
rect 32126 0 32182 160
rect 32402 0 32458 160
rect 32678 0 32734 160
rect 32954 0 33010 160
rect 33230 0 33286 160
rect 33506 0 33562 160
rect 33782 0 33838 160
rect 34058 0 34114 160
rect 34334 0 34390 160
rect 34610 0 34666 160
rect 34886 0 34942 160
rect 35162 0 35218 160
rect 35438 0 35494 160
rect 35714 0 35770 160
rect 35990 0 36046 160
rect 36266 0 36322 160
rect 36542 0 36598 160
rect 36818 0 36874 160
rect 37094 0 37150 160
rect 37370 0 37426 160
rect 37646 0 37702 160
rect 37922 0 37978 160
rect 38198 0 38254 160
rect 38474 0 38530 160
rect 38750 0 38806 160
rect 39026 0 39082 160
rect 39302 0 39358 160
rect 39578 0 39634 160
<< obsm2 >>
rect 20 90584 5298 90640
rect 5466 90584 5574 90640
rect 5742 90584 5850 90640
rect 6018 90584 6126 90640
rect 6294 90584 6402 90640
rect 6570 90584 6678 90640
rect 6846 90584 6954 90640
rect 7122 90584 7230 90640
rect 7398 90584 7506 90640
rect 7674 90584 7782 90640
rect 7950 90584 8058 90640
rect 8226 90584 8334 90640
rect 8502 90584 8610 90640
rect 8778 90584 8886 90640
rect 9054 90584 9162 90640
rect 9330 90584 9438 90640
rect 9606 90584 9714 90640
rect 9882 90584 9990 90640
rect 10158 90584 10266 90640
rect 10434 90584 10542 90640
rect 10710 90584 10818 90640
rect 10986 90584 11094 90640
rect 11262 90584 11370 90640
rect 11538 90584 11646 90640
rect 11814 90584 11922 90640
rect 12090 90584 12198 90640
rect 12366 90584 12474 90640
rect 12642 90584 12750 90640
rect 12918 90584 13026 90640
rect 13194 90584 13302 90640
rect 13470 90584 13578 90640
rect 13746 90584 13854 90640
rect 14022 90584 14130 90640
rect 14298 90584 14406 90640
rect 14574 90584 14682 90640
rect 14850 90584 14958 90640
rect 15126 90584 15234 90640
rect 15402 90584 15510 90640
rect 15678 90584 15786 90640
rect 15954 90584 16062 90640
rect 16230 90584 16338 90640
rect 16506 90584 16614 90640
rect 16782 90584 16890 90640
rect 17058 90584 17166 90640
rect 17334 90584 17442 90640
rect 17610 90584 17718 90640
rect 17886 90584 17994 90640
rect 18162 90584 18270 90640
rect 18438 90584 18546 90640
rect 18714 90584 18822 90640
rect 18990 90584 19098 90640
rect 19266 90584 19374 90640
rect 19542 90584 19650 90640
rect 19818 90584 19926 90640
rect 20094 90584 20202 90640
rect 20370 90584 20478 90640
rect 20646 90584 20754 90640
rect 20922 90584 21030 90640
rect 21198 90584 21306 90640
rect 21474 90584 21582 90640
rect 21750 90584 21858 90640
rect 22026 90584 22134 90640
rect 22302 90584 22410 90640
rect 22578 90584 22686 90640
rect 22854 90584 22962 90640
rect 23130 90584 23238 90640
rect 23406 90584 23514 90640
rect 23682 90584 23790 90640
rect 23958 90584 24066 90640
rect 24234 90584 24342 90640
rect 24510 90584 24618 90640
rect 24786 90584 24894 90640
rect 25062 90584 25170 90640
rect 25338 90584 25446 90640
rect 25614 90584 25722 90640
rect 25890 90584 25998 90640
rect 26166 90584 26274 90640
rect 26442 90584 26550 90640
rect 26718 90584 26826 90640
rect 26994 90584 27102 90640
rect 27270 90584 27378 90640
rect 27546 90584 27654 90640
rect 27822 90584 27930 90640
rect 28098 90584 28206 90640
rect 28374 90584 28482 90640
rect 28650 90584 28758 90640
rect 28926 90584 29034 90640
rect 29202 90584 29310 90640
rect 29478 90584 29586 90640
rect 29754 90584 29862 90640
rect 30030 90584 30138 90640
rect 30306 90584 30414 90640
rect 30582 90584 30690 90640
rect 30858 90584 30966 90640
rect 31134 90584 31242 90640
rect 31410 90584 31518 90640
rect 31686 90584 31794 90640
rect 31962 90584 32070 90640
rect 32238 90584 32346 90640
rect 32514 90584 32622 90640
rect 32790 90584 32898 90640
rect 33066 90584 33174 90640
rect 33342 90584 33450 90640
rect 33618 90584 33726 90640
rect 33894 90584 34002 90640
rect 34170 90584 34278 90640
rect 34446 90584 34554 90640
rect 34722 90584 34830 90640
rect 34998 90584 35106 90640
rect 35274 90584 35382 90640
rect 35550 90584 35658 90640
rect 35826 90584 35934 90640
rect 36102 90584 36210 90640
rect 36378 90584 36486 90640
rect 36654 90584 36762 90640
rect 36930 90584 37038 90640
rect 37206 90584 37314 90640
rect 37482 90584 37590 90640
rect 37758 90584 37866 90640
rect 38034 90584 38142 90640
rect 38310 90584 38418 90640
rect 38586 90584 38694 90640
rect 38862 90584 38970 90640
rect 39138 90584 39246 90640
rect 39414 90584 39522 90640
rect 39690 90584 44876 90640
rect 20 216 44876 90584
rect 20 54 5298 216
rect 5466 54 5574 216
rect 5742 54 5850 216
rect 6018 54 6126 216
rect 6294 54 6402 216
rect 6570 54 6678 216
rect 6846 54 6954 216
rect 7122 54 7230 216
rect 7398 54 7506 216
rect 7674 54 7782 216
rect 7950 54 8058 216
rect 8226 54 8334 216
rect 8502 54 8610 216
rect 8778 54 8886 216
rect 9054 54 9162 216
rect 9330 54 9438 216
rect 9606 54 9714 216
rect 9882 54 9990 216
rect 10158 54 10266 216
rect 10434 54 10542 216
rect 10710 54 10818 216
rect 10986 54 11094 216
rect 11262 54 11370 216
rect 11538 54 11646 216
rect 11814 54 11922 216
rect 12090 54 12198 216
rect 12366 54 12474 216
rect 12642 54 12750 216
rect 12918 54 13026 216
rect 13194 54 13302 216
rect 13470 54 13578 216
rect 13746 54 13854 216
rect 14022 54 14130 216
rect 14298 54 14406 216
rect 14574 54 14682 216
rect 14850 54 14958 216
rect 15126 54 15234 216
rect 15402 54 15510 216
rect 15678 54 15786 216
rect 15954 54 16062 216
rect 16230 54 16338 216
rect 16506 54 16614 216
rect 16782 54 16890 216
rect 17058 54 17166 216
rect 17334 54 17442 216
rect 17610 54 17718 216
rect 17886 54 17994 216
rect 18162 54 18270 216
rect 18438 54 18546 216
rect 18714 54 18822 216
rect 18990 54 19098 216
rect 19266 54 19374 216
rect 19542 54 19650 216
rect 19818 54 19926 216
rect 20094 54 20202 216
rect 20370 54 20478 216
rect 20646 54 20754 216
rect 20922 54 21030 216
rect 21198 54 21306 216
rect 21474 54 21582 216
rect 21750 54 21858 216
rect 22026 54 22134 216
rect 22302 54 22410 216
rect 22578 54 22686 216
rect 22854 54 22962 216
rect 23130 54 23238 216
rect 23406 54 23514 216
rect 23682 54 23790 216
rect 23958 54 24066 216
rect 24234 54 24342 216
rect 24510 54 24618 216
rect 24786 54 24894 216
rect 25062 54 25170 216
rect 25338 54 25446 216
rect 25614 54 25722 216
rect 25890 54 25998 216
rect 26166 54 26274 216
rect 26442 54 26550 216
rect 26718 54 26826 216
rect 26994 54 27102 216
rect 27270 54 27378 216
rect 27546 54 27654 216
rect 27822 54 27930 216
rect 28098 54 28206 216
rect 28374 54 28482 216
rect 28650 54 28758 216
rect 28926 54 29034 216
rect 29202 54 29310 216
rect 29478 54 29586 216
rect 29754 54 29862 216
rect 30030 54 30138 216
rect 30306 54 30414 216
rect 30582 54 30690 216
rect 30858 54 30966 216
rect 31134 54 31242 216
rect 31410 54 31518 216
rect 31686 54 31794 216
rect 31962 54 32070 216
rect 32238 54 32346 216
rect 32514 54 32622 216
rect 32790 54 32898 216
rect 33066 54 33174 216
rect 33342 54 33450 216
rect 33618 54 33726 216
rect 33894 54 34002 216
rect 34170 54 34278 216
rect 34446 54 34554 216
rect 34722 54 34830 216
rect 34998 54 35106 216
rect 35274 54 35382 216
rect 35550 54 35658 216
rect 35826 54 35934 216
rect 36102 54 36210 216
rect 36378 54 36486 216
rect 36654 54 36762 216
rect 36930 54 37038 216
rect 37206 54 37314 216
rect 37482 54 37590 216
rect 37758 54 37866 216
rect 38034 54 38142 216
rect 38310 54 38418 216
rect 38586 54 38694 216
rect 38862 54 38970 216
rect 39138 54 39246 216
rect 39414 54 39522 216
rect 39690 54 44876 216
<< metal3 >>
rect 0 85144 160 85264
rect 0 84872 160 84992
rect 0 84600 160 84720
rect 0 84328 160 84448
rect 0 84056 160 84176
rect 0 83784 160 83904
rect 0 83512 160 83632
rect 0 83240 160 83360
rect 0 82968 160 83088
rect 0 82696 160 82816
rect 0 82424 160 82544
rect 0 82152 160 82272
rect 0 81880 160 82000
rect 0 81608 160 81728
rect 0 81336 160 81456
rect 0 81064 160 81184
rect 0 80792 160 80912
rect 0 80520 160 80640
rect 0 80248 160 80368
rect 0 79976 160 80096
rect 0 79704 160 79824
rect 0 79432 160 79552
rect 0 79160 160 79280
rect 0 78888 160 79008
rect 0 78616 160 78736
rect 0 78344 160 78464
rect 0 78072 160 78192
rect 0 77800 160 77920
rect 0 77528 160 77648
rect 0 77256 160 77376
rect 0 76984 160 77104
rect 0 76712 160 76832
rect 0 76440 160 76560
rect 0 76168 160 76288
rect 0 75896 160 76016
rect 0 75624 160 75744
rect 0 75352 160 75472
rect 0 75080 160 75200
rect 0 74808 160 74928
rect 0 74536 160 74656
rect 0 74264 160 74384
rect 0 73992 160 74112
rect 0 73720 160 73840
rect 0 73448 160 73568
rect 0 73176 160 73296
rect 0 72904 160 73024
rect 0 72632 160 72752
rect 0 72360 160 72480
rect 0 72088 160 72208
rect 0 71816 160 71936
rect 0 71544 160 71664
rect 0 71272 160 71392
rect 0 71000 160 71120
rect 0 70728 160 70848
rect 0 70456 160 70576
rect 0 70184 160 70304
rect 0 69912 160 70032
rect 0 69640 160 69760
rect 0 69368 160 69488
rect 0 69096 160 69216
rect 0 68824 160 68944
rect 0 68552 160 68672
rect 0 68280 160 68400
rect 0 68008 160 68128
rect 0 67736 160 67856
rect 0 67464 160 67584
rect 0 67192 160 67312
rect 0 66920 160 67040
rect 0 66648 160 66768
rect 0 66376 160 66496
rect 0 66104 160 66224
rect 0 65832 160 65952
rect 0 65560 160 65680
rect 0 65288 160 65408
rect 0 65016 160 65136
rect 0 64744 160 64864
rect 0 64472 160 64592
rect 0 64200 160 64320
rect 0 63928 160 64048
rect 0 63656 160 63776
rect 0 63384 160 63504
rect 0 63112 160 63232
rect 0 62840 160 62960
rect 0 62568 160 62688
rect 0 62296 160 62416
rect 0 62024 160 62144
rect 0 61752 160 61872
rect 0 61480 160 61600
rect 0 61208 160 61328
rect 0 60936 160 61056
rect 0 60664 160 60784
rect 0 60392 160 60512
rect 0 60120 160 60240
rect 0 59848 160 59968
rect 0 59576 160 59696
rect 0 59304 160 59424
rect 0 59032 160 59152
rect 0 58760 160 58880
rect 0 58488 160 58608
rect 0 58216 160 58336
rect 0 57944 160 58064
rect 0 57672 160 57792
rect 0 57400 160 57520
rect 0 57128 160 57248
rect 0 56856 160 56976
rect 0 56584 160 56704
rect 0 56312 160 56432
rect 0 56040 160 56160
rect 0 55768 160 55888
rect 0 55496 160 55616
rect 0 55224 160 55344
rect 0 54952 160 55072
rect 0 54680 160 54800
rect 0 54408 160 54528
rect 0 54136 160 54256
rect 0 53864 160 53984
rect 0 53592 160 53712
rect 0 53320 160 53440
rect 0 53048 160 53168
rect 0 52776 160 52896
rect 0 52504 160 52624
rect 0 52232 160 52352
rect 0 51960 160 52080
rect 0 51688 160 51808
rect 0 51416 160 51536
rect 0 51144 160 51264
rect 0 50872 160 50992
rect 0 50600 160 50720
rect 44840 85144 45000 85264
rect 44840 84872 45000 84992
rect 44840 84600 45000 84720
rect 44840 84328 45000 84448
rect 44840 84056 45000 84176
rect 44840 83784 45000 83904
rect 44840 83512 45000 83632
rect 44840 83240 45000 83360
rect 44840 82968 45000 83088
rect 44840 82696 45000 82816
rect 44840 82424 45000 82544
rect 44840 82152 45000 82272
rect 44840 81880 45000 82000
rect 44840 81608 45000 81728
rect 44840 81336 45000 81456
rect 44840 81064 45000 81184
rect 44840 80792 45000 80912
rect 44840 80520 45000 80640
rect 44840 80248 45000 80368
rect 44840 79976 45000 80096
rect 44840 79704 45000 79824
rect 44840 79432 45000 79552
rect 44840 79160 45000 79280
rect 44840 78888 45000 79008
rect 44840 78616 45000 78736
rect 44840 78344 45000 78464
rect 44840 78072 45000 78192
rect 44840 77800 45000 77920
rect 44840 77528 45000 77648
rect 44840 77256 45000 77376
rect 44840 76984 45000 77104
rect 44840 76712 45000 76832
rect 44840 76440 45000 76560
rect 44840 76168 45000 76288
rect 44840 75896 45000 76016
rect 44840 75624 45000 75744
rect 44840 75352 45000 75472
rect 44840 75080 45000 75200
rect 44840 74808 45000 74928
rect 44840 74536 45000 74656
rect 44840 74264 45000 74384
rect 44840 73992 45000 74112
rect 44840 73720 45000 73840
rect 44840 73448 45000 73568
rect 44840 73176 45000 73296
rect 44840 72904 45000 73024
rect 44840 72632 45000 72752
rect 44840 72360 45000 72480
rect 44840 72088 45000 72208
rect 44840 71816 45000 71936
rect 44840 71544 45000 71664
rect 44840 71272 45000 71392
rect 44840 71000 45000 71120
rect 44840 70728 45000 70848
rect 44840 70456 45000 70576
rect 44840 70184 45000 70304
rect 44840 69912 45000 70032
rect 44840 69640 45000 69760
rect 44840 69368 45000 69488
rect 44840 69096 45000 69216
rect 44840 68824 45000 68944
rect 44840 68552 45000 68672
rect 44840 68280 45000 68400
rect 44840 68008 45000 68128
rect 44840 67736 45000 67856
rect 44840 67464 45000 67584
rect 44840 67192 45000 67312
rect 44840 66920 45000 67040
rect 44840 66648 45000 66768
rect 44840 66376 45000 66496
rect 44840 66104 45000 66224
rect 44840 65832 45000 65952
rect 44840 65560 45000 65680
rect 44840 65288 45000 65408
rect 44840 65016 45000 65136
rect 44840 64744 45000 64864
rect 44840 64472 45000 64592
rect 44840 64200 45000 64320
rect 44840 63928 45000 64048
rect 44840 63656 45000 63776
rect 44840 63384 45000 63504
rect 44840 63112 45000 63232
rect 44840 62840 45000 62960
rect 44840 62568 45000 62688
rect 44840 62296 45000 62416
rect 44840 62024 45000 62144
rect 44840 61752 45000 61872
rect 44840 61480 45000 61600
rect 44840 61208 45000 61328
rect 44840 60936 45000 61056
rect 44840 60664 45000 60784
rect 44840 60392 45000 60512
rect 44840 60120 45000 60240
rect 44840 59848 45000 59968
rect 44840 59576 45000 59696
rect 44840 59304 45000 59424
rect 44840 59032 45000 59152
rect 44840 58760 45000 58880
rect 44840 58488 45000 58608
rect 44840 58216 45000 58336
rect 44840 57944 45000 58064
rect 44840 57672 45000 57792
rect 44840 57400 45000 57520
rect 44840 57128 45000 57248
rect 44840 56856 45000 56976
rect 44840 56584 45000 56704
rect 44840 56312 45000 56432
rect 44840 56040 45000 56160
rect 44840 55768 45000 55888
rect 44840 55496 45000 55616
rect 44840 55224 45000 55344
rect 44840 54952 45000 55072
rect 44840 54680 45000 54800
rect 44840 54408 45000 54528
rect 44840 54136 45000 54256
rect 44840 53864 45000 53984
rect 44840 53592 45000 53712
rect 44840 53320 45000 53440
rect 44840 53048 45000 53168
rect 44840 52776 45000 52896
rect 44840 52504 45000 52624
rect 44840 52232 45000 52352
rect 44840 51960 45000 52080
rect 44840 51688 45000 51808
rect 44840 51416 45000 51536
rect 44840 51144 45000 51264
rect 44840 50872 45000 50992
rect 44840 50600 45000 50720
rect 0 39176 160 39296
rect 0 38904 160 39024
rect 0 38632 160 38752
rect 0 38360 160 38480
rect 0 38088 160 38208
rect 0 37816 160 37936
rect 0 37544 160 37664
rect 0 37272 160 37392
rect 0 37000 160 37120
rect 0 36728 160 36848
rect 0 36456 160 36576
rect 0 36184 160 36304
rect 0 35912 160 36032
rect 0 35640 160 35760
rect 0 35368 160 35488
rect 0 35096 160 35216
rect 0 34824 160 34944
rect 0 34552 160 34672
rect 0 34280 160 34400
rect 0 34008 160 34128
rect 0 33736 160 33856
rect 0 33464 160 33584
rect 0 33192 160 33312
rect 0 32920 160 33040
rect 0 32648 160 32768
rect 0 32376 160 32496
rect 0 32104 160 32224
rect 0 31832 160 31952
rect 0 31560 160 31680
rect 0 31288 160 31408
rect 0 31016 160 31136
rect 0 30744 160 30864
rect 0 30472 160 30592
rect 0 30200 160 30320
rect 0 29928 160 30048
rect 0 29656 160 29776
rect 0 29384 160 29504
rect 0 29112 160 29232
rect 0 28840 160 28960
rect 0 28568 160 28688
rect 0 28296 160 28416
rect 0 28024 160 28144
rect 0 27752 160 27872
rect 0 27480 160 27600
rect 0 27208 160 27328
rect 0 26936 160 27056
rect 0 26664 160 26784
rect 0 26392 160 26512
rect 0 26120 160 26240
rect 0 25848 160 25968
rect 0 25576 160 25696
rect 0 25304 160 25424
rect 0 25032 160 25152
rect 0 24760 160 24880
rect 0 24488 160 24608
rect 0 24216 160 24336
rect 0 23944 160 24064
rect 0 23672 160 23792
rect 0 23400 160 23520
rect 0 23128 160 23248
rect 0 22856 160 22976
rect 0 22584 160 22704
rect 0 22312 160 22432
rect 0 22040 160 22160
rect 0 21768 160 21888
rect 0 21496 160 21616
rect 0 21224 160 21344
rect 0 20952 160 21072
rect 0 20680 160 20800
rect 0 20408 160 20528
rect 0 20136 160 20256
rect 0 19864 160 19984
rect 0 19592 160 19712
rect 0 19320 160 19440
rect 0 19048 160 19168
rect 0 18776 160 18896
rect 0 18504 160 18624
rect 0 18232 160 18352
rect 0 17960 160 18080
rect 0 17688 160 17808
rect 0 17416 160 17536
rect 0 17144 160 17264
rect 0 16872 160 16992
rect 0 16600 160 16720
rect 0 16328 160 16448
rect 0 16056 160 16176
rect 0 15784 160 15904
rect 0 15512 160 15632
rect 0 15240 160 15360
rect 0 14968 160 15088
rect 0 14696 160 14816
rect 0 14424 160 14544
rect 0 14152 160 14272
rect 0 13880 160 14000
rect 0 13608 160 13728
rect 0 13336 160 13456
rect 0 13064 160 13184
rect 0 12792 160 12912
rect 0 12520 160 12640
rect 0 12248 160 12368
rect 0 11976 160 12096
rect 0 11704 160 11824
rect 0 11432 160 11552
rect 0 11160 160 11280
rect 0 10888 160 11008
rect 0 10616 160 10736
rect 0 10344 160 10464
rect 0 10072 160 10192
rect 0 9800 160 9920
rect 0 9528 160 9648
rect 0 9256 160 9376
rect 0 8984 160 9104
rect 0 8712 160 8832
rect 0 8440 160 8560
rect 0 8168 160 8288
rect 0 7896 160 8016
rect 0 7624 160 7744
rect 0 7352 160 7472
rect 0 7080 160 7200
rect 0 6808 160 6928
rect 0 6536 160 6656
rect 0 6264 160 6384
rect 0 5992 160 6112
rect 0 5720 160 5840
rect 0 5448 160 5568
rect 0 5176 160 5296
rect 0 4904 160 5024
rect 0 4632 160 4752
rect 44840 39176 45000 39296
rect 44840 38904 45000 39024
rect 44840 38632 45000 38752
rect 44840 38360 45000 38480
rect 44840 38088 45000 38208
rect 44840 37816 45000 37936
rect 44840 37544 45000 37664
rect 44840 37272 45000 37392
rect 44840 37000 45000 37120
rect 44840 36728 45000 36848
rect 44840 36456 45000 36576
rect 44840 36184 45000 36304
rect 44840 35912 45000 36032
rect 44840 35640 45000 35760
rect 44840 35368 45000 35488
rect 44840 35096 45000 35216
rect 44840 34824 45000 34944
rect 44840 34552 45000 34672
rect 44840 34280 45000 34400
rect 44840 34008 45000 34128
rect 44840 33736 45000 33856
rect 44840 33464 45000 33584
rect 44840 33192 45000 33312
rect 44840 32920 45000 33040
rect 44840 32648 45000 32768
rect 44840 32376 45000 32496
rect 44840 32104 45000 32224
rect 44840 31832 45000 31952
rect 44840 31560 45000 31680
rect 44840 31288 45000 31408
rect 44840 31016 45000 31136
rect 44840 30744 45000 30864
rect 44840 30472 45000 30592
rect 44840 30200 45000 30320
rect 44840 29928 45000 30048
rect 44840 29656 45000 29776
rect 44840 29384 45000 29504
rect 44840 29112 45000 29232
rect 44840 28840 45000 28960
rect 44840 28568 45000 28688
rect 44840 28296 45000 28416
rect 44840 28024 45000 28144
rect 44840 27752 45000 27872
rect 44840 27480 45000 27600
rect 44840 27208 45000 27328
rect 44840 26936 45000 27056
rect 44840 26664 45000 26784
rect 44840 26392 45000 26512
rect 44840 26120 45000 26240
rect 44840 25848 45000 25968
rect 44840 25576 45000 25696
rect 44840 25304 45000 25424
rect 44840 25032 45000 25152
rect 44840 24760 45000 24880
rect 44840 24488 45000 24608
rect 44840 24216 45000 24336
rect 44840 23944 45000 24064
rect 44840 23672 45000 23792
rect 44840 23400 45000 23520
rect 44840 23128 45000 23248
rect 44840 22856 45000 22976
rect 44840 22584 45000 22704
rect 44840 22312 45000 22432
rect 44840 22040 45000 22160
rect 44840 21768 45000 21888
rect 44840 21496 45000 21616
rect 44840 21224 45000 21344
rect 44840 20952 45000 21072
rect 44840 20680 45000 20800
rect 44840 20408 45000 20528
rect 44840 20136 45000 20256
rect 44840 19864 45000 19984
rect 44840 19592 45000 19712
rect 44840 19320 45000 19440
rect 44840 19048 45000 19168
rect 44840 18776 45000 18896
rect 44840 18504 45000 18624
rect 44840 18232 45000 18352
rect 44840 17960 45000 18080
rect 44840 17688 45000 17808
rect 44840 17416 45000 17536
rect 44840 17144 45000 17264
rect 44840 16872 45000 16992
rect 44840 16600 45000 16720
rect 44840 16328 45000 16448
rect 44840 16056 45000 16176
rect 44840 15784 45000 15904
rect 44840 15512 45000 15632
rect 44840 15240 45000 15360
rect 44840 14968 45000 15088
rect 44840 14696 45000 14816
rect 44840 14424 45000 14544
rect 44840 14152 45000 14272
rect 44840 13880 45000 14000
rect 44840 13608 45000 13728
rect 44840 13336 45000 13456
rect 44840 13064 45000 13184
rect 44840 12792 45000 12912
rect 44840 12520 45000 12640
rect 44840 12248 45000 12368
rect 44840 11976 45000 12096
rect 44840 11704 45000 11824
rect 44840 11432 45000 11552
rect 44840 11160 45000 11280
rect 44840 10888 45000 11008
rect 44840 10616 45000 10736
rect 44840 10344 45000 10464
rect 44840 10072 45000 10192
rect 44840 9800 45000 9920
rect 44840 9528 45000 9648
rect 44840 9256 45000 9376
rect 44840 8984 45000 9104
rect 44840 8712 45000 8832
rect 44840 8440 45000 8560
rect 44840 8168 45000 8288
rect 44840 7896 45000 8016
rect 44840 7624 45000 7744
rect 44840 7352 45000 7472
rect 44840 7080 45000 7200
rect 44840 6808 45000 6928
rect 44840 6536 45000 6656
rect 44840 6264 45000 6384
rect 44840 5992 45000 6112
rect 44840 5720 45000 5840
rect 44840 5448 45000 5568
rect 44840 5176 45000 5296
rect 44840 4904 45000 5024
rect 44840 4632 45000 4752
<< obsm3 >>
rect 160 85344 44840 89453
rect 240 50520 44760 85344
rect 160 39376 44840 50520
rect 240 4552 44760 39376
rect 160 851 44840 4552
<< metal4 >>
rect 4208 1040 4528 89264
rect 19568 1040 19888 89264
rect 34928 1040 35248 89264
<< obsm4 >>
rect 795 89344 42629 89453
rect 795 960 4128 89344
rect 4608 960 19488 89344
rect 19968 960 34848 89344
rect 35328 960 42629 89344
rect 795 851 42629 960
<< labels >>
rlabel metal3 s 44840 63656 45000 63776 6 Tile_X0Y0_E1BEG[0]
port 1 nsew signal output
rlabel metal3 s 44840 63928 45000 64048 6 Tile_X0Y0_E1BEG[1]
port 2 nsew signal output
rlabel metal3 s 44840 64200 45000 64320 6 Tile_X0Y0_E1BEG[2]
port 3 nsew signal output
rlabel metal3 s 44840 64472 45000 64592 6 Tile_X0Y0_E1BEG[3]
port 4 nsew signal output
rlabel metal3 s 0 63656 160 63776 6 Tile_X0Y0_E1END[0]
port 5 nsew signal input
rlabel metal3 s 0 63928 160 64048 6 Tile_X0Y0_E1END[1]
port 6 nsew signal input
rlabel metal3 s 0 64200 160 64320 6 Tile_X0Y0_E1END[2]
port 7 nsew signal input
rlabel metal3 s 0 64472 160 64592 6 Tile_X0Y0_E1END[3]
port 8 nsew signal input
rlabel metal3 s 44840 64744 45000 64864 6 Tile_X0Y0_E2BEG[0]
port 9 nsew signal output
rlabel metal3 s 44840 65016 45000 65136 6 Tile_X0Y0_E2BEG[1]
port 10 nsew signal output
rlabel metal3 s 44840 65288 45000 65408 6 Tile_X0Y0_E2BEG[2]
port 11 nsew signal output
rlabel metal3 s 44840 65560 45000 65680 6 Tile_X0Y0_E2BEG[3]
port 12 nsew signal output
rlabel metal3 s 44840 65832 45000 65952 6 Tile_X0Y0_E2BEG[4]
port 13 nsew signal output
rlabel metal3 s 44840 66104 45000 66224 6 Tile_X0Y0_E2BEG[5]
port 14 nsew signal output
rlabel metal3 s 44840 66376 45000 66496 6 Tile_X0Y0_E2BEG[6]
port 15 nsew signal output
rlabel metal3 s 44840 66648 45000 66768 6 Tile_X0Y0_E2BEG[7]
port 16 nsew signal output
rlabel metal3 s 44840 66920 45000 67040 6 Tile_X0Y0_E2BEGb[0]
port 17 nsew signal output
rlabel metal3 s 44840 67192 45000 67312 6 Tile_X0Y0_E2BEGb[1]
port 18 nsew signal output
rlabel metal3 s 44840 67464 45000 67584 6 Tile_X0Y0_E2BEGb[2]
port 19 nsew signal output
rlabel metal3 s 44840 67736 45000 67856 6 Tile_X0Y0_E2BEGb[3]
port 20 nsew signal output
rlabel metal3 s 44840 68008 45000 68128 6 Tile_X0Y0_E2BEGb[4]
port 21 nsew signal output
rlabel metal3 s 44840 68280 45000 68400 6 Tile_X0Y0_E2BEGb[5]
port 22 nsew signal output
rlabel metal3 s 44840 68552 45000 68672 6 Tile_X0Y0_E2BEGb[6]
port 23 nsew signal output
rlabel metal3 s 44840 68824 45000 68944 6 Tile_X0Y0_E2BEGb[7]
port 24 nsew signal output
rlabel metal3 s 0 66920 160 67040 6 Tile_X0Y0_E2END[0]
port 25 nsew signal input
rlabel metal3 s 0 67192 160 67312 6 Tile_X0Y0_E2END[1]
port 26 nsew signal input
rlabel metal3 s 0 67464 160 67584 6 Tile_X0Y0_E2END[2]
port 27 nsew signal input
rlabel metal3 s 0 67736 160 67856 6 Tile_X0Y0_E2END[3]
port 28 nsew signal input
rlabel metal3 s 0 68008 160 68128 6 Tile_X0Y0_E2END[4]
port 29 nsew signal input
rlabel metal3 s 0 68280 160 68400 6 Tile_X0Y0_E2END[5]
port 30 nsew signal input
rlabel metal3 s 0 68552 160 68672 6 Tile_X0Y0_E2END[6]
port 31 nsew signal input
rlabel metal3 s 0 68824 160 68944 6 Tile_X0Y0_E2END[7]
port 32 nsew signal input
rlabel metal3 s 0 64744 160 64864 6 Tile_X0Y0_E2MID[0]
port 33 nsew signal input
rlabel metal3 s 0 65016 160 65136 6 Tile_X0Y0_E2MID[1]
port 34 nsew signal input
rlabel metal3 s 0 65288 160 65408 6 Tile_X0Y0_E2MID[2]
port 35 nsew signal input
rlabel metal3 s 0 65560 160 65680 6 Tile_X0Y0_E2MID[3]
port 36 nsew signal input
rlabel metal3 s 0 65832 160 65952 6 Tile_X0Y0_E2MID[4]
port 37 nsew signal input
rlabel metal3 s 0 66104 160 66224 6 Tile_X0Y0_E2MID[5]
port 38 nsew signal input
rlabel metal3 s 0 66376 160 66496 6 Tile_X0Y0_E2MID[6]
port 39 nsew signal input
rlabel metal3 s 0 66648 160 66768 6 Tile_X0Y0_E2MID[7]
port 40 nsew signal input
rlabel metal3 s 44840 73448 45000 73568 6 Tile_X0Y0_E6BEG[0]
port 41 nsew signal output
rlabel metal3 s 44840 76168 45000 76288 6 Tile_X0Y0_E6BEG[10]
port 42 nsew signal output
rlabel metal3 s 44840 76440 45000 76560 6 Tile_X0Y0_E6BEG[11]
port 43 nsew signal output
rlabel metal3 s 44840 73720 45000 73840 6 Tile_X0Y0_E6BEG[1]
port 44 nsew signal output
rlabel metal3 s 44840 73992 45000 74112 6 Tile_X0Y0_E6BEG[2]
port 45 nsew signal output
rlabel metal3 s 44840 74264 45000 74384 6 Tile_X0Y0_E6BEG[3]
port 46 nsew signal output
rlabel metal3 s 44840 74536 45000 74656 6 Tile_X0Y0_E6BEG[4]
port 47 nsew signal output
rlabel metal3 s 44840 74808 45000 74928 6 Tile_X0Y0_E6BEG[5]
port 48 nsew signal output
rlabel metal3 s 44840 75080 45000 75200 6 Tile_X0Y0_E6BEG[6]
port 49 nsew signal output
rlabel metal3 s 44840 75352 45000 75472 6 Tile_X0Y0_E6BEG[7]
port 50 nsew signal output
rlabel metal3 s 44840 75624 45000 75744 6 Tile_X0Y0_E6BEG[8]
port 51 nsew signal output
rlabel metal3 s 44840 75896 45000 76016 6 Tile_X0Y0_E6BEG[9]
port 52 nsew signal output
rlabel metal3 s 0 73448 160 73568 6 Tile_X0Y0_E6END[0]
port 53 nsew signal input
rlabel metal3 s 0 76168 160 76288 6 Tile_X0Y0_E6END[10]
port 54 nsew signal input
rlabel metal3 s 0 76440 160 76560 6 Tile_X0Y0_E6END[11]
port 55 nsew signal input
rlabel metal3 s 0 73720 160 73840 6 Tile_X0Y0_E6END[1]
port 56 nsew signal input
rlabel metal3 s 0 73992 160 74112 6 Tile_X0Y0_E6END[2]
port 57 nsew signal input
rlabel metal3 s 0 74264 160 74384 6 Tile_X0Y0_E6END[3]
port 58 nsew signal input
rlabel metal3 s 0 74536 160 74656 6 Tile_X0Y0_E6END[4]
port 59 nsew signal input
rlabel metal3 s 0 74808 160 74928 6 Tile_X0Y0_E6END[5]
port 60 nsew signal input
rlabel metal3 s 0 75080 160 75200 6 Tile_X0Y0_E6END[6]
port 61 nsew signal input
rlabel metal3 s 0 75352 160 75472 6 Tile_X0Y0_E6END[7]
port 62 nsew signal input
rlabel metal3 s 0 75624 160 75744 6 Tile_X0Y0_E6END[8]
port 63 nsew signal input
rlabel metal3 s 0 75896 160 76016 6 Tile_X0Y0_E6END[9]
port 64 nsew signal input
rlabel metal3 s 44840 69096 45000 69216 6 Tile_X0Y0_EE4BEG[0]
port 65 nsew signal output
rlabel metal3 s 44840 71816 45000 71936 6 Tile_X0Y0_EE4BEG[10]
port 66 nsew signal output
rlabel metal3 s 44840 72088 45000 72208 6 Tile_X0Y0_EE4BEG[11]
port 67 nsew signal output
rlabel metal3 s 44840 72360 45000 72480 6 Tile_X0Y0_EE4BEG[12]
port 68 nsew signal output
rlabel metal3 s 44840 72632 45000 72752 6 Tile_X0Y0_EE4BEG[13]
port 69 nsew signal output
rlabel metal3 s 44840 72904 45000 73024 6 Tile_X0Y0_EE4BEG[14]
port 70 nsew signal output
rlabel metal3 s 44840 73176 45000 73296 6 Tile_X0Y0_EE4BEG[15]
port 71 nsew signal output
rlabel metal3 s 44840 69368 45000 69488 6 Tile_X0Y0_EE4BEG[1]
port 72 nsew signal output
rlabel metal3 s 44840 69640 45000 69760 6 Tile_X0Y0_EE4BEG[2]
port 73 nsew signal output
rlabel metal3 s 44840 69912 45000 70032 6 Tile_X0Y0_EE4BEG[3]
port 74 nsew signal output
rlabel metal3 s 44840 70184 45000 70304 6 Tile_X0Y0_EE4BEG[4]
port 75 nsew signal output
rlabel metal3 s 44840 70456 45000 70576 6 Tile_X0Y0_EE4BEG[5]
port 76 nsew signal output
rlabel metal3 s 44840 70728 45000 70848 6 Tile_X0Y0_EE4BEG[6]
port 77 nsew signal output
rlabel metal3 s 44840 71000 45000 71120 6 Tile_X0Y0_EE4BEG[7]
port 78 nsew signal output
rlabel metal3 s 44840 71272 45000 71392 6 Tile_X0Y0_EE4BEG[8]
port 79 nsew signal output
rlabel metal3 s 44840 71544 45000 71664 6 Tile_X0Y0_EE4BEG[9]
port 80 nsew signal output
rlabel metal3 s 0 69096 160 69216 6 Tile_X0Y0_EE4END[0]
port 81 nsew signal input
rlabel metal3 s 0 71816 160 71936 6 Tile_X0Y0_EE4END[10]
port 82 nsew signal input
rlabel metal3 s 0 72088 160 72208 6 Tile_X0Y0_EE4END[11]
port 83 nsew signal input
rlabel metal3 s 0 72360 160 72480 6 Tile_X0Y0_EE4END[12]
port 84 nsew signal input
rlabel metal3 s 0 72632 160 72752 6 Tile_X0Y0_EE4END[13]
port 85 nsew signal input
rlabel metal3 s 0 72904 160 73024 6 Tile_X0Y0_EE4END[14]
port 86 nsew signal input
rlabel metal3 s 0 73176 160 73296 6 Tile_X0Y0_EE4END[15]
port 87 nsew signal input
rlabel metal3 s 0 69368 160 69488 6 Tile_X0Y0_EE4END[1]
port 88 nsew signal input
rlabel metal3 s 0 69640 160 69760 6 Tile_X0Y0_EE4END[2]
port 89 nsew signal input
rlabel metal3 s 0 69912 160 70032 6 Tile_X0Y0_EE4END[3]
port 90 nsew signal input
rlabel metal3 s 0 70184 160 70304 6 Tile_X0Y0_EE4END[4]
port 91 nsew signal input
rlabel metal3 s 0 70456 160 70576 6 Tile_X0Y0_EE4END[5]
port 92 nsew signal input
rlabel metal3 s 0 70728 160 70848 6 Tile_X0Y0_EE4END[6]
port 93 nsew signal input
rlabel metal3 s 0 71000 160 71120 6 Tile_X0Y0_EE4END[7]
port 94 nsew signal input
rlabel metal3 s 0 71272 160 71392 6 Tile_X0Y0_EE4END[8]
port 95 nsew signal input
rlabel metal3 s 0 71544 160 71664 6 Tile_X0Y0_EE4END[9]
port 96 nsew signal input
rlabel metal3 s 0 76712 160 76832 6 Tile_X0Y0_FrameData[0]
port 97 nsew signal input
rlabel metal3 s 0 79432 160 79552 6 Tile_X0Y0_FrameData[10]
port 98 nsew signal input
rlabel metal3 s 0 79704 160 79824 6 Tile_X0Y0_FrameData[11]
port 99 nsew signal input
rlabel metal3 s 0 79976 160 80096 6 Tile_X0Y0_FrameData[12]
port 100 nsew signal input
rlabel metal3 s 0 80248 160 80368 6 Tile_X0Y0_FrameData[13]
port 101 nsew signal input
rlabel metal3 s 0 80520 160 80640 6 Tile_X0Y0_FrameData[14]
port 102 nsew signal input
rlabel metal3 s 0 80792 160 80912 6 Tile_X0Y0_FrameData[15]
port 103 nsew signal input
rlabel metal3 s 0 81064 160 81184 6 Tile_X0Y0_FrameData[16]
port 104 nsew signal input
rlabel metal3 s 0 81336 160 81456 6 Tile_X0Y0_FrameData[17]
port 105 nsew signal input
rlabel metal3 s 0 81608 160 81728 6 Tile_X0Y0_FrameData[18]
port 106 nsew signal input
rlabel metal3 s 0 81880 160 82000 6 Tile_X0Y0_FrameData[19]
port 107 nsew signal input
rlabel metal3 s 0 76984 160 77104 6 Tile_X0Y0_FrameData[1]
port 108 nsew signal input
rlabel metal3 s 0 82152 160 82272 6 Tile_X0Y0_FrameData[20]
port 109 nsew signal input
rlabel metal3 s 0 82424 160 82544 6 Tile_X0Y0_FrameData[21]
port 110 nsew signal input
rlabel metal3 s 0 82696 160 82816 6 Tile_X0Y0_FrameData[22]
port 111 nsew signal input
rlabel metal3 s 0 82968 160 83088 6 Tile_X0Y0_FrameData[23]
port 112 nsew signal input
rlabel metal3 s 0 83240 160 83360 6 Tile_X0Y0_FrameData[24]
port 113 nsew signal input
rlabel metal3 s 0 83512 160 83632 6 Tile_X0Y0_FrameData[25]
port 114 nsew signal input
rlabel metal3 s 0 83784 160 83904 6 Tile_X0Y0_FrameData[26]
port 115 nsew signal input
rlabel metal3 s 0 84056 160 84176 6 Tile_X0Y0_FrameData[27]
port 116 nsew signal input
rlabel metal3 s 0 84328 160 84448 6 Tile_X0Y0_FrameData[28]
port 117 nsew signal input
rlabel metal3 s 0 84600 160 84720 6 Tile_X0Y0_FrameData[29]
port 118 nsew signal input
rlabel metal3 s 0 77256 160 77376 6 Tile_X0Y0_FrameData[2]
port 119 nsew signal input
rlabel metal3 s 0 84872 160 84992 6 Tile_X0Y0_FrameData[30]
port 120 nsew signal input
rlabel metal3 s 0 85144 160 85264 6 Tile_X0Y0_FrameData[31]
port 121 nsew signal input
rlabel metal3 s 0 77528 160 77648 6 Tile_X0Y0_FrameData[3]
port 122 nsew signal input
rlabel metal3 s 0 77800 160 77920 6 Tile_X0Y0_FrameData[4]
port 123 nsew signal input
rlabel metal3 s 0 78072 160 78192 6 Tile_X0Y0_FrameData[5]
port 124 nsew signal input
rlabel metal3 s 0 78344 160 78464 6 Tile_X0Y0_FrameData[6]
port 125 nsew signal input
rlabel metal3 s 0 78616 160 78736 6 Tile_X0Y0_FrameData[7]
port 126 nsew signal input
rlabel metal3 s 0 78888 160 79008 6 Tile_X0Y0_FrameData[8]
port 127 nsew signal input
rlabel metal3 s 0 79160 160 79280 6 Tile_X0Y0_FrameData[9]
port 128 nsew signal input
rlabel metal3 s 44840 76712 45000 76832 6 Tile_X0Y0_FrameData_O[0]
port 129 nsew signal output
rlabel metal3 s 44840 79432 45000 79552 6 Tile_X0Y0_FrameData_O[10]
port 130 nsew signal output
rlabel metal3 s 44840 79704 45000 79824 6 Tile_X0Y0_FrameData_O[11]
port 131 nsew signal output
rlabel metal3 s 44840 79976 45000 80096 6 Tile_X0Y0_FrameData_O[12]
port 132 nsew signal output
rlabel metal3 s 44840 80248 45000 80368 6 Tile_X0Y0_FrameData_O[13]
port 133 nsew signal output
rlabel metal3 s 44840 80520 45000 80640 6 Tile_X0Y0_FrameData_O[14]
port 134 nsew signal output
rlabel metal3 s 44840 80792 45000 80912 6 Tile_X0Y0_FrameData_O[15]
port 135 nsew signal output
rlabel metal3 s 44840 81064 45000 81184 6 Tile_X0Y0_FrameData_O[16]
port 136 nsew signal output
rlabel metal3 s 44840 81336 45000 81456 6 Tile_X0Y0_FrameData_O[17]
port 137 nsew signal output
rlabel metal3 s 44840 81608 45000 81728 6 Tile_X0Y0_FrameData_O[18]
port 138 nsew signal output
rlabel metal3 s 44840 81880 45000 82000 6 Tile_X0Y0_FrameData_O[19]
port 139 nsew signal output
rlabel metal3 s 44840 76984 45000 77104 6 Tile_X0Y0_FrameData_O[1]
port 140 nsew signal output
rlabel metal3 s 44840 82152 45000 82272 6 Tile_X0Y0_FrameData_O[20]
port 141 nsew signal output
rlabel metal3 s 44840 82424 45000 82544 6 Tile_X0Y0_FrameData_O[21]
port 142 nsew signal output
rlabel metal3 s 44840 82696 45000 82816 6 Tile_X0Y0_FrameData_O[22]
port 143 nsew signal output
rlabel metal3 s 44840 82968 45000 83088 6 Tile_X0Y0_FrameData_O[23]
port 144 nsew signal output
rlabel metal3 s 44840 83240 45000 83360 6 Tile_X0Y0_FrameData_O[24]
port 145 nsew signal output
rlabel metal3 s 44840 83512 45000 83632 6 Tile_X0Y0_FrameData_O[25]
port 146 nsew signal output
rlabel metal3 s 44840 83784 45000 83904 6 Tile_X0Y0_FrameData_O[26]
port 147 nsew signal output
rlabel metal3 s 44840 84056 45000 84176 6 Tile_X0Y0_FrameData_O[27]
port 148 nsew signal output
rlabel metal3 s 44840 84328 45000 84448 6 Tile_X0Y0_FrameData_O[28]
port 149 nsew signal output
rlabel metal3 s 44840 84600 45000 84720 6 Tile_X0Y0_FrameData_O[29]
port 150 nsew signal output
rlabel metal3 s 44840 77256 45000 77376 6 Tile_X0Y0_FrameData_O[2]
port 151 nsew signal output
rlabel metal3 s 44840 84872 45000 84992 6 Tile_X0Y0_FrameData_O[30]
port 152 nsew signal output
rlabel metal3 s 44840 85144 45000 85264 6 Tile_X0Y0_FrameData_O[31]
port 153 nsew signal output
rlabel metal3 s 44840 77528 45000 77648 6 Tile_X0Y0_FrameData_O[3]
port 154 nsew signal output
rlabel metal3 s 44840 77800 45000 77920 6 Tile_X0Y0_FrameData_O[4]
port 155 nsew signal output
rlabel metal3 s 44840 78072 45000 78192 6 Tile_X0Y0_FrameData_O[5]
port 156 nsew signal output
rlabel metal3 s 44840 78344 45000 78464 6 Tile_X0Y0_FrameData_O[6]
port 157 nsew signal output
rlabel metal3 s 44840 78616 45000 78736 6 Tile_X0Y0_FrameData_O[7]
port 158 nsew signal output
rlabel metal3 s 44840 78888 45000 79008 6 Tile_X0Y0_FrameData_O[8]
port 159 nsew signal output
rlabel metal3 s 44840 79160 45000 79280 6 Tile_X0Y0_FrameData_O[9]
port 160 nsew signal output
rlabel metal2 s 34334 90640 34390 90800 6 Tile_X0Y0_FrameStrobe_O[0]
port 161 nsew signal output
rlabel metal2 s 37094 90640 37150 90800 6 Tile_X0Y0_FrameStrobe_O[10]
port 162 nsew signal output
rlabel metal2 s 37370 90640 37426 90800 6 Tile_X0Y0_FrameStrobe_O[11]
port 163 nsew signal output
rlabel metal2 s 37646 90640 37702 90800 6 Tile_X0Y0_FrameStrobe_O[12]
port 164 nsew signal output
rlabel metal2 s 37922 90640 37978 90800 6 Tile_X0Y0_FrameStrobe_O[13]
port 165 nsew signal output
rlabel metal2 s 38198 90640 38254 90800 6 Tile_X0Y0_FrameStrobe_O[14]
port 166 nsew signal output
rlabel metal2 s 38474 90640 38530 90800 6 Tile_X0Y0_FrameStrobe_O[15]
port 167 nsew signal output
rlabel metal2 s 38750 90640 38806 90800 6 Tile_X0Y0_FrameStrobe_O[16]
port 168 nsew signal output
rlabel metal2 s 39026 90640 39082 90800 6 Tile_X0Y0_FrameStrobe_O[17]
port 169 nsew signal output
rlabel metal2 s 39302 90640 39358 90800 6 Tile_X0Y0_FrameStrobe_O[18]
port 170 nsew signal output
rlabel metal2 s 39578 90640 39634 90800 6 Tile_X0Y0_FrameStrobe_O[19]
port 171 nsew signal output
rlabel metal2 s 34610 90640 34666 90800 6 Tile_X0Y0_FrameStrobe_O[1]
port 172 nsew signal output
rlabel metal2 s 34886 90640 34942 90800 6 Tile_X0Y0_FrameStrobe_O[2]
port 173 nsew signal output
rlabel metal2 s 35162 90640 35218 90800 6 Tile_X0Y0_FrameStrobe_O[3]
port 174 nsew signal output
rlabel metal2 s 35438 90640 35494 90800 6 Tile_X0Y0_FrameStrobe_O[4]
port 175 nsew signal output
rlabel metal2 s 35714 90640 35770 90800 6 Tile_X0Y0_FrameStrobe_O[5]
port 176 nsew signal output
rlabel metal2 s 35990 90640 36046 90800 6 Tile_X0Y0_FrameStrobe_O[6]
port 177 nsew signal output
rlabel metal2 s 36266 90640 36322 90800 6 Tile_X0Y0_FrameStrobe_O[7]
port 178 nsew signal output
rlabel metal2 s 36542 90640 36598 90800 6 Tile_X0Y0_FrameStrobe_O[8]
port 179 nsew signal output
rlabel metal2 s 36818 90640 36874 90800 6 Tile_X0Y0_FrameStrobe_O[9]
port 180 nsew signal output
rlabel metal2 s 5354 90640 5410 90800 6 Tile_X0Y0_N1BEG[0]
port 181 nsew signal output
rlabel metal2 s 5630 90640 5686 90800 6 Tile_X0Y0_N1BEG[1]
port 182 nsew signal output
rlabel metal2 s 5906 90640 5962 90800 6 Tile_X0Y0_N1BEG[2]
port 183 nsew signal output
rlabel metal2 s 6182 90640 6238 90800 6 Tile_X0Y0_N1BEG[3]
port 184 nsew signal output
rlabel metal2 s 6458 90640 6514 90800 6 Tile_X0Y0_N2BEG[0]
port 185 nsew signal output
rlabel metal2 s 6734 90640 6790 90800 6 Tile_X0Y0_N2BEG[1]
port 186 nsew signal output
rlabel metal2 s 7010 90640 7066 90800 6 Tile_X0Y0_N2BEG[2]
port 187 nsew signal output
rlabel metal2 s 7286 90640 7342 90800 6 Tile_X0Y0_N2BEG[3]
port 188 nsew signal output
rlabel metal2 s 7562 90640 7618 90800 6 Tile_X0Y0_N2BEG[4]
port 189 nsew signal output
rlabel metal2 s 7838 90640 7894 90800 6 Tile_X0Y0_N2BEG[5]
port 190 nsew signal output
rlabel metal2 s 8114 90640 8170 90800 6 Tile_X0Y0_N2BEG[6]
port 191 nsew signal output
rlabel metal2 s 8390 90640 8446 90800 6 Tile_X0Y0_N2BEG[7]
port 192 nsew signal output
rlabel metal2 s 8666 90640 8722 90800 6 Tile_X0Y0_N2BEGb[0]
port 193 nsew signal output
rlabel metal2 s 8942 90640 8998 90800 6 Tile_X0Y0_N2BEGb[1]
port 194 nsew signal output
rlabel metal2 s 9218 90640 9274 90800 6 Tile_X0Y0_N2BEGb[2]
port 195 nsew signal output
rlabel metal2 s 9494 90640 9550 90800 6 Tile_X0Y0_N2BEGb[3]
port 196 nsew signal output
rlabel metal2 s 9770 90640 9826 90800 6 Tile_X0Y0_N2BEGb[4]
port 197 nsew signal output
rlabel metal2 s 10046 90640 10102 90800 6 Tile_X0Y0_N2BEGb[5]
port 198 nsew signal output
rlabel metal2 s 10322 90640 10378 90800 6 Tile_X0Y0_N2BEGb[6]
port 199 nsew signal output
rlabel metal2 s 10598 90640 10654 90800 6 Tile_X0Y0_N2BEGb[7]
port 200 nsew signal output
rlabel metal2 s 10874 90640 10930 90800 6 Tile_X0Y0_N4BEG[0]
port 201 nsew signal output
rlabel metal2 s 13634 90640 13690 90800 6 Tile_X0Y0_N4BEG[10]
port 202 nsew signal output
rlabel metal2 s 13910 90640 13966 90800 6 Tile_X0Y0_N4BEG[11]
port 203 nsew signal output
rlabel metal2 s 14186 90640 14242 90800 6 Tile_X0Y0_N4BEG[12]
port 204 nsew signal output
rlabel metal2 s 14462 90640 14518 90800 6 Tile_X0Y0_N4BEG[13]
port 205 nsew signal output
rlabel metal2 s 14738 90640 14794 90800 6 Tile_X0Y0_N4BEG[14]
port 206 nsew signal output
rlabel metal2 s 15014 90640 15070 90800 6 Tile_X0Y0_N4BEG[15]
port 207 nsew signal output
rlabel metal2 s 11150 90640 11206 90800 6 Tile_X0Y0_N4BEG[1]
port 208 nsew signal output
rlabel metal2 s 11426 90640 11482 90800 6 Tile_X0Y0_N4BEG[2]
port 209 nsew signal output
rlabel metal2 s 11702 90640 11758 90800 6 Tile_X0Y0_N4BEG[3]
port 210 nsew signal output
rlabel metal2 s 11978 90640 12034 90800 6 Tile_X0Y0_N4BEG[4]
port 211 nsew signal output
rlabel metal2 s 12254 90640 12310 90800 6 Tile_X0Y0_N4BEG[5]
port 212 nsew signal output
rlabel metal2 s 12530 90640 12586 90800 6 Tile_X0Y0_N4BEG[6]
port 213 nsew signal output
rlabel metal2 s 12806 90640 12862 90800 6 Tile_X0Y0_N4BEG[7]
port 214 nsew signal output
rlabel metal2 s 13082 90640 13138 90800 6 Tile_X0Y0_N4BEG[8]
port 215 nsew signal output
rlabel metal2 s 13358 90640 13414 90800 6 Tile_X0Y0_N4BEG[9]
port 216 nsew signal output
rlabel metal2 s 15290 90640 15346 90800 6 Tile_X0Y0_NN4BEG[0]
port 217 nsew signal output
rlabel metal2 s 18050 90640 18106 90800 6 Tile_X0Y0_NN4BEG[10]
port 218 nsew signal output
rlabel metal2 s 18326 90640 18382 90800 6 Tile_X0Y0_NN4BEG[11]
port 219 nsew signal output
rlabel metal2 s 18602 90640 18658 90800 6 Tile_X0Y0_NN4BEG[12]
port 220 nsew signal output
rlabel metal2 s 18878 90640 18934 90800 6 Tile_X0Y0_NN4BEG[13]
port 221 nsew signal output
rlabel metal2 s 19154 90640 19210 90800 6 Tile_X0Y0_NN4BEG[14]
port 222 nsew signal output
rlabel metal2 s 19430 90640 19486 90800 6 Tile_X0Y0_NN4BEG[15]
port 223 nsew signal output
rlabel metal2 s 15566 90640 15622 90800 6 Tile_X0Y0_NN4BEG[1]
port 224 nsew signal output
rlabel metal2 s 15842 90640 15898 90800 6 Tile_X0Y0_NN4BEG[2]
port 225 nsew signal output
rlabel metal2 s 16118 90640 16174 90800 6 Tile_X0Y0_NN4BEG[3]
port 226 nsew signal output
rlabel metal2 s 16394 90640 16450 90800 6 Tile_X0Y0_NN4BEG[4]
port 227 nsew signal output
rlabel metal2 s 16670 90640 16726 90800 6 Tile_X0Y0_NN4BEG[5]
port 228 nsew signal output
rlabel metal2 s 16946 90640 17002 90800 6 Tile_X0Y0_NN4BEG[6]
port 229 nsew signal output
rlabel metal2 s 17222 90640 17278 90800 6 Tile_X0Y0_NN4BEG[7]
port 230 nsew signal output
rlabel metal2 s 17498 90640 17554 90800 6 Tile_X0Y0_NN4BEG[8]
port 231 nsew signal output
rlabel metal2 s 17774 90640 17830 90800 6 Tile_X0Y0_NN4BEG[9]
port 232 nsew signal output
rlabel metal2 s 19706 90640 19762 90800 6 Tile_X0Y0_S1END[0]
port 233 nsew signal input
rlabel metal2 s 19982 90640 20038 90800 6 Tile_X0Y0_S1END[1]
port 234 nsew signal input
rlabel metal2 s 20258 90640 20314 90800 6 Tile_X0Y0_S1END[2]
port 235 nsew signal input
rlabel metal2 s 20534 90640 20590 90800 6 Tile_X0Y0_S1END[3]
port 236 nsew signal input
rlabel metal2 s 20810 90640 20866 90800 6 Tile_X0Y0_S2END[0]
port 237 nsew signal input
rlabel metal2 s 21086 90640 21142 90800 6 Tile_X0Y0_S2END[1]
port 238 nsew signal input
rlabel metal2 s 21362 90640 21418 90800 6 Tile_X0Y0_S2END[2]
port 239 nsew signal input
rlabel metal2 s 21638 90640 21694 90800 6 Tile_X0Y0_S2END[3]
port 240 nsew signal input
rlabel metal2 s 21914 90640 21970 90800 6 Tile_X0Y0_S2END[4]
port 241 nsew signal input
rlabel metal2 s 22190 90640 22246 90800 6 Tile_X0Y0_S2END[5]
port 242 nsew signal input
rlabel metal2 s 22466 90640 22522 90800 6 Tile_X0Y0_S2END[6]
port 243 nsew signal input
rlabel metal2 s 22742 90640 22798 90800 6 Tile_X0Y0_S2END[7]
port 244 nsew signal input
rlabel metal2 s 23018 90640 23074 90800 6 Tile_X0Y0_S2MID[0]
port 245 nsew signal input
rlabel metal2 s 23294 90640 23350 90800 6 Tile_X0Y0_S2MID[1]
port 246 nsew signal input
rlabel metal2 s 23570 90640 23626 90800 6 Tile_X0Y0_S2MID[2]
port 247 nsew signal input
rlabel metal2 s 23846 90640 23902 90800 6 Tile_X0Y0_S2MID[3]
port 248 nsew signal input
rlabel metal2 s 24122 90640 24178 90800 6 Tile_X0Y0_S2MID[4]
port 249 nsew signal input
rlabel metal2 s 24398 90640 24454 90800 6 Tile_X0Y0_S2MID[5]
port 250 nsew signal input
rlabel metal2 s 24674 90640 24730 90800 6 Tile_X0Y0_S2MID[6]
port 251 nsew signal input
rlabel metal2 s 24950 90640 25006 90800 6 Tile_X0Y0_S2MID[7]
port 252 nsew signal input
rlabel metal2 s 25226 90640 25282 90800 6 Tile_X0Y0_S4END[0]
port 253 nsew signal input
rlabel metal2 s 27986 90640 28042 90800 6 Tile_X0Y0_S4END[10]
port 254 nsew signal input
rlabel metal2 s 28262 90640 28318 90800 6 Tile_X0Y0_S4END[11]
port 255 nsew signal input
rlabel metal2 s 28538 90640 28594 90800 6 Tile_X0Y0_S4END[12]
port 256 nsew signal input
rlabel metal2 s 28814 90640 28870 90800 6 Tile_X0Y0_S4END[13]
port 257 nsew signal input
rlabel metal2 s 29090 90640 29146 90800 6 Tile_X0Y0_S4END[14]
port 258 nsew signal input
rlabel metal2 s 29366 90640 29422 90800 6 Tile_X0Y0_S4END[15]
port 259 nsew signal input
rlabel metal2 s 25502 90640 25558 90800 6 Tile_X0Y0_S4END[1]
port 260 nsew signal input
rlabel metal2 s 25778 90640 25834 90800 6 Tile_X0Y0_S4END[2]
port 261 nsew signal input
rlabel metal2 s 26054 90640 26110 90800 6 Tile_X0Y0_S4END[3]
port 262 nsew signal input
rlabel metal2 s 26330 90640 26386 90800 6 Tile_X0Y0_S4END[4]
port 263 nsew signal input
rlabel metal2 s 26606 90640 26662 90800 6 Tile_X0Y0_S4END[5]
port 264 nsew signal input
rlabel metal2 s 26882 90640 26938 90800 6 Tile_X0Y0_S4END[6]
port 265 nsew signal input
rlabel metal2 s 27158 90640 27214 90800 6 Tile_X0Y0_S4END[7]
port 266 nsew signal input
rlabel metal2 s 27434 90640 27490 90800 6 Tile_X0Y0_S4END[8]
port 267 nsew signal input
rlabel metal2 s 27710 90640 27766 90800 6 Tile_X0Y0_S4END[9]
port 268 nsew signal input
rlabel metal2 s 29642 90640 29698 90800 6 Tile_X0Y0_SS4END[0]
port 269 nsew signal input
rlabel metal2 s 32402 90640 32458 90800 6 Tile_X0Y0_SS4END[10]
port 270 nsew signal input
rlabel metal2 s 32678 90640 32734 90800 6 Tile_X0Y0_SS4END[11]
port 271 nsew signal input
rlabel metal2 s 32954 90640 33010 90800 6 Tile_X0Y0_SS4END[12]
port 272 nsew signal input
rlabel metal2 s 33230 90640 33286 90800 6 Tile_X0Y0_SS4END[13]
port 273 nsew signal input
rlabel metal2 s 33506 90640 33562 90800 6 Tile_X0Y0_SS4END[14]
port 274 nsew signal input
rlabel metal2 s 33782 90640 33838 90800 6 Tile_X0Y0_SS4END[15]
port 275 nsew signal input
rlabel metal2 s 29918 90640 29974 90800 6 Tile_X0Y0_SS4END[1]
port 276 nsew signal input
rlabel metal2 s 30194 90640 30250 90800 6 Tile_X0Y0_SS4END[2]
port 277 nsew signal input
rlabel metal2 s 30470 90640 30526 90800 6 Tile_X0Y0_SS4END[3]
port 278 nsew signal input
rlabel metal2 s 30746 90640 30802 90800 6 Tile_X0Y0_SS4END[4]
port 279 nsew signal input
rlabel metal2 s 31022 90640 31078 90800 6 Tile_X0Y0_SS4END[5]
port 280 nsew signal input
rlabel metal2 s 31298 90640 31354 90800 6 Tile_X0Y0_SS4END[6]
port 281 nsew signal input
rlabel metal2 s 31574 90640 31630 90800 6 Tile_X0Y0_SS4END[7]
port 282 nsew signal input
rlabel metal2 s 31850 90640 31906 90800 6 Tile_X0Y0_SS4END[8]
port 283 nsew signal input
rlabel metal2 s 32126 90640 32182 90800 6 Tile_X0Y0_SS4END[9]
port 284 nsew signal input
rlabel metal2 s 34058 90640 34114 90800 6 Tile_X0Y0_UserCLKo
port 285 nsew signal output
rlabel metal3 s 0 50600 160 50720 6 Tile_X0Y0_W1BEG[0]
port 286 nsew signal output
rlabel metal3 s 0 50872 160 50992 6 Tile_X0Y0_W1BEG[1]
port 287 nsew signal output
rlabel metal3 s 0 51144 160 51264 6 Tile_X0Y0_W1BEG[2]
port 288 nsew signal output
rlabel metal3 s 0 51416 160 51536 6 Tile_X0Y0_W1BEG[3]
port 289 nsew signal output
rlabel metal3 s 44840 50600 45000 50720 6 Tile_X0Y0_W1END[0]
port 290 nsew signal input
rlabel metal3 s 44840 50872 45000 50992 6 Tile_X0Y0_W1END[1]
port 291 nsew signal input
rlabel metal3 s 44840 51144 45000 51264 6 Tile_X0Y0_W1END[2]
port 292 nsew signal input
rlabel metal3 s 44840 51416 45000 51536 6 Tile_X0Y0_W1END[3]
port 293 nsew signal input
rlabel metal3 s 0 51688 160 51808 6 Tile_X0Y0_W2BEG[0]
port 294 nsew signal output
rlabel metal3 s 0 51960 160 52080 6 Tile_X0Y0_W2BEG[1]
port 295 nsew signal output
rlabel metal3 s 0 52232 160 52352 6 Tile_X0Y0_W2BEG[2]
port 296 nsew signal output
rlabel metal3 s 0 52504 160 52624 6 Tile_X0Y0_W2BEG[3]
port 297 nsew signal output
rlabel metal3 s 0 52776 160 52896 6 Tile_X0Y0_W2BEG[4]
port 298 nsew signal output
rlabel metal3 s 0 53048 160 53168 6 Tile_X0Y0_W2BEG[5]
port 299 nsew signal output
rlabel metal3 s 0 53320 160 53440 6 Tile_X0Y0_W2BEG[6]
port 300 nsew signal output
rlabel metal3 s 0 53592 160 53712 6 Tile_X0Y0_W2BEG[7]
port 301 nsew signal output
rlabel metal3 s 0 53864 160 53984 6 Tile_X0Y0_W2BEGb[0]
port 302 nsew signal output
rlabel metal3 s 0 54136 160 54256 6 Tile_X0Y0_W2BEGb[1]
port 303 nsew signal output
rlabel metal3 s 0 54408 160 54528 6 Tile_X0Y0_W2BEGb[2]
port 304 nsew signal output
rlabel metal3 s 0 54680 160 54800 6 Tile_X0Y0_W2BEGb[3]
port 305 nsew signal output
rlabel metal3 s 0 54952 160 55072 6 Tile_X0Y0_W2BEGb[4]
port 306 nsew signal output
rlabel metal3 s 0 55224 160 55344 6 Tile_X0Y0_W2BEGb[5]
port 307 nsew signal output
rlabel metal3 s 0 55496 160 55616 6 Tile_X0Y0_W2BEGb[6]
port 308 nsew signal output
rlabel metal3 s 0 55768 160 55888 6 Tile_X0Y0_W2BEGb[7]
port 309 nsew signal output
rlabel metal3 s 44840 53864 45000 53984 6 Tile_X0Y0_W2END[0]
port 310 nsew signal input
rlabel metal3 s 44840 54136 45000 54256 6 Tile_X0Y0_W2END[1]
port 311 nsew signal input
rlabel metal3 s 44840 54408 45000 54528 6 Tile_X0Y0_W2END[2]
port 312 nsew signal input
rlabel metal3 s 44840 54680 45000 54800 6 Tile_X0Y0_W2END[3]
port 313 nsew signal input
rlabel metal3 s 44840 54952 45000 55072 6 Tile_X0Y0_W2END[4]
port 314 nsew signal input
rlabel metal3 s 44840 55224 45000 55344 6 Tile_X0Y0_W2END[5]
port 315 nsew signal input
rlabel metal3 s 44840 55496 45000 55616 6 Tile_X0Y0_W2END[6]
port 316 nsew signal input
rlabel metal3 s 44840 55768 45000 55888 6 Tile_X0Y0_W2END[7]
port 317 nsew signal input
rlabel metal3 s 44840 51688 45000 51808 6 Tile_X0Y0_W2MID[0]
port 318 nsew signal input
rlabel metal3 s 44840 51960 45000 52080 6 Tile_X0Y0_W2MID[1]
port 319 nsew signal input
rlabel metal3 s 44840 52232 45000 52352 6 Tile_X0Y0_W2MID[2]
port 320 nsew signal input
rlabel metal3 s 44840 52504 45000 52624 6 Tile_X0Y0_W2MID[3]
port 321 nsew signal input
rlabel metal3 s 44840 52776 45000 52896 6 Tile_X0Y0_W2MID[4]
port 322 nsew signal input
rlabel metal3 s 44840 53048 45000 53168 6 Tile_X0Y0_W2MID[5]
port 323 nsew signal input
rlabel metal3 s 44840 53320 45000 53440 6 Tile_X0Y0_W2MID[6]
port 324 nsew signal input
rlabel metal3 s 44840 53592 45000 53712 6 Tile_X0Y0_W2MID[7]
port 325 nsew signal input
rlabel metal3 s 0 60392 160 60512 6 Tile_X0Y0_W6BEG[0]
port 326 nsew signal output
rlabel metal3 s 0 63112 160 63232 6 Tile_X0Y0_W6BEG[10]
port 327 nsew signal output
rlabel metal3 s 0 63384 160 63504 6 Tile_X0Y0_W6BEG[11]
port 328 nsew signal output
rlabel metal3 s 0 60664 160 60784 6 Tile_X0Y0_W6BEG[1]
port 329 nsew signal output
rlabel metal3 s 0 60936 160 61056 6 Tile_X0Y0_W6BEG[2]
port 330 nsew signal output
rlabel metal3 s 0 61208 160 61328 6 Tile_X0Y0_W6BEG[3]
port 331 nsew signal output
rlabel metal3 s 0 61480 160 61600 6 Tile_X0Y0_W6BEG[4]
port 332 nsew signal output
rlabel metal3 s 0 61752 160 61872 6 Tile_X0Y0_W6BEG[5]
port 333 nsew signal output
rlabel metal3 s 0 62024 160 62144 6 Tile_X0Y0_W6BEG[6]
port 334 nsew signal output
rlabel metal3 s 0 62296 160 62416 6 Tile_X0Y0_W6BEG[7]
port 335 nsew signal output
rlabel metal3 s 0 62568 160 62688 6 Tile_X0Y0_W6BEG[8]
port 336 nsew signal output
rlabel metal3 s 0 62840 160 62960 6 Tile_X0Y0_W6BEG[9]
port 337 nsew signal output
rlabel metal3 s 44840 60392 45000 60512 6 Tile_X0Y0_W6END[0]
port 338 nsew signal input
rlabel metal3 s 44840 63112 45000 63232 6 Tile_X0Y0_W6END[10]
port 339 nsew signal input
rlabel metal3 s 44840 63384 45000 63504 6 Tile_X0Y0_W6END[11]
port 340 nsew signal input
rlabel metal3 s 44840 60664 45000 60784 6 Tile_X0Y0_W6END[1]
port 341 nsew signal input
rlabel metal3 s 44840 60936 45000 61056 6 Tile_X0Y0_W6END[2]
port 342 nsew signal input
rlabel metal3 s 44840 61208 45000 61328 6 Tile_X0Y0_W6END[3]
port 343 nsew signal input
rlabel metal3 s 44840 61480 45000 61600 6 Tile_X0Y0_W6END[4]
port 344 nsew signal input
rlabel metal3 s 44840 61752 45000 61872 6 Tile_X0Y0_W6END[5]
port 345 nsew signal input
rlabel metal3 s 44840 62024 45000 62144 6 Tile_X0Y0_W6END[6]
port 346 nsew signal input
rlabel metal3 s 44840 62296 45000 62416 6 Tile_X0Y0_W6END[7]
port 347 nsew signal input
rlabel metal3 s 44840 62568 45000 62688 6 Tile_X0Y0_W6END[8]
port 348 nsew signal input
rlabel metal3 s 44840 62840 45000 62960 6 Tile_X0Y0_W6END[9]
port 349 nsew signal input
rlabel metal3 s 0 56040 160 56160 6 Tile_X0Y0_WW4BEG[0]
port 350 nsew signal output
rlabel metal3 s 0 58760 160 58880 6 Tile_X0Y0_WW4BEG[10]
port 351 nsew signal output
rlabel metal3 s 0 59032 160 59152 6 Tile_X0Y0_WW4BEG[11]
port 352 nsew signal output
rlabel metal3 s 0 59304 160 59424 6 Tile_X0Y0_WW4BEG[12]
port 353 nsew signal output
rlabel metal3 s 0 59576 160 59696 6 Tile_X0Y0_WW4BEG[13]
port 354 nsew signal output
rlabel metal3 s 0 59848 160 59968 6 Tile_X0Y0_WW4BEG[14]
port 355 nsew signal output
rlabel metal3 s 0 60120 160 60240 6 Tile_X0Y0_WW4BEG[15]
port 356 nsew signal output
rlabel metal3 s 0 56312 160 56432 6 Tile_X0Y0_WW4BEG[1]
port 357 nsew signal output
rlabel metal3 s 0 56584 160 56704 6 Tile_X0Y0_WW4BEG[2]
port 358 nsew signal output
rlabel metal3 s 0 56856 160 56976 6 Tile_X0Y0_WW4BEG[3]
port 359 nsew signal output
rlabel metal3 s 0 57128 160 57248 6 Tile_X0Y0_WW4BEG[4]
port 360 nsew signal output
rlabel metal3 s 0 57400 160 57520 6 Tile_X0Y0_WW4BEG[5]
port 361 nsew signal output
rlabel metal3 s 0 57672 160 57792 6 Tile_X0Y0_WW4BEG[6]
port 362 nsew signal output
rlabel metal3 s 0 57944 160 58064 6 Tile_X0Y0_WW4BEG[7]
port 363 nsew signal output
rlabel metal3 s 0 58216 160 58336 6 Tile_X0Y0_WW4BEG[8]
port 364 nsew signal output
rlabel metal3 s 0 58488 160 58608 6 Tile_X0Y0_WW4BEG[9]
port 365 nsew signal output
rlabel metal3 s 44840 56040 45000 56160 6 Tile_X0Y0_WW4END[0]
port 366 nsew signal input
rlabel metal3 s 44840 58760 45000 58880 6 Tile_X0Y0_WW4END[10]
port 367 nsew signal input
rlabel metal3 s 44840 59032 45000 59152 6 Tile_X0Y0_WW4END[11]
port 368 nsew signal input
rlabel metal3 s 44840 59304 45000 59424 6 Tile_X0Y0_WW4END[12]
port 369 nsew signal input
rlabel metal3 s 44840 59576 45000 59696 6 Tile_X0Y0_WW4END[13]
port 370 nsew signal input
rlabel metal3 s 44840 59848 45000 59968 6 Tile_X0Y0_WW4END[14]
port 371 nsew signal input
rlabel metal3 s 44840 60120 45000 60240 6 Tile_X0Y0_WW4END[15]
port 372 nsew signal input
rlabel metal3 s 44840 56312 45000 56432 6 Tile_X0Y0_WW4END[1]
port 373 nsew signal input
rlabel metal3 s 44840 56584 45000 56704 6 Tile_X0Y0_WW4END[2]
port 374 nsew signal input
rlabel metal3 s 44840 56856 45000 56976 6 Tile_X0Y0_WW4END[3]
port 375 nsew signal input
rlabel metal3 s 44840 57128 45000 57248 6 Tile_X0Y0_WW4END[4]
port 376 nsew signal input
rlabel metal3 s 44840 57400 45000 57520 6 Tile_X0Y0_WW4END[5]
port 377 nsew signal input
rlabel metal3 s 44840 57672 45000 57792 6 Tile_X0Y0_WW4END[6]
port 378 nsew signal input
rlabel metal3 s 44840 57944 45000 58064 6 Tile_X0Y0_WW4END[7]
port 379 nsew signal input
rlabel metal3 s 44840 58216 45000 58336 6 Tile_X0Y0_WW4END[8]
port 380 nsew signal input
rlabel metal3 s 44840 58488 45000 58608 6 Tile_X0Y0_WW4END[9]
port 381 nsew signal input
rlabel metal3 s 44840 17688 45000 17808 6 Tile_X0Y1_E1BEG[0]
port 382 nsew signal output
rlabel metal3 s 44840 17960 45000 18080 6 Tile_X0Y1_E1BEG[1]
port 383 nsew signal output
rlabel metal3 s 44840 18232 45000 18352 6 Tile_X0Y1_E1BEG[2]
port 384 nsew signal output
rlabel metal3 s 44840 18504 45000 18624 6 Tile_X0Y1_E1BEG[3]
port 385 nsew signal output
rlabel metal3 s 0 17688 160 17808 6 Tile_X0Y1_E1END[0]
port 386 nsew signal input
rlabel metal3 s 0 17960 160 18080 6 Tile_X0Y1_E1END[1]
port 387 nsew signal input
rlabel metal3 s 0 18232 160 18352 6 Tile_X0Y1_E1END[2]
port 388 nsew signal input
rlabel metal3 s 0 18504 160 18624 6 Tile_X0Y1_E1END[3]
port 389 nsew signal input
rlabel metal3 s 44840 18776 45000 18896 6 Tile_X0Y1_E2BEG[0]
port 390 nsew signal output
rlabel metal3 s 44840 19048 45000 19168 6 Tile_X0Y1_E2BEG[1]
port 391 nsew signal output
rlabel metal3 s 44840 19320 45000 19440 6 Tile_X0Y1_E2BEG[2]
port 392 nsew signal output
rlabel metal3 s 44840 19592 45000 19712 6 Tile_X0Y1_E2BEG[3]
port 393 nsew signal output
rlabel metal3 s 44840 19864 45000 19984 6 Tile_X0Y1_E2BEG[4]
port 394 nsew signal output
rlabel metal3 s 44840 20136 45000 20256 6 Tile_X0Y1_E2BEG[5]
port 395 nsew signal output
rlabel metal3 s 44840 20408 45000 20528 6 Tile_X0Y1_E2BEG[6]
port 396 nsew signal output
rlabel metal3 s 44840 20680 45000 20800 6 Tile_X0Y1_E2BEG[7]
port 397 nsew signal output
rlabel metal3 s 44840 20952 45000 21072 6 Tile_X0Y1_E2BEGb[0]
port 398 nsew signal output
rlabel metal3 s 44840 21224 45000 21344 6 Tile_X0Y1_E2BEGb[1]
port 399 nsew signal output
rlabel metal3 s 44840 21496 45000 21616 6 Tile_X0Y1_E2BEGb[2]
port 400 nsew signal output
rlabel metal3 s 44840 21768 45000 21888 6 Tile_X0Y1_E2BEGb[3]
port 401 nsew signal output
rlabel metal3 s 44840 22040 45000 22160 6 Tile_X0Y1_E2BEGb[4]
port 402 nsew signal output
rlabel metal3 s 44840 22312 45000 22432 6 Tile_X0Y1_E2BEGb[5]
port 403 nsew signal output
rlabel metal3 s 44840 22584 45000 22704 6 Tile_X0Y1_E2BEGb[6]
port 404 nsew signal output
rlabel metal3 s 44840 22856 45000 22976 6 Tile_X0Y1_E2BEGb[7]
port 405 nsew signal output
rlabel metal3 s 0 20952 160 21072 6 Tile_X0Y1_E2END[0]
port 406 nsew signal input
rlabel metal3 s 0 21224 160 21344 6 Tile_X0Y1_E2END[1]
port 407 nsew signal input
rlabel metal3 s 0 21496 160 21616 6 Tile_X0Y1_E2END[2]
port 408 nsew signal input
rlabel metal3 s 0 21768 160 21888 6 Tile_X0Y1_E2END[3]
port 409 nsew signal input
rlabel metal3 s 0 22040 160 22160 6 Tile_X0Y1_E2END[4]
port 410 nsew signal input
rlabel metal3 s 0 22312 160 22432 6 Tile_X0Y1_E2END[5]
port 411 nsew signal input
rlabel metal3 s 0 22584 160 22704 6 Tile_X0Y1_E2END[6]
port 412 nsew signal input
rlabel metal3 s 0 22856 160 22976 6 Tile_X0Y1_E2END[7]
port 413 nsew signal input
rlabel metal3 s 0 18776 160 18896 6 Tile_X0Y1_E2MID[0]
port 414 nsew signal input
rlabel metal3 s 0 19048 160 19168 6 Tile_X0Y1_E2MID[1]
port 415 nsew signal input
rlabel metal3 s 0 19320 160 19440 6 Tile_X0Y1_E2MID[2]
port 416 nsew signal input
rlabel metal3 s 0 19592 160 19712 6 Tile_X0Y1_E2MID[3]
port 417 nsew signal input
rlabel metal3 s 0 19864 160 19984 6 Tile_X0Y1_E2MID[4]
port 418 nsew signal input
rlabel metal3 s 0 20136 160 20256 6 Tile_X0Y1_E2MID[5]
port 419 nsew signal input
rlabel metal3 s 0 20408 160 20528 6 Tile_X0Y1_E2MID[6]
port 420 nsew signal input
rlabel metal3 s 0 20680 160 20800 6 Tile_X0Y1_E2MID[7]
port 421 nsew signal input
rlabel metal3 s 44840 27480 45000 27600 6 Tile_X0Y1_E6BEG[0]
port 422 nsew signal output
rlabel metal3 s 44840 30200 45000 30320 6 Tile_X0Y1_E6BEG[10]
port 423 nsew signal output
rlabel metal3 s 44840 30472 45000 30592 6 Tile_X0Y1_E6BEG[11]
port 424 nsew signal output
rlabel metal3 s 44840 27752 45000 27872 6 Tile_X0Y1_E6BEG[1]
port 425 nsew signal output
rlabel metal3 s 44840 28024 45000 28144 6 Tile_X0Y1_E6BEG[2]
port 426 nsew signal output
rlabel metal3 s 44840 28296 45000 28416 6 Tile_X0Y1_E6BEG[3]
port 427 nsew signal output
rlabel metal3 s 44840 28568 45000 28688 6 Tile_X0Y1_E6BEG[4]
port 428 nsew signal output
rlabel metal3 s 44840 28840 45000 28960 6 Tile_X0Y1_E6BEG[5]
port 429 nsew signal output
rlabel metal3 s 44840 29112 45000 29232 6 Tile_X0Y1_E6BEG[6]
port 430 nsew signal output
rlabel metal3 s 44840 29384 45000 29504 6 Tile_X0Y1_E6BEG[7]
port 431 nsew signal output
rlabel metal3 s 44840 29656 45000 29776 6 Tile_X0Y1_E6BEG[8]
port 432 nsew signal output
rlabel metal3 s 44840 29928 45000 30048 6 Tile_X0Y1_E6BEG[9]
port 433 nsew signal output
rlabel metal3 s 0 27480 160 27600 6 Tile_X0Y1_E6END[0]
port 434 nsew signal input
rlabel metal3 s 0 30200 160 30320 6 Tile_X0Y1_E6END[10]
port 435 nsew signal input
rlabel metal3 s 0 30472 160 30592 6 Tile_X0Y1_E6END[11]
port 436 nsew signal input
rlabel metal3 s 0 27752 160 27872 6 Tile_X0Y1_E6END[1]
port 437 nsew signal input
rlabel metal3 s 0 28024 160 28144 6 Tile_X0Y1_E6END[2]
port 438 nsew signal input
rlabel metal3 s 0 28296 160 28416 6 Tile_X0Y1_E6END[3]
port 439 nsew signal input
rlabel metal3 s 0 28568 160 28688 6 Tile_X0Y1_E6END[4]
port 440 nsew signal input
rlabel metal3 s 0 28840 160 28960 6 Tile_X0Y1_E6END[5]
port 441 nsew signal input
rlabel metal3 s 0 29112 160 29232 6 Tile_X0Y1_E6END[6]
port 442 nsew signal input
rlabel metal3 s 0 29384 160 29504 6 Tile_X0Y1_E6END[7]
port 443 nsew signal input
rlabel metal3 s 0 29656 160 29776 6 Tile_X0Y1_E6END[8]
port 444 nsew signal input
rlabel metal3 s 0 29928 160 30048 6 Tile_X0Y1_E6END[9]
port 445 nsew signal input
rlabel metal3 s 44840 23128 45000 23248 6 Tile_X0Y1_EE4BEG[0]
port 446 nsew signal output
rlabel metal3 s 44840 25848 45000 25968 6 Tile_X0Y1_EE4BEG[10]
port 447 nsew signal output
rlabel metal3 s 44840 26120 45000 26240 6 Tile_X0Y1_EE4BEG[11]
port 448 nsew signal output
rlabel metal3 s 44840 26392 45000 26512 6 Tile_X0Y1_EE4BEG[12]
port 449 nsew signal output
rlabel metal3 s 44840 26664 45000 26784 6 Tile_X0Y1_EE4BEG[13]
port 450 nsew signal output
rlabel metal3 s 44840 26936 45000 27056 6 Tile_X0Y1_EE4BEG[14]
port 451 nsew signal output
rlabel metal3 s 44840 27208 45000 27328 6 Tile_X0Y1_EE4BEG[15]
port 452 nsew signal output
rlabel metal3 s 44840 23400 45000 23520 6 Tile_X0Y1_EE4BEG[1]
port 453 nsew signal output
rlabel metal3 s 44840 23672 45000 23792 6 Tile_X0Y1_EE4BEG[2]
port 454 nsew signal output
rlabel metal3 s 44840 23944 45000 24064 6 Tile_X0Y1_EE4BEG[3]
port 455 nsew signal output
rlabel metal3 s 44840 24216 45000 24336 6 Tile_X0Y1_EE4BEG[4]
port 456 nsew signal output
rlabel metal3 s 44840 24488 45000 24608 6 Tile_X0Y1_EE4BEG[5]
port 457 nsew signal output
rlabel metal3 s 44840 24760 45000 24880 6 Tile_X0Y1_EE4BEG[6]
port 458 nsew signal output
rlabel metal3 s 44840 25032 45000 25152 6 Tile_X0Y1_EE4BEG[7]
port 459 nsew signal output
rlabel metal3 s 44840 25304 45000 25424 6 Tile_X0Y1_EE4BEG[8]
port 460 nsew signal output
rlabel metal3 s 44840 25576 45000 25696 6 Tile_X0Y1_EE4BEG[9]
port 461 nsew signal output
rlabel metal3 s 0 23128 160 23248 6 Tile_X0Y1_EE4END[0]
port 462 nsew signal input
rlabel metal3 s 0 25848 160 25968 6 Tile_X0Y1_EE4END[10]
port 463 nsew signal input
rlabel metal3 s 0 26120 160 26240 6 Tile_X0Y1_EE4END[11]
port 464 nsew signal input
rlabel metal3 s 0 26392 160 26512 6 Tile_X0Y1_EE4END[12]
port 465 nsew signal input
rlabel metal3 s 0 26664 160 26784 6 Tile_X0Y1_EE4END[13]
port 466 nsew signal input
rlabel metal3 s 0 26936 160 27056 6 Tile_X0Y1_EE4END[14]
port 467 nsew signal input
rlabel metal3 s 0 27208 160 27328 6 Tile_X0Y1_EE4END[15]
port 468 nsew signal input
rlabel metal3 s 0 23400 160 23520 6 Tile_X0Y1_EE4END[1]
port 469 nsew signal input
rlabel metal3 s 0 23672 160 23792 6 Tile_X0Y1_EE4END[2]
port 470 nsew signal input
rlabel metal3 s 0 23944 160 24064 6 Tile_X0Y1_EE4END[3]
port 471 nsew signal input
rlabel metal3 s 0 24216 160 24336 6 Tile_X0Y1_EE4END[4]
port 472 nsew signal input
rlabel metal3 s 0 24488 160 24608 6 Tile_X0Y1_EE4END[5]
port 473 nsew signal input
rlabel metal3 s 0 24760 160 24880 6 Tile_X0Y1_EE4END[6]
port 474 nsew signal input
rlabel metal3 s 0 25032 160 25152 6 Tile_X0Y1_EE4END[7]
port 475 nsew signal input
rlabel metal3 s 0 25304 160 25424 6 Tile_X0Y1_EE4END[8]
port 476 nsew signal input
rlabel metal3 s 0 25576 160 25696 6 Tile_X0Y1_EE4END[9]
port 477 nsew signal input
rlabel metal3 s 0 30744 160 30864 6 Tile_X0Y1_FrameData[0]
port 478 nsew signal input
rlabel metal3 s 0 33464 160 33584 6 Tile_X0Y1_FrameData[10]
port 479 nsew signal input
rlabel metal3 s 0 33736 160 33856 6 Tile_X0Y1_FrameData[11]
port 480 nsew signal input
rlabel metal3 s 0 34008 160 34128 6 Tile_X0Y1_FrameData[12]
port 481 nsew signal input
rlabel metal3 s 0 34280 160 34400 6 Tile_X0Y1_FrameData[13]
port 482 nsew signal input
rlabel metal3 s 0 34552 160 34672 6 Tile_X0Y1_FrameData[14]
port 483 nsew signal input
rlabel metal3 s 0 34824 160 34944 6 Tile_X0Y1_FrameData[15]
port 484 nsew signal input
rlabel metal3 s 0 35096 160 35216 6 Tile_X0Y1_FrameData[16]
port 485 nsew signal input
rlabel metal3 s 0 35368 160 35488 6 Tile_X0Y1_FrameData[17]
port 486 nsew signal input
rlabel metal3 s 0 35640 160 35760 6 Tile_X0Y1_FrameData[18]
port 487 nsew signal input
rlabel metal3 s 0 35912 160 36032 6 Tile_X0Y1_FrameData[19]
port 488 nsew signal input
rlabel metal3 s 0 31016 160 31136 6 Tile_X0Y1_FrameData[1]
port 489 nsew signal input
rlabel metal3 s 0 36184 160 36304 6 Tile_X0Y1_FrameData[20]
port 490 nsew signal input
rlabel metal3 s 0 36456 160 36576 6 Tile_X0Y1_FrameData[21]
port 491 nsew signal input
rlabel metal3 s 0 36728 160 36848 6 Tile_X0Y1_FrameData[22]
port 492 nsew signal input
rlabel metal3 s 0 37000 160 37120 6 Tile_X0Y1_FrameData[23]
port 493 nsew signal input
rlabel metal3 s 0 37272 160 37392 6 Tile_X0Y1_FrameData[24]
port 494 nsew signal input
rlabel metal3 s 0 37544 160 37664 6 Tile_X0Y1_FrameData[25]
port 495 nsew signal input
rlabel metal3 s 0 37816 160 37936 6 Tile_X0Y1_FrameData[26]
port 496 nsew signal input
rlabel metal3 s 0 38088 160 38208 6 Tile_X0Y1_FrameData[27]
port 497 nsew signal input
rlabel metal3 s 0 38360 160 38480 6 Tile_X0Y1_FrameData[28]
port 498 nsew signal input
rlabel metal3 s 0 38632 160 38752 6 Tile_X0Y1_FrameData[29]
port 499 nsew signal input
rlabel metal3 s 0 31288 160 31408 6 Tile_X0Y1_FrameData[2]
port 500 nsew signal input
rlabel metal3 s 0 38904 160 39024 6 Tile_X0Y1_FrameData[30]
port 501 nsew signal input
rlabel metal3 s 0 39176 160 39296 6 Tile_X0Y1_FrameData[31]
port 502 nsew signal input
rlabel metal3 s 0 31560 160 31680 6 Tile_X0Y1_FrameData[3]
port 503 nsew signal input
rlabel metal3 s 0 31832 160 31952 6 Tile_X0Y1_FrameData[4]
port 504 nsew signal input
rlabel metal3 s 0 32104 160 32224 6 Tile_X0Y1_FrameData[5]
port 505 nsew signal input
rlabel metal3 s 0 32376 160 32496 6 Tile_X0Y1_FrameData[6]
port 506 nsew signal input
rlabel metal3 s 0 32648 160 32768 6 Tile_X0Y1_FrameData[7]
port 507 nsew signal input
rlabel metal3 s 0 32920 160 33040 6 Tile_X0Y1_FrameData[8]
port 508 nsew signal input
rlabel metal3 s 0 33192 160 33312 6 Tile_X0Y1_FrameData[9]
port 509 nsew signal input
rlabel metal3 s 44840 30744 45000 30864 6 Tile_X0Y1_FrameData_O[0]
port 510 nsew signal output
rlabel metal3 s 44840 33464 45000 33584 6 Tile_X0Y1_FrameData_O[10]
port 511 nsew signal output
rlabel metal3 s 44840 33736 45000 33856 6 Tile_X0Y1_FrameData_O[11]
port 512 nsew signal output
rlabel metal3 s 44840 34008 45000 34128 6 Tile_X0Y1_FrameData_O[12]
port 513 nsew signal output
rlabel metal3 s 44840 34280 45000 34400 6 Tile_X0Y1_FrameData_O[13]
port 514 nsew signal output
rlabel metal3 s 44840 34552 45000 34672 6 Tile_X0Y1_FrameData_O[14]
port 515 nsew signal output
rlabel metal3 s 44840 34824 45000 34944 6 Tile_X0Y1_FrameData_O[15]
port 516 nsew signal output
rlabel metal3 s 44840 35096 45000 35216 6 Tile_X0Y1_FrameData_O[16]
port 517 nsew signal output
rlabel metal3 s 44840 35368 45000 35488 6 Tile_X0Y1_FrameData_O[17]
port 518 nsew signal output
rlabel metal3 s 44840 35640 45000 35760 6 Tile_X0Y1_FrameData_O[18]
port 519 nsew signal output
rlabel metal3 s 44840 35912 45000 36032 6 Tile_X0Y1_FrameData_O[19]
port 520 nsew signal output
rlabel metal3 s 44840 31016 45000 31136 6 Tile_X0Y1_FrameData_O[1]
port 521 nsew signal output
rlabel metal3 s 44840 36184 45000 36304 6 Tile_X0Y1_FrameData_O[20]
port 522 nsew signal output
rlabel metal3 s 44840 36456 45000 36576 6 Tile_X0Y1_FrameData_O[21]
port 523 nsew signal output
rlabel metal3 s 44840 36728 45000 36848 6 Tile_X0Y1_FrameData_O[22]
port 524 nsew signal output
rlabel metal3 s 44840 37000 45000 37120 6 Tile_X0Y1_FrameData_O[23]
port 525 nsew signal output
rlabel metal3 s 44840 37272 45000 37392 6 Tile_X0Y1_FrameData_O[24]
port 526 nsew signal output
rlabel metal3 s 44840 37544 45000 37664 6 Tile_X0Y1_FrameData_O[25]
port 527 nsew signal output
rlabel metal3 s 44840 37816 45000 37936 6 Tile_X0Y1_FrameData_O[26]
port 528 nsew signal output
rlabel metal3 s 44840 38088 45000 38208 6 Tile_X0Y1_FrameData_O[27]
port 529 nsew signal output
rlabel metal3 s 44840 38360 45000 38480 6 Tile_X0Y1_FrameData_O[28]
port 530 nsew signal output
rlabel metal3 s 44840 38632 45000 38752 6 Tile_X0Y1_FrameData_O[29]
port 531 nsew signal output
rlabel metal3 s 44840 31288 45000 31408 6 Tile_X0Y1_FrameData_O[2]
port 532 nsew signal output
rlabel metal3 s 44840 38904 45000 39024 6 Tile_X0Y1_FrameData_O[30]
port 533 nsew signal output
rlabel metal3 s 44840 39176 45000 39296 6 Tile_X0Y1_FrameData_O[31]
port 534 nsew signal output
rlabel metal3 s 44840 31560 45000 31680 6 Tile_X0Y1_FrameData_O[3]
port 535 nsew signal output
rlabel metal3 s 44840 31832 45000 31952 6 Tile_X0Y1_FrameData_O[4]
port 536 nsew signal output
rlabel metal3 s 44840 32104 45000 32224 6 Tile_X0Y1_FrameData_O[5]
port 537 nsew signal output
rlabel metal3 s 44840 32376 45000 32496 6 Tile_X0Y1_FrameData_O[6]
port 538 nsew signal output
rlabel metal3 s 44840 32648 45000 32768 6 Tile_X0Y1_FrameData_O[7]
port 539 nsew signal output
rlabel metal3 s 44840 32920 45000 33040 6 Tile_X0Y1_FrameData_O[8]
port 540 nsew signal output
rlabel metal3 s 44840 33192 45000 33312 6 Tile_X0Y1_FrameData_O[9]
port 541 nsew signal output
rlabel metal2 s 34334 0 34390 160 6 Tile_X0Y1_FrameStrobe[0]
port 542 nsew signal input
rlabel metal2 s 37094 0 37150 160 6 Tile_X0Y1_FrameStrobe[10]
port 543 nsew signal input
rlabel metal2 s 37370 0 37426 160 6 Tile_X0Y1_FrameStrobe[11]
port 544 nsew signal input
rlabel metal2 s 37646 0 37702 160 6 Tile_X0Y1_FrameStrobe[12]
port 545 nsew signal input
rlabel metal2 s 37922 0 37978 160 6 Tile_X0Y1_FrameStrobe[13]
port 546 nsew signal input
rlabel metal2 s 38198 0 38254 160 6 Tile_X0Y1_FrameStrobe[14]
port 547 nsew signal input
rlabel metal2 s 38474 0 38530 160 6 Tile_X0Y1_FrameStrobe[15]
port 548 nsew signal input
rlabel metal2 s 38750 0 38806 160 6 Tile_X0Y1_FrameStrobe[16]
port 549 nsew signal input
rlabel metal2 s 39026 0 39082 160 6 Tile_X0Y1_FrameStrobe[17]
port 550 nsew signal input
rlabel metal2 s 39302 0 39358 160 6 Tile_X0Y1_FrameStrobe[18]
port 551 nsew signal input
rlabel metal2 s 39578 0 39634 160 6 Tile_X0Y1_FrameStrobe[19]
port 552 nsew signal input
rlabel metal2 s 34610 0 34666 160 6 Tile_X0Y1_FrameStrobe[1]
port 553 nsew signal input
rlabel metal2 s 34886 0 34942 160 6 Tile_X0Y1_FrameStrobe[2]
port 554 nsew signal input
rlabel metal2 s 35162 0 35218 160 6 Tile_X0Y1_FrameStrobe[3]
port 555 nsew signal input
rlabel metal2 s 35438 0 35494 160 6 Tile_X0Y1_FrameStrobe[4]
port 556 nsew signal input
rlabel metal2 s 35714 0 35770 160 6 Tile_X0Y1_FrameStrobe[5]
port 557 nsew signal input
rlabel metal2 s 35990 0 36046 160 6 Tile_X0Y1_FrameStrobe[6]
port 558 nsew signal input
rlabel metal2 s 36266 0 36322 160 6 Tile_X0Y1_FrameStrobe[7]
port 559 nsew signal input
rlabel metal2 s 36542 0 36598 160 6 Tile_X0Y1_FrameStrobe[8]
port 560 nsew signal input
rlabel metal2 s 36818 0 36874 160 6 Tile_X0Y1_FrameStrobe[9]
port 561 nsew signal input
rlabel metal2 s 5354 0 5410 160 6 Tile_X0Y1_N1END[0]
port 562 nsew signal input
rlabel metal2 s 5630 0 5686 160 6 Tile_X0Y1_N1END[1]
port 563 nsew signal input
rlabel metal2 s 5906 0 5962 160 6 Tile_X0Y1_N1END[2]
port 564 nsew signal input
rlabel metal2 s 6182 0 6238 160 6 Tile_X0Y1_N1END[3]
port 565 nsew signal input
rlabel metal2 s 8666 0 8722 160 6 Tile_X0Y1_N2END[0]
port 566 nsew signal input
rlabel metal2 s 8942 0 8998 160 6 Tile_X0Y1_N2END[1]
port 567 nsew signal input
rlabel metal2 s 9218 0 9274 160 6 Tile_X0Y1_N2END[2]
port 568 nsew signal input
rlabel metal2 s 9494 0 9550 160 6 Tile_X0Y1_N2END[3]
port 569 nsew signal input
rlabel metal2 s 9770 0 9826 160 6 Tile_X0Y1_N2END[4]
port 570 nsew signal input
rlabel metal2 s 10046 0 10102 160 6 Tile_X0Y1_N2END[5]
port 571 nsew signal input
rlabel metal2 s 10322 0 10378 160 6 Tile_X0Y1_N2END[6]
port 572 nsew signal input
rlabel metal2 s 10598 0 10654 160 6 Tile_X0Y1_N2END[7]
port 573 nsew signal input
rlabel metal2 s 6458 0 6514 160 6 Tile_X0Y1_N2MID[0]
port 574 nsew signal input
rlabel metal2 s 6734 0 6790 160 6 Tile_X0Y1_N2MID[1]
port 575 nsew signal input
rlabel metal2 s 7010 0 7066 160 6 Tile_X0Y1_N2MID[2]
port 576 nsew signal input
rlabel metal2 s 7286 0 7342 160 6 Tile_X0Y1_N2MID[3]
port 577 nsew signal input
rlabel metal2 s 7562 0 7618 160 6 Tile_X0Y1_N2MID[4]
port 578 nsew signal input
rlabel metal2 s 7838 0 7894 160 6 Tile_X0Y1_N2MID[5]
port 579 nsew signal input
rlabel metal2 s 8114 0 8170 160 6 Tile_X0Y1_N2MID[6]
port 580 nsew signal input
rlabel metal2 s 8390 0 8446 160 6 Tile_X0Y1_N2MID[7]
port 581 nsew signal input
rlabel metal2 s 10874 0 10930 160 6 Tile_X0Y1_N4END[0]
port 582 nsew signal input
rlabel metal2 s 13634 0 13690 160 6 Tile_X0Y1_N4END[10]
port 583 nsew signal input
rlabel metal2 s 13910 0 13966 160 6 Tile_X0Y1_N4END[11]
port 584 nsew signal input
rlabel metal2 s 14186 0 14242 160 6 Tile_X0Y1_N4END[12]
port 585 nsew signal input
rlabel metal2 s 14462 0 14518 160 6 Tile_X0Y1_N4END[13]
port 586 nsew signal input
rlabel metal2 s 14738 0 14794 160 6 Tile_X0Y1_N4END[14]
port 587 nsew signal input
rlabel metal2 s 15014 0 15070 160 6 Tile_X0Y1_N4END[15]
port 588 nsew signal input
rlabel metal2 s 11150 0 11206 160 6 Tile_X0Y1_N4END[1]
port 589 nsew signal input
rlabel metal2 s 11426 0 11482 160 6 Tile_X0Y1_N4END[2]
port 590 nsew signal input
rlabel metal2 s 11702 0 11758 160 6 Tile_X0Y1_N4END[3]
port 591 nsew signal input
rlabel metal2 s 11978 0 12034 160 6 Tile_X0Y1_N4END[4]
port 592 nsew signal input
rlabel metal2 s 12254 0 12310 160 6 Tile_X0Y1_N4END[5]
port 593 nsew signal input
rlabel metal2 s 12530 0 12586 160 6 Tile_X0Y1_N4END[6]
port 594 nsew signal input
rlabel metal2 s 12806 0 12862 160 6 Tile_X0Y1_N4END[7]
port 595 nsew signal input
rlabel metal2 s 13082 0 13138 160 6 Tile_X0Y1_N4END[8]
port 596 nsew signal input
rlabel metal2 s 13358 0 13414 160 6 Tile_X0Y1_N4END[9]
port 597 nsew signal input
rlabel metal2 s 15290 0 15346 160 6 Tile_X0Y1_NN4END[0]
port 598 nsew signal input
rlabel metal2 s 18050 0 18106 160 6 Tile_X0Y1_NN4END[10]
port 599 nsew signal input
rlabel metal2 s 18326 0 18382 160 6 Tile_X0Y1_NN4END[11]
port 600 nsew signal input
rlabel metal2 s 18602 0 18658 160 6 Tile_X0Y1_NN4END[12]
port 601 nsew signal input
rlabel metal2 s 18878 0 18934 160 6 Tile_X0Y1_NN4END[13]
port 602 nsew signal input
rlabel metal2 s 19154 0 19210 160 6 Tile_X0Y1_NN4END[14]
port 603 nsew signal input
rlabel metal2 s 19430 0 19486 160 6 Tile_X0Y1_NN4END[15]
port 604 nsew signal input
rlabel metal2 s 15566 0 15622 160 6 Tile_X0Y1_NN4END[1]
port 605 nsew signal input
rlabel metal2 s 15842 0 15898 160 6 Tile_X0Y1_NN4END[2]
port 606 nsew signal input
rlabel metal2 s 16118 0 16174 160 6 Tile_X0Y1_NN4END[3]
port 607 nsew signal input
rlabel metal2 s 16394 0 16450 160 6 Tile_X0Y1_NN4END[4]
port 608 nsew signal input
rlabel metal2 s 16670 0 16726 160 6 Tile_X0Y1_NN4END[5]
port 609 nsew signal input
rlabel metal2 s 16946 0 17002 160 6 Tile_X0Y1_NN4END[6]
port 610 nsew signal input
rlabel metal2 s 17222 0 17278 160 6 Tile_X0Y1_NN4END[7]
port 611 nsew signal input
rlabel metal2 s 17498 0 17554 160 6 Tile_X0Y1_NN4END[8]
port 612 nsew signal input
rlabel metal2 s 17774 0 17830 160 6 Tile_X0Y1_NN4END[9]
port 613 nsew signal input
rlabel metal2 s 19706 0 19762 160 6 Tile_X0Y1_S1BEG[0]
port 614 nsew signal output
rlabel metal2 s 19982 0 20038 160 6 Tile_X0Y1_S1BEG[1]
port 615 nsew signal output
rlabel metal2 s 20258 0 20314 160 6 Tile_X0Y1_S1BEG[2]
port 616 nsew signal output
rlabel metal2 s 20534 0 20590 160 6 Tile_X0Y1_S1BEG[3]
port 617 nsew signal output
rlabel metal2 s 23018 0 23074 160 6 Tile_X0Y1_S2BEG[0]
port 618 nsew signal output
rlabel metal2 s 23294 0 23350 160 6 Tile_X0Y1_S2BEG[1]
port 619 nsew signal output
rlabel metal2 s 23570 0 23626 160 6 Tile_X0Y1_S2BEG[2]
port 620 nsew signal output
rlabel metal2 s 23846 0 23902 160 6 Tile_X0Y1_S2BEG[3]
port 621 nsew signal output
rlabel metal2 s 24122 0 24178 160 6 Tile_X0Y1_S2BEG[4]
port 622 nsew signal output
rlabel metal2 s 24398 0 24454 160 6 Tile_X0Y1_S2BEG[5]
port 623 nsew signal output
rlabel metal2 s 24674 0 24730 160 6 Tile_X0Y1_S2BEG[6]
port 624 nsew signal output
rlabel metal2 s 24950 0 25006 160 6 Tile_X0Y1_S2BEG[7]
port 625 nsew signal output
rlabel metal2 s 20810 0 20866 160 6 Tile_X0Y1_S2BEGb[0]
port 626 nsew signal output
rlabel metal2 s 21086 0 21142 160 6 Tile_X0Y1_S2BEGb[1]
port 627 nsew signal output
rlabel metal2 s 21362 0 21418 160 6 Tile_X0Y1_S2BEGb[2]
port 628 nsew signal output
rlabel metal2 s 21638 0 21694 160 6 Tile_X0Y1_S2BEGb[3]
port 629 nsew signal output
rlabel metal2 s 21914 0 21970 160 6 Tile_X0Y1_S2BEGb[4]
port 630 nsew signal output
rlabel metal2 s 22190 0 22246 160 6 Tile_X0Y1_S2BEGb[5]
port 631 nsew signal output
rlabel metal2 s 22466 0 22522 160 6 Tile_X0Y1_S2BEGb[6]
port 632 nsew signal output
rlabel metal2 s 22742 0 22798 160 6 Tile_X0Y1_S2BEGb[7]
port 633 nsew signal output
rlabel metal2 s 25226 0 25282 160 6 Tile_X0Y1_S4BEG[0]
port 634 nsew signal output
rlabel metal2 s 27986 0 28042 160 6 Tile_X0Y1_S4BEG[10]
port 635 nsew signal output
rlabel metal2 s 28262 0 28318 160 6 Tile_X0Y1_S4BEG[11]
port 636 nsew signal output
rlabel metal2 s 28538 0 28594 160 6 Tile_X0Y1_S4BEG[12]
port 637 nsew signal output
rlabel metal2 s 28814 0 28870 160 6 Tile_X0Y1_S4BEG[13]
port 638 nsew signal output
rlabel metal2 s 29090 0 29146 160 6 Tile_X0Y1_S4BEG[14]
port 639 nsew signal output
rlabel metal2 s 29366 0 29422 160 6 Tile_X0Y1_S4BEG[15]
port 640 nsew signal output
rlabel metal2 s 25502 0 25558 160 6 Tile_X0Y1_S4BEG[1]
port 641 nsew signal output
rlabel metal2 s 25778 0 25834 160 6 Tile_X0Y1_S4BEG[2]
port 642 nsew signal output
rlabel metal2 s 26054 0 26110 160 6 Tile_X0Y1_S4BEG[3]
port 643 nsew signal output
rlabel metal2 s 26330 0 26386 160 6 Tile_X0Y1_S4BEG[4]
port 644 nsew signal output
rlabel metal2 s 26606 0 26662 160 6 Tile_X0Y1_S4BEG[5]
port 645 nsew signal output
rlabel metal2 s 26882 0 26938 160 6 Tile_X0Y1_S4BEG[6]
port 646 nsew signal output
rlabel metal2 s 27158 0 27214 160 6 Tile_X0Y1_S4BEG[7]
port 647 nsew signal output
rlabel metal2 s 27434 0 27490 160 6 Tile_X0Y1_S4BEG[8]
port 648 nsew signal output
rlabel metal2 s 27710 0 27766 160 6 Tile_X0Y1_S4BEG[9]
port 649 nsew signal output
rlabel metal2 s 29642 0 29698 160 6 Tile_X0Y1_SS4BEG[0]
port 650 nsew signal output
rlabel metal2 s 32402 0 32458 160 6 Tile_X0Y1_SS4BEG[10]
port 651 nsew signal output
rlabel metal2 s 32678 0 32734 160 6 Tile_X0Y1_SS4BEG[11]
port 652 nsew signal output
rlabel metal2 s 32954 0 33010 160 6 Tile_X0Y1_SS4BEG[12]
port 653 nsew signal output
rlabel metal2 s 33230 0 33286 160 6 Tile_X0Y1_SS4BEG[13]
port 654 nsew signal output
rlabel metal2 s 33506 0 33562 160 6 Tile_X0Y1_SS4BEG[14]
port 655 nsew signal output
rlabel metal2 s 33782 0 33838 160 6 Tile_X0Y1_SS4BEG[15]
port 656 nsew signal output
rlabel metal2 s 29918 0 29974 160 6 Tile_X0Y1_SS4BEG[1]
port 657 nsew signal output
rlabel metal2 s 30194 0 30250 160 6 Tile_X0Y1_SS4BEG[2]
port 658 nsew signal output
rlabel metal2 s 30470 0 30526 160 6 Tile_X0Y1_SS4BEG[3]
port 659 nsew signal output
rlabel metal2 s 30746 0 30802 160 6 Tile_X0Y1_SS4BEG[4]
port 660 nsew signal output
rlabel metal2 s 31022 0 31078 160 6 Tile_X0Y1_SS4BEG[5]
port 661 nsew signal output
rlabel metal2 s 31298 0 31354 160 6 Tile_X0Y1_SS4BEG[6]
port 662 nsew signal output
rlabel metal2 s 31574 0 31630 160 6 Tile_X0Y1_SS4BEG[7]
port 663 nsew signal output
rlabel metal2 s 31850 0 31906 160 6 Tile_X0Y1_SS4BEG[8]
port 664 nsew signal output
rlabel metal2 s 32126 0 32182 160 6 Tile_X0Y1_SS4BEG[9]
port 665 nsew signal output
rlabel metal2 s 34058 0 34114 160 6 Tile_X0Y1_UserCLK
port 666 nsew signal input
rlabel metal3 s 0 4632 160 4752 6 Tile_X0Y1_W1BEG[0]
port 667 nsew signal output
rlabel metal3 s 0 4904 160 5024 6 Tile_X0Y1_W1BEG[1]
port 668 nsew signal output
rlabel metal3 s 0 5176 160 5296 6 Tile_X0Y1_W1BEG[2]
port 669 nsew signal output
rlabel metal3 s 0 5448 160 5568 6 Tile_X0Y1_W1BEG[3]
port 670 nsew signal output
rlabel metal3 s 44840 4632 45000 4752 6 Tile_X0Y1_W1END[0]
port 671 nsew signal input
rlabel metal3 s 44840 4904 45000 5024 6 Tile_X0Y1_W1END[1]
port 672 nsew signal input
rlabel metal3 s 44840 5176 45000 5296 6 Tile_X0Y1_W1END[2]
port 673 nsew signal input
rlabel metal3 s 44840 5448 45000 5568 6 Tile_X0Y1_W1END[3]
port 674 nsew signal input
rlabel metal3 s 0 5720 160 5840 6 Tile_X0Y1_W2BEG[0]
port 675 nsew signal output
rlabel metal3 s 0 5992 160 6112 6 Tile_X0Y1_W2BEG[1]
port 676 nsew signal output
rlabel metal3 s 0 6264 160 6384 6 Tile_X0Y1_W2BEG[2]
port 677 nsew signal output
rlabel metal3 s 0 6536 160 6656 6 Tile_X0Y1_W2BEG[3]
port 678 nsew signal output
rlabel metal3 s 0 6808 160 6928 6 Tile_X0Y1_W2BEG[4]
port 679 nsew signal output
rlabel metal3 s 0 7080 160 7200 6 Tile_X0Y1_W2BEG[5]
port 680 nsew signal output
rlabel metal3 s 0 7352 160 7472 6 Tile_X0Y1_W2BEG[6]
port 681 nsew signal output
rlabel metal3 s 0 7624 160 7744 6 Tile_X0Y1_W2BEG[7]
port 682 nsew signal output
rlabel metal3 s 0 7896 160 8016 6 Tile_X0Y1_W2BEGb[0]
port 683 nsew signal output
rlabel metal3 s 0 8168 160 8288 6 Tile_X0Y1_W2BEGb[1]
port 684 nsew signal output
rlabel metal3 s 0 8440 160 8560 6 Tile_X0Y1_W2BEGb[2]
port 685 nsew signal output
rlabel metal3 s 0 8712 160 8832 6 Tile_X0Y1_W2BEGb[3]
port 686 nsew signal output
rlabel metal3 s 0 8984 160 9104 6 Tile_X0Y1_W2BEGb[4]
port 687 nsew signal output
rlabel metal3 s 0 9256 160 9376 6 Tile_X0Y1_W2BEGb[5]
port 688 nsew signal output
rlabel metal3 s 0 9528 160 9648 6 Tile_X0Y1_W2BEGb[6]
port 689 nsew signal output
rlabel metal3 s 0 9800 160 9920 6 Tile_X0Y1_W2BEGb[7]
port 690 nsew signal output
rlabel metal3 s 44840 7896 45000 8016 6 Tile_X0Y1_W2END[0]
port 691 nsew signal input
rlabel metal3 s 44840 8168 45000 8288 6 Tile_X0Y1_W2END[1]
port 692 nsew signal input
rlabel metal3 s 44840 8440 45000 8560 6 Tile_X0Y1_W2END[2]
port 693 nsew signal input
rlabel metal3 s 44840 8712 45000 8832 6 Tile_X0Y1_W2END[3]
port 694 nsew signal input
rlabel metal3 s 44840 8984 45000 9104 6 Tile_X0Y1_W2END[4]
port 695 nsew signal input
rlabel metal3 s 44840 9256 45000 9376 6 Tile_X0Y1_W2END[5]
port 696 nsew signal input
rlabel metal3 s 44840 9528 45000 9648 6 Tile_X0Y1_W2END[6]
port 697 nsew signal input
rlabel metal3 s 44840 9800 45000 9920 6 Tile_X0Y1_W2END[7]
port 698 nsew signal input
rlabel metal3 s 44840 5720 45000 5840 6 Tile_X0Y1_W2MID[0]
port 699 nsew signal input
rlabel metal3 s 44840 5992 45000 6112 6 Tile_X0Y1_W2MID[1]
port 700 nsew signal input
rlabel metal3 s 44840 6264 45000 6384 6 Tile_X0Y1_W2MID[2]
port 701 nsew signal input
rlabel metal3 s 44840 6536 45000 6656 6 Tile_X0Y1_W2MID[3]
port 702 nsew signal input
rlabel metal3 s 44840 6808 45000 6928 6 Tile_X0Y1_W2MID[4]
port 703 nsew signal input
rlabel metal3 s 44840 7080 45000 7200 6 Tile_X0Y1_W2MID[5]
port 704 nsew signal input
rlabel metal3 s 44840 7352 45000 7472 6 Tile_X0Y1_W2MID[6]
port 705 nsew signal input
rlabel metal3 s 44840 7624 45000 7744 6 Tile_X0Y1_W2MID[7]
port 706 nsew signal input
rlabel metal3 s 0 14424 160 14544 6 Tile_X0Y1_W6BEG[0]
port 707 nsew signal output
rlabel metal3 s 0 17144 160 17264 6 Tile_X0Y1_W6BEG[10]
port 708 nsew signal output
rlabel metal3 s 0 17416 160 17536 6 Tile_X0Y1_W6BEG[11]
port 709 nsew signal output
rlabel metal3 s 0 14696 160 14816 6 Tile_X0Y1_W6BEG[1]
port 710 nsew signal output
rlabel metal3 s 0 14968 160 15088 6 Tile_X0Y1_W6BEG[2]
port 711 nsew signal output
rlabel metal3 s 0 15240 160 15360 6 Tile_X0Y1_W6BEG[3]
port 712 nsew signal output
rlabel metal3 s 0 15512 160 15632 6 Tile_X0Y1_W6BEG[4]
port 713 nsew signal output
rlabel metal3 s 0 15784 160 15904 6 Tile_X0Y1_W6BEG[5]
port 714 nsew signal output
rlabel metal3 s 0 16056 160 16176 6 Tile_X0Y1_W6BEG[6]
port 715 nsew signal output
rlabel metal3 s 0 16328 160 16448 6 Tile_X0Y1_W6BEG[7]
port 716 nsew signal output
rlabel metal3 s 0 16600 160 16720 6 Tile_X0Y1_W6BEG[8]
port 717 nsew signal output
rlabel metal3 s 0 16872 160 16992 6 Tile_X0Y1_W6BEG[9]
port 718 nsew signal output
rlabel metal3 s 44840 14424 45000 14544 6 Tile_X0Y1_W6END[0]
port 719 nsew signal input
rlabel metal3 s 44840 17144 45000 17264 6 Tile_X0Y1_W6END[10]
port 720 nsew signal input
rlabel metal3 s 44840 17416 45000 17536 6 Tile_X0Y1_W6END[11]
port 721 nsew signal input
rlabel metal3 s 44840 14696 45000 14816 6 Tile_X0Y1_W6END[1]
port 722 nsew signal input
rlabel metal3 s 44840 14968 45000 15088 6 Tile_X0Y1_W6END[2]
port 723 nsew signal input
rlabel metal3 s 44840 15240 45000 15360 6 Tile_X0Y1_W6END[3]
port 724 nsew signal input
rlabel metal3 s 44840 15512 45000 15632 6 Tile_X0Y1_W6END[4]
port 725 nsew signal input
rlabel metal3 s 44840 15784 45000 15904 6 Tile_X0Y1_W6END[5]
port 726 nsew signal input
rlabel metal3 s 44840 16056 45000 16176 6 Tile_X0Y1_W6END[6]
port 727 nsew signal input
rlabel metal3 s 44840 16328 45000 16448 6 Tile_X0Y1_W6END[7]
port 728 nsew signal input
rlabel metal3 s 44840 16600 45000 16720 6 Tile_X0Y1_W6END[8]
port 729 nsew signal input
rlabel metal3 s 44840 16872 45000 16992 6 Tile_X0Y1_W6END[9]
port 730 nsew signal input
rlabel metal3 s 0 10072 160 10192 6 Tile_X0Y1_WW4BEG[0]
port 731 nsew signal output
rlabel metal3 s 0 12792 160 12912 6 Tile_X0Y1_WW4BEG[10]
port 732 nsew signal output
rlabel metal3 s 0 13064 160 13184 6 Tile_X0Y1_WW4BEG[11]
port 733 nsew signal output
rlabel metal3 s 0 13336 160 13456 6 Tile_X0Y1_WW4BEG[12]
port 734 nsew signal output
rlabel metal3 s 0 13608 160 13728 6 Tile_X0Y1_WW4BEG[13]
port 735 nsew signal output
rlabel metal3 s 0 13880 160 14000 6 Tile_X0Y1_WW4BEG[14]
port 736 nsew signal output
rlabel metal3 s 0 14152 160 14272 6 Tile_X0Y1_WW4BEG[15]
port 737 nsew signal output
rlabel metal3 s 0 10344 160 10464 6 Tile_X0Y1_WW4BEG[1]
port 738 nsew signal output
rlabel metal3 s 0 10616 160 10736 6 Tile_X0Y1_WW4BEG[2]
port 739 nsew signal output
rlabel metal3 s 0 10888 160 11008 6 Tile_X0Y1_WW4BEG[3]
port 740 nsew signal output
rlabel metal3 s 0 11160 160 11280 6 Tile_X0Y1_WW4BEG[4]
port 741 nsew signal output
rlabel metal3 s 0 11432 160 11552 6 Tile_X0Y1_WW4BEG[5]
port 742 nsew signal output
rlabel metal3 s 0 11704 160 11824 6 Tile_X0Y1_WW4BEG[6]
port 743 nsew signal output
rlabel metal3 s 0 11976 160 12096 6 Tile_X0Y1_WW4BEG[7]
port 744 nsew signal output
rlabel metal3 s 0 12248 160 12368 6 Tile_X0Y1_WW4BEG[8]
port 745 nsew signal output
rlabel metal3 s 0 12520 160 12640 6 Tile_X0Y1_WW4BEG[9]
port 746 nsew signal output
rlabel metal3 s 44840 10072 45000 10192 6 Tile_X0Y1_WW4END[0]
port 747 nsew signal input
rlabel metal3 s 44840 12792 45000 12912 6 Tile_X0Y1_WW4END[10]
port 748 nsew signal input
rlabel metal3 s 44840 13064 45000 13184 6 Tile_X0Y1_WW4END[11]
port 749 nsew signal input
rlabel metal3 s 44840 13336 45000 13456 6 Tile_X0Y1_WW4END[12]
port 750 nsew signal input
rlabel metal3 s 44840 13608 45000 13728 6 Tile_X0Y1_WW4END[13]
port 751 nsew signal input
rlabel metal3 s 44840 13880 45000 14000 6 Tile_X0Y1_WW4END[14]
port 752 nsew signal input
rlabel metal3 s 44840 14152 45000 14272 6 Tile_X0Y1_WW4END[15]
port 753 nsew signal input
rlabel metal3 s 44840 10344 45000 10464 6 Tile_X0Y1_WW4END[1]
port 754 nsew signal input
rlabel metal3 s 44840 10616 45000 10736 6 Tile_X0Y1_WW4END[2]
port 755 nsew signal input
rlabel metal3 s 44840 10888 45000 11008 6 Tile_X0Y1_WW4END[3]
port 756 nsew signal input
rlabel metal3 s 44840 11160 45000 11280 6 Tile_X0Y1_WW4END[4]
port 757 nsew signal input
rlabel metal3 s 44840 11432 45000 11552 6 Tile_X0Y1_WW4END[5]
port 758 nsew signal input
rlabel metal3 s 44840 11704 45000 11824 6 Tile_X0Y1_WW4END[6]
port 759 nsew signal input
rlabel metal3 s 44840 11976 45000 12096 6 Tile_X0Y1_WW4END[7]
port 760 nsew signal input
rlabel metal3 s 44840 12248 45000 12368 6 Tile_X0Y1_WW4END[8]
port 761 nsew signal input
rlabel metal3 s 44840 12520 45000 12640 6 Tile_X0Y1_WW4END[9]
port 762 nsew signal input
rlabel metal4 s 19568 1040 19888 89264 6 VGND
port 763 nsew ground bidirectional
rlabel metal4 s 4208 1040 4528 89264 6 VPWR
port 764 nsew power bidirectional
rlabel metal4 s 34928 1040 35248 89264 6 VPWR
port 764 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 45000 90800
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13985226
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/DSP/runs/24_12_05_16_33/results/signoff/DSP.magic.gds
string GDS_START 1116864
<< end >>

