magic
tech sky130A
magscale 1 2
timestamp 1733529900
<< viali >>
rect 1593 8585 1627 8619
rect 2421 8585 2455 8619
rect 3985 8585 4019 8619
rect 4813 8585 4847 8619
rect 6009 8585 6043 8619
rect 6377 8585 6411 8619
rect 7389 8585 7423 8619
rect 8217 8585 8251 8619
rect 9597 8585 9631 8619
rect 10793 8585 10827 8619
rect 10977 8585 11011 8619
rect 11989 8585 12023 8619
rect 13185 8585 13219 8619
rect 13369 8585 13403 8619
rect 14381 8585 14415 8619
rect 15393 8585 15427 8619
rect 17233 8585 17267 8619
rect 17785 8585 17819 8619
rect 19441 8585 19475 8619
rect 20361 8585 20395 8619
rect 21557 8585 21591 8619
rect 22753 8585 22787 8619
rect 23949 8585 23983 8619
rect 6929 8517 6963 8551
rect 7297 8517 7331 8551
rect 16773 8517 16807 8551
rect 1501 8449 1535 8483
rect 2237 8449 2271 8483
rect 3801 8449 3835 8483
rect 4629 8449 4663 8483
rect 5825 8449 5859 8483
rect 6561 8449 6595 8483
rect 7573 8449 7607 8483
rect 8125 8449 8159 8483
rect 9413 8449 9447 8483
rect 10609 8449 10643 8483
rect 11161 8449 11195 8483
rect 11805 8449 11839 8483
rect 13001 8449 13035 8483
rect 13553 8449 13587 8483
rect 14197 8449 14231 8483
rect 15301 8449 15335 8483
rect 17417 8449 17451 8483
rect 17693 8449 17727 8483
rect 19349 8449 19383 8483
rect 20177 8449 20211 8483
rect 21373 8449 21407 8483
rect 22569 8449 22603 8483
rect 23121 8449 23155 8483
rect 23673 8449 23707 8483
rect 23765 8449 23799 8483
rect 16957 8313 16991 8347
rect 22937 8313 22971 8347
rect 23489 8313 23523 8347
rect 6101 8041 6135 8075
rect 7297 8041 7331 8075
rect 11161 8041 11195 8075
rect 13645 8041 13679 8075
rect 17233 8041 17267 8075
rect 22753 8041 22787 8075
rect 23489 8041 23523 8075
rect 24133 8041 24167 8075
rect 13369 7973 13403 8007
rect 16957 7973 16991 8007
rect 6285 7837 6319 7871
rect 7481 7837 7515 7871
rect 11069 7837 11103 7871
rect 11345 7837 11379 7871
rect 13553 7837 13587 7871
rect 13829 7837 13863 7871
rect 17141 7837 17175 7871
rect 17417 7837 17451 7871
rect 22937 7837 22971 7871
rect 23213 7837 23247 7871
rect 23673 7837 23707 7871
rect 23857 7769 23891 7803
rect 10885 7701 10919 7735
rect 23029 7701 23063 7735
rect 6377 7497 6411 7531
rect 7389 7497 7423 7531
rect 24041 7497 24075 7531
rect 6561 7361 6595 7395
rect 7573 7361 7607 7395
rect 7941 7361 7975 7395
rect 24225 7361 24259 7395
rect 6929 7157 6963 7191
rect 14473 5865 14507 5899
rect 19441 5797 19475 5831
rect 14657 5661 14691 5695
rect 19257 5661 19291 5695
rect 19901 5593 19935 5627
rect 19993 5525 20027 5559
rect 11897 5321 11931 5355
rect 12173 5321 12207 5355
rect 14657 5321 14691 5355
rect 14933 5321 14967 5355
rect 19441 5321 19475 5355
rect 12081 5185 12115 5219
rect 12357 5185 12391 5219
rect 14841 5185 14875 5219
rect 15117 5185 15151 5219
rect 19625 5185 19659 5219
rect 12173 4777 12207 4811
rect 19809 4777 19843 4811
rect 12357 4573 12391 4607
rect 19993 4573 20027 4607
rect 8585 4097 8619 4131
rect 8861 4097 8895 4131
rect 9689 4097 9723 4131
rect 24317 4097 24351 4131
rect 8401 3961 8435 3995
rect 8677 3961 8711 3995
rect 9505 3961 9539 3995
rect 24133 3893 24167 3927
rect 8953 3689 8987 3723
rect 9781 3689 9815 3723
rect 23397 3689 23431 3723
rect 23673 3689 23707 3723
rect 23765 3689 23799 3723
rect 20269 3621 20303 3655
rect 9137 3485 9171 3519
rect 9965 3485 9999 3519
rect 10241 3485 10275 3519
rect 20085 3485 20119 3519
rect 23213 3485 23247 3519
rect 23489 3485 23523 3519
rect 23949 3485 23983 3519
rect 24225 3485 24259 3519
rect 9505 3417 9539 3451
rect 10057 3349 10091 3383
rect 24041 3349 24075 3383
rect 2421 3145 2455 3179
rect 20361 3145 20395 3179
rect 22937 3145 22971 3179
rect 23581 3145 23615 3179
rect 1593 3009 1627 3043
rect 1869 3009 1903 3043
rect 2145 3009 2179 3043
rect 2237 3009 2271 3043
rect 20085 3009 20119 3043
rect 20545 3009 20579 3043
rect 22661 3009 22695 3043
rect 22753 3009 22787 3043
rect 23213 3009 23247 3043
rect 23489 3009 23523 3043
rect 23765 3009 23799 3043
rect 24041 3009 24075 3043
rect 24317 3009 24351 3043
rect 20269 2873 20303 2907
rect 23857 2873 23891 2907
rect 1409 2805 1443 2839
rect 1685 2805 1719 2839
rect 1961 2805 1995 2839
rect 22477 2805 22511 2839
rect 23029 2805 23063 2839
rect 23305 2805 23339 2839
rect 24133 2805 24167 2839
rect 9689 2601 9723 2635
rect 11253 2601 11287 2635
rect 17141 2601 17175 2635
rect 17877 2601 17911 2635
rect 19257 2601 19291 2635
rect 20361 2601 20395 2635
rect 21097 2601 21131 2635
rect 22109 2601 22143 2635
rect 23029 2601 23063 2635
rect 23305 2601 23339 2635
rect 23765 2601 23799 2635
rect 1593 2533 1627 2567
rect 2145 2533 2179 2567
rect 12633 2533 12667 2567
rect 17509 2533 17543 2567
rect 20913 2533 20947 2567
rect 22661 2533 22695 2567
rect 23857 2533 23891 2567
rect 1409 2397 1443 2431
rect 1869 2397 1903 2431
rect 1961 2397 1995 2431
rect 2421 2397 2455 2431
rect 2697 2397 2731 2431
rect 4905 2397 4939 2431
rect 5181 2397 5215 2431
rect 5457 2397 5491 2431
rect 6377 2397 6411 2431
rect 9873 2397 9907 2431
rect 10977 2397 11011 2431
rect 11437 2397 11471 2431
rect 11713 2397 11747 2431
rect 11989 2397 12023 2431
rect 12817 2397 12851 2431
rect 13185 2397 13219 2431
rect 13461 2397 13495 2431
rect 15117 2397 15151 2431
rect 15393 2397 15427 2431
rect 15945 2397 15979 2431
rect 16497 2397 16531 2431
rect 16773 2397 16807 2431
rect 17049 2397 17083 2431
rect 17325 2397 17359 2431
rect 17693 2397 17727 2431
rect 18061 2397 18095 2431
rect 18337 2397 18371 2431
rect 18613 2397 18647 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 19717 2397 19751 2431
rect 19993 2397 20027 2431
rect 20269 2397 20303 2431
rect 20545 2397 20579 2431
rect 20729 2397 20763 2431
rect 21281 2397 21315 2431
rect 21557 2397 21591 2431
rect 21833 2397 21867 2431
rect 21925 2397 21959 2431
rect 22385 2397 22419 2431
rect 22477 2397 22511 2431
rect 22937 2397 22971 2431
rect 23213 2397 23247 2431
rect 23489 2397 23523 2431
rect 23581 2397 23615 2431
rect 24041 2397 24075 2431
rect 1685 2261 1719 2295
rect 2237 2261 2271 2295
rect 2513 2261 2547 2295
rect 4721 2261 4755 2295
rect 4997 2261 5031 2295
rect 5273 2261 5307 2295
rect 6561 2261 6595 2295
rect 10793 2261 10827 2295
rect 11529 2261 11563 2295
rect 11805 2261 11839 2295
rect 13001 2261 13035 2295
rect 13277 2261 13311 2295
rect 14933 2261 14967 2295
rect 15209 2261 15243 2295
rect 16129 2261 16163 2295
rect 16313 2261 16347 2295
rect 16589 2261 16623 2295
rect 16865 2261 16899 2295
rect 18153 2261 18187 2295
rect 18429 2261 18463 2295
rect 18705 2261 18739 2295
rect 19533 2261 19567 2295
rect 19809 2261 19843 2295
rect 20085 2261 20119 2295
rect 21373 2261 21407 2295
rect 21649 2261 21683 2295
rect 22201 2261 22235 2295
rect 22753 2261 22787 2295
rect 1777 2057 1811 2091
rect 3433 2057 3467 2091
rect 4261 2057 4295 2091
rect 4537 2057 4571 2091
rect 5457 2057 5491 2091
rect 6653 2057 6687 2091
rect 6929 2057 6963 2091
rect 7573 2057 7607 2091
rect 8125 2057 8159 2091
rect 8953 2057 8987 2091
rect 17417 2057 17451 2091
rect 17693 2057 17727 2091
rect 21097 2057 21131 2091
rect 21833 2057 21867 2091
rect 22109 2057 22143 2091
rect 22661 2057 22695 2091
rect 23489 2057 23523 2091
rect 24041 2057 24075 2091
rect 24317 2057 24351 2091
rect 10425 1989 10459 2023
rect 11989 1989 12023 2023
rect 15853 1989 15887 2023
rect 16957 1989 16991 2023
rect 18061 1989 18095 2023
rect 18613 1989 18647 2023
rect 20269 1989 20303 2023
rect 21005 1989 21039 2023
rect 1593 1921 1627 1955
rect 2053 1921 2087 1955
rect 2145 1921 2179 1955
rect 2789 1921 2823 1955
rect 3065 1921 3099 1955
rect 3341 1921 3375 1955
rect 3617 1921 3651 1955
rect 3893 1921 3927 1955
rect 4169 1921 4203 1955
rect 4445 1921 4479 1955
rect 4721 1921 4755 1955
rect 5181 1921 5215 1955
rect 5641 1921 5675 1955
rect 5917 1921 5951 1955
rect 6193 1921 6227 1955
rect 6469 1921 6503 1955
rect 6745 1921 6779 1955
rect 7205 1921 7239 1955
rect 7481 1921 7515 1955
rect 7757 1921 7791 1955
rect 8033 1921 8067 1955
rect 8309 1921 8343 1955
rect 8585 1921 8619 1955
rect 8861 1921 8895 1955
rect 9137 1921 9171 1955
rect 9413 1921 9447 1955
rect 9689 1921 9723 1955
rect 9965 1921 9999 1955
rect 10241 1921 10275 1955
rect 10977 1921 11011 1955
rect 11529 1921 11563 1955
rect 12633 1921 12667 1955
rect 12817 1921 12851 1955
rect 13645 1921 13679 1955
rect 14013 1921 14047 1955
rect 14289 1921 14323 1955
rect 14473 1921 14507 1955
rect 14841 1921 14875 1955
rect 15393 1921 15427 1955
rect 15669 1921 15703 1955
rect 16497 1921 16531 1955
rect 17601 1921 17635 1955
rect 17877 1921 17911 1955
rect 19165 1921 19199 1955
rect 19717 1921 19751 1955
rect 21649 1921 21683 1955
rect 22017 1921 22051 1955
rect 22293 1921 22327 1955
rect 22569 1921 22603 1955
rect 22845 1921 22879 1955
rect 22937 1921 22971 1955
rect 23397 1921 23431 1955
rect 23673 1921 23707 1955
rect 23949 1921 23983 1955
rect 24225 1921 24259 1955
rect 24501 1921 24535 1955
rect 2605 1785 2639 1819
rect 3985 1785 4019 1819
rect 7021 1785 7055 1819
rect 7849 1785 7883 1819
rect 8401 1785 8435 1819
rect 9229 1785 9263 1819
rect 9505 1785 9539 1819
rect 12449 1785 12483 1819
rect 13461 1785 13495 1819
rect 13829 1785 13863 1819
rect 15485 1785 15519 1819
rect 19349 1785 19383 1819
rect 20453 1785 20487 1819
rect 22385 1785 22419 1819
rect 23121 1785 23155 1819
rect 23213 1785 23247 1819
rect 23765 1785 23799 1819
rect 1869 1717 1903 1751
rect 2329 1717 2363 1751
rect 2881 1717 2915 1751
rect 3157 1717 3191 1751
rect 3709 1717 3743 1751
rect 4997 1717 5031 1751
rect 5733 1717 5767 1751
rect 6009 1717 6043 1751
rect 7297 1717 7331 1751
rect 8677 1717 8711 1751
rect 9781 1717 9815 1751
rect 10057 1717 10091 1751
rect 10517 1717 10551 1751
rect 11069 1717 11103 1751
rect 11713 1717 11747 1751
rect 12081 1717 12115 1751
rect 12909 1717 12943 1751
rect 14105 1717 14139 1751
rect 14657 1717 14691 1751
rect 15025 1717 15059 1751
rect 15209 1717 15243 1751
rect 15945 1717 15979 1751
rect 16313 1717 16347 1751
rect 17049 1717 17083 1751
rect 18153 1717 18187 1751
rect 18705 1717 18739 1751
rect 19809 1717 19843 1751
rect 21465 1717 21499 1751
rect 2881 1513 2915 1547
rect 14289 1513 14323 1547
rect 15393 1513 15427 1547
rect 15945 1513 15979 1547
rect 16865 1513 16899 1547
rect 17417 1513 17451 1547
rect 18521 1513 18555 1547
rect 18889 1513 18923 1547
rect 20545 1513 20579 1547
rect 21833 1513 21867 1547
rect 22109 1513 22143 1547
rect 22661 1513 22695 1547
rect 3157 1445 3191 1479
rect 4353 1445 4387 1479
rect 7113 1445 7147 1479
rect 8309 1445 8343 1479
rect 11069 1377 11103 1411
rect 19625 1377 19659 1411
rect 20177 1377 20211 1411
rect 1501 1309 1535 1343
rect 1961 1309 1995 1343
rect 2237 1309 2271 1343
rect 2513 1309 2547 1343
rect 2789 1309 2823 1343
rect 3065 1309 3099 1343
rect 3341 1309 3375 1343
rect 3617 1309 3651 1343
rect 3801 1309 3835 1343
rect 4077 1309 4111 1343
rect 4537 1309 4571 1343
rect 4629 1309 4663 1343
rect 5089 1309 5123 1343
rect 5181 1309 5215 1343
rect 5641 1309 5675 1343
rect 5733 1309 5767 1343
rect 6193 1309 6227 1343
rect 6377 1309 6411 1343
rect 6837 1309 6871 1343
rect 6929 1309 6963 1343
rect 7389 1309 7423 1343
rect 7665 1309 7699 1343
rect 7757 1309 7791 1343
rect 8217 1309 8251 1343
rect 8493 1309 8527 1343
rect 8769 1309 8803 1343
rect 9229 1309 9263 1343
rect 9505 1309 9539 1343
rect 9597 1309 9631 1343
rect 9965 1309 9999 1343
rect 10333 1309 10367 1343
rect 11713 1309 11747 1343
rect 11805 1309 11839 1343
rect 12909 1309 12943 1343
rect 13277 1309 13311 1343
rect 14657 1309 14691 1343
rect 15853 1309 15887 1343
rect 16497 1309 16531 1343
rect 16773 1309 16807 1343
rect 19073 1309 19107 1343
rect 21649 1309 21683 1343
rect 22017 1309 22051 1343
rect 22293 1309 22327 1343
rect 22569 1309 22603 1343
rect 22845 1309 22879 1343
rect 22937 1309 22971 1343
rect 23397 1309 23431 1343
rect 23489 1309 23523 1343
rect 23765 1309 23799 1343
rect 24225 1309 24259 1343
rect 10793 1241 10827 1275
rect 12265 1241 12299 1275
rect 14197 1241 14231 1275
rect 15301 1241 15335 1275
rect 17325 1241 17359 1275
rect 17877 1241 17911 1275
rect 18429 1241 18463 1275
rect 19349 1241 19383 1275
rect 19901 1241 19935 1275
rect 20453 1241 20487 1275
rect 1685 1173 1719 1207
rect 1777 1173 1811 1207
rect 2053 1173 2087 1207
rect 2329 1173 2363 1207
rect 2605 1173 2639 1207
rect 3433 1173 3467 1207
rect 3985 1173 4019 1207
rect 4261 1173 4295 1207
rect 4813 1173 4847 1207
rect 4905 1173 4939 1207
rect 5365 1173 5399 1207
rect 5457 1173 5491 1207
rect 5917 1173 5951 1207
rect 6009 1173 6043 1207
rect 6561 1173 6595 1207
rect 6653 1173 6687 1207
rect 7205 1173 7239 1207
rect 7481 1173 7515 1207
rect 7941 1173 7975 1207
rect 8033 1173 8067 1207
rect 8585 1173 8619 1207
rect 9045 1173 9079 1207
rect 9321 1173 9355 1207
rect 9781 1173 9815 1207
rect 10149 1173 10183 1207
rect 10517 1173 10551 1207
rect 11529 1173 11563 1207
rect 11989 1173 12023 1207
rect 12357 1173 12391 1207
rect 13093 1173 13127 1207
rect 13461 1173 13495 1207
rect 14841 1173 14875 1207
rect 16313 1173 16347 1207
rect 17969 1173 18003 1207
rect 21097 1173 21131 1207
rect 21465 1173 21499 1207
rect 22385 1173 22419 1207
rect 23121 1173 23155 1207
rect 23213 1173 23247 1207
rect 23673 1173 23707 1207
rect 23949 1173 23983 1207
rect 24041 1173 24075 1207
<< metal1 >>
rect 1104 8730 25000 8752
rect 1104 8678 6884 8730
rect 6936 8678 6948 8730
rect 7000 8678 7012 8730
rect 7064 8678 7076 8730
rect 7128 8678 7140 8730
rect 7192 8678 12818 8730
rect 12870 8678 12882 8730
rect 12934 8678 12946 8730
rect 12998 8678 13010 8730
rect 13062 8678 13074 8730
rect 13126 8678 18752 8730
rect 18804 8678 18816 8730
rect 18868 8678 18880 8730
rect 18932 8678 18944 8730
rect 18996 8678 19008 8730
rect 19060 8678 24686 8730
rect 24738 8678 24750 8730
rect 24802 8678 24814 8730
rect 24866 8678 24878 8730
rect 24930 8678 24942 8730
rect 24994 8678 25000 8730
rect 1104 8656 25000 8678
rect 1210 8576 1216 8628
rect 1268 8616 1274 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1268 8588 1593 8616
rect 1268 8576 1274 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 1581 8579 1639 8585
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 2409 8619 2467 8625
rect 2409 8616 2421 8619
rect 2188 8588 2421 8616
rect 2188 8576 2194 8588
rect 2409 8585 2421 8588
rect 2455 8585 2467 8619
rect 2409 8579 2467 8585
rect 3326 8576 3332 8628
rect 3384 8616 3390 8628
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3384 8588 3985 8616
rect 3384 8576 3390 8588
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 3973 8579 4031 8585
rect 4522 8576 4528 8628
rect 4580 8616 4586 8628
rect 4801 8619 4859 8625
rect 4801 8616 4813 8619
rect 4580 8588 4813 8616
rect 4580 8576 4586 8588
rect 4801 8585 4813 8588
rect 4847 8585 4859 8619
rect 4801 8579 4859 8585
rect 5718 8576 5724 8628
rect 5776 8616 5782 8628
rect 5997 8619 6055 8625
rect 5997 8616 6009 8619
rect 5776 8588 6009 8616
rect 5776 8576 5782 8588
rect 5997 8585 6009 8588
rect 6043 8585 6055 8619
rect 5997 8579 6055 8585
rect 6365 8619 6423 8625
rect 6365 8585 6377 8619
rect 6411 8585 6423 8619
rect 7377 8619 7435 8625
rect 7377 8616 7389 8619
rect 6365 8579 6423 8585
rect 6932 8588 7389 8616
rect 1486 8440 1492 8492
rect 1544 8440 1550 8492
rect 2222 8440 2228 8492
rect 2280 8440 2286 8492
rect 3786 8440 3792 8492
rect 3844 8440 3850 8492
rect 4614 8440 4620 8492
rect 4672 8440 4678 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6380 8480 6408 8579
rect 6932 8557 6960 8588
rect 7377 8585 7389 8588
rect 7423 8585 7435 8619
rect 7377 8579 7435 8585
rect 8202 8576 8208 8628
rect 8260 8576 8266 8628
rect 9306 8576 9312 8628
rect 9364 8616 9370 8628
rect 9585 8619 9643 8625
rect 9585 8616 9597 8619
rect 9364 8588 9597 8616
rect 9364 8576 9370 8588
rect 9585 8585 9597 8588
rect 9631 8585 9643 8619
rect 9585 8579 9643 8585
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 10781 8619 10839 8625
rect 10781 8616 10793 8619
rect 10560 8588 10793 8616
rect 10560 8576 10566 8588
rect 10781 8585 10793 8588
rect 10827 8585 10839 8619
rect 10781 8579 10839 8585
rect 10965 8619 11023 8625
rect 10965 8585 10977 8619
rect 11011 8585 11023 8619
rect 10965 8579 11023 8585
rect 6917 8551 6975 8557
rect 6917 8517 6929 8551
rect 6963 8517 6975 8551
rect 6917 8511 6975 8517
rect 7282 8508 7288 8560
rect 7340 8508 7346 8560
rect 5859 8452 6408 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6546 8440 6552 8492
rect 6604 8440 6610 8492
rect 7558 8440 7564 8492
rect 7616 8440 7622 8492
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8480 8171 8483
rect 8294 8480 8300 8492
rect 8159 8452 8300 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 9490 8480 9496 8492
rect 9447 8452 9496 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8480 10655 8483
rect 10980 8480 11008 8579
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 11977 8619 12035 8625
rect 11977 8616 11989 8619
rect 11756 8588 11989 8616
rect 11756 8576 11762 8588
rect 11977 8585 11989 8588
rect 12023 8585 12035 8619
rect 11977 8579 12035 8585
rect 13170 8576 13176 8628
rect 13228 8576 13234 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8585 13415 8619
rect 13357 8579 13415 8585
rect 10643 8452 11008 8480
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 11146 8440 11152 8492
rect 11204 8440 11210 8492
rect 11790 8440 11796 8492
rect 11848 8440 11854 8492
rect 12989 8483 13047 8489
rect 12989 8449 13001 8483
rect 13035 8480 13047 8483
rect 13372 8480 13400 8579
rect 14090 8576 14096 8628
rect 14148 8616 14154 8628
rect 14369 8619 14427 8625
rect 14369 8616 14381 8619
rect 14148 8588 14381 8616
rect 14148 8576 14154 8588
rect 14369 8585 14381 8588
rect 14415 8585 14427 8619
rect 14369 8579 14427 8585
rect 15378 8576 15384 8628
rect 15436 8576 15442 8628
rect 17221 8619 17279 8625
rect 17221 8616 17233 8619
rect 16776 8588 17233 8616
rect 16776 8557 16804 8588
rect 17221 8585 17233 8588
rect 17267 8585 17279 8619
rect 17221 8579 17279 8585
rect 17770 8576 17776 8628
rect 17828 8576 17834 8628
rect 19150 8576 19156 8628
rect 19208 8616 19214 8628
rect 19429 8619 19487 8625
rect 19429 8616 19441 8619
rect 19208 8588 19441 8616
rect 19208 8576 19214 8588
rect 19429 8585 19441 8588
rect 19475 8585 19487 8619
rect 19429 8579 19487 8585
rect 20070 8576 20076 8628
rect 20128 8616 20134 8628
rect 20349 8619 20407 8625
rect 20349 8616 20361 8619
rect 20128 8588 20361 8616
rect 20128 8576 20134 8588
rect 20349 8585 20361 8588
rect 20395 8585 20407 8619
rect 20349 8579 20407 8585
rect 21266 8576 21272 8628
rect 21324 8616 21330 8628
rect 21545 8619 21603 8625
rect 21545 8616 21557 8619
rect 21324 8588 21557 8616
rect 21324 8576 21330 8588
rect 21545 8585 21557 8588
rect 21591 8585 21603 8619
rect 21545 8579 21603 8585
rect 22462 8576 22468 8628
rect 22520 8616 22526 8628
rect 22741 8619 22799 8625
rect 22741 8616 22753 8619
rect 22520 8588 22753 8616
rect 22520 8576 22526 8588
rect 22741 8585 22753 8588
rect 22787 8585 22799 8619
rect 22741 8579 22799 8585
rect 23658 8576 23664 8628
rect 23716 8616 23722 8628
rect 23937 8619 23995 8625
rect 23937 8616 23949 8619
rect 23716 8588 23949 8616
rect 23716 8576 23722 8588
rect 23937 8585 23949 8588
rect 23983 8585 23995 8619
rect 23937 8579 23995 8585
rect 16761 8551 16819 8557
rect 16761 8517 16773 8551
rect 16807 8517 16819 8551
rect 16761 8511 16819 8517
rect 22066 8520 23612 8548
rect 13035 8452 13400 8480
rect 13035 8449 13047 8452
rect 12989 8443 13047 8449
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 14182 8440 14188 8492
rect 14240 8440 14246 8492
rect 15289 8483 15347 8489
rect 15289 8449 15301 8483
rect 15335 8449 15347 8483
rect 15289 8443 15347 8449
rect 15304 8412 15332 8443
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17678 8440 17684 8492
rect 17736 8440 17742 8492
rect 19150 8440 19156 8492
rect 19208 8480 19214 8492
rect 19337 8483 19395 8489
rect 19337 8480 19349 8483
rect 19208 8452 19349 8480
rect 19208 8440 19214 8452
rect 19337 8449 19349 8452
rect 19383 8449 19395 8483
rect 19337 8443 19395 8449
rect 20165 8483 20223 8489
rect 20165 8449 20177 8483
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 21361 8483 21419 8489
rect 21361 8449 21373 8483
rect 21407 8480 21419 8483
rect 22066 8480 22094 8520
rect 23584 8492 23612 8520
rect 21407 8452 22094 8480
rect 21407 8449 21419 8452
rect 21361 8443 21419 8449
rect 20180 8412 20208 8443
rect 22554 8440 22560 8492
rect 22612 8440 22618 8492
rect 23106 8440 23112 8492
rect 23164 8440 23170 8492
rect 23566 8440 23572 8492
rect 23624 8440 23630 8492
rect 23658 8440 23664 8492
rect 23716 8440 23722 8492
rect 23753 8483 23811 8489
rect 23753 8449 23765 8483
rect 23799 8449 23811 8483
rect 23753 8443 23811 8449
rect 22094 8412 22100 8424
rect 15304 8384 18736 8412
rect 20180 8384 22100 8412
rect 16482 8304 16488 8356
rect 16540 8344 16546 8356
rect 16945 8347 17003 8353
rect 16945 8344 16957 8347
rect 16540 8316 16957 8344
rect 16540 8304 16546 8316
rect 16945 8313 16957 8316
rect 16991 8313 17003 8347
rect 18708 8344 18736 8384
rect 22094 8372 22100 8384
rect 22152 8372 22158 8424
rect 23768 8412 23796 8443
rect 23492 8384 23796 8412
rect 23492 8353 23520 8384
rect 22925 8347 22983 8353
rect 22925 8344 22937 8347
rect 18708 8316 22937 8344
rect 16945 8307 17003 8313
rect 22925 8313 22937 8316
rect 22971 8313 22983 8347
rect 22925 8307 22983 8313
rect 23477 8347 23535 8353
rect 23477 8313 23489 8347
rect 23523 8313 23535 8347
rect 23477 8307 23535 8313
rect 1104 8186 24840 8208
rect 1104 8134 3917 8186
rect 3969 8134 3981 8186
rect 4033 8134 4045 8186
rect 4097 8134 4109 8186
rect 4161 8134 4173 8186
rect 4225 8134 9851 8186
rect 9903 8134 9915 8186
rect 9967 8134 9979 8186
rect 10031 8134 10043 8186
rect 10095 8134 10107 8186
rect 10159 8134 15785 8186
rect 15837 8134 15849 8186
rect 15901 8134 15913 8186
rect 15965 8134 15977 8186
rect 16029 8134 16041 8186
rect 16093 8134 21719 8186
rect 21771 8134 21783 8186
rect 21835 8134 21847 8186
rect 21899 8134 21911 8186
rect 21963 8134 21975 8186
rect 22027 8134 24840 8186
rect 1104 8112 24840 8134
rect 6089 8075 6147 8081
rect 6089 8041 6101 8075
rect 6135 8072 6147 8075
rect 6546 8072 6552 8084
rect 6135 8044 6552 8072
rect 6135 8041 6147 8044
rect 6089 8035 6147 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 7285 8075 7343 8081
rect 7285 8041 7297 8075
rect 7331 8072 7343 8075
rect 7558 8072 7564 8084
rect 7331 8044 7564 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 11146 8032 11152 8084
rect 11204 8032 11210 8084
rect 13538 8032 13544 8084
rect 13596 8072 13602 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13596 8044 13645 8072
rect 13596 8032 13602 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 17221 8075 17279 8081
rect 17221 8041 17233 8075
rect 17267 8072 17279 8075
rect 17402 8072 17408 8084
rect 17267 8044 17408 8072
rect 17267 8041 17279 8044
rect 17221 8035 17279 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 22741 8075 22799 8081
rect 22741 8041 22753 8075
rect 22787 8072 22799 8075
rect 23106 8072 23112 8084
rect 22787 8044 23112 8072
rect 22787 8041 22799 8044
rect 22741 8035 22799 8041
rect 23106 8032 23112 8044
rect 23164 8032 23170 8084
rect 23477 8075 23535 8081
rect 23477 8041 23489 8075
rect 23523 8072 23535 8075
rect 23658 8072 23664 8084
rect 23523 8044 23664 8072
rect 23523 8041 23535 8044
rect 23477 8035 23535 8041
rect 23658 8032 23664 8044
rect 23716 8032 23722 8084
rect 24121 8075 24179 8081
rect 24121 8041 24133 8075
rect 24167 8072 24179 8075
rect 24486 8072 24492 8084
rect 24167 8044 24492 8072
rect 24167 8041 24179 8044
rect 24121 8035 24179 8041
rect 24486 8032 24492 8044
rect 24544 8032 24550 8084
rect 13357 8007 13415 8013
rect 13357 7973 13369 8007
rect 13403 7973 13415 8007
rect 13357 7967 13415 7973
rect 16945 8007 17003 8013
rect 16945 7973 16957 8007
rect 16991 7973 17003 8007
rect 16945 7967 17003 7973
rect 13372 7936 13400 7967
rect 16960 7936 16988 7967
rect 23842 7936 23848 7948
rect 13372 7908 13860 7936
rect 16960 7908 17448 7936
rect 6270 7828 6276 7880
rect 6328 7828 6334 7880
rect 7466 7828 7472 7880
rect 7524 7828 7530 7880
rect 11054 7828 11060 7880
rect 11112 7828 11118 7880
rect 13832 7877 13860 7908
rect 17420 7877 17448 7908
rect 22066 7908 23848 7936
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 13817 7871 13875 7877
rect 13817 7837 13829 7871
rect 13863 7837 13875 7871
rect 13817 7831 13875 7837
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7837 17187 7871
rect 17129 7831 17187 7837
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7837 17463 7871
rect 17405 7831 17463 7837
rect 11348 7800 11376 7831
rect 10888 7772 11376 7800
rect 10888 7741 10916 7772
rect 10873 7735 10931 7741
rect 10873 7701 10885 7735
rect 10919 7701 10931 7735
rect 13556 7732 13584 7831
rect 17144 7800 17172 7831
rect 22066 7800 22094 7908
rect 23842 7896 23848 7908
rect 23900 7896 23906 7948
rect 22925 7871 22983 7877
rect 22925 7837 22937 7871
rect 22971 7868 22983 7871
rect 23201 7871 23259 7877
rect 22971 7840 23060 7868
rect 22971 7837 22983 7840
rect 22925 7831 22983 7837
rect 17144 7772 22094 7800
rect 22186 7732 22192 7744
rect 13556 7704 22192 7732
rect 10873 7695 10931 7701
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 23032 7741 23060 7840
rect 23201 7837 23213 7871
rect 23247 7837 23259 7871
rect 23201 7831 23259 7837
rect 23017 7735 23075 7741
rect 23017 7701 23029 7735
rect 23063 7701 23075 7735
rect 23216 7732 23244 7831
rect 23658 7828 23664 7880
rect 23716 7828 23722 7880
rect 23845 7803 23903 7809
rect 23845 7769 23857 7803
rect 23891 7800 23903 7803
rect 23934 7800 23940 7812
rect 23891 7772 23940 7800
rect 23891 7769 23903 7772
rect 23845 7763 23903 7769
rect 23934 7760 23940 7772
rect 23992 7760 23998 7812
rect 24394 7732 24400 7744
rect 23216 7704 24400 7732
rect 23017 7695 23075 7701
rect 24394 7692 24400 7704
rect 24452 7692 24458 7744
rect 1104 7642 25000 7664
rect 1104 7590 6884 7642
rect 6936 7590 6948 7642
rect 7000 7590 7012 7642
rect 7064 7590 7076 7642
rect 7128 7590 7140 7642
rect 7192 7590 12818 7642
rect 12870 7590 12882 7642
rect 12934 7590 12946 7642
rect 12998 7590 13010 7642
rect 13062 7590 13074 7642
rect 13126 7590 18752 7642
rect 18804 7590 18816 7642
rect 18868 7590 18880 7642
rect 18932 7590 18944 7642
rect 18996 7590 19008 7642
rect 19060 7590 24686 7642
rect 24738 7590 24750 7642
rect 24802 7590 24814 7642
rect 24866 7590 24878 7642
rect 24930 7590 24942 7642
rect 24994 7590 25000 7642
rect 1104 7568 25000 7590
rect 6270 7488 6276 7540
rect 6328 7528 6334 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 6328 7500 6377 7528
rect 6328 7488 6334 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 7377 7531 7435 7537
rect 7377 7497 7389 7531
rect 7423 7528 7435 7531
rect 7466 7528 7472 7540
rect 7423 7500 7472 7528
rect 7423 7497 7435 7500
rect 7377 7491 7435 7497
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 23382 7528 23388 7540
rect 11112 7500 23388 7528
rect 11112 7488 11118 7500
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 23658 7488 23664 7540
rect 23716 7528 23722 7540
rect 24029 7531 24087 7537
rect 24029 7528 24041 7531
rect 23716 7500 24041 7528
rect 23716 7488 23722 7500
rect 24029 7497 24041 7500
rect 24075 7497 24087 7531
rect 24029 7491 24087 7497
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7392 6607 7395
rect 7561 7395 7619 7401
rect 6595 7364 6960 7392
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 6932 7197 6960 7364
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7607 7364 7941 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 7929 7361 7941 7364
rect 7975 7392 7987 7395
rect 23014 7392 23020 7404
rect 7975 7364 23020 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 23014 7352 23020 7364
rect 23072 7352 23078 7404
rect 23198 7352 23204 7404
rect 23256 7392 23262 7404
rect 24213 7395 24271 7401
rect 24213 7392 24225 7395
rect 23256 7364 24225 7392
rect 23256 7352 23262 7364
rect 24213 7361 24225 7364
rect 24259 7361 24271 7395
rect 24213 7355 24271 7361
rect 6917 7191 6975 7197
rect 6917 7157 6929 7191
rect 6963 7188 6975 7191
rect 8202 7188 8208 7200
rect 6963 7160 8208 7188
rect 6963 7157 6975 7160
rect 6917 7151 6975 7157
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 1104 7098 24840 7120
rect 1104 7046 3917 7098
rect 3969 7046 3981 7098
rect 4033 7046 4045 7098
rect 4097 7046 4109 7098
rect 4161 7046 4173 7098
rect 4225 7046 9851 7098
rect 9903 7046 9915 7098
rect 9967 7046 9979 7098
rect 10031 7046 10043 7098
rect 10095 7046 10107 7098
rect 10159 7046 15785 7098
rect 15837 7046 15849 7098
rect 15901 7046 15913 7098
rect 15965 7046 15977 7098
rect 16029 7046 16041 7098
rect 16093 7046 21719 7098
rect 21771 7046 21783 7098
rect 21835 7046 21847 7098
rect 21899 7046 21911 7098
rect 21963 7046 21975 7098
rect 22027 7046 24840 7098
rect 1104 7024 24840 7046
rect 1104 6554 25000 6576
rect 1104 6502 6884 6554
rect 6936 6502 6948 6554
rect 7000 6502 7012 6554
rect 7064 6502 7076 6554
rect 7128 6502 7140 6554
rect 7192 6502 12818 6554
rect 12870 6502 12882 6554
rect 12934 6502 12946 6554
rect 12998 6502 13010 6554
rect 13062 6502 13074 6554
rect 13126 6502 18752 6554
rect 18804 6502 18816 6554
rect 18868 6502 18880 6554
rect 18932 6502 18944 6554
rect 18996 6502 19008 6554
rect 19060 6502 24686 6554
rect 24738 6502 24750 6554
rect 24802 6502 24814 6554
rect 24866 6502 24878 6554
rect 24930 6502 24942 6554
rect 24994 6502 25000 6554
rect 1104 6480 25000 6502
rect 1104 6010 24840 6032
rect 1104 5958 3917 6010
rect 3969 5958 3981 6010
rect 4033 5958 4045 6010
rect 4097 5958 4109 6010
rect 4161 5958 4173 6010
rect 4225 5958 9851 6010
rect 9903 5958 9915 6010
rect 9967 5958 9979 6010
rect 10031 5958 10043 6010
rect 10095 5958 10107 6010
rect 10159 5958 15785 6010
rect 15837 5958 15849 6010
rect 15901 5958 15913 6010
rect 15965 5958 15977 6010
rect 16029 5958 16041 6010
rect 16093 5958 21719 6010
rect 21771 5958 21783 6010
rect 21835 5958 21847 6010
rect 21899 5958 21911 6010
rect 21963 5958 21975 6010
rect 22027 5958 24840 6010
rect 1104 5936 24840 5958
rect 14182 5856 14188 5908
rect 14240 5896 14246 5908
rect 14461 5899 14519 5905
rect 14461 5896 14473 5899
rect 14240 5868 14473 5896
rect 14240 5856 14246 5868
rect 14461 5865 14473 5868
rect 14507 5865 14519 5899
rect 14461 5859 14519 5865
rect 19429 5831 19487 5837
rect 19429 5828 19441 5831
rect 2746 5800 19441 5828
rect 2222 5720 2228 5772
rect 2280 5760 2286 5772
rect 2746 5760 2774 5800
rect 19429 5797 19441 5800
rect 19475 5797 19487 5831
rect 19429 5791 19487 5797
rect 2280 5732 2774 5760
rect 2280 5720 2286 5732
rect 14642 5652 14648 5704
rect 14700 5652 14706 5704
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5692 19303 5695
rect 19426 5692 19432 5704
rect 19291 5664 19432 5692
rect 19291 5661 19303 5664
rect 19245 5655 19303 5661
rect 19426 5652 19432 5664
rect 19484 5652 19490 5704
rect 19889 5627 19947 5633
rect 2746 5596 19564 5624
rect 1486 5516 1492 5568
rect 1544 5556 1550 5568
rect 2746 5556 2774 5596
rect 1544 5528 2774 5556
rect 19536 5556 19564 5596
rect 19889 5593 19901 5627
rect 19935 5624 19947 5627
rect 19935 5596 22094 5624
rect 19935 5593 19947 5596
rect 19889 5587 19947 5593
rect 19981 5559 20039 5565
rect 19981 5556 19993 5559
rect 19536 5528 19993 5556
rect 1544 5516 1550 5528
rect 19981 5525 19993 5528
rect 20027 5525 20039 5559
rect 22066 5556 22094 5596
rect 22462 5556 22468 5568
rect 22066 5528 22468 5556
rect 19981 5519 20039 5525
rect 22462 5516 22468 5528
rect 22520 5516 22526 5568
rect 1104 5466 25000 5488
rect 1104 5414 6884 5466
rect 6936 5414 6948 5466
rect 7000 5414 7012 5466
rect 7064 5414 7076 5466
rect 7128 5414 7140 5466
rect 7192 5414 12818 5466
rect 12870 5414 12882 5466
rect 12934 5414 12946 5466
rect 12998 5414 13010 5466
rect 13062 5414 13074 5466
rect 13126 5414 18752 5466
rect 18804 5414 18816 5466
rect 18868 5414 18880 5466
rect 18932 5414 18944 5466
rect 18996 5414 19008 5466
rect 19060 5414 24686 5466
rect 24738 5414 24750 5466
rect 24802 5414 24814 5466
rect 24866 5414 24878 5466
rect 24930 5414 24942 5466
rect 24994 5414 25000 5466
rect 1104 5392 25000 5414
rect 11790 5312 11796 5364
rect 11848 5352 11854 5364
rect 11885 5355 11943 5361
rect 11885 5352 11897 5355
rect 11848 5324 11897 5352
rect 11848 5312 11854 5324
rect 11885 5321 11897 5324
rect 11931 5321 11943 5355
rect 11885 5315 11943 5321
rect 12161 5355 12219 5361
rect 12161 5321 12173 5355
rect 12207 5321 12219 5355
rect 12161 5315 12219 5321
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5216 12127 5219
rect 12176 5216 12204 5315
rect 14642 5312 14648 5364
rect 14700 5312 14706 5364
rect 14921 5355 14979 5361
rect 14921 5321 14933 5355
rect 14967 5321 14979 5355
rect 14921 5315 14979 5321
rect 12115 5188 12204 5216
rect 12115 5185 12127 5188
rect 12069 5179 12127 5185
rect 12342 5176 12348 5228
rect 12400 5176 12406 5228
rect 14829 5219 14887 5225
rect 14829 5185 14841 5219
rect 14875 5216 14887 5219
rect 14936 5216 14964 5315
rect 19426 5312 19432 5364
rect 19484 5312 19490 5364
rect 14875 5188 14964 5216
rect 15105 5219 15163 5225
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 15105 5185 15117 5219
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 15120 5148 15148 5179
rect 19610 5176 19616 5228
rect 19668 5176 19674 5228
rect 20714 5148 20720 5160
rect 15120 5120 20720 5148
rect 20714 5108 20720 5120
rect 20772 5108 20778 5160
rect 1104 4922 24840 4944
rect 1104 4870 3917 4922
rect 3969 4870 3981 4922
rect 4033 4870 4045 4922
rect 4097 4870 4109 4922
rect 4161 4870 4173 4922
rect 4225 4870 9851 4922
rect 9903 4870 9915 4922
rect 9967 4870 9979 4922
rect 10031 4870 10043 4922
rect 10095 4870 10107 4922
rect 10159 4870 15785 4922
rect 15837 4870 15849 4922
rect 15901 4870 15913 4922
rect 15965 4870 15977 4922
rect 16029 4870 16041 4922
rect 16093 4870 21719 4922
rect 21771 4870 21783 4922
rect 21835 4870 21847 4922
rect 21899 4870 21911 4922
rect 21963 4870 21975 4922
rect 22027 4870 24840 4922
rect 1104 4848 24840 4870
rect 12161 4811 12219 4817
rect 12161 4777 12173 4811
rect 12207 4808 12219 4811
rect 12342 4808 12348 4820
rect 12207 4780 12348 4808
rect 12207 4777 12219 4780
rect 12161 4771 12219 4777
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 19610 4768 19616 4820
rect 19668 4808 19674 4820
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 19668 4780 19809 4808
rect 19668 4768 19674 4780
rect 19797 4777 19809 4780
rect 19843 4777 19855 4811
rect 19797 4771 19855 4777
rect 12360 4613 12480 4620
rect 12345 4607 12480 4613
rect 12345 4573 12357 4607
rect 12391 4592 12480 4607
rect 12391 4573 12403 4592
rect 12345 4567 12403 4573
rect 12452 4536 12480 4592
rect 19981 4607 20039 4613
rect 19981 4573 19993 4607
rect 20027 4604 20039 4607
rect 20990 4604 20996 4616
rect 20027 4576 20996 4604
rect 20027 4573 20039 4576
rect 19981 4567 20039 4573
rect 20990 4564 20996 4576
rect 21048 4564 21054 4616
rect 23658 4536 23664 4548
rect 12452 4508 23664 4536
rect 23658 4496 23664 4508
rect 23716 4496 23722 4548
rect 1104 4378 25000 4400
rect 1104 4326 6884 4378
rect 6936 4326 6948 4378
rect 7000 4326 7012 4378
rect 7064 4326 7076 4378
rect 7128 4326 7140 4378
rect 7192 4326 12818 4378
rect 12870 4326 12882 4378
rect 12934 4326 12946 4378
rect 12998 4326 13010 4378
rect 13062 4326 13074 4378
rect 13126 4326 18752 4378
rect 18804 4326 18816 4378
rect 18868 4326 18880 4378
rect 18932 4326 18944 4378
rect 18996 4326 19008 4378
rect 19060 4326 24686 4378
rect 24738 4326 24750 4378
rect 24802 4326 24814 4378
rect 24866 4326 24878 4378
rect 24930 4326 24942 4378
rect 24994 4326 25000 4378
rect 1104 4304 25000 4326
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4128 8631 4131
rect 8619 4100 8708 4128
rect 8619 4097 8631 4100
rect 8573 4091 8631 4097
rect 8294 4020 8300 4072
rect 8352 4020 8358 4072
rect 8312 3992 8340 4020
rect 8680 4001 8708 4100
rect 8846 4088 8852 4140
rect 8904 4088 8910 4140
rect 9674 4088 9680 4140
rect 9732 4088 9738 4140
rect 24302 4088 24308 4140
rect 24360 4088 24366 4140
rect 8389 3995 8447 4001
rect 8389 3992 8401 3995
rect 8312 3964 8401 3992
rect 8389 3961 8401 3964
rect 8435 3961 8447 3995
rect 8389 3955 8447 3961
rect 8665 3995 8723 4001
rect 8665 3961 8677 3995
rect 8711 3961 8723 3995
rect 8665 3955 8723 3961
rect 9490 3952 9496 4004
rect 9548 3952 9554 4004
rect 24118 3884 24124 3936
rect 24176 3884 24182 3936
rect 1104 3834 24840 3856
rect 1104 3782 3917 3834
rect 3969 3782 3981 3834
rect 4033 3782 4045 3834
rect 4097 3782 4109 3834
rect 4161 3782 4173 3834
rect 4225 3782 9851 3834
rect 9903 3782 9915 3834
rect 9967 3782 9979 3834
rect 10031 3782 10043 3834
rect 10095 3782 10107 3834
rect 10159 3782 15785 3834
rect 15837 3782 15849 3834
rect 15901 3782 15913 3834
rect 15965 3782 15977 3834
rect 16029 3782 16041 3834
rect 16093 3782 21719 3834
rect 21771 3782 21783 3834
rect 21835 3782 21847 3834
rect 21899 3782 21911 3834
rect 21963 3782 21975 3834
rect 22027 3782 24840 3834
rect 1104 3760 24840 3782
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 8904 3692 8953 3720
rect 8904 3680 8910 3692
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 8941 3683 8999 3689
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 9769 3723 9827 3729
rect 9769 3720 9781 3723
rect 9732 3692 9781 3720
rect 9732 3680 9738 3692
rect 9769 3689 9781 3692
rect 9815 3689 9827 3723
rect 9769 3683 9827 3689
rect 23382 3680 23388 3732
rect 23440 3680 23446 3732
rect 23658 3680 23664 3732
rect 23716 3680 23722 3732
rect 23753 3723 23811 3729
rect 23753 3689 23765 3723
rect 23799 3720 23811 3723
rect 24302 3720 24308 3732
rect 23799 3692 24308 3720
rect 23799 3689 23811 3692
rect 23753 3683 23811 3689
rect 24302 3680 24308 3692
rect 24360 3680 24366 3732
rect 3786 3612 3792 3664
rect 3844 3652 3850 3664
rect 20257 3655 20315 3661
rect 20257 3652 20269 3655
rect 3844 3624 20269 3652
rect 3844 3612 3850 3624
rect 20257 3621 20269 3624
rect 20303 3621 20315 3655
rect 20257 3615 20315 3621
rect 23474 3612 23480 3664
rect 23532 3652 23538 3664
rect 25314 3652 25320 3664
rect 23532 3624 25320 3652
rect 23532 3612 23538 3624
rect 25314 3612 25320 3624
rect 25372 3612 25378 3664
rect 23106 3544 23112 3596
rect 23164 3584 23170 3596
rect 24578 3584 24584 3596
rect 23164 3556 24584 3584
rect 23164 3544 23170 3556
rect 24578 3544 24584 3556
rect 24636 3544 24642 3596
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10229 3519 10287 3525
rect 9999 3488 10088 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 9140 3448 9168 3479
rect 9490 3448 9496 3460
rect 9140 3420 9496 3448
rect 9490 3408 9496 3420
rect 9548 3408 9554 3460
rect 10060 3389 10088 3488
rect 10229 3485 10241 3519
rect 10275 3516 10287 3519
rect 13906 3516 13912 3528
rect 10275 3488 13912 3516
rect 10275 3485 10287 3488
rect 10229 3479 10287 3485
rect 13906 3476 13912 3488
rect 13964 3476 13970 3528
rect 20070 3476 20076 3528
rect 20128 3476 20134 3528
rect 22646 3476 22652 3528
rect 22704 3516 22710 3528
rect 23201 3519 23259 3525
rect 23201 3516 23213 3519
rect 22704 3488 23213 3516
rect 22704 3476 22710 3488
rect 23201 3485 23213 3488
rect 23247 3485 23259 3519
rect 23201 3479 23259 3485
rect 23477 3519 23535 3525
rect 23477 3485 23489 3519
rect 23523 3485 23535 3519
rect 23477 3479 23535 3485
rect 23937 3519 23995 3525
rect 23937 3485 23949 3519
rect 23983 3485 23995 3519
rect 23937 3479 23995 3485
rect 24213 3519 24271 3525
rect 24213 3485 24225 3519
rect 24259 3516 24271 3519
rect 24486 3516 24492 3528
rect 24259 3488 24492 3516
rect 24259 3485 24271 3488
rect 24213 3479 24271 3485
rect 22830 3408 22836 3460
rect 22888 3448 22894 3460
rect 23492 3448 23520 3479
rect 22888 3420 23520 3448
rect 23952 3448 23980 3479
rect 24486 3476 24492 3488
rect 24544 3476 24550 3528
rect 25590 3448 25596 3460
rect 23952 3420 25596 3448
rect 22888 3408 22894 3420
rect 25590 3408 25596 3420
rect 25648 3408 25654 3460
rect 10045 3383 10103 3389
rect 10045 3349 10057 3383
rect 10091 3349 10103 3383
rect 10045 3343 10103 3349
rect 23750 3340 23756 3392
rect 23808 3380 23814 3392
rect 24029 3383 24087 3389
rect 24029 3380 24041 3383
rect 23808 3352 24041 3380
rect 23808 3340 23814 3352
rect 24029 3349 24041 3352
rect 24075 3349 24087 3383
rect 24029 3343 24087 3349
rect 1104 3290 25000 3312
rect 1104 3238 6884 3290
rect 6936 3238 6948 3290
rect 7000 3238 7012 3290
rect 7064 3238 7076 3290
rect 7128 3238 7140 3290
rect 7192 3238 12818 3290
rect 12870 3238 12882 3290
rect 12934 3238 12946 3290
rect 12998 3238 13010 3290
rect 13062 3238 13074 3290
rect 13126 3238 18752 3290
rect 18804 3238 18816 3290
rect 18868 3238 18880 3290
rect 18932 3238 18944 3290
rect 18996 3238 19008 3290
rect 19060 3238 24686 3290
rect 24738 3238 24750 3290
rect 24802 3238 24814 3290
rect 24866 3238 24878 3290
rect 24930 3238 24942 3290
rect 24994 3238 25000 3290
rect 1104 3216 25000 3238
rect 2409 3179 2467 3185
rect 2409 3145 2421 3179
rect 2455 3145 2467 3179
rect 2409 3139 2467 3145
rect 750 3068 756 3120
rect 808 3108 814 3120
rect 808 3080 2176 3108
rect 808 3068 814 3080
rect 198 3000 204 3052
rect 256 3040 262 3052
rect 2148 3049 2176 3080
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 256 3012 1593 3040
rect 256 3000 262 3012
rect 1581 3009 1593 3012
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3009 2191 3043
rect 2133 3003 2191 3009
rect 474 2932 480 2984
rect 532 2972 538 2984
rect 1872 2972 1900 3003
rect 2222 3000 2228 3052
rect 2280 3000 2286 3052
rect 532 2944 1900 2972
rect 2424 2972 2452 3139
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 4672 3148 12434 3176
rect 4672 3136 4678 3148
rect 12406 2972 12434 3148
rect 20070 3136 20076 3188
rect 20128 3176 20134 3188
rect 20349 3179 20407 3185
rect 20349 3176 20361 3179
rect 20128 3148 20361 3176
rect 20128 3136 20134 3148
rect 20349 3145 20361 3148
rect 20395 3145 20407 3179
rect 20349 3139 20407 3145
rect 20714 3136 20720 3188
rect 20772 3176 20778 3188
rect 22925 3179 22983 3185
rect 22925 3176 22937 3179
rect 20772 3148 22937 3176
rect 20772 3136 20778 3148
rect 22925 3145 22937 3148
rect 22971 3145 22983 3179
rect 22925 3139 22983 3145
rect 23569 3179 23627 3185
rect 23569 3145 23581 3179
rect 23615 3176 23627 3179
rect 24210 3176 24216 3188
rect 23615 3148 24216 3176
rect 23615 3145 23627 3148
rect 23569 3139 23627 3145
rect 24210 3136 24216 3148
rect 24268 3136 24274 3188
rect 23290 3068 23296 3120
rect 23348 3108 23354 3120
rect 23348 3080 24072 3108
rect 23348 3068 23354 3080
rect 20070 3000 20076 3052
rect 20128 3000 20134 3052
rect 20533 3043 20591 3049
rect 20533 3009 20545 3043
rect 20579 3040 20591 3043
rect 21082 3040 21088 3052
rect 20579 3012 21088 3040
rect 20579 3009 20591 3012
rect 20533 3003 20591 3009
rect 21082 3000 21088 3012
rect 21140 3000 21146 3052
rect 22649 3043 22707 3049
rect 22649 3009 22661 3043
rect 22695 3009 22707 3043
rect 22649 3003 22707 3009
rect 22741 3043 22799 3049
rect 22741 3009 22753 3043
rect 22787 3040 22799 3043
rect 22922 3040 22928 3052
rect 22787 3012 22928 3040
rect 22787 3009 22799 3012
rect 22741 3003 22799 3009
rect 22664 2972 22692 3003
rect 22922 3000 22928 3012
rect 22980 3000 22986 3052
rect 23106 3000 23112 3052
rect 23164 3040 23170 3052
rect 23201 3043 23259 3049
rect 23201 3040 23213 3043
rect 23164 3012 23213 3040
rect 23164 3000 23170 3012
rect 23201 3009 23213 3012
rect 23247 3009 23259 3043
rect 23201 3003 23259 3009
rect 23474 3000 23480 3052
rect 23532 3000 23538 3052
rect 23658 3000 23664 3052
rect 23716 3040 23722 3052
rect 24044 3049 24072 3080
rect 23753 3043 23811 3049
rect 23753 3040 23765 3043
rect 23716 3012 23765 3040
rect 23716 3000 23722 3012
rect 23753 3009 23765 3012
rect 23799 3009 23811 3043
rect 23753 3003 23811 3009
rect 24029 3043 24087 3049
rect 24029 3009 24041 3043
rect 24075 3009 24087 3043
rect 24029 3003 24087 3009
rect 24305 3043 24363 3049
rect 24305 3009 24317 3043
rect 24351 3009 24363 3043
rect 24305 3003 24363 3009
rect 2424 2944 9536 2972
rect 12406 2944 20300 2972
rect 22664 2944 23520 2972
rect 532 2932 538 2944
rect 9398 2904 9404 2916
rect 1964 2876 9404 2904
rect 1397 2839 1455 2845
rect 1397 2805 1409 2839
rect 1443 2836 1455 2839
rect 1578 2836 1584 2848
rect 1443 2808 1584 2836
rect 1443 2805 1455 2808
rect 1397 2799 1455 2805
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 1670 2796 1676 2848
rect 1728 2796 1734 2848
rect 1964 2845 1992 2876
rect 9398 2864 9404 2876
rect 9456 2864 9462 2916
rect 9508 2904 9536 2944
rect 13446 2904 13452 2916
rect 9508 2876 13452 2904
rect 13446 2864 13452 2876
rect 13504 2864 13510 2916
rect 20272 2913 20300 2944
rect 20257 2907 20315 2913
rect 20257 2873 20269 2907
rect 20303 2873 20315 2907
rect 20257 2867 20315 2873
rect 20438 2864 20444 2916
rect 20496 2904 20502 2916
rect 22278 2904 22284 2916
rect 20496 2876 22284 2904
rect 20496 2864 20502 2876
rect 22278 2864 22284 2876
rect 22336 2864 22342 2916
rect 1949 2839 2007 2845
rect 1949 2805 1961 2839
rect 1995 2805 2007 2839
rect 1949 2799 2007 2805
rect 9306 2796 9312 2848
rect 9364 2836 9370 2848
rect 12618 2836 12624 2848
rect 9364 2808 12624 2836
rect 9364 2796 9370 2808
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 19426 2796 19432 2848
rect 19484 2836 19490 2848
rect 22465 2839 22523 2845
rect 22465 2836 22477 2839
rect 19484 2808 22477 2836
rect 19484 2796 19490 2808
rect 22465 2805 22477 2808
rect 22511 2805 22523 2839
rect 22465 2799 22523 2805
rect 23014 2796 23020 2848
rect 23072 2796 23078 2848
rect 23198 2796 23204 2848
rect 23256 2836 23262 2848
rect 23293 2839 23351 2845
rect 23293 2836 23305 2839
rect 23256 2808 23305 2836
rect 23256 2796 23262 2808
rect 23293 2805 23305 2808
rect 23339 2805 23351 2839
rect 23492 2836 23520 2944
rect 23845 2907 23903 2913
rect 23845 2873 23857 2907
rect 23891 2873 23903 2907
rect 23845 2867 23903 2873
rect 23860 2836 23888 2867
rect 23934 2864 23940 2916
rect 23992 2864 23998 2916
rect 24026 2864 24032 2916
rect 24084 2904 24090 2916
rect 24320 2904 24348 3003
rect 24084 2876 24348 2904
rect 24084 2864 24090 2876
rect 23492 2808 23888 2836
rect 23952 2836 23980 2864
rect 24121 2839 24179 2845
rect 24121 2836 24133 2839
rect 23952 2808 24133 2836
rect 23293 2799 23351 2805
rect 24121 2805 24133 2808
rect 24167 2805 24179 2839
rect 24121 2799 24179 2805
rect 1104 2746 24840 2768
rect 1104 2694 3917 2746
rect 3969 2694 3981 2746
rect 4033 2694 4045 2746
rect 4097 2694 4109 2746
rect 4161 2694 4173 2746
rect 4225 2694 9851 2746
rect 9903 2694 9915 2746
rect 9967 2694 9979 2746
rect 10031 2694 10043 2746
rect 10095 2694 10107 2746
rect 10159 2694 15785 2746
rect 15837 2694 15849 2746
rect 15901 2694 15913 2746
rect 15965 2694 15977 2746
rect 16029 2694 16041 2746
rect 16093 2694 21719 2746
rect 21771 2694 21783 2746
rect 21835 2694 21847 2746
rect 21899 2694 21911 2746
rect 21963 2694 21975 2746
rect 22027 2694 24840 2746
rect 1104 2672 24840 2694
rect 1670 2592 1676 2644
rect 1728 2592 1734 2644
rect 2038 2592 2044 2644
rect 2096 2632 2102 2644
rect 9030 2632 9036 2644
rect 2096 2604 9036 2632
rect 2096 2592 2102 2604
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 9677 2635 9735 2641
rect 9677 2632 9689 2635
rect 9600 2604 9689 2632
rect 1486 2524 1492 2576
rect 1544 2564 1550 2576
rect 1581 2567 1639 2573
rect 1581 2564 1593 2567
rect 1544 2536 1593 2564
rect 1544 2524 1550 2536
rect 1581 2533 1593 2536
rect 1627 2533 1639 2567
rect 1581 2527 1639 2533
rect 1688 2496 1716 2592
rect 2133 2567 2191 2573
rect 2133 2533 2145 2567
rect 2179 2564 2191 2567
rect 9306 2564 9312 2576
rect 2179 2536 9312 2564
rect 2179 2533 2191 2536
rect 2133 2527 2191 2533
rect 9306 2524 9312 2536
rect 9364 2524 9370 2576
rect 1688 2468 2452 2496
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1360 2400 1409 2428
rect 1360 2388 1366 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1578 2388 1584 2440
rect 1636 2428 1642 2440
rect 2424 2437 2452 2468
rect 3142 2456 3148 2508
rect 3200 2496 3206 2508
rect 3200 2468 8294 2496
rect 3200 2456 3206 2468
rect 1857 2431 1915 2437
rect 1857 2428 1869 2431
rect 1636 2400 1869 2428
rect 1636 2388 1642 2400
rect 1857 2397 1869 2400
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 1486 2320 1492 2372
rect 1544 2360 1550 2372
rect 1964 2360 1992 2391
rect 2682 2388 2688 2440
rect 2740 2388 2746 2440
rect 4614 2388 4620 2440
rect 4672 2428 4678 2440
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 4672 2400 4905 2428
rect 4672 2388 4678 2400
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 5166 2388 5172 2440
rect 5224 2388 5230 2440
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 6362 2388 6368 2440
rect 6420 2388 6426 2440
rect 8266 2428 8294 2468
rect 9214 2456 9220 2508
rect 9272 2496 9278 2508
rect 9600 2496 9628 2604
rect 9677 2601 9689 2604
rect 9723 2601 9735 2635
rect 9677 2595 9735 2601
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 17129 2635 17187 2641
rect 11287 2604 17080 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 12621 2567 12679 2573
rect 12621 2533 12633 2567
rect 12667 2533 12679 2567
rect 17052 2564 17080 2604
rect 17129 2601 17141 2635
rect 17175 2632 17187 2635
rect 17175 2604 17632 2632
rect 17175 2601 17187 2604
rect 17129 2595 17187 2601
rect 17218 2564 17224 2576
rect 17052 2536 17224 2564
rect 12621 2527 12679 2533
rect 9272 2468 9628 2496
rect 9272 2456 9278 2468
rect 9950 2456 9956 2508
rect 10008 2496 10014 2508
rect 12636 2496 12664 2527
rect 17218 2524 17224 2536
rect 17276 2524 17282 2576
rect 17497 2567 17555 2573
rect 17497 2533 17509 2567
rect 17543 2533 17555 2567
rect 17604 2564 17632 2604
rect 17678 2592 17684 2644
rect 17736 2632 17742 2644
rect 17865 2635 17923 2641
rect 17865 2632 17877 2635
rect 17736 2604 17877 2632
rect 17736 2592 17742 2604
rect 17865 2601 17877 2604
rect 17911 2601 17923 2635
rect 17865 2595 17923 2601
rect 19150 2592 19156 2644
rect 19208 2632 19214 2644
rect 19245 2635 19303 2641
rect 19245 2632 19257 2635
rect 19208 2604 19257 2632
rect 19208 2592 19214 2604
rect 19245 2601 19257 2604
rect 19291 2601 19303 2635
rect 19245 2595 19303 2601
rect 20070 2592 20076 2644
rect 20128 2632 20134 2644
rect 20349 2635 20407 2641
rect 20349 2632 20361 2635
rect 20128 2604 20361 2632
rect 20128 2592 20134 2604
rect 20349 2601 20361 2604
rect 20395 2601 20407 2635
rect 20349 2595 20407 2601
rect 21082 2592 21088 2644
rect 21140 2592 21146 2644
rect 22094 2592 22100 2644
rect 22152 2592 22158 2644
rect 22186 2592 22192 2644
rect 22244 2592 22250 2644
rect 22554 2592 22560 2644
rect 22612 2632 22618 2644
rect 23017 2635 23075 2641
rect 23017 2632 23029 2635
rect 22612 2604 23029 2632
rect 22612 2592 22618 2604
rect 23017 2601 23029 2604
rect 23063 2601 23075 2635
rect 23017 2595 23075 2601
rect 23290 2592 23296 2644
rect 23348 2592 23354 2644
rect 23753 2635 23811 2641
rect 23753 2601 23765 2635
rect 23799 2632 23811 2635
rect 23934 2632 23940 2644
rect 23799 2604 23940 2632
rect 23799 2601 23811 2604
rect 23753 2595 23811 2601
rect 23934 2592 23940 2604
rect 23992 2592 23998 2644
rect 24394 2592 24400 2644
rect 24452 2592 24458 2644
rect 19334 2564 19340 2576
rect 17604 2536 19340 2564
rect 17497 2527 17555 2533
rect 10008 2468 11744 2496
rect 12636 2468 13216 2496
rect 10008 2456 10014 2468
rect 8266 2400 9812 2428
rect 8846 2360 8852 2372
rect 1544 2332 1992 2360
rect 2516 2332 8852 2360
rect 1544 2320 1550 2332
rect 1670 2252 1676 2304
rect 1728 2252 1734 2304
rect 2222 2252 2228 2304
rect 2280 2252 2286 2304
rect 2516 2301 2544 2332
rect 8846 2320 8852 2332
rect 8904 2320 8910 2372
rect 9784 2360 9812 2400
rect 9858 2388 9864 2440
rect 9916 2388 9922 2440
rect 10962 2388 10968 2440
rect 11020 2388 11026 2440
rect 11716 2437 11744 2468
rect 11425 2431 11483 2437
rect 11425 2397 11437 2431
rect 11471 2397 11483 2431
rect 11425 2391 11483 2397
rect 11701 2431 11759 2437
rect 11701 2397 11713 2431
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 10318 2360 10324 2372
rect 9784 2332 10324 2360
rect 10318 2320 10324 2332
rect 10376 2320 10382 2372
rect 11440 2360 11468 2391
rect 11974 2388 11980 2440
rect 12032 2388 12038 2440
rect 12526 2388 12532 2440
rect 12584 2428 12590 2440
rect 13188 2437 13216 2468
rect 13262 2456 13268 2508
rect 13320 2496 13326 2508
rect 13320 2468 15424 2496
rect 13320 2456 13326 2468
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12584 2400 12817 2428
rect 12584 2388 12590 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 13446 2388 13452 2440
rect 13504 2388 13510 2440
rect 15102 2388 15108 2440
rect 15160 2388 15166 2440
rect 15396 2437 15424 2468
rect 15470 2456 15476 2508
rect 15528 2496 15534 2508
rect 17512 2496 17540 2527
rect 19334 2524 19340 2536
rect 19392 2524 19398 2576
rect 19610 2524 19616 2576
rect 19668 2564 19674 2576
rect 20901 2567 20959 2573
rect 20901 2564 20913 2567
rect 19668 2536 20913 2564
rect 19668 2524 19674 2536
rect 20901 2533 20913 2536
rect 20947 2533 20959 2567
rect 22204 2564 22232 2592
rect 22649 2567 22707 2573
rect 22649 2564 22661 2567
rect 22204 2536 22661 2564
rect 20901 2527 20959 2533
rect 22649 2533 22661 2536
rect 22695 2533 22707 2567
rect 22649 2527 22707 2533
rect 22830 2524 22836 2576
rect 22888 2564 22894 2576
rect 23845 2567 23903 2573
rect 23845 2564 23857 2567
rect 22888 2536 23857 2564
rect 22888 2524 22894 2536
rect 23845 2533 23857 2536
rect 23891 2533 23903 2567
rect 23845 2527 23903 2533
rect 20622 2496 20628 2508
rect 15528 2468 16804 2496
rect 17512 2468 18368 2496
rect 15528 2456 15534 2468
rect 15381 2431 15439 2437
rect 15381 2397 15393 2431
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 15933 2431 15991 2437
rect 15933 2397 15945 2431
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 16485 2431 16543 2437
rect 16485 2397 16497 2431
rect 16531 2428 16543 2431
rect 16666 2428 16672 2440
rect 16531 2400 16672 2428
rect 16531 2397 16543 2400
rect 16485 2391 16543 2397
rect 13722 2360 13728 2372
rect 10796 2332 11468 2360
rect 13004 2332 13728 2360
rect 2501 2295 2559 2301
rect 2501 2261 2513 2295
rect 2547 2261 2559 2295
rect 2501 2255 2559 2261
rect 4706 2252 4712 2304
rect 4764 2252 4770 2304
rect 4798 2252 4804 2304
rect 4856 2292 4862 2304
rect 4985 2295 5043 2301
rect 4985 2292 4997 2295
rect 4856 2264 4997 2292
rect 4856 2252 4862 2264
rect 4985 2261 4997 2264
rect 5031 2261 5043 2295
rect 4985 2255 5043 2261
rect 5074 2252 5080 2304
rect 5132 2292 5138 2304
rect 5261 2295 5319 2301
rect 5261 2292 5273 2295
rect 5132 2264 5273 2292
rect 5132 2252 5138 2264
rect 5261 2261 5273 2264
rect 5307 2261 5319 2295
rect 5261 2255 5319 2261
rect 6546 2252 6552 2304
rect 6604 2252 6610 2304
rect 6730 2252 6736 2304
rect 6788 2292 6794 2304
rect 9214 2292 9220 2304
rect 6788 2264 9220 2292
rect 6788 2252 6794 2264
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 10796 2301 10824 2332
rect 10781 2295 10839 2301
rect 10781 2261 10793 2295
rect 10827 2261 10839 2295
rect 10781 2255 10839 2261
rect 11514 2252 11520 2304
rect 11572 2252 11578 2304
rect 11698 2252 11704 2304
rect 11756 2292 11762 2304
rect 13004 2301 13032 2332
rect 13722 2320 13728 2332
rect 13780 2320 13786 2372
rect 15948 2360 15976 2391
rect 16666 2388 16672 2400
rect 16724 2388 16730 2440
rect 16776 2437 16804 2468
rect 16761 2431 16819 2437
rect 16761 2397 16773 2431
rect 16807 2397 16819 2431
rect 16761 2391 16819 2397
rect 16850 2388 16856 2440
rect 16908 2428 16914 2440
rect 18340 2437 18368 2468
rect 19628 2468 20628 2496
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 16908 2400 17049 2428
rect 16908 2388 16914 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17313 2431 17371 2437
rect 17313 2397 17325 2431
rect 17359 2397 17371 2431
rect 17313 2391 17371 2397
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 18325 2431 18383 2437
rect 18325 2397 18337 2431
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 17328 2360 17356 2391
rect 14936 2332 15976 2360
rect 16868 2332 17356 2360
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11756 2264 11805 2292
rect 11756 2252 11762 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 12989 2295 13047 2301
rect 12989 2261 13001 2295
rect 13035 2261 13047 2295
rect 12989 2255 13047 2261
rect 13262 2252 13268 2304
rect 13320 2252 13326 2304
rect 14936 2301 14964 2332
rect 14921 2295 14979 2301
rect 14921 2261 14933 2295
rect 14967 2261 14979 2295
rect 14921 2255 14979 2261
rect 15194 2252 15200 2304
rect 15252 2252 15258 2304
rect 15378 2252 15384 2304
rect 15436 2292 15442 2304
rect 16117 2295 16175 2301
rect 16117 2292 16129 2295
rect 15436 2264 16129 2292
rect 15436 2252 15442 2264
rect 16117 2261 16129 2264
rect 16163 2261 16175 2295
rect 16117 2255 16175 2261
rect 16301 2295 16359 2301
rect 16301 2261 16313 2295
rect 16347 2292 16359 2295
rect 16482 2292 16488 2304
rect 16347 2264 16488 2292
rect 16347 2261 16359 2264
rect 16301 2255 16359 2261
rect 16482 2252 16488 2264
rect 16540 2252 16546 2304
rect 16574 2252 16580 2304
rect 16632 2252 16638 2304
rect 16868 2301 16896 2332
rect 16853 2295 16911 2301
rect 16853 2261 16865 2295
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 17126 2252 17132 2304
rect 17184 2292 17190 2304
rect 17696 2292 17724 2391
rect 18064 2360 18092 2391
rect 18414 2388 18420 2440
rect 18472 2428 18478 2440
rect 18601 2431 18659 2437
rect 18601 2428 18613 2431
rect 18472 2400 18613 2428
rect 18472 2388 18478 2400
rect 18601 2397 18613 2400
rect 18647 2397 18659 2431
rect 18601 2391 18659 2397
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2428 18935 2431
rect 19150 2428 19156 2440
rect 18923 2400 19156 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 19150 2388 19156 2400
rect 19208 2388 19214 2440
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 19628 2360 19656 2468
rect 20622 2456 20628 2468
rect 20680 2456 20686 2508
rect 21634 2456 21640 2508
rect 21692 2496 21698 2508
rect 23382 2496 23388 2508
rect 21692 2468 21956 2496
rect 21692 2456 21698 2468
rect 19705 2431 19763 2437
rect 19705 2397 19717 2431
rect 19751 2428 19763 2431
rect 19886 2428 19892 2440
rect 19751 2400 19892 2428
rect 19751 2397 19763 2400
rect 19705 2391 19763 2397
rect 19886 2388 19892 2400
rect 19944 2388 19950 2440
rect 19978 2388 19984 2440
rect 20036 2388 20042 2440
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 20533 2431 20591 2437
rect 20533 2397 20545 2431
rect 20579 2397 20591 2431
rect 20533 2391 20591 2397
rect 20272 2360 20300 2391
rect 18064 2332 19656 2360
rect 19812 2332 20300 2360
rect 20548 2360 20576 2391
rect 20714 2388 20720 2440
rect 20772 2388 20778 2440
rect 21174 2388 21180 2440
rect 21232 2428 21238 2440
rect 21269 2431 21327 2437
rect 21269 2428 21281 2431
rect 21232 2400 21281 2428
rect 21232 2388 21238 2400
rect 21269 2397 21281 2400
rect 21315 2397 21327 2431
rect 21269 2391 21327 2397
rect 21545 2431 21603 2437
rect 21545 2397 21557 2431
rect 21591 2397 21603 2431
rect 21545 2391 21603 2397
rect 21560 2360 21588 2391
rect 21818 2388 21824 2440
rect 21876 2388 21882 2440
rect 21928 2437 21956 2468
rect 22296 2468 23388 2496
rect 21913 2431 21971 2437
rect 21913 2397 21925 2431
rect 21959 2397 21971 2431
rect 21913 2391 21971 2397
rect 22002 2360 22008 2372
rect 20548 2332 21404 2360
rect 21560 2332 22008 2360
rect 17184 2264 17724 2292
rect 17184 2252 17190 2264
rect 18138 2252 18144 2304
rect 18196 2252 18202 2304
rect 18414 2252 18420 2304
rect 18472 2252 18478 2304
rect 18506 2252 18512 2304
rect 18564 2292 18570 2304
rect 18693 2295 18751 2301
rect 18693 2292 18705 2295
rect 18564 2264 18705 2292
rect 18564 2252 18570 2264
rect 18693 2261 18705 2264
rect 18739 2261 18751 2295
rect 18693 2255 18751 2261
rect 19518 2252 19524 2304
rect 19576 2252 19582 2304
rect 19812 2301 19840 2332
rect 19797 2295 19855 2301
rect 19797 2261 19809 2295
rect 19843 2261 19855 2295
rect 19797 2255 19855 2261
rect 20070 2252 20076 2304
rect 20128 2252 20134 2304
rect 21376 2301 21404 2332
rect 22002 2320 22008 2332
rect 22060 2320 22066 2372
rect 21361 2295 21419 2301
rect 21361 2261 21373 2295
rect 21407 2261 21419 2295
rect 21361 2255 21419 2261
rect 21450 2252 21456 2304
rect 21508 2292 21514 2304
rect 21637 2295 21695 2301
rect 21637 2292 21649 2295
rect 21508 2264 21649 2292
rect 21508 2252 21514 2264
rect 21637 2261 21649 2264
rect 21683 2261 21695 2295
rect 21637 2255 21695 2261
rect 22189 2295 22247 2301
rect 22189 2261 22201 2295
rect 22235 2292 22247 2295
rect 22296 2292 22324 2468
rect 23382 2456 23388 2468
rect 23440 2456 23446 2508
rect 23934 2456 23940 2508
rect 23992 2496 23998 2508
rect 24412 2496 24440 2592
rect 23992 2468 24440 2496
rect 23992 2456 23998 2468
rect 22370 2388 22376 2440
rect 22428 2388 22434 2440
rect 22465 2431 22523 2437
rect 22465 2397 22477 2431
rect 22511 2428 22523 2431
rect 22830 2428 22836 2440
rect 22511 2400 22836 2428
rect 22511 2397 22523 2400
rect 22465 2391 22523 2397
rect 22830 2388 22836 2400
rect 22888 2388 22894 2440
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 22235 2264 22324 2292
rect 22235 2261 22247 2264
rect 22189 2255 22247 2261
rect 22738 2252 22744 2304
rect 22796 2252 22802 2304
rect 22940 2292 22968 2391
rect 23198 2388 23204 2440
rect 23256 2388 23262 2440
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 23492 2360 23520 2391
rect 23566 2388 23572 2440
rect 23624 2388 23630 2440
rect 24029 2431 24087 2437
rect 24029 2397 24041 2431
rect 24075 2428 24087 2431
rect 24302 2428 24308 2440
rect 24075 2400 24308 2428
rect 24075 2397 24087 2400
rect 24029 2391 24087 2397
rect 24302 2388 24308 2400
rect 24360 2388 24366 2440
rect 23750 2360 23756 2372
rect 23492 2332 23756 2360
rect 23750 2320 23756 2332
rect 23808 2320 23814 2372
rect 25038 2292 25044 2304
rect 22940 2264 25044 2292
rect 25038 2252 25044 2264
rect 25096 2252 25102 2304
rect 1104 2202 25000 2224
rect 1104 2150 6884 2202
rect 6936 2150 6948 2202
rect 7000 2150 7012 2202
rect 7064 2150 7076 2202
rect 7128 2150 7140 2202
rect 7192 2150 12818 2202
rect 12870 2150 12882 2202
rect 12934 2150 12946 2202
rect 12998 2150 13010 2202
rect 13062 2150 13074 2202
rect 13126 2150 18752 2202
rect 18804 2150 18816 2202
rect 18868 2150 18880 2202
rect 18932 2150 18944 2202
rect 18996 2150 19008 2202
rect 19060 2150 24686 2202
rect 24738 2150 24750 2202
rect 24802 2150 24814 2202
rect 24866 2150 24878 2202
rect 24930 2150 24942 2202
rect 24994 2150 25000 2202
rect 1104 2128 25000 2150
rect 1670 2048 1676 2100
rect 1728 2048 1734 2100
rect 1765 2091 1823 2097
rect 1765 2057 1777 2091
rect 1811 2088 1823 2091
rect 3421 2091 3479 2097
rect 1811 2060 3280 2088
rect 1811 2057 1823 2060
rect 1765 2051 1823 2057
rect 1578 1912 1584 1964
rect 1636 1912 1642 1964
rect 1688 1884 1716 2048
rect 2222 2020 2228 2032
rect 2056 1992 2228 2020
rect 2056 1961 2084 1992
rect 2222 1980 2228 1992
rect 2280 1980 2286 2032
rect 3142 1980 3148 2032
rect 3200 1980 3206 2032
rect 2041 1955 2099 1961
rect 2041 1921 2053 1955
rect 2087 1921 2099 1955
rect 2041 1915 2099 1921
rect 2133 1955 2191 1961
rect 2133 1921 2145 1955
rect 2179 1921 2191 1955
rect 2682 1952 2688 1964
rect 2133 1915 2191 1921
rect 2240 1924 2688 1952
rect 2148 1884 2176 1915
rect 1688 1856 2176 1884
rect 1026 1776 1032 1828
rect 1084 1816 1090 1828
rect 2240 1816 2268 1924
rect 2682 1912 2688 1924
rect 2740 1912 2746 1964
rect 2774 1912 2780 1964
rect 2832 1912 2838 1964
rect 3050 1912 3056 1964
rect 3108 1912 3114 1964
rect 3160 1884 3188 1980
rect 1084 1788 2268 1816
rect 2332 1856 3188 1884
rect 3252 1884 3280 2060
rect 3421 2057 3433 2091
rect 3467 2057 3479 2091
rect 3421 2051 3479 2057
rect 3329 1955 3387 1961
rect 3329 1921 3341 1955
rect 3375 1952 3387 1955
rect 3436 1952 3464 2051
rect 4246 2048 4252 2100
rect 4304 2048 4310 2100
rect 4525 2091 4583 2097
rect 4525 2057 4537 2091
rect 4571 2057 4583 2091
rect 4525 2051 4583 2057
rect 4540 2020 4568 2051
rect 4706 2048 4712 2100
rect 4764 2088 4770 2100
rect 5445 2091 5503 2097
rect 4764 2060 5304 2088
rect 4764 2048 4770 2060
rect 4540 1992 5212 2020
rect 3375 1924 3464 1952
rect 3375 1921 3387 1924
rect 3329 1915 3387 1921
rect 3602 1912 3608 1964
rect 3660 1912 3666 1964
rect 3878 1912 3884 1964
rect 3936 1912 3942 1964
rect 4157 1955 4215 1961
rect 4157 1921 4169 1955
rect 4203 1952 4215 1955
rect 4338 1952 4344 1964
rect 4203 1924 4344 1952
rect 4203 1921 4215 1924
rect 4157 1915 4215 1921
rect 4338 1912 4344 1924
rect 4396 1912 4402 1964
rect 4430 1912 4436 1964
rect 4488 1912 4494 1964
rect 5184 1961 5212 1992
rect 4709 1955 4767 1961
rect 4709 1952 4721 1955
rect 4540 1924 4721 1952
rect 4540 1884 4568 1924
rect 4709 1921 4721 1924
rect 4755 1921 4767 1955
rect 4709 1915 4767 1921
rect 5169 1955 5227 1961
rect 5169 1921 5181 1955
rect 5215 1921 5227 1955
rect 5276 1952 5304 2060
rect 5445 2057 5457 2091
rect 5491 2057 5503 2091
rect 5445 2051 5503 2057
rect 5460 2020 5488 2051
rect 6638 2048 6644 2100
rect 6696 2048 6702 2100
rect 6917 2091 6975 2097
rect 6917 2057 6929 2091
rect 6963 2088 6975 2091
rect 7374 2088 7380 2100
rect 6963 2060 7380 2088
rect 6963 2057 6975 2060
rect 6917 2051 6975 2057
rect 7374 2048 7380 2060
rect 7432 2048 7438 2100
rect 7561 2091 7619 2097
rect 7561 2057 7573 2091
rect 7607 2088 7619 2091
rect 7926 2088 7932 2100
rect 7607 2060 7932 2088
rect 7607 2057 7619 2060
rect 7561 2051 7619 2057
rect 7926 2048 7932 2060
rect 7984 2048 7990 2100
rect 8110 2048 8116 2100
rect 8168 2048 8174 2100
rect 8938 2048 8944 2100
rect 8996 2048 9002 2100
rect 9214 2048 9220 2100
rect 9272 2088 9278 2100
rect 9674 2088 9680 2100
rect 9272 2060 9680 2088
rect 9272 2048 9278 2060
rect 9674 2048 9680 2060
rect 9732 2048 9738 2100
rect 9784 2060 11100 2088
rect 7282 2020 7288 2032
rect 5460 1992 6224 2020
rect 5629 1955 5687 1961
rect 5629 1952 5641 1955
rect 5276 1924 5641 1952
rect 5169 1915 5227 1921
rect 5629 1921 5641 1924
rect 5675 1921 5687 1955
rect 5629 1915 5687 1921
rect 5902 1912 5908 1964
rect 5960 1912 5966 1964
rect 6196 1961 6224 1992
rect 6748 1992 7288 2020
rect 6181 1955 6239 1961
rect 6181 1921 6193 1955
rect 6227 1921 6239 1955
rect 6181 1915 6239 1921
rect 6454 1912 6460 1964
rect 6512 1912 6518 1964
rect 6748 1961 6776 1992
rect 7282 1980 7288 1992
rect 7340 1980 7346 2032
rect 9784 2020 9812 2060
rect 10413 2023 10471 2029
rect 10413 2020 10425 2023
rect 7392 1992 9812 2020
rect 9876 1992 10425 2020
rect 6733 1955 6791 1961
rect 6733 1921 6745 1955
rect 6779 1921 6791 1955
rect 6733 1915 6791 1921
rect 6822 1912 6828 1964
rect 6880 1912 6886 1964
rect 7193 1955 7251 1961
rect 7193 1952 7205 1955
rect 6932 1924 7205 1952
rect 6840 1884 6868 1912
rect 3252 1856 3832 1884
rect 1084 1776 1090 1788
rect 1857 1751 1915 1757
rect 1857 1717 1869 1751
rect 1903 1748 1915 1751
rect 2038 1748 2044 1760
rect 1903 1720 2044 1748
rect 1903 1717 1915 1720
rect 1857 1711 1915 1717
rect 2038 1708 2044 1720
rect 2096 1708 2102 1760
rect 2332 1757 2360 1856
rect 2593 1819 2651 1825
rect 2593 1785 2605 1819
rect 2639 1816 2651 1819
rect 3510 1816 3516 1828
rect 2639 1788 3516 1816
rect 2639 1785 2651 1788
rect 2593 1779 2651 1785
rect 3510 1776 3516 1788
rect 3568 1776 3574 1828
rect 2317 1751 2375 1757
rect 2317 1717 2329 1751
rect 2363 1717 2375 1751
rect 2317 1711 2375 1717
rect 2682 1708 2688 1760
rect 2740 1748 2746 1760
rect 2869 1751 2927 1757
rect 2869 1748 2881 1751
rect 2740 1720 2881 1748
rect 2740 1708 2746 1720
rect 2869 1717 2881 1720
rect 2915 1717 2927 1751
rect 2869 1711 2927 1717
rect 2958 1708 2964 1760
rect 3016 1748 3022 1760
rect 3145 1751 3203 1757
rect 3145 1748 3157 1751
rect 3016 1720 3157 1748
rect 3016 1708 3022 1720
rect 3145 1717 3157 1720
rect 3191 1717 3203 1751
rect 3145 1711 3203 1717
rect 3234 1708 3240 1760
rect 3292 1748 3298 1760
rect 3697 1751 3755 1757
rect 3697 1748 3709 1751
rect 3292 1720 3709 1748
rect 3292 1708 3298 1720
rect 3697 1717 3709 1720
rect 3743 1717 3755 1751
rect 3804 1748 3832 1856
rect 3988 1856 4568 1884
rect 4816 1856 6868 1884
rect 3988 1825 4016 1856
rect 3973 1819 4031 1825
rect 3973 1785 3985 1819
rect 4019 1785 4031 1819
rect 4816 1816 4844 1856
rect 3973 1779 4031 1785
rect 4632 1788 4844 1816
rect 4632 1748 4660 1788
rect 5626 1776 5632 1828
rect 5684 1816 5690 1828
rect 6932 1816 6960 1924
rect 7193 1921 7205 1924
rect 7239 1921 7251 1955
rect 7392 1952 7420 1992
rect 9876 1964 9904 1992
rect 10413 1989 10425 1992
rect 10459 1989 10471 2023
rect 10413 1983 10471 1989
rect 7193 1915 7251 1921
rect 7300 1924 7420 1952
rect 5684 1788 6960 1816
rect 5684 1776 5690 1788
rect 7006 1776 7012 1828
rect 7064 1776 7070 1828
rect 7300 1816 7328 1924
rect 7466 1912 7472 1964
rect 7524 1912 7530 1964
rect 7745 1955 7803 1961
rect 7745 1952 7757 1955
rect 7576 1924 7757 1952
rect 7576 1896 7604 1924
rect 7745 1921 7757 1924
rect 7791 1921 7803 1955
rect 7745 1915 7803 1921
rect 7834 1912 7840 1964
rect 7892 1952 7898 1964
rect 7892 1924 7972 1952
rect 7892 1912 7898 1924
rect 7558 1844 7564 1896
rect 7616 1844 7622 1896
rect 7208 1788 7328 1816
rect 3804 1720 4660 1748
rect 3697 1711 3755 1717
rect 4706 1708 4712 1760
rect 4764 1748 4770 1760
rect 4985 1751 5043 1757
rect 4985 1748 4997 1751
rect 4764 1720 4997 1748
rect 4764 1708 4770 1720
rect 4985 1717 4997 1720
rect 5031 1717 5043 1751
rect 4985 1711 5043 1717
rect 5534 1708 5540 1760
rect 5592 1748 5598 1760
rect 5721 1751 5779 1757
rect 5721 1748 5733 1751
rect 5592 1720 5733 1748
rect 5592 1708 5598 1720
rect 5721 1717 5733 1720
rect 5767 1717 5779 1751
rect 5721 1711 5779 1717
rect 5997 1751 6055 1757
rect 5997 1717 6009 1751
rect 6043 1748 6055 1751
rect 7208 1748 7236 1788
rect 7834 1776 7840 1828
rect 7892 1776 7898 1828
rect 7944 1816 7972 1924
rect 8018 1912 8024 1964
rect 8076 1912 8082 1964
rect 8294 1912 8300 1964
rect 8352 1912 8358 1964
rect 8570 1912 8576 1964
rect 8628 1912 8634 1964
rect 8846 1912 8852 1964
rect 8904 1912 8910 1964
rect 9122 1912 9128 1964
rect 9180 1912 9186 1964
rect 9398 1912 9404 1964
rect 9456 1912 9462 1964
rect 9677 1955 9735 1961
rect 9677 1921 9689 1955
rect 9723 1952 9735 1955
rect 9766 1952 9772 1964
rect 9723 1924 9772 1952
rect 9723 1921 9735 1924
rect 9677 1915 9735 1921
rect 9766 1912 9772 1924
rect 9824 1912 9830 1964
rect 9858 1912 9864 1964
rect 9916 1912 9922 1964
rect 9953 1955 10011 1961
rect 9953 1921 9965 1955
rect 9999 1921 10011 1955
rect 9953 1915 10011 1921
rect 10229 1955 10287 1961
rect 10229 1921 10241 1955
rect 10275 1921 10287 1955
rect 10229 1915 10287 1921
rect 9968 1884 9996 1915
rect 9232 1856 9996 1884
rect 9232 1825 9260 1856
rect 8389 1819 8447 1825
rect 8389 1816 8401 1819
rect 7944 1788 8401 1816
rect 8389 1785 8401 1788
rect 8435 1785 8447 1819
rect 9217 1819 9275 1825
rect 8389 1779 8447 1785
rect 8588 1788 9168 1816
rect 6043 1720 7236 1748
rect 7285 1751 7343 1757
rect 6043 1717 6055 1720
rect 5997 1711 6055 1717
rect 7285 1717 7297 1751
rect 7331 1748 7343 1751
rect 8588 1748 8616 1788
rect 7331 1720 8616 1748
rect 7331 1717 7343 1720
rect 7285 1711 7343 1717
rect 8662 1708 8668 1760
rect 8720 1708 8726 1760
rect 9140 1748 9168 1788
rect 9217 1785 9229 1819
rect 9263 1785 9275 1819
rect 9217 1779 9275 1785
rect 9398 1776 9404 1828
rect 9456 1776 9462 1828
rect 9493 1819 9551 1825
rect 9493 1785 9505 1819
rect 9539 1816 9551 1819
rect 10244 1816 10272 1915
rect 10318 1912 10324 1964
rect 10376 1952 10382 1964
rect 10965 1955 11023 1961
rect 10965 1952 10977 1955
rect 10376 1924 10977 1952
rect 10376 1912 10382 1924
rect 10965 1921 10977 1924
rect 11011 1921 11023 1955
rect 11072 1952 11100 2060
rect 11514 2048 11520 2100
rect 11572 2048 11578 2100
rect 12250 2048 12256 2100
rect 12308 2088 12314 2100
rect 13170 2088 13176 2100
rect 12308 2060 13176 2088
rect 12308 2048 12314 2060
rect 13170 2048 13176 2060
rect 13228 2048 13234 2100
rect 13262 2048 13268 2100
rect 13320 2048 13326 2100
rect 13722 2048 13728 2100
rect 13780 2088 13786 2100
rect 13780 2060 14504 2088
rect 13780 2048 13786 2060
rect 11532 2020 11560 2048
rect 11977 2023 12035 2029
rect 11977 2020 11989 2023
rect 11532 1992 11989 2020
rect 11977 1989 11989 1992
rect 12023 1989 12035 2023
rect 13280 2020 13308 2048
rect 13280 1992 14044 2020
rect 11977 1983 12035 1989
rect 11517 1955 11575 1961
rect 11517 1952 11529 1955
rect 11072 1924 11529 1952
rect 10965 1915 11023 1921
rect 11517 1921 11529 1924
rect 11563 1921 11575 1955
rect 11517 1915 11575 1921
rect 12618 1912 12624 1964
rect 12676 1912 12682 1964
rect 12802 1912 12808 1964
rect 12860 1912 12866 1964
rect 13630 1912 13636 1964
rect 13688 1912 13694 1964
rect 14016 1961 14044 1992
rect 14108 1992 14412 2020
rect 14108 1964 14136 1992
rect 14001 1955 14059 1961
rect 14001 1921 14013 1955
rect 14047 1921 14059 1955
rect 14001 1915 14059 1921
rect 14090 1912 14096 1964
rect 14148 1912 14154 1964
rect 14277 1955 14335 1961
rect 14277 1921 14289 1955
rect 14323 1921 14335 1955
rect 14277 1915 14335 1921
rect 13354 1884 13360 1896
rect 9539 1788 10272 1816
rect 10428 1856 13360 1884
rect 9539 1785 9551 1788
rect 9493 1779 9551 1785
rect 9416 1748 9444 1776
rect 9140 1720 9444 1748
rect 9769 1751 9827 1757
rect 9769 1717 9781 1751
rect 9815 1748 9827 1751
rect 9858 1748 9864 1760
rect 9815 1720 9864 1748
rect 9815 1717 9827 1720
rect 9769 1711 9827 1717
rect 9858 1708 9864 1720
rect 9916 1708 9922 1760
rect 10045 1751 10103 1757
rect 10045 1717 10057 1751
rect 10091 1748 10103 1751
rect 10428 1748 10456 1856
rect 13354 1844 13360 1856
rect 13412 1844 13418 1896
rect 14292 1884 14320 1915
rect 13464 1856 14320 1884
rect 14384 1884 14412 1992
rect 14476 1961 14504 2060
rect 15194 2048 15200 2100
rect 15252 2088 15258 2100
rect 15252 2060 15884 2088
rect 15252 2048 15258 2060
rect 15856 2029 15884 2060
rect 16574 2048 16580 2100
rect 16632 2048 16638 2100
rect 16666 2048 16672 2100
rect 16724 2088 16730 2100
rect 17405 2091 17463 2097
rect 17405 2088 17417 2091
rect 16724 2060 17417 2088
rect 16724 2048 16730 2060
rect 17405 2057 17417 2060
rect 17451 2057 17463 2091
rect 17405 2051 17463 2057
rect 17681 2091 17739 2097
rect 17681 2057 17693 2091
rect 17727 2088 17739 2091
rect 17727 2060 18092 2088
rect 17727 2057 17739 2060
rect 17681 2051 17739 2057
rect 15841 2023 15899 2029
rect 14752 1992 15424 2020
rect 14461 1955 14519 1961
rect 14461 1921 14473 1955
rect 14507 1921 14519 1955
rect 14461 1915 14519 1921
rect 14752 1884 14780 1992
rect 14829 1955 14887 1961
rect 14829 1921 14841 1955
rect 14875 1921 14887 1955
rect 14829 1915 14887 1921
rect 14384 1856 14780 1884
rect 11882 1816 11888 1828
rect 11716 1788 11888 1816
rect 10091 1720 10456 1748
rect 10091 1717 10103 1720
rect 10045 1711 10103 1717
rect 10502 1708 10508 1760
rect 10560 1708 10566 1760
rect 11054 1708 11060 1760
rect 11112 1708 11118 1760
rect 11716 1757 11744 1788
rect 11882 1776 11888 1788
rect 11940 1776 11946 1828
rect 13464 1825 13492 1856
rect 12437 1819 12495 1825
rect 12437 1785 12449 1819
rect 12483 1816 12495 1819
rect 13449 1819 13507 1825
rect 12483 1788 13400 1816
rect 12483 1785 12495 1788
rect 12437 1779 12495 1785
rect 11701 1751 11759 1757
rect 11701 1717 11713 1751
rect 11747 1717 11759 1751
rect 11701 1711 11759 1717
rect 11790 1708 11796 1760
rect 11848 1748 11854 1760
rect 12069 1751 12127 1757
rect 12069 1748 12081 1751
rect 11848 1720 12081 1748
rect 11848 1708 11854 1720
rect 12069 1717 12081 1720
rect 12115 1717 12127 1751
rect 12069 1711 12127 1717
rect 12618 1708 12624 1760
rect 12676 1748 12682 1760
rect 12897 1751 12955 1757
rect 12897 1748 12909 1751
rect 12676 1720 12909 1748
rect 12676 1708 12682 1720
rect 12897 1717 12909 1720
rect 12943 1717 12955 1751
rect 13372 1748 13400 1788
rect 13449 1785 13461 1819
rect 13495 1785 13507 1819
rect 13449 1779 13507 1785
rect 13817 1819 13875 1825
rect 13817 1785 13829 1819
rect 13863 1816 13875 1819
rect 14844 1816 14872 1915
rect 15102 1912 15108 1964
rect 15160 1912 15166 1964
rect 15396 1961 15424 1992
rect 15841 1989 15853 2023
rect 15887 1989 15899 2023
rect 16592 2020 16620 2048
rect 18064 2029 18092 2060
rect 18138 2048 18144 2100
rect 18196 2048 18202 2100
rect 18414 2048 18420 2100
rect 18472 2088 18478 2100
rect 18472 2060 19104 2088
rect 18472 2048 18478 2060
rect 16945 2023 17003 2029
rect 16945 2020 16957 2023
rect 16592 1992 16957 2020
rect 15841 1983 15899 1989
rect 16945 1989 16957 1992
rect 16991 1989 17003 2023
rect 16945 1983 17003 1989
rect 18049 2023 18107 2029
rect 18049 1989 18061 2023
rect 18095 1989 18107 2023
rect 18156 2020 18184 2048
rect 18601 2023 18659 2029
rect 18601 2020 18613 2023
rect 18156 1992 18613 2020
rect 18049 1983 18107 1989
rect 18601 1989 18613 1992
rect 18647 1989 18659 2023
rect 19076 2020 19104 2060
rect 19518 2048 19524 2100
rect 19576 2048 19582 2100
rect 19794 2048 19800 2100
rect 19852 2088 19858 2100
rect 21085 2091 21143 2097
rect 21085 2088 21097 2091
rect 19852 2060 21097 2088
rect 19852 2048 19858 2060
rect 21085 2057 21097 2060
rect 21131 2057 21143 2091
rect 21085 2051 21143 2057
rect 21450 2048 21456 2100
rect 21508 2048 21514 2100
rect 21818 2048 21824 2100
rect 21876 2048 21882 2100
rect 22097 2091 22155 2097
rect 22097 2057 22109 2091
rect 22143 2057 22155 2091
rect 22097 2051 22155 2057
rect 19536 2020 19564 2048
rect 20257 2023 20315 2029
rect 20257 2020 20269 2023
rect 19076 1992 19288 2020
rect 19536 1992 20269 2020
rect 18601 1983 18659 1989
rect 15381 1955 15439 1961
rect 15381 1921 15393 1955
rect 15427 1921 15439 1955
rect 15381 1915 15439 1921
rect 15654 1912 15660 1964
rect 15712 1912 15718 1964
rect 16206 1912 16212 1964
rect 16264 1952 16270 1964
rect 16485 1955 16543 1961
rect 16485 1952 16497 1955
rect 16264 1924 16497 1952
rect 16264 1912 16270 1924
rect 16485 1921 16497 1924
rect 16531 1921 16543 1955
rect 17589 1955 17647 1961
rect 17589 1952 17601 1955
rect 16485 1915 16543 1921
rect 16592 1924 17601 1952
rect 13863 1788 14872 1816
rect 15120 1816 15148 1912
rect 15286 1844 15292 1896
rect 15344 1884 15350 1896
rect 16592 1884 16620 1924
rect 17589 1921 17601 1924
rect 17635 1921 17647 1955
rect 17589 1915 17647 1921
rect 17865 1955 17923 1961
rect 17865 1921 17877 1955
rect 17911 1921 17923 1955
rect 17865 1915 17923 1921
rect 19153 1955 19211 1961
rect 19153 1921 19165 1955
rect 19199 1921 19211 1955
rect 19260 1952 19288 1992
rect 20257 1989 20269 1992
rect 20303 1989 20315 2023
rect 20257 1983 20315 1989
rect 20993 2023 21051 2029
rect 20993 1989 21005 2023
rect 21039 2020 21051 2023
rect 21468 2020 21496 2048
rect 21039 1992 21496 2020
rect 21039 1989 21051 1992
rect 20993 1983 21051 1989
rect 21542 1980 21548 2032
rect 21600 2020 21606 2032
rect 22112 2020 22140 2051
rect 22370 2048 22376 2100
rect 22428 2088 22434 2100
rect 22649 2091 22707 2097
rect 22649 2088 22661 2091
rect 22428 2060 22661 2088
rect 22428 2048 22434 2060
rect 22649 2057 22661 2060
rect 22695 2057 22707 2091
rect 22649 2051 22707 2057
rect 22738 2048 22744 2100
rect 22796 2088 22802 2100
rect 22796 2060 23152 2088
rect 22796 2048 22802 2060
rect 22462 2020 22468 2032
rect 21600 1992 22048 2020
rect 22112 1992 22468 2020
rect 21600 1980 21606 1992
rect 19705 1955 19763 1961
rect 19705 1952 19717 1955
rect 19260 1924 19717 1952
rect 19153 1915 19211 1921
rect 19705 1921 19717 1924
rect 19751 1921 19763 1955
rect 19705 1915 19763 1921
rect 15344 1856 16620 1884
rect 15344 1844 15350 1856
rect 16942 1844 16948 1896
rect 17000 1884 17006 1896
rect 17880 1884 17908 1915
rect 18966 1884 18972 1896
rect 17000 1856 17908 1884
rect 18340 1856 18972 1884
rect 17000 1844 17006 1856
rect 15473 1819 15531 1825
rect 15473 1816 15485 1819
rect 15120 1788 15485 1816
rect 13863 1785 13875 1788
rect 13817 1779 13875 1785
rect 15473 1785 15485 1788
rect 15519 1785 15531 1819
rect 15473 1779 15531 1785
rect 16482 1776 16488 1828
rect 16540 1816 16546 1828
rect 18340 1816 18368 1856
rect 18966 1844 18972 1856
rect 19024 1844 19030 1896
rect 19168 1884 19196 1915
rect 20070 1912 20076 1964
rect 20128 1912 20134 1964
rect 21637 1955 21695 1961
rect 21637 1921 21649 1955
rect 21683 1952 21695 1955
rect 21726 1952 21732 1964
rect 21683 1924 21732 1952
rect 21683 1921 21695 1924
rect 21637 1915 21695 1921
rect 21726 1912 21732 1924
rect 21784 1912 21790 1964
rect 22020 1961 22048 1992
rect 22462 1980 22468 1992
rect 22520 1980 22526 2032
rect 23124 2020 23152 2060
rect 23198 2048 23204 2100
rect 23256 2088 23262 2100
rect 23477 2091 23535 2097
rect 23477 2088 23489 2091
rect 23256 2060 23489 2088
rect 23256 2048 23262 2060
rect 23477 2057 23489 2060
rect 23523 2057 23535 2091
rect 23477 2051 23535 2057
rect 24026 2048 24032 2100
rect 24084 2048 24090 2100
rect 24302 2048 24308 2100
rect 24360 2048 24366 2100
rect 22664 1992 22968 2020
rect 23124 1992 23980 2020
rect 22005 1955 22063 1961
rect 22005 1921 22017 1955
rect 22051 1921 22063 1955
rect 22005 1915 22063 1921
rect 22278 1912 22284 1964
rect 22336 1912 22342 1964
rect 22557 1955 22615 1961
rect 22557 1921 22569 1955
rect 22603 1921 22615 1955
rect 22557 1915 22615 1921
rect 20088 1884 20116 1912
rect 19168 1856 20116 1884
rect 20622 1844 20628 1896
rect 20680 1884 20686 1896
rect 22572 1884 22600 1915
rect 20680 1856 22600 1884
rect 20680 1844 20686 1856
rect 16540 1788 18368 1816
rect 16540 1776 16546 1788
rect 19334 1776 19340 1828
rect 19392 1776 19398 1828
rect 20438 1776 20444 1828
rect 20496 1776 20502 1828
rect 21174 1776 21180 1828
rect 21232 1816 21238 1828
rect 22373 1819 22431 1825
rect 22373 1816 22385 1819
rect 21232 1788 22385 1816
rect 21232 1776 21238 1788
rect 22373 1785 22385 1788
rect 22419 1785 22431 1819
rect 22373 1779 22431 1785
rect 13998 1748 14004 1760
rect 13372 1720 14004 1748
rect 12897 1711 12955 1717
rect 13998 1708 14004 1720
rect 14056 1708 14062 1760
rect 14090 1708 14096 1760
rect 14148 1708 14154 1760
rect 14274 1708 14280 1760
rect 14332 1748 14338 1760
rect 14645 1751 14703 1757
rect 14645 1748 14657 1751
rect 14332 1720 14657 1748
rect 14332 1708 14338 1720
rect 14645 1717 14657 1720
rect 14691 1717 14703 1751
rect 14645 1711 14703 1717
rect 14734 1708 14740 1760
rect 14792 1748 14798 1760
rect 15013 1751 15071 1757
rect 15013 1748 15025 1751
rect 14792 1720 15025 1748
rect 14792 1708 14798 1720
rect 15013 1717 15025 1720
rect 15059 1717 15071 1751
rect 15013 1711 15071 1717
rect 15194 1708 15200 1760
rect 15252 1708 15258 1760
rect 15654 1708 15660 1760
rect 15712 1748 15718 1760
rect 15933 1751 15991 1757
rect 15933 1748 15945 1751
rect 15712 1720 15945 1748
rect 15712 1708 15718 1720
rect 15933 1717 15945 1720
rect 15979 1717 15991 1751
rect 15933 1711 15991 1717
rect 16301 1751 16359 1757
rect 16301 1717 16313 1751
rect 16347 1748 16359 1751
rect 16574 1748 16580 1760
rect 16347 1720 16580 1748
rect 16347 1717 16359 1720
rect 16301 1711 16359 1717
rect 16574 1708 16580 1720
rect 16632 1708 16638 1760
rect 16758 1708 16764 1760
rect 16816 1748 16822 1760
rect 17037 1751 17095 1757
rect 17037 1748 17049 1751
rect 16816 1720 17049 1748
rect 16816 1708 16822 1720
rect 17037 1717 17049 1720
rect 17083 1717 17095 1751
rect 17037 1711 17095 1717
rect 17954 1708 17960 1760
rect 18012 1748 18018 1760
rect 18141 1751 18199 1757
rect 18141 1748 18153 1751
rect 18012 1720 18153 1748
rect 18012 1708 18018 1720
rect 18141 1717 18153 1720
rect 18187 1717 18199 1751
rect 18141 1711 18199 1717
rect 18230 1708 18236 1760
rect 18288 1748 18294 1760
rect 18693 1751 18751 1757
rect 18693 1748 18705 1751
rect 18288 1720 18705 1748
rect 18288 1708 18294 1720
rect 18693 1717 18705 1720
rect 18739 1717 18751 1751
rect 18693 1711 18751 1717
rect 19702 1708 19708 1760
rect 19760 1748 19766 1760
rect 19797 1751 19855 1757
rect 19797 1748 19809 1751
rect 19760 1720 19809 1748
rect 19760 1708 19766 1720
rect 19797 1717 19809 1720
rect 19843 1717 19855 1751
rect 19797 1711 19855 1717
rect 19886 1708 19892 1760
rect 19944 1748 19950 1760
rect 21453 1751 21511 1757
rect 21453 1748 21465 1751
rect 19944 1720 21465 1748
rect 19944 1708 19950 1720
rect 21453 1717 21465 1720
rect 21499 1717 21511 1751
rect 21453 1711 21511 1717
rect 21542 1708 21548 1760
rect 21600 1748 21606 1760
rect 22664 1748 22692 1992
rect 22940 1961 22968 1992
rect 22833 1955 22891 1961
rect 22833 1921 22845 1955
rect 22879 1921 22891 1955
rect 22833 1915 22891 1921
rect 22925 1955 22983 1961
rect 22925 1921 22937 1955
rect 22971 1921 22983 1955
rect 22925 1915 22983 1921
rect 22848 1884 22876 1915
rect 23014 1912 23020 1964
rect 23072 1952 23078 1964
rect 23952 1961 23980 1992
rect 23385 1955 23443 1961
rect 23385 1952 23397 1955
rect 23072 1924 23397 1952
rect 23072 1912 23078 1924
rect 23385 1921 23397 1924
rect 23431 1921 23443 1955
rect 23385 1915 23443 1921
rect 23661 1955 23719 1961
rect 23661 1921 23673 1955
rect 23707 1952 23719 1955
rect 23937 1955 23995 1961
rect 23707 1924 23796 1952
rect 23707 1921 23719 1924
rect 23661 1915 23719 1921
rect 22848 1856 23244 1884
rect 23106 1776 23112 1828
rect 23164 1776 23170 1828
rect 23216 1825 23244 1856
rect 23768 1825 23796 1924
rect 23937 1921 23949 1955
rect 23983 1921 23995 1955
rect 23937 1915 23995 1921
rect 24210 1912 24216 1964
rect 24268 1912 24274 1964
rect 24394 1912 24400 1964
rect 24452 1952 24458 1964
rect 24489 1955 24547 1961
rect 24489 1952 24501 1955
rect 24452 1924 24501 1952
rect 24452 1912 24458 1924
rect 24489 1921 24501 1924
rect 24535 1921 24547 1955
rect 24489 1915 24547 1921
rect 23201 1819 23259 1825
rect 23201 1785 23213 1819
rect 23247 1785 23259 1819
rect 23201 1779 23259 1785
rect 23753 1819 23811 1825
rect 23753 1785 23765 1819
rect 23799 1785 23811 1819
rect 23753 1779 23811 1785
rect 21600 1720 22692 1748
rect 21600 1708 21606 1720
rect 1104 1658 24840 1680
rect 1104 1606 3917 1658
rect 3969 1606 3981 1658
rect 4033 1606 4045 1658
rect 4097 1606 4109 1658
rect 4161 1606 4173 1658
rect 4225 1606 9851 1658
rect 9903 1606 9915 1658
rect 9967 1606 9979 1658
rect 10031 1606 10043 1658
rect 10095 1606 10107 1658
rect 10159 1606 15785 1658
rect 15837 1606 15849 1658
rect 15901 1606 15913 1658
rect 15965 1606 15977 1658
rect 16029 1606 16041 1658
rect 16093 1606 21719 1658
rect 21771 1606 21783 1658
rect 21835 1606 21847 1658
rect 21899 1606 21911 1658
rect 21963 1606 21975 1658
rect 22027 1606 24840 1658
rect 1104 1584 24840 1606
rect 2682 1504 2688 1556
rect 2740 1504 2746 1556
rect 2869 1547 2927 1553
rect 2869 1513 2881 1547
rect 2915 1544 2927 1547
rect 4430 1544 4436 1556
rect 2915 1516 4436 1544
rect 2915 1513 2927 1516
rect 2869 1507 2927 1513
rect 4430 1504 4436 1516
rect 4488 1504 4494 1556
rect 4522 1504 4528 1556
rect 4580 1544 4586 1556
rect 6730 1544 6736 1556
rect 4580 1516 6736 1544
rect 4580 1504 4586 1516
rect 6730 1504 6736 1516
rect 6788 1504 6794 1556
rect 7006 1504 7012 1556
rect 7064 1544 7070 1556
rect 7558 1544 7564 1556
rect 7064 1516 7564 1544
rect 7064 1504 7070 1516
rect 7558 1504 7564 1516
rect 7616 1504 7622 1556
rect 7926 1504 7932 1556
rect 7984 1544 7990 1556
rect 7984 1516 12434 1544
rect 7984 1504 7990 1516
rect 2700 1408 2728 1504
rect 3145 1479 3203 1485
rect 3145 1445 3157 1479
rect 3191 1445 3203 1479
rect 3145 1439 3203 1445
rect 4341 1479 4399 1485
rect 4341 1445 4353 1479
rect 4387 1476 4399 1479
rect 7101 1479 7159 1485
rect 4387 1448 5580 1476
rect 4387 1445 4399 1448
rect 4341 1439 4399 1445
rect 2240 1380 2728 1408
rect 3160 1408 3188 1439
rect 4798 1408 4804 1420
rect 3160 1380 3464 1408
rect 1486 1300 1492 1352
rect 1544 1300 1550 1352
rect 1946 1300 1952 1352
rect 2004 1300 2010 1352
rect 2240 1349 2268 1380
rect 2225 1343 2283 1349
rect 2225 1309 2237 1343
rect 2271 1309 2283 1343
rect 2225 1303 2283 1309
rect 2501 1343 2559 1349
rect 2501 1309 2513 1343
rect 2547 1309 2559 1343
rect 2501 1303 2559 1309
rect 2777 1343 2835 1349
rect 2777 1309 2789 1343
rect 2823 1340 2835 1343
rect 2958 1340 2964 1352
rect 2823 1312 2964 1340
rect 2823 1309 2835 1312
rect 2777 1303 2835 1309
rect 2516 1272 2544 1303
rect 2958 1300 2964 1312
rect 3016 1300 3022 1352
rect 3053 1343 3111 1349
rect 3053 1309 3065 1343
rect 3099 1340 3111 1343
rect 3234 1340 3240 1352
rect 3099 1312 3240 1340
rect 3099 1309 3111 1312
rect 3053 1303 3111 1309
rect 3234 1300 3240 1312
rect 3292 1300 3298 1352
rect 3326 1300 3332 1352
rect 3384 1300 3390 1352
rect 3436 1340 3464 1380
rect 4448 1380 4804 1408
rect 3605 1343 3663 1349
rect 3605 1340 3617 1343
rect 3436 1312 3617 1340
rect 3605 1309 3617 1312
rect 3651 1309 3663 1343
rect 3605 1303 3663 1309
rect 3789 1343 3847 1349
rect 3789 1309 3801 1343
rect 3835 1309 3847 1343
rect 3789 1303 3847 1309
rect 4065 1343 4123 1349
rect 4065 1309 4077 1343
rect 4111 1340 4123 1343
rect 4448 1340 4476 1380
rect 4798 1368 4804 1380
rect 4856 1368 4862 1420
rect 5552 1408 5580 1448
rect 7101 1445 7113 1479
rect 7147 1476 7159 1479
rect 7466 1476 7472 1488
rect 7147 1448 7472 1476
rect 7147 1445 7159 1448
rect 7101 1439 7159 1445
rect 7466 1436 7472 1448
rect 7524 1436 7530 1488
rect 8018 1476 8024 1488
rect 7576 1448 8024 1476
rect 7576 1408 7604 1448
rect 8018 1436 8024 1448
rect 8076 1436 8082 1488
rect 8297 1479 8355 1485
rect 8297 1445 8309 1479
rect 8343 1476 8355 1479
rect 8343 1448 9628 1476
rect 8343 1445 8355 1448
rect 8297 1439 8355 1445
rect 8846 1408 8852 1420
rect 5552 1380 7604 1408
rect 7668 1380 7972 1408
rect 4111 1312 4476 1340
rect 4111 1309 4123 1312
rect 4065 1303 4123 1309
rect 3804 1272 3832 1303
rect 4522 1300 4528 1352
rect 4580 1300 4586 1352
rect 4617 1343 4675 1349
rect 4617 1309 4629 1343
rect 4663 1340 4675 1343
rect 4982 1340 4988 1352
rect 4663 1312 4988 1340
rect 4663 1309 4675 1312
rect 4617 1303 4675 1309
rect 4982 1300 4988 1312
rect 5040 1300 5046 1352
rect 5074 1300 5080 1352
rect 5132 1300 5138 1352
rect 5169 1343 5227 1349
rect 5169 1309 5181 1343
rect 5215 1340 5227 1343
rect 5534 1340 5540 1352
rect 5215 1312 5540 1340
rect 5215 1309 5227 1312
rect 5169 1303 5227 1309
rect 5534 1300 5540 1312
rect 5592 1300 5598 1352
rect 5629 1343 5687 1349
rect 5629 1309 5641 1343
rect 5675 1309 5687 1343
rect 5629 1303 5687 1309
rect 4430 1272 4436 1284
rect 2056 1244 2544 1272
rect 3436 1244 3832 1272
rect 4264 1244 4436 1272
rect 1670 1164 1676 1216
rect 1728 1164 1734 1216
rect 1762 1164 1768 1216
rect 1820 1164 1826 1216
rect 2056 1213 2084 1244
rect 2041 1207 2099 1213
rect 2041 1173 2053 1207
rect 2087 1173 2099 1207
rect 2041 1167 2099 1173
rect 2314 1164 2320 1216
rect 2372 1164 2378 1216
rect 2590 1164 2596 1216
rect 2648 1164 2654 1216
rect 3436 1213 3464 1244
rect 3421 1207 3479 1213
rect 3421 1173 3433 1207
rect 3467 1173 3479 1207
rect 3421 1167 3479 1173
rect 3973 1207 4031 1213
rect 3973 1173 3985 1207
rect 4019 1204 4031 1207
rect 4154 1204 4160 1216
rect 4019 1176 4160 1204
rect 4019 1173 4031 1176
rect 3973 1167 4031 1173
rect 4154 1164 4160 1176
rect 4212 1164 4218 1216
rect 4264 1213 4292 1244
rect 4430 1232 4436 1244
rect 4488 1232 4494 1284
rect 5644 1272 5672 1303
rect 5718 1300 5724 1352
rect 5776 1300 5782 1352
rect 6178 1300 6184 1352
rect 6236 1300 6242 1352
rect 6365 1343 6423 1349
rect 6365 1309 6377 1343
rect 6411 1340 6423 1343
rect 6730 1340 6736 1352
rect 6411 1312 6736 1340
rect 6411 1309 6423 1312
rect 6365 1303 6423 1309
rect 6730 1300 6736 1312
rect 6788 1300 6794 1352
rect 6825 1343 6883 1349
rect 6825 1309 6837 1343
rect 6871 1309 6883 1343
rect 6825 1303 6883 1309
rect 6840 1272 6868 1303
rect 6914 1300 6920 1352
rect 6972 1300 6978 1352
rect 7668 1349 7696 1380
rect 7377 1343 7435 1349
rect 7377 1309 7389 1343
rect 7423 1309 7435 1343
rect 7377 1303 7435 1309
rect 7653 1343 7711 1349
rect 7653 1309 7665 1343
rect 7699 1309 7711 1343
rect 7653 1303 7711 1309
rect 4908 1244 5672 1272
rect 6012 1244 6868 1272
rect 7392 1272 7420 1303
rect 7742 1300 7748 1352
rect 7800 1300 7806 1352
rect 7834 1300 7840 1352
rect 7892 1300 7898 1352
rect 7852 1272 7880 1300
rect 7392 1244 7880 1272
rect 7944 1272 7972 1380
rect 8220 1380 8852 1408
rect 8220 1349 8248 1380
rect 8846 1368 8852 1380
rect 8904 1368 8910 1420
rect 9306 1408 9312 1420
rect 9232 1380 9312 1408
rect 8205 1343 8263 1349
rect 8205 1309 8217 1343
rect 8251 1309 8263 1343
rect 8205 1303 8263 1309
rect 8481 1343 8539 1349
rect 8481 1309 8493 1343
rect 8527 1340 8539 1343
rect 8662 1340 8668 1352
rect 8527 1312 8668 1340
rect 8527 1309 8539 1312
rect 8481 1303 8539 1309
rect 8662 1300 8668 1312
rect 8720 1300 8726 1352
rect 8757 1343 8815 1349
rect 8757 1309 8769 1343
rect 8803 1340 8815 1343
rect 9030 1340 9036 1352
rect 8803 1312 9036 1340
rect 8803 1309 8815 1312
rect 8757 1303 8815 1309
rect 9030 1300 9036 1312
rect 9088 1300 9094 1352
rect 9232 1349 9260 1380
rect 9306 1368 9312 1380
rect 9364 1368 9370 1420
rect 9600 1349 9628 1448
rect 11054 1368 11060 1420
rect 11112 1368 11118 1420
rect 12406 1408 12434 1516
rect 13354 1504 13360 1556
rect 13412 1504 13418 1556
rect 13814 1504 13820 1556
rect 13872 1544 13878 1556
rect 14277 1547 14335 1553
rect 14277 1544 14289 1547
rect 13872 1516 14289 1544
rect 13872 1504 13878 1516
rect 14277 1513 14289 1516
rect 14323 1513 14335 1547
rect 14277 1507 14335 1513
rect 15102 1504 15108 1556
rect 15160 1544 15166 1556
rect 15381 1547 15439 1553
rect 15381 1544 15393 1547
rect 15160 1516 15393 1544
rect 15160 1504 15166 1516
rect 15381 1513 15393 1516
rect 15427 1513 15439 1547
rect 15381 1507 15439 1513
rect 15933 1547 15991 1553
rect 15933 1513 15945 1547
rect 15979 1513 15991 1547
rect 15933 1507 15991 1513
rect 13372 1408 13400 1504
rect 14090 1436 14096 1488
rect 14148 1476 14154 1488
rect 14148 1448 15056 1476
rect 14148 1436 14154 1448
rect 12406 1380 12572 1408
rect 13372 1380 14964 1408
rect 9217 1343 9275 1349
rect 9217 1309 9229 1343
rect 9263 1309 9275 1343
rect 9493 1343 9551 1349
rect 9493 1336 9505 1343
rect 9217 1303 9275 1309
rect 9416 1309 9505 1336
rect 9539 1309 9551 1343
rect 9416 1308 9551 1309
rect 8294 1272 8300 1284
rect 7944 1244 8300 1272
rect 4249 1207 4307 1213
rect 4249 1173 4261 1207
rect 4295 1173 4307 1207
rect 4249 1167 4307 1173
rect 4798 1164 4804 1216
rect 4856 1164 4862 1216
rect 4908 1213 4936 1244
rect 4893 1207 4951 1213
rect 4893 1173 4905 1207
rect 4939 1173 4951 1207
rect 4893 1167 4951 1173
rect 5350 1164 5356 1216
rect 5408 1164 5414 1216
rect 5442 1164 5448 1216
rect 5500 1164 5506 1216
rect 5810 1164 5816 1216
rect 5868 1204 5874 1216
rect 6012 1213 6040 1244
rect 8294 1232 8300 1244
rect 8352 1232 8358 1284
rect 9416 1272 9444 1308
rect 9493 1303 9551 1308
rect 9585 1343 9643 1349
rect 9585 1309 9597 1343
rect 9631 1309 9643 1343
rect 9585 1303 9643 1309
rect 9674 1300 9680 1352
rect 9732 1340 9738 1352
rect 9953 1343 10011 1349
rect 9953 1340 9965 1343
rect 9732 1312 9965 1340
rect 9732 1300 9738 1312
rect 9953 1309 9965 1312
rect 9999 1309 10011 1343
rect 10321 1343 10379 1349
rect 10321 1340 10333 1343
rect 9953 1303 10011 1309
rect 10060 1312 10333 1340
rect 10060 1272 10088 1312
rect 10321 1309 10333 1312
rect 10367 1309 10379 1343
rect 10321 1303 10379 1309
rect 11698 1300 11704 1352
rect 11756 1300 11762 1352
rect 11793 1343 11851 1349
rect 11793 1309 11805 1343
rect 11839 1309 11851 1343
rect 12434 1340 12440 1352
rect 11793 1303 11851 1309
rect 11992 1312 12440 1340
rect 10686 1272 10692 1284
rect 8588 1244 9444 1272
rect 9692 1244 10088 1272
rect 10152 1244 10692 1272
rect 5905 1207 5963 1213
rect 5905 1204 5917 1207
rect 5868 1176 5917 1204
rect 5868 1164 5874 1176
rect 5905 1173 5917 1176
rect 5951 1173 5963 1207
rect 5905 1167 5963 1173
rect 5997 1207 6055 1213
rect 5997 1173 6009 1207
rect 6043 1173 6055 1207
rect 5997 1167 6055 1173
rect 6546 1164 6552 1216
rect 6604 1164 6610 1216
rect 6638 1164 6644 1216
rect 6696 1164 6702 1216
rect 7193 1207 7251 1213
rect 7193 1173 7205 1207
rect 7239 1204 7251 1207
rect 7374 1204 7380 1216
rect 7239 1176 7380 1204
rect 7239 1173 7251 1176
rect 7193 1167 7251 1173
rect 7374 1164 7380 1176
rect 7432 1164 7438 1216
rect 7469 1207 7527 1213
rect 7469 1173 7481 1207
rect 7515 1204 7527 1207
rect 7742 1204 7748 1216
rect 7515 1176 7748 1204
rect 7515 1173 7527 1176
rect 7469 1167 7527 1173
rect 7742 1164 7748 1176
rect 7800 1164 7806 1216
rect 7834 1164 7840 1216
rect 7892 1204 7898 1216
rect 7929 1207 7987 1213
rect 7929 1204 7941 1207
rect 7892 1176 7941 1204
rect 7892 1164 7898 1176
rect 7929 1173 7941 1176
rect 7975 1173 7987 1207
rect 7929 1167 7987 1173
rect 8018 1164 8024 1216
rect 8076 1164 8082 1216
rect 8588 1213 8616 1244
rect 8573 1207 8631 1213
rect 8573 1173 8585 1207
rect 8619 1173 8631 1207
rect 8573 1167 8631 1173
rect 9033 1207 9091 1213
rect 9033 1173 9045 1207
rect 9079 1204 9091 1207
rect 9214 1204 9220 1216
rect 9079 1176 9220 1204
rect 9079 1173 9091 1176
rect 9033 1167 9091 1173
rect 9214 1164 9220 1176
rect 9272 1164 9278 1216
rect 9306 1164 9312 1216
rect 9364 1164 9370 1216
rect 9398 1164 9404 1216
rect 9456 1204 9462 1216
rect 9692 1204 9720 1244
rect 9456 1176 9720 1204
rect 9769 1207 9827 1213
rect 9456 1164 9462 1176
rect 9769 1173 9781 1207
rect 9815 1204 9827 1207
rect 10042 1204 10048 1216
rect 9815 1176 10048 1204
rect 9815 1173 9827 1176
rect 9769 1167 9827 1173
rect 10042 1164 10048 1176
rect 10100 1164 10106 1216
rect 10152 1213 10180 1244
rect 10686 1232 10692 1244
rect 10744 1232 10750 1284
rect 10778 1232 10784 1284
rect 10836 1232 10842 1284
rect 11808 1272 11836 1303
rect 11624 1244 11836 1272
rect 11624 1216 11652 1244
rect 10137 1207 10195 1213
rect 10137 1173 10149 1207
rect 10183 1173 10195 1207
rect 10137 1167 10195 1173
rect 10505 1207 10563 1213
rect 10505 1173 10517 1207
rect 10551 1204 10563 1207
rect 11146 1204 11152 1216
rect 10551 1176 11152 1204
rect 10551 1173 10563 1176
rect 10505 1167 10563 1173
rect 11146 1164 11152 1176
rect 11204 1164 11210 1216
rect 11514 1164 11520 1216
rect 11572 1164 11578 1216
rect 11606 1164 11612 1216
rect 11664 1164 11670 1216
rect 11992 1213 12020 1312
rect 12434 1300 12440 1312
rect 12492 1300 12498 1352
rect 12253 1275 12311 1281
rect 12253 1272 12265 1275
rect 12084 1244 12265 1272
rect 12084 1216 12112 1244
rect 12253 1241 12265 1244
rect 12299 1241 12311 1275
rect 12544 1272 12572 1380
rect 12894 1300 12900 1352
rect 12952 1300 12958 1352
rect 13262 1300 13268 1352
rect 13320 1300 13326 1352
rect 14645 1343 14703 1349
rect 14645 1340 14657 1343
rect 13372 1312 14657 1340
rect 13372 1272 13400 1312
rect 14645 1309 14657 1312
rect 14691 1309 14703 1343
rect 14645 1303 14703 1309
rect 12544 1244 13400 1272
rect 12253 1235 12311 1241
rect 14182 1232 14188 1284
rect 14240 1232 14246 1284
rect 11977 1207 12035 1213
rect 11977 1173 11989 1207
rect 12023 1173 12035 1207
rect 11977 1167 12035 1173
rect 12066 1164 12072 1216
rect 12124 1164 12130 1216
rect 12342 1164 12348 1216
rect 12400 1164 12406 1216
rect 13078 1164 13084 1216
rect 13136 1164 13142 1216
rect 13446 1164 13452 1216
rect 13504 1164 13510 1216
rect 13998 1164 14004 1216
rect 14056 1204 14062 1216
rect 14829 1207 14887 1213
rect 14829 1204 14841 1207
rect 14056 1176 14841 1204
rect 14056 1164 14062 1176
rect 14829 1173 14841 1176
rect 14875 1173 14887 1207
rect 14936 1204 14964 1380
rect 15028 1272 15056 1448
rect 15102 1368 15108 1420
rect 15160 1408 15166 1420
rect 15948 1408 15976 1507
rect 16114 1504 16120 1556
rect 16172 1544 16178 1556
rect 16853 1547 16911 1553
rect 16853 1544 16865 1547
rect 16172 1516 16865 1544
rect 16172 1504 16178 1516
rect 16853 1513 16865 1516
rect 16899 1513 16911 1547
rect 16853 1507 16911 1513
rect 17405 1547 17463 1553
rect 17405 1513 17417 1547
rect 17451 1513 17463 1547
rect 18509 1547 18567 1553
rect 18509 1544 18521 1547
rect 17405 1507 17463 1513
rect 17512 1516 18521 1544
rect 17420 1476 17448 1507
rect 16132 1448 17448 1476
rect 16132 1420 16160 1448
rect 15160 1380 15976 1408
rect 15160 1368 15166 1380
rect 16114 1368 16120 1420
rect 16172 1368 16178 1420
rect 16224 1380 16896 1408
rect 15194 1300 15200 1352
rect 15252 1340 15258 1352
rect 15841 1343 15899 1349
rect 15841 1340 15853 1343
rect 15252 1312 15853 1340
rect 15252 1300 15258 1312
rect 15841 1309 15853 1312
rect 15887 1309 15899 1343
rect 15841 1303 15899 1309
rect 15289 1275 15347 1281
rect 15289 1272 15301 1275
rect 15028 1244 15301 1272
rect 15289 1241 15301 1244
rect 15335 1241 15347 1275
rect 15289 1235 15347 1241
rect 16224 1204 16252 1380
rect 16298 1300 16304 1352
rect 16356 1340 16362 1352
rect 16485 1343 16543 1349
rect 16485 1340 16497 1343
rect 16356 1312 16497 1340
rect 16356 1300 16362 1312
rect 16485 1309 16497 1312
rect 16531 1309 16543 1343
rect 16485 1303 16543 1309
rect 16574 1300 16580 1352
rect 16632 1340 16638 1352
rect 16761 1343 16819 1349
rect 16761 1340 16773 1343
rect 16632 1312 16773 1340
rect 16632 1300 16638 1312
rect 16761 1309 16773 1312
rect 16807 1309 16819 1343
rect 16868 1340 16896 1380
rect 17034 1368 17040 1420
rect 17092 1408 17098 1420
rect 17512 1408 17540 1516
rect 18509 1513 18521 1516
rect 18555 1513 18567 1547
rect 18509 1507 18567 1513
rect 18877 1547 18935 1553
rect 18877 1513 18889 1547
rect 18923 1544 18935 1547
rect 19150 1544 19156 1556
rect 18923 1516 19156 1544
rect 18923 1513 18935 1516
rect 18877 1507 18935 1513
rect 19150 1504 19156 1516
rect 19208 1504 19214 1556
rect 20533 1547 20591 1553
rect 20533 1513 20545 1547
rect 20579 1513 20591 1547
rect 20533 1507 20591 1513
rect 17586 1436 17592 1488
rect 17644 1476 17650 1488
rect 17644 1448 18644 1476
rect 17644 1436 17650 1448
rect 17092 1380 17540 1408
rect 18616 1408 18644 1448
rect 18690 1436 18696 1488
rect 18748 1476 18754 1488
rect 20548 1476 20576 1507
rect 20714 1504 20720 1556
rect 20772 1504 20778 1556
rect 21634 1504 21640 1556
rect 21692 1544 21698 1556
rect 21821 1547 21879 1553
rect 21821 1544 21833 1547
rect 21692 1516 21833 1544
rect 21692 1504 21698 1516
rect 21821 1513 21833 1516
rect 21867 1513 21879 1547
rect 22097 1547 22155 1553
rect 22097 1544 22109 1547
rect 21821 1507 21879 1513
rect 21928 1516 22109 1544
rect 18748 1448 20576 1476
rect 20732 1476 20760 1504
rect 21928 1476 21956 1516
rect 22097 1513 22109 1516
rect 22143 1513 22155 1547
rect 22097 1507 22155 1513
rect 22186 1504 22192 1556
rect 22244 1544 22250 1556
rect 22649 1547 22707 1553
rect 22649 1544 22661 1547
rect 22244 1516 22661 1544
rect 22244 1504 22250 1516
rect 22649 1513 22661 1516
rect 22695 1513 22707 1547
rect 22649 1507 22707 1513
rect 20732 1448 21956 1476
rect 18748 1436 18754 1448
rect 22002 1436 22008 1488
rect 22060 1476 22066 1488
rect 22060 1448 23520 1476
rect 22060 1436 22066 1448
rect 19613 1411 19671 1417
rect 19613 1408 19625 1411
rect 18616 1380 19625 1408
rect 17092 1368 17098 1380
rect 19613 1377 19625 1380
rect 19659 1377 19671 1411
rect 20165 1411 20223 1417
rect 20165 1408 20177 1411
rect 19613 1371 19671 1377
rect 19720 1380 20177 1408
rect 16868 1312 17448 1340
rect 16761 1303 16819 1309
rect 16942 1272 16948 1284
rect 16316 1244 16948 1272
rect 16316 1213 16344 1244
rect 16942 1232 16948 1244
rect 17000 1232 17006 1284
rect 17218 1232 17224 1284
rect 17276 1272 17282 1284
rect 17313 1275 17371 1281
rect 17313 1272 17325 1275
rect 17276 1244 17325 1272
rect 17276 1232 17282 1244
rect 17313 1241 17325 1244
rect 17359 1241 17371 1275
rect 17420 1272 17448 1312
rect 17770 1300 17776 1352
rect 17828 1340 17834 1352
rect 17828 1312 18552 1340
rect 17828 1300 17834 1312
rect 17865 1275 17923 1281
rect 17865 1272 17877 1275
rect 17420 1244 17877 1272
rect 17313 1235 17371 1241
rect 17865 1241 17877 1244
rect 17911 1241 17923 1275
rect 17865 1235 17923 1241
rect 18046 1232 18052 1284
rect 18104 1272 18110 1284
rect 18417 1275 18475 1281
rect 18417 1272 18429 1275
rect 18104 1244 18429 1272
rect 18104 1232 18110 1244
rect 18417 1241 18429 1244
rect 18463 1241 18475 1275
rect 18524 1272 18552 1312
rect 18598 1300 18604 1352
rect 18656 1340 18662 1352
rect 19061 1343 19119 1349
rect 19061 1340 19073 1343
rect 18656 1312 19073 1340
rect 18656 1300 18662 1312
rect 19061 1309 19073 1312
rect 19107 1309 19119 1343
rect 19720 1340 19748 1380
rect 20165 1377 20177 1380
rect 20211 1377 20223 1411
rect 20165 1371 20223 1377
rect 21637 1343 21695 1349
rect 21637 1340 21649 1343
rect 19061 1303 19119 1309
rect 19168 1312 19748 1340
rect 20916 1312 21649 1340
rect 19168 1272 19196 1312
rect 18524 1244 19196 1272
rect 18417 1235 18475 1241
rect 19334 1232 19340 1284
rect 19392 1232 19398 1284
rect 19426 1232 19432 1284
rect 19484 1272 19490 1284
rect 19889 1275 19947 1281
rect 19889 1272 19901 1275
rect 19484 1244 19901 1272
rect 19484 1232 19490 1244
rect 19889 1241 19901 1244
rect 19935 1241 19947 1275
rect 19889 1235 19947 1241
rect 20441 1275 20499 1281
rect 20441 1241 20453 1275
rect 20487 1241 20499 1275
rect 20441 1235 20499 1241
rect 14936 1176 16252 1204
rect 16301 1207 16359 1213
rect 14829 1167 14887 1173
rect 16301 1173 16313 1207
rect 16347 1173 16359 1207
rect 16301 1167 16359 1173
rect 16390 1164 16396 1216
rect 16448 1204 16454 1216
rect 17957 1207 18015 1213
rect 17957 1204 17969 1207
rect 16448 1176 17969 1204
rect 16448 1164 16454 1176
rect 17957 1173 17969 1176
rect 18003 1173 18015 1207
rect 17957 1167 18015 1173
rect 18506 1164 18512 1216
rect 18564 1204 18570 1216
rect 20456 1204 20484 1235
rect 18564 1176 20484 1204
rect 18564 1164 18570 1176
rect 20806 1164 20812 1216
rect 20864 1204 20870 1216
rect 20916 1204 20944 1312
rect 21637 1309 21649 1312
rect 21683 1309 21695 1343
rect 21637 1303 21695 1309
rect 22005 1343 22063 1349
rect 22005 1309 22017 1343
rect 22051 1309 22063 1343
rect 22005 1303 22063 1309
rect 20990 1232 20996 1284
rect 21048 1272 21054 1284
rect 22020 1272 22048 1303
rect 22278 1300 22284 1352
rect 22336 1300 22342 1352
rect 22554 1300 22560 1352
rect 22612 1300 22618 1352
rect 22738 1300 22744 1352
rect 22796 1340 22802 1352
rect 22833 1343 22891 1349
rect 22833 1340 22845 1343
rect 22796 1312 22845 1340
rect 22796 1300 22802 1312
rect 22833 1309 22845 1312
rect 22879 1309 22891 1343
rect 22833 1303 22891 1309
rect 22925 1343 22983 1349
rect 22925 1309 22937 1343
rect 22971 1340 22983 1343
rect 23014 1340 23020 1352
rect 22971 1312 23020 1340
rect 22971 1309 22983 1312
rect 22925 1303 22983 1309
rect 23014 1300 23020 1312
rect 23072 1300 23078 1352
rect 23382 1300 23388 1352
rect 23440 1300 23446 1352
rect 23492 1349 23520 1448
rect 23750 1436 23756 1488
rect 23808 1476 23814 1488
rect 24026 1476 24032 1488
rect 23808 1448 24032 1476
rect 23808 1436 23814 1448
rect 24026 1436 24032 1448
rect 24084 1436 24090 1488
rect 23477 1343 23535 1349
rect 23477 1309 23489 1343
rect 23523 1309 23535 1343
rect 23477 1303 23535 1309
rect 23750 1300 23756 1352
rect 23808 1300 23814 1352
rect 23934 1300 23940 1352
rect 23992 1300 23998 1352
rect 24210 1300 24216 1352
rect 24268 1300 24274 1352
rect 23952 1272 23980 1300
rect 21048 1244 21588 1272
rect 22020 1244 23244 1272
rect 23952 1244 24072 1272
rect 21048 1232 21054 1244
rect 21085 1207 21143 1213
rect 21085 1204 21097 1207
rect 20864 1176 21097 1204
rect 20864 1164 20870 1176
rect 21085 1173 21097 1176
rect 21131 1173 21143 1207
rect 21085 1167 21143 1173
rect 21450 1164 21456 1216
rect 21508 1164 21514 1216
rect 21560 1204 21588 1244
rect 22373 1207 22431 1213
rect 22373 1204 22385 1207
rect 21560 1176 22385 1204
rect 22373 1173 22385 1176
rect 22419 1173 22431 1207
rect 22373 1167 22431 1173
rect 23106 1164 23112 1216
rect 23164 1164 23170 1216
rect 23216 1213 23244 1244
rect 23201 1207 23259 1213
rect 23201 1173 23213 1207
rect 23247 1173 23259 1207
rect 23201 1167 23259 1173
rect 23474 1164 23480 1216
rect 23532 1204 23538 1216
rect 23661 1207 23719 1213
rect 23661 1204 23673 1207
rect 23532 1176 23673 1204
rect 23532 1164 23538 1176
rect 23661 1173 23673 1176
rect 23707 1173 23719 1207
rect 23661 1167 23719 1173
rect 23934 1164 23940 1216
rect 23992 1164 23998 1216
rect 24044 1213 24072 1244
rect 24029 1207 24087 1213
rect 24029 1173 24041 1207
rect 24075 1173 24087 1207
rect 24029 1167 24087 1173
rect 1104 1114 25000 1136
rect 1104 1062 6884 1114
rect 6936 1062 6948 1114
rect 7000 1062 7012 1114
rect 7064 1062 7076 1114
rect 7128 1062 7140 1114
rect 7192 1062 12818 1114
rect 12870 1062 12882 1114
rect 12934 1062 12946 1114
rect 12998 1062 13010 1114
rect 13062 1062 13074 1114
rect 13126 1062 18752 1114
rect 18804 1062 18816 1114
rect 18868 1062 18880 1114
rect 18932 1062 18944 1114
rect 18996 1062 19008 1114
rect 19060 1062 24686 1114
rect 24738 1062 24750 1114
rect 24802 1062 24814 1114
rect 24866 1062 24878 1114
rect 24930 1062 24942 1114
rect 24994 1062 25000 1114
rect 1104 1040 25000 1062
rect 4982 960 4988 1012
rect 5040 1000 5046 1012
rect 5534 1000 5540 1012
rect 5040 972 5540 1000
rect 5040 960 5046 972
rect 5534 960 5540 972
rect 5592 960 5598 1012
rect 6178 960 6184 1012
rect 6236 960 6242 1012
rect 7374 960 7380 1012
rect 7432 1000 7438 1012
rect 10778 1000 10784 1012
rect 7432 972 10784 1000
rect 7432 960 7438 972
rect 10778 960 10784 972
rect 10836 960 10842 1012
rect 11514 960 11520 1012
rect 11572 1000 11578 1012
rect 11572 972 12434 1000
rect 11572 960 11578 972
rect 1762 892 1768 944
rect 1820 932 1826 944
rect 1820 904 2774 932
rect 1820 892 1826 904
rect 2746 796 2774 904
rect 3510 892 3516 944
rect 3568 932 3574 944
rect 6196 932 6224 960
rect 3568 904 6224 932
rect 3568 892 3574 904
rect 8018 892 8024 944
rect 8076 932 8082 944
rect 9766 932 9772 944
rect 8076 904 9772 932
rect 8076 892 8082 904
rect 9766 892 9772 904
rect 9824 892 9830 944
rect 12250 892 12256 944
rect 12308 892 12314 944
rect 5442 824 5448 876
rect 5500 864 5506 876
rect 9398 864 9404 876
rect 5500 836 9404 864
rect 5500 824 5506 836
rect 9398 824 9404 836
rect 9456 824 9462 876
rect 9490 824 9496 876
rect 9548 864 9554 876
rect 12268 864 12296 892
rect 9548 836 12296 864
rect 12406 864 12434 972
rect 18046 960 18052 1012
rect 18104 960 18110 1012
rect 18322 960 18328 1012
rect 18380 960 18386 1012
rect 18506 960 18512 1012
rect 18564 1000 18570 1012
rect 19702 1000 19708 1012
rect 18564 972 19708 1000
rect 18564 960 18570 972
rect 19702 960 19708 972
rect 19760 960 19766 1012
rect 20622 960 20628 1012
rect 20680 1000 20686 1012
rect 22554 1000 22560 1012
rect 20680 972 22560 1000
rect 20680 960 20686 972
rect 22554 960 22560 972
rect 22612 960 22618 1012
rect 23934 960 23940 1012
rect 23992 960 23998 1012
rect 18064 864 18092 960
rect 18340 932 18368 960
rect 21450 932 21456 944
rect 18340 904 21456 932
rect 21450 892 21456 904
rect 21508 892 21514 944
rect 23952 932 23980 960
rect 21652 904 23980 932
rect 21652 864 21680 904
rect 23014 864 23020 876
rect 12406 836 18092 864
rect 21560 836 21680 864
rect 22066 836 23020 864
rect 9548 824 9554 836
rect 5626 796 5632 808
rect 2746 768 5632 796
rect 5626 756 5632 768
rect 5684 756 5690 808
rect 6638 756 6644 808
rect 6696 796 6702 808
rect 14182 796 14188 808
rect 6696 768 14188 796
rect 6696 756 6702 768
rect 14182 756 14188 768
rect 14240 756 14246 808
rect 21560 796 21588 836
rect 16960 768 21588 796
rect 1946 688 1952 740
rect 2004 728 2010 740
rect 2682 728 2688 740
rect 2004 700 2688 728
rect 2004 688 2010 700
rect 2682 688 2688 700
rect 2740 688 2746 740
rect 3326 688 3332 740
rect 3384 728 3390 740
rect 4062 728 4068 740
rect 3384 700 4068 728
rect 3384 688 3390 700
rect 4062 688 4068 700
rect 4120 688 4126 740
rect 4522 688 4528 740
rect 4580 728 4586 740
rect 5442 728 5448 740
rect 4580 700 5448 728
rect 4580 688 4586 700
rect 5442 688 5448 700
rect 5500 688 5506 740
rect 6730 688 6736 740
rect 6788 728 6794 740
rect 7374 728 7380 740
rect 6788 700 7380 728
rect 6788 688 6794 700
rect 7374 688 7380 700
rect 7432 688 7438 740
rect 7466 688 7472 740
rect 7524 688 7530 740
rect 9030 688 9036 740
rect 9088 728 9094 740
rect 9674 728 9680 740
rect 9088 700 9680 728
rect 9088 688 9094 700
rect 9674 688 9680 700
rect 9732 688 9738 740
rect 16850 728 16856 740
rect 9784 700 16856 728
rect 1486 620 1492 672
rect 1544 660 1550 672
rect 2406 660 2412 672
rect 1544 632 2412 660
rect 1544 620 1550 632
rect 2406 620 2412 632
rect 2464 620 2470 672
rect 4706 620 4712 672
rect 4764 620 4770 672
rect 5718 620 5724 672
rect 5776 660 5782 672
rect 6822 660 6828 672
rect 5776 632 6828 660
rect 5776 620 5782 632
rect 6822 620 6828 632
rect 6880 620 6886 672
rect 7484 660 7512 688
rect 9784 660 9812 700
rect 16850 688 16856 700
rect 16908 688 16914 740
rect 7484 632 9812 660
rect 12434 620 12440 672
rect 12492 660 12498 672
rect 12894 660 12900 672
rect 12492 632 12900 660
rect 12492 620 12498 632
rect 12894 620 12900 632
rect 12952 620 12958 672
rect 13262 620 13268 672
rect 13320 620 13326 672
rect 13906 620 13912 672
rect 13964 660 13970 672
rect 16960 660 16988 768
rect 21634 756 21640 808
rect 21692 796 21698 808
rect 22066 796 22094 836
rect 23014 824 23020 836
rect 23072 824 23078 876
rect 21692 768 22094 796
rect 21692 756 21698 768
rect 23474 756 23480 808
rect 23532 796 23538 808
rect 24210 796 24216 808
rect 23532 768 24216 796
rect 23532 756 23538 768
rect 24210 756 24216 768
rect 24268 756 24274 808
rect 21082 688 21088 740
rect 21140 728 21146 740
rect 22738 728 22744 740
rect 21140 700 22744 728
rect 21140 688 21146 700
rect 22738 688 22744 700
rect 22796 688 22802 740
rect 13964 632 16988 660
rect 13964 620 13970 632
rect 22002 620 22008 672
rect 22060 660 22066 672
rect 23750 660 23756 672
rect 22060 632 23756 660
rect 22060 620 22066 632
rect 23750 620 23756 632
rect 23808 620 23814 672
rect 2314 552 2320 604
rect 2372 552 2378 604
rect 4724 592 4752 620
rect 12066 592 12072 604
rect 4724 564 12072 592
rect 12066 552 12072 564
rect 12124 552 12130 604
rect 2332 388 2360 552
rect 4246 484 4252 536
rect 4304 524 4310 536
rect 11606 524 11612 536
rect 4304 496 11612 524
rect 4304 484 4310 496
rect 11606 484 11612 496
rect 11664 484 11670 536
rect 11974 484 11980 536
rect 12032 484 12038 536
rect 2590 416 2596 468
rect 2648 456 2654 468
rect 6730 456 6736 468
rect 2648 428 6736 456
rect 2648 416 2654 428
rect 6730 416 6736 428
rect 6788 416 6794 468
rect 7742 416 7748 468
rect 7800 456 7806 468
rect 11992 456 12020 484
rect 7800 428 12020 456
rect 7800 416 7806 428
rect 13280 388 13308 620
rect 19242 484 19248 536
rect 19300 524 19306 536
rect 20438 524 20444 536
rect 19300 496 20444 524
rect 19300 484 19306 496
rect 20438 484 20444 496
rect 20496 484 20502 536
rect 21174 416 21180 468
rect 21232 456 21238 468
rect 21634 456 21640 468
rect 21232 428 21640 456
rect 21232 416 21238 428
rect 21634 416 21640 428
rect 21692 416 21698 468
rect 2332 360 13308 388
rect 7834 280 7840 332
rect 7892 320 7898 332
rect 7892 292 12434 320
rect 7892 280 7898 292
rect 4798 212 4804 264
rect 4856 252 4862 264
rect 8938 252 8944 264
rect 4856 224 8944 252
rect 4856 212 4862 224
rect 8938 212 8944 224
rect 8996 212 9002 264
rect 12406 252 12434 292
rect 15470 252 15476 264
rect 12406 224 15476 252
rect 15470 212 15476 224
rect 15528 212 15534 264
<< via1 >>
rect 6884 8678 6936 8730
rect 6948 8678 7000 8730
rect 7012 8678 7064 8730
rect 7076 8678 7128 8730
rect 7140 8678 7192 8730
rect 12818 8678 12870 8730
rect 12882 8678 12934 8730
rect 12946 8678 12998 8730
rect 13010 8678 13062 8730
rect 13074 8678 13126 8730
rect 18752 8678 18804 8730
rect 18816 8678 18868 8730
rect 18880 8678 18932 8730
rect 18944 8678 18996 8730
rect 19008 8678 19060 8730
rect 24686 8678 24738 8730
rect 24750 8678 24802 8730
rect 24814 8678 24866 8730
rect 24878 8678 24930 8730
rect 24942 8678 24994 8730
rect 1216 8576 1268 8628
rect 2136 8576 2188 8628
rect 3332 8576 3384 8628
rect 4528 8576 4580 8628
rect 5724 8576 5776 8628
rect 1492 8483 1544 8492
rect 1492 8449 1501 8483
rect 1501 8449 1535 8483
rect 1535 8449 1544 8483
rect 1492 8440 1544 8449
rect 2228 8483 2280 8492
rect 2228 8449 2237 8483
rect 2237 8449 2271 8483
rect 2271 8449 2280 8483
rect 2228 8440 2280 8449
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 4620 8483 4672 8492
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 4620 8440 4672 8449
rect 8208 8619 8260 8628
rect 8208 8585 8217 8619
rect 8217 8585 8251 8619
rect 8251 8585 8260 8619
rect 8208 8576 8260 8585
rect 9312 8576 9364 8628
rect 10508 8576 10560 8628
rect 7288 8551 7340 8560
rect 7288 8517 7297 8551
rect 7297 8517 7331 8551
rect 7331 8517 7340 8551
rect 7288 8508 7340 8517
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 8300 8440 8352 8492
rect 9496 8440 9548 8492
rect 11704 8576 11756 8628
rect 13176 8619 13228 8628
rect 13176 8585 13185 8619
rect 13185 8585 13219 8619
rect 13219 8585 13228 8619
rect 13176 8576 13228 8585
rect 11152 8483 11204 8492
rect 11152 8449 11161 8483
rect 11161 8449 11195 8483
rect 11195 8449 11204 8483
rect 11152 8440 11204 8449
rect 11796 8483 11848 8492
rect 11796 8449 11805 8483
rect 11805 8449 11839 8483
rect 11839 8449 11848 8483
rect 11796 8440 11848 8449
rect 14096 8576 14148 8628
rect 15384 8619 15436 8628
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 17776 8619 17828 8628
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 19156 8576 19208 8628
rect 20076 8576 20128 8628
rect 21272 8576 21324 8628
rect 22468 8576 22520 8628
rect 23664 8576 23716 8628
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 17684 8483 17736 8492
rect 17684 8449 17693 8483
rect 17693 8449 17727 8483
rect 17727 8449 17736 8483
rect 17684 8440 17736 8449
rect 19156 8440 19208 8492
rect 22560 8483 22612 8492
rect 22560 8449 22569 8483
rect 22569 8449 22603 8483
rect 22603 8449 22612 8483
rect 22560 8440 22612 8449
rect 23112 8483 23164 8492
rect 23112 8449 23121 8483
rect 23121 8449 23155 8483
rect 23155 8449 23164 8483
rect 23112 8440 23164 8449
rect 23572 8440 23624 8492
rect 23664 8483 23716 8492
rect 23664 8449 23673 8483
rect 23673 8449 23707 8483
rect 23707 8449 23716 8483
rect 23664 8440 23716 8449
rect 16488 8304 16540 8356
rect 22100 8372 22152 8424
rect 3917 8134 3969 8186
rect 3981 8134 4033 8186
rect 4045 8134 4097 8186
rect 4109 8134 4161 8186
rect 4173 8134 4225 8186
rect 9851 8134 9903 8186
rect 9915 8134 9967 8186
rect 9979 8134 10031 8186
rect 10043 8134 10095 8186
rect 10107 8134 10159 8186
rect 15785 8134 15837 8186
rect 15849 8134 15901 8186
rect 15913 8134 15965 8186
rect 15977 8134 16029 8186
rect 16041 8134 16093 8186
rect 21719 8134 21771 8186
rect 21783 8134 21835 8186
rect 21847 8134 21899 8186
rect 21911 8134 21963 8186
rect 21975 8134 22027 8186
rect 6552 8032 6604 8084
rect 7564 8032 7616 8084
rect 11152 8075 11204 8084
rect 11152 8041 11161 8075
rect 11161 8041 11195 8075
rect 11195 8041 11204 8075
rect 11152 8032 11204 8041
rect 13544 8032 13596 8084
rect 17408 8032 17460 8084
rect 23112 8032 23164 8084
rect 23664 8032 23716 8084
rect 24492 8032 24544 8084
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 6276 7828 6328 7837
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 11060 7871 11112 7880
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 23848 7896 23900 7948
rect 22192 7692 22244 7744
rect 23664 7871 23716 7880
rect 23664 7837 23673 7871
rect 23673 7837 23707 7871
rect 23707 7837 23716 7871
rect 23664 7828 23716 7837
rect 23940 7760 23992 7812
rect 24400 7692 24452 7744
rect 6884 7590 6936 7642
rect 6948 7590 7000 7642
rect 7012 7590 7064 7642
rect 7076 7590 7128 7642
rect 7140 7590 7192 7642
rect 12818 7590 12870 7642
rect 12882 7590 12934 7642
rect 12946 7590 12998 7642
rect 13010 7590 13062 7642
rect 13074 7590 13126 7642
rect 18752 7590 18804 7642
rect 18816 7590 18868 7642
rect 18880 7590 18932 7642
rect 18944 7590 18996 7642
rect 19008 7590 19060 7642
rect 24686 7590 24738 7642
rect 24750 7590 24802 7642
rect 24814 7590 24866 7642
rect 24878 7590 24930 7642
rect 24942 7590 24994 7642
rect 6276 7488 6328 7540
rect 7472 7488 7524 7540
rect 11060 7488 11112 7540
rect 23388 7488 23440 7540
rect 23664 7488 23716 7540
rect 23020 7352 23072 7404
rect 23204 7352 23256 7404
rect 8208 7148 8260 7200
rect 3917 7046 3969 7098
rect 3981 7046 4033 7098
rect 4045 7046 4097 7098
rect 4109 7046 4161 7098
rect 4173 7046 4225 7098
rect 9851 7046 9903 7098
rect 9915 7046 9967 7098
rect 9979 7046 10031 7098
rect 10043 7046 10095 7098
rect 10107 7046 10159 7098
rect 15785 7046 15837 7098
rect 15849 7046 15901 7098
rect 15913 7046 15965 7098
rect 15977 7046 16029 7098
rect 16041 7046 16093 7098
rect 21719 7046 21771 7098
rect 21783 7046 21835 7098
rect 21847 7046 21899 7098
rect 21911 7046 21963 7098
rect 21975 7046 22027 7098
rect 6884 6502 6936 6554
rect 6948 6502 7000 6554
rect 7012 6502 7064 6554
rect 7076 6502 7128 6554
rect 7140 6502 7192 6554
rect 12818 6502 12870 6554
rect 12882 6502 12934 6554
rect 12946 6502 12998 6554
rect 13010 6502 13062 6554
rect 13074 6502 13126 6554
rect 18752 6502 18804 6554
rect 18816 6502 18868 6554
rect 18880 6502 18932 6554
rect 18944 6502 18996 6554
rect 19008 6502 19060 6554
rect 24686 6502 24738 6554
rect 24750 6502 24802 6554
rect 24814 6502 24866 6554
rect 24878 6502 24930 6554
rect 24942 6502 24994 6554
rect 3917 5958 3969 6010
rect 3981 5958 4033 6010
rect 4045 5958 4097 6010
rect 4109 5958 4161 6010
rect 4173 5958 4225 6010
rect 9851 5958 9903 6010
rect 9915 5958 9967 6010
rect 9979 5958 10031 6010
rect 10043 5958 10095 6010
rect 10107 5958 10159 6010
rect 15785 5958 15837 6010
rect 15849 5958 15901 6010
rect 15913 5958 15965 6010
rect 15977 5958 16029 6010
rect 16041 5958 16093 6010
rect 21719 5958 21771 6010
rect 21783 5958 21835 6010
rect 21847 5958 21899 6010
rect 21911 5958 21963 6010
rect 21975 5958 22027 6010
rect 14188 5856 14240 5908
rect 2228 5720 2280 5772
rect 14648 5695 14700 5704
rect 14648 5661 14657 5695
rect 14657 5661 14691 5695
rect 14691 5661 14700 5695
rect 14648 5652 14700 5661
rect 19432 5652 19484 5704
rect 1492 5516 1544 5568
rect 22468 5516 22520 5568
rect 6884 5414 6936 5466
rect 6948 5414 7000 5466
rect 7012 5414 7064 5466
rect 7076 5414 7128 5466
rect 7140 5414 7192 5466
rect 12818 5414 12870 5466
rect 12882 5414 12934 5466
rect 12946 5414 12998 5466
rect 13010 5414 13062 5466
rect 13074 5414 13126 5466
rect 18752 5414 18804 5466
rect 18816 5414 18868 5466
rect 18880 5414 18932 5466
rect 18944 5414 18996 5466
rect 19008 5414 19060 5466
rect 24686 5414 24738 5466
rect 24750 5414 24802 5466
rect 24814 5414 24866 5466
rect 24878 5414 24930 5466
rect 24942 5414 24994 5466
rect 11796 5312 11848 5364
rect 14648 5355 14700 5364
rect 14648 5321 14657 5355
rect 14657 5321 14691 5355
rect 14691 5321 14700 5355
rect 14648 5312 14700 5321
rect 12348 5219 12400 5228
rect 12348 5185 12357 5219
rect 12357 5185 12391 5219
rect 12391 5185 12400 5219
rect 12348 5176 12400 5185
rect 19432 5355 19484 5364
rect 19432 5321 19441 5355
rect 19441 5321 19475 5355
rect 19475 5321 19484 5355
rect 19432 5312 19484 5321
rect 19616 5219 19668 5228
rect 19616 5185 19625 5219
rect 19625 5185 19659 5219
rect 19659 5185 19668 5219
rect 19616 5176 19668 5185
rect 20720 5108 20772 5160
rect 3917 4870 3969 4922
rect 3981 4870 4033 4922
rect 4045 4870 4097 4922
rect 4109 4870 4161 4922
rect 4173 4870 4225 4922
rect 9851 4870 9903 4922
rect 9915 4870 9967 4922
rect 9979 4870 10031 4922
rect 10043 4870 10095 4922
rect 10107 4870 10159 4922
rect 15785 4870 15837 4922
rect 15849 4870 15901 4922
rect 15913 4870 15965 4922
rect 15977 4870 16029 4922
rect 16041 4870 16093 4922
rect 21719 4870 21771 4922
rect 21783 4870 21835 4922
rect 21847 4870 21899 4922
rect 21911 4870 21963 4922
rect 21975 4870 22027 4922
rect 12348 4768 12400 4820
rect 19616 4768 19668 4820
rect 20996 4564 21048 4616
rect 23664 4496 23716 4548
rect 6884 4326 6936 4378
rect 6948 4326 7000 4378
rect 7012 4326 7064 4378
rect 7076 4326 7128 4378
rect 7140 4326 7192 4378
rect 12818 4326 12870 4378
rect 12882 4326 12934 4378
rect 12946 4326 12998 4378
rect 13010 4326 13062 4378
rect 13074 4326 13126 4378
rect 18752 4326 18804 4378
rect 18816 4326 18868 4378
rect 18880 4326 18932 4378
rect 18944 4326 18996 4378
rect 19008 4326 19060 4378
rect 24686 4326 24738 4378
rect 24750 4326 24802 4378
rect 24814 4326 24866 4378
rect 24878 4326 24930 4378
rect 24942 4326 24994 4378
rect 8300 4020 8352 4072
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 9680 4131 9732 4140
rect 9680 4097 9689 4131
rect 9689 4097 9723 4131
rect 9723 4097 9732 4131
rect 9680 4088 9732 4097
rect 24308 4131 24360 4140
rect 24308 4097 24317 4131
rect 24317 4097 24351 4131
rect 24351 4097 24360 4131
rect 24308 4088 24360 4097
rect 9496 3995 9548 4004
rect 9496 3961 9505 3995
rect 9505 3961 9539 3995
rect 9539 3961 9548 3995
rect 9496 3952 9548 3961
rect 24124 3927 24176 3936
rect 24124 3893 24133 3927
rect 24133 3893 24167 3927
rect 24167 3893 24176 3927
rect 24124 3884 24176 3893
rect 3917 3782 3969 3834
rect 3981 3782 4033 3834
rect 4045 3782 4097 3834
rect 4109 3782 4161 3834
rect 4173 3782 4225 3834
rect 9851 3782 9903 3834
rect 9915 3782 9967 3834
rect 9979 3782 10031 3834
rect 10043 3782 10095 3834
rect 10107 3782 10159 3834
rect 15785 3782 15837 3834
rect 15849 3782 15901 3834
rect 15913 3782 15965 3834
rect 15977 3782 16029 3834
rect 16041 3782 16093 3834
rect 21719 3782 21771 3834
rect 21783 3782 21835 3834
rect 21847 3782 21899 3834
rect 21911 3782 21963 3834
rect 21975 3782 22027 3834
rect 8852 3680 8904 3732
rect 9680 3680 9732 3732
rect 23388 3723 23440 3732
rect 23388 3689 23397 3723
rect 23397 3689 23431 3723
rect 23431 3689 23440 3723
rect 23388 3680 23440 3689
rect 23664 3723 23716 3732
rect 23664 3689 23673 3723
rect 23673 3689 23707 3723
rect 23707 3689 23716 3723
rect 23664 3680 23716 3689
rect 24308 3680 24360 3732
rect 3792 3612 3844 3664
rect 23480 3612 23532 3664
rect 25320 3612 25372 3664
rect 23112 3544 23164 3596
rect 24584 3544 24636 3596
rect 9496 3451 9548 3460
rect 9496 3417 9505 3451
rect 9505 3417 9539 3451
rect 9539 3417 9548 3451
rect 9496 3408 9548 3417
rect 13912 3476 13964 3528
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 22652 3476 22704 3528
rect 22836 3408 22888 3460
rect 24492 3476 24544 3528
rect 25596 3408 25648 3460
rect 23756 3340 23808 3392
rect 6884 3238 6936 3290
rect 6948 3238 7000 3290
rect 7012 3238 7064 3290
rect 7076 3238 7128 3290
rect 7140 3238 7192 3290
rect 12818 3238 12870 3290
rect 12882 3238 12934 3290
rect 12946 3238 12998 3290
rect 13010 3238 13062 3290
rect 13074 3238 13126 3290
rect 18752 3238 18804 3290
rect 18816 3238 18868 3290
rect 18880 3238 18932 3290
rect 18944 3238 18996 3290
rect 19008 3238 19060 3290
rect 24686 3238 24738 3290
rect 24750 3238 24802 3290
rect 24814 3238 24866 3290
rect 24878 3238 24930 3290
rect 24942 3238 24994 3290
rect 756 3068 808 3120
rect 204 3000 256 3052
rect 480 2932 532 2984
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 4620 3136 4672 3188
rect 20076 3136 20128 3188
rect 20720 3136 20772 3188
rect 24216 3136 24268 3188
rect 23296 3068 23348 3120
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 21088 3000 21140 3052
rect 22928 3000 22980 3052
rect 23112 3000 23164 3052
rect 23480 3043 23532 3052
rect 23480 3009 23489 3043
rect 23489 3009 23523 3043
rect 23523 3009 23532 3043
rect 23480 3000 23532 3009
rect 23664 3000 23716 3052
rect 1584 2796 1636 2848
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 9404 2864 9456 2916
rect 13452 2864 13504 2916
rect 20444 2864 20496 2916
rect 22284 2864 22336 2916
rect 9312 2796 9364 2848
rect 12624 2796 12676 2848
rect 19432 2796 19484 2848
rect 23020 2839 23072 2848
rect 23020 2805 23029 2839
rect 23029 2805 23063 2839
rect 23063 2805 23072 2839
rect 23020 2796 23072 2805
rect 23204 2796 23256 2848
rect 23940 2864 23992 2916
rect 24032 2864 24084 2916
rect 3917 2694 3969 2746
rect 3981 2694 4033 2746
rect 4045 2694 4097 2746
rect 4109 2694 4161 2746
rect 4173 2694 4225 2746
rect 9851 2694 9903 2746
rect 9915 2694 9967 2746
rect 9979 2694 10031 2746
rect 10043 2694 10095 2746
rect 10107 2694 10159 2746
rect 15785 2694 15837 2746
rect 15849 2694 15901 2746
rect 15913 2694 15965 2746
rect 15977 2694 16029 2746
rect 16041 2694 16093 2746
rect 21719 2694 21771 2746
rect 21783 2694 21835 2746
rect 21847 2694 21899 2746
rect 21911 2694 21963 2746
rect 21975 2694 22027 2746
rect 1676 2592 1728 2644
rect 2044 2592 2096 2644
rect 9036 2592 9088 2644
rect 1492 2524 1544 2576
rect 9312 2524 9364 2576
rect 1308 2388 1360 2440
rect 1584 2388 1636 2440
rect 3148 2456 3200 2508
rect 1492 2320 1544 2372
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 4620 2388 4672 2440
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 6368 2388 6420 2397
rect 9220 2456 9272 2508
rect 9956 2456 10008 2508
rect 17224 2524 17276 2576
rect 17684 2592 17736 2644
rect 19156 2592 19208 2644
rect 20076 2592 20128 2644
rect 21088 2635 21140 2644
rect 21088 2601 21097 2635
rect 21097 2601 21131 2635
rect 21131 2601 21140 2635
rect 21088 2592 21140 2601
rect 22100 2635 22152 2644
rect 22100 2601 22109 2635
rect 22109 2601 22143 2635
rect 22143 2601 22152 2635
rect 22100 2592 22152 2601
rect 22192 2592 22244 2644
rect 22560 2592 22612 2644
rect 23296 2635 23348 2644
rect 23296 2601 23305 2635
rect 23305 2601 23339 2635
rect 23339 2601 23348 2635
rect 23296 2592 23348 2601
rect 23940 2592 23992 2644
rect 24400 2592 24452 2644
rect 1676 2295 1728 2304
rect 1676 2261 1685 2295
rect 1685 2261 1719 2295
rect 1719 2261 1728 2295
rect 1676 2252 1728 2261
rect 2228 2295 2280 2304
rect 2228 2261 2237 2295
rect 2237 2261 2271 2295
rect 2271 2261 2280 2295
rect 2228 2252 2280 2261
rect 8852 2320 8904 2372
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 10324 2320 10376 2372
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12532 2388 12584 2440
rect 13268 2456 13320 2508
rect 13452 2431 13504 2440
rect 13452 2397 13461 2431
rect 13461 2397 13495 2431
rect 13495 2397 13504 2431
rect 13452 2388 13504 2397
rect 15108 2431 15160 2440
rect 15108 2397 15117 2431
rect 15117 2397 15151 2431
rect 15151 2397 15160 2431
rect 15108 2388 15160 2397
rect 15476 2456 15528 2508
rect 19340 2524 19392 2576
rect 19616 2524 19668 2576
rect 22836 2524 22888 2576
rect 4712 2295 4764 2304
rect 4712 2261 4721 2295
rect 4721 2261 4755 2295
rect 4755 2261 4764 2295
rect 4712 2252 4764 2261
rect 4804 2252 4856 2304
rect 5080 2252 5132 2304
rect 6552 2295 6604 2304
rect 6552 2261 6561 2295
rect 6561 2261 6595 2295
rect 6595 2261 6604 2295
rect 6552 2252 6604 2261
rect 6736 2252 6788 2304
rect 9220 2252 9272 2304
rect 11520 2295 11572 2304
rect 11520 2261 11529 2295
rect 11529 2261 11563 2295
rect 11563 2261 11572 2295
rect 11520 2252 11572 2261
rect 11704 2252 11756 2304
rect 13728 2320 13780 2372
rect 16672 2388 16724 2440
rect 16856 2388 16908 2440
rect 13268 2295 13320 2304
rect 13268 2261 13277 2295
rect 13277 2261 13311 2295
rect 13311 2261 13320 2295
rect 13268 2252 13320 2261
rect 15200 2295 15252 2304
rect 15200 2261 15209 2295
rect 15209 2261 15243 2295
rect 15243 2261 15252 2295
rect 15200 2252 15252 2261
rect 15384 2252 15436 2304
rect 16488 2252 16540 2304
rect 16580 2295 16632 2304
rect 16580 2261 16589 2295
rect 16589 2261 16623 2295
rect 16623 2261 16632 2295
rect 16580 2252 16632 2261
rect 17132 2252 17184 2304
rect 18420 2388 18472 2440
rect 19156 2388 19208 2440
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 20628 2456 20680 2508
rect 21640 2456 21692 2508
rect 19892 2388 19944 2440
rect 19984 2431 20036 2440
rect 19984 2397 19993 2431
rect 19993 2397 20027 2431
rect 20027 2397 20036 2431
rect 19984 2388 20036 2397
rect 20720 2431 20772 2440
rect 20720 2397 20729 2431
rect 20729 2397 20763 2431
rect 20763 2397 20772 2431
rect 20720 2388 20772 2397
rect 21180 2388 21232 2440
rect 21824 2431 21876 2440
rect 21824 2397 21833 2431
rect 21833 2397 21867 2431
rect 21867 2397 21876 2431
rect 21824 2388 21876 2397
rect 18144 2295 18196 2304
rect 18144 2261 18153 2295
rect 18153 2261 18187 2295
rect 18187 2261 18196 2295
rect 18144 2252 18196 2261
rect 18420 2295 18472 2304
rect 18420 2261 18429 2295
rect 18429 2261 18463 2295
rect 18463 2261 18472 2295
rect 18420 2252 18472 2261
rect 18512 2252 18564 2304
rect 19524 2295 19576 2304
rect 19524 2261 19533 2295
rect 19533 2261 19567 2295
rect 19567 2261 19576 2295
rect 19524 2252 19576 2261
rect 20076 2295 20128 2304
rect 20076 2261 20085 2295
rect 20085 2261 20119 2295
rect 20119 2261 20128 2295
rect 20076 2252 20128 2261
rect 22008 2320 22060 2372
rect 21456 2252 21508 2304
rect 23388 2456 23440 2508
rect 23940 2456 23992 2508
rect 22376 2431 22428 2440
rect 22376 2397 22385 2431
rect 22385 2397 22419 2431
rect 22419 2397 22428 2431
rect 22376 2388 22428 2397
rect 22836 2388 22888 2440
rect 22744 2295 22796 2304
rect 22744 2261 22753 2295
rect 22753 2261 22787 2295
rect 22787 2261 22796 2295
rect 22744 2252 22796 2261
rect 23204 2431 23256 2440
rect 23204 2397 23213 2431
rect 23213 2397 23247 2431
rect 23247 2397 23256 2431
rect 23204 2388 23256 2397
rect 23572 2431 23624 2440
rect 23572 2397 23581 2431
rect 23581 2397 23615 2431
rect 23615 2397 23624 2431
rect 23572 2388 23624 2397
rect 24308 2388 24360 2440
rect 23756 2320 23808 2372
rect 25044 2252 25096 2304
rect 6884 2150 6936 2202
rect 6948 2150 7000 2202
rect 7012 2150 7064 2202
rect 7076 2150 7128 2202
rect 7140 2150 7192 2202
rect 12818 2150 12870 2202
rect 12882 2150 12934 2202
rect 12946 2150 12998 2202
rect 13010 2150 13062 2202
rect 13074 2150 13126 2202
rect 18752 2150 18804 2202
rect 18816 2150 18868 2202
rect 18880 2150 18932 2202
rect 18944 2150 18996 2202
rect 19008 2150 19060 2202
rect 24686 2150 24738 2202
rect 24750 2150 24802 2202
rect 24814 2150 24866 2202
rect 24878 2150 24930 2202
rect 24942 2150 24994 2202
rect 1676 2048 1728 2100
rect 1584 1955 1636 1964
rect 1584 1921 1593 1955
rect 1593 1921 1627 1955
rect 1627 1921 1636 1955
rect 1584 1912 1636 1921
rect 2228 1980 2280 2032
rect 3148 1980 3200 2032
rect 1032 1776 1084 1828
rect 2688 1912 2740 1964
rect 2780 1955 2832 1964
rect 2780 1921 2789 1955
rect 2789 1921 2823 1955
rect 2823 1921 2832 1955
rect 2780 1912 2832 1921
rect 3056 1955 3108 1964
rect 3056 1921 3065 1955
rect 3065 1921 3099 1955
rect 3099 1921 3108 1955
rect 3056 1912 3108 1921
rect 4252 2091 4304 2100
rect 4252 2057 4261 2091
rect 4261 2057 4295 2091
rect 4295 2057 4304 2091
rect 4252 2048 4304 2057
rect 4712 2048 4764 2100
rect 3608 1955 3660 1964
rect 3608 1921 3617 1955
rect 3617 1921 3651 1955
rect 3651 1921 3660 1955
rect 3608 1912 3660 1921
rect 3884 1955 3936 1964
rect 3884 1921 3893 1955
rect 3893 1921 3927 1955
rect 3927 1921 3936 1955
rect 3884 1912 3936 1921
rect 4344 1912 4396 1964
rect 4436 1955 4488 1964
rect 4436 1921 4445 1955
rect 4445 1921 4479 1955
rect 4479 1921 4488 1955
rect 4436 1912 4488 1921
rect 6644 2091 6696 2100
rect 6644 2057 6653 2091
rect 6653 2057 6687 2091
rect 6687 2057 6696 2091
rect 6644 2048 6696 2057
rect 7380 2048 7432 2100
rect 7932 2048 7984 2100
rect 8116 2091 8168 2100
rect 8116 2057 8125 2091
rect 8125 2057 8159 2091
rect 8159 2057 8168 2091
rect 8116 2048 8168 2057
rect 8944 2091 8996 2100
rect 8944 2057 8953 2091
rect 8953 2057 8987 2091
rect 8987 2057 8996 2091
rect 8944 2048 8996 2057
rect 9220 2048 9272 2100
rect 9680 2048 9732 2100
rect 5908 1955 5960 1964
rect 5908 1921 5917 1955
rect 5917 1921 5951 1955
rect 5951 1921 5960 1955
rect 5908 1912 5960 1921
rect 6460 1955 6512 1964
rect 6460 1921 6469 1955
rect 6469 1921 6503 1955
rect 6503 1921 6512 1955
rect 6460 1912 6512 1921
rect 7288 1980 7340 2032
rect 6828 1912 6880 1964
rect 2044 1708 2096 1760
rect 3516 1776 3568 1828
rect 2688 1708 2740 1760
rect 2964 1708 3016 1760
rect 3240 1708 3292 1760
rect 5632 1776 5684 1828
rect 7012 1819 7064 1828
rect 7012 1785 7021 1819
rect 7021 1785 7055 1819
rect 7055 1785 7064 1819
rect 7012 1776 7064 1785
rect 7472 1955 7524 1964
rect 7472 1921 7481 1955
rect 7481 1921 7515 1955
rect 7515 1921 7524 1955
rect 7472 1912 7524 1921
rect 7840 1912 7892 1964
rect 7564 1844 7616 1896
rect 4712 1708 4764 1760
rect 5540 1708 5592 1760
rect 7840 1819 7892 1828
rect 7840 1785 7849 1819
rect 7849 1785 7883 1819
rect 7883 1785 7892 1819
rect 7840 1776 7892 1785
rect 8024 1955 8076 1964
rect 8024 1921 8033 1955
rect 8033 1921 8067 1955
rect 8067 1921 8076 1955
rect 8024 1912 8076 1921
rect 8300 1955 8352 1964
rect 8300 1921 8309 1955
rect 8309 1921 8343 1955
rect 8343 1921 8352 1955
rect 8300 1912 8352 1921
rect 8576 1955 8628 1964
rect 8576 1921 8585 1955
rect 8585 1921 8619 1955
rect 8619 1921 8628 1955
rect 8576 1912 8628 1921
rect 8852 1955 8904 1964
rect 8852 1921 8861 1955
rect 8861 1921 8895 1955
rect 8895 1921 8904 1955
rect 8852 1912 8904 1921
rect 9128 1955 9180 1964
rect 9128 1921 9137 1955
rect 9137 1921 9171 1955
rect 9171 1921 9180 1955
rect 9128 1912 9180 1921
rect 9404 1955 9456 1964
rect 9404 1921 9413 1955
rect 9413 1921 9447 1955
rect 9447 1921 9456 1955
rect 9404 1912 9456 1921
rect 9772 1912 9824 1964
rect 9864 1912 9916 1964
rect 8668 1751 8720 1760
rect 8668 1717 8677 1751
rect 8677 1717 8711 1751
rect 8711 1717 8720 1751
rect 8668 1708 8720 1717
rect 9404 1776 9456 1828
rect 10324 1912 10376 1964
rect 11520 2048 11572 2100
rect 12256 2048 12308 2100
rect 13176 2048 13228 2100
rect 13268 2048 13320 2100
rect 13728 2048 13780 2100
rect 12624 1955 12676 1964
rect 12624 1921 12633 1955
rect 12633 1921 12667 1955
rect 12667 1921 12676 1955
rect 12624 1912 12676 1921
rect 12808 1955 12860 1964
rect 12808 1921 12817 1955
rect 12817 1921 12851 1955
rect 12851 1921 12860 1955
rect 12808 1912 12860 1921
rect 13636 1955 13688 1964
rect 13636 1921 13645 1955
rect 13645 1921 13679 1955
rect 13679 1921 13688 1955
rect 13636 1912 13688 1921
rect 14096 1912 14148 1964
rect 9864 1708 9916 1760
rect 13360 1844 13412 1896
rect 15200 2048 15252 2100
rect 16580 2048 16632 2100
rect 16672 2048 16724 2100
rect 10508 1751 10560 1760
rect 10508 1717 10517 1751
rect 10517 1717 10551 1751
rect 10551 1717 10560 1751
rect 10508 1708 10560 1717
rect 11060 1751 11112 1760
rect 11060 1717 11069 1751
rect 11069 1717 11103 1751
rect 11103 1717 11112 1751
rect 11060 1708 11112 1717
rect 11888 1776 11940 1828
rect 11796 1708 11848 1760
rect 12624 1708 12676 1760
rect 15108 1912 15160 1964
rect 18144 2048 18196 2100
rect 18420 2048 18472 2100
rect 19524 2048 19576 2100
rect 19800 2048 19852 2100
rect 21456 2048 21508 2100
rect 21824 2091 21876 2100
rect 21824 2057 21833 2091
rect 21833 2057 21867 2091
rect 21867 2057 21876 2091
rect 21824 2048 21876 2057
rect 15660 1955 15712 1964
rect 15660 1921 15669 1955
rect 15669 1921 15703 1955
rect 15703 1921 15712 1955
rect 15660 1912 15712 1921
rect 16212 1912 16264 1964
rect 15292 1844 15344 1896
rect 21548 1980 21600 2032
rect 22376 2048 22428 2100
rect 22744 2048 22796 2100
rect 16948 1844 17000 1896
rect 16488 1776 16540 1828
rect 18972 1844 19024 1896
rect 20076 1912 20128 1964
rect 21732 1912 21784 1964
rect 22468 1980 22520 2032
rect 23204 2048 23256 2100
rect 24032 2091 24084 2100
rect 24032 2057 24041 2091
rect 24041 2057 24075 2091
rect 24075 2057 24084 2091
rect 24032 2048 24084 2057
rect 24308 2091 24360 2100
rect 24308 2057 24317 2091
rect 24317 2057 24351 2091
rect 24351 2057 24360 2091
rect 24308 2048 24360 2057
rect 22284 1955 22336 1964
rect 22284 1921 22293 1955
rect 22293 1921 22327 1955
rect 22327 1921 22336 1955
rect 22284 1912 22336 1921
rect 20628 1844 20680 1896
rect 19340 1819 19392 1828
rect 19340 1785 19349 1819
rect 19349 1785 19383 1819
rect 19383 1785 19392 1819
rect 19340 1776 19392 1785
rect 20444 1819 20496 1828
rect 20444 1785 20453 1819
rect 20453 1785 20487 1819
rect 20487 1785 20496 1819
rect 20444 1776 20496 1785
rect 21180 1776 21232 1828
rect 14004 1708 14056 1760
rect 14096 1751 14148 1760
rect 14096 1717 14105 1751
rect 14105 1717 14139 1751
rect 14139 1717 14148 1751
rect 14096 1708 14148 1717
rect 14280 1708 14332 1760
rect 14740 1708 14792 1760
rect 15200 1751 15252 1760
rect 15200 1717 15209 1751
rect 15209 1717 15243 1751
rect 15243 1717 15252 1751
rect 15200 1708 15252 1717
rect 15660 1708 15712 1760
rect 16580 1708 16632 1760
rect 16764 1708 16816 1760
rect 17960 1708 18012 1760
rect 18236 1708 18288 1760
rect 19708 1708 19760 1760
rect 19892 1708 19944 1760
rect 21548 1708 21600 1760
rect 23020 1912 23072 1964
rect 23112 1819 23164 1828
rect 23112 1785 23121 1819
rect 23121 1785 23155 1819
rect 23155 1785 23164 1819
rect 23112 1776 23164 1785
rect 24216 1955 24268 1964
rect 24216 1921 24225 1955
rect 24225 1921 24259 1955
rect 24259 1921 24268 1955
rect 24216 1912 24268 1921
rect 24400 1912 24452 1964
rect 3917 1606 3969 1658
rect 3981 1606 4033 1658
rect 4045 1606 4097 1658
rect 4109 1606 4161 1658
rect 4173 1606 4225 1658
rect 9851 1606 9903 1658
rect 9915 1606 9967 1658
rect 9979 1606 10031 1658
rect 10043 1606 10095 1658
rect 10107 1606 10159 1658
rect 15785 1606 15837 1658
rect 15849 1606 15901 1658
rect 15913 1606 15965 1658
rect 15977 1606 16029 1658
rect 16041 1606 16093 1658
rect 21719 1606 21771 1658
rect 21783 1606 21835 1658
rect 21847 1606 21899 1658
rect 21911 1606 21963 1658
rect 21975 1606 22027 1658
rect 2688 1504 2740 1556
rect 4436 1504 4488 1556
rect 4528 1504 4580 1556
rect 6736 1504 6788 1556
rect 7012 1504 7064 1556
rect 7564 1504 7616 1556
rect 7932 1504 7984 1556
rect 1492 1343 1544 1352
rect 1492 1309 1501 1343
rect 1501 1309 1535 1343
rect 1535 1309 1544 1343
rect 1492 1300 1544 1309
rect 1952 1343 2004 1352
rect 1952 1309 1961 1343
rect 1961 1309 1995 1343
rect 1995 1309 2004 1343
rect 1952 1300 2004 1309
rect 2964 1300 3016 1352
rect 3240 1300 3292 1352
rect 3332 1343 3384 1352
rect 3332 1309 3341 1343
rect 3341 1309 3375 1343
rect 3375 1309 3384 1343
rect 3332 1300 3384 1309
rect 4804 1368 4856 1420
rect 7472 1436 7524 1488
rect 8024 1436 8076 1488
rect 4528 1343 4580 1352
rect 4528 1309 4537 1343
rect 4537 1309 4571 1343
rect 4571 1309 4580 1343
rect 4528 1300 4580 1309
rect 4988 1300 5040 1352
rect 5080 1343 5132 1352
rect 5080 1309 5089 1343
rect 5089 1309 5123 1343
rect 5123 1309 5132 1343
rect 5080 1300 5132 1309
rect 5540 1300 5592 1352
rect 1676 1207 1728 1216
rect 1676 1173 1685 1207
rect 1685 1173 1719 1207
rect 1719 1173 1728 1207
rect 1676 1164 1728 1173
rect 1768 1207 1820 1216
rect 1768 1173 1777 1207
rect 1777 1173 1811 1207
rect 1811 1173 1820 1207
rect 1768 1164 1820 1173
rect 2320 1207 2372 1216
rect 2320 1173 2329 1207
rect 2329 1173 2363 1207
rect 2363 1173 2372 1207
rect 2320 1164 2372 1173
rect 2596 1207 2648 1216
rect 2596 1173 2605 1207
rect 2605 1173 2639 1207
rect 2639 1173 2648 1207
rect 2596 1164 2648 1173
rect 4160 1164 4212 1216
rect 4436 1232 4488 1284
rect 5724 1343 5776 1352
rect 5724 1309 5733 1343
rect 5733 1309 5767 1343
rect 5767 1309 5776 1343
rect 5724 1300 5776 1309
rect 6184 1343 6236 1352
rect 6184 1309 6193 1343
rect 6193 1309 6227 1343
rect 6227 1309 6236 1343
rect 6184 1300 6236 1309
rect 6736 1300 6788 1352
rect 6920 1343 6972 1352
rect 6920 1309 6929 1343
rect 6929 1309 6963 1343
rect 6963 1309 6972 1343
rect 6920 1300 6972 1309
rect 7748 1343 7800 1352
rect 7748 1309 7757 1343
rect 7757 1309 7791 1343
rect 7791 1309 7800 1343
rect 7748 1300 7800 1309
rect 7840 1300 7892 1352
rect 8852 1368 8904 1420
rect 8668 1300 8720 1352
rect 9036 1300 9088 1352
rect 9312 1368 9364 1420
rect 11060 1411 11112 1420
rect 11060 1377 11069 1411
rect 11069 1377 11103 1411
rect 11103 1377 11112 1411
rect 11060 1368 11112 1377
rect 13360 1504 13412 1556
rect 13820 1504 13872 1556
rect 15108 1504 15160 1556
rect 14096 1436 14148 1488
rect 4804 1207 4856 1216
rect 4804 1173 4813 1207
rect 4813 1173 4847 1207
rect 4847 1173 4856 1207
rect 4804 1164 4856 1173
rect 5356 1207 5408 1216
rect 5356 1173 5365 1207
rect 5365 1173 5399 1207
rect 5399 1173 5408 1207
rect 5356 1164 5408 1173
rect 5448 1207 5500 1216
rect 5448 1173 5457 1207
rect 5457 1173 5491 1207
rect 5491 1173 5500 1207
rect 5448 1164 5500 1173
rect 5816 1164 5868 1216
rect 8300 1232 8352 1284
rect 9680 1300 9732 1352
rect 11704 1343 11756 1352
rect 11704 1309 11713 1343
rect 11713 1309 11747 1343
rect 11747 1309 11756 1343
rect 11704 1300 11756 1309
rect 6552 1207 6604 1216
rect 6552 1173 6561 1207
rect 6561 1173 6595 1207
rect 6595 1173 6604 1207
rect 6552 1164 6604 1173
rect 6644 1207 6696 1216
rect 6644 1173 6653 1207
rect 6653 1173 6687 1207
rect 6687 1173 6696 1207
rect 6644 1164 6696 1173
rect 7380 1164 7432 1216
rect 7748 1164 7800 1216
rect 7840 1164 7892 1216
rect 8024 1207 8076 1216
rect 8024 1173 8033 1207
rect 8033 1173 8067 1207
rect 8067 1173 8076 1207
rect 8024 1164 8076 1173
rect 9220 1164 9272 1216
rect 9312 1207 9364 1216
rect 9312 1173 9321 1207
rect 9321 1173 9355 1207
rect 9355 1173 9364 1207
rect 9312 1164 9364 1173
rect 9404 1164 9456 1216
rect 10048 1164 10100 1216
rect 10692 1232 10744 1284
rect 10784 1275 10836 1284
rect 10784 1241 10793 1275
rect 10793 1241 10827 1275
rect 10827 1241 10836 1275
rect 10784 1232 10836 1241
rect 11152 1164 11204 1216
rect 11520 1207 11572 1216
rect 11520 1173 11529 1207
rect 11529 1173 11563 1207
rect 11563 1173 11572 1207
rect 11520 1164 11572 1173
rect 11612 1164 11664 1216
rect 12440 1300 12492 1352
rect 12900 1343 12952 1352
rect 12900 1309 12909 1343
rect 12909 1309 12943 1343
rect 12943 1309 12952 1343
rect 12900 1300 12952 1309
rect 13268 1343 13320 1352
rect 13268 1309 13277 1343
rect 13277 1309 13311 1343
rect 13311 1309 13320 1343
rect 13268 1300 13320 1309
rect 14188 1275 14240 1284
rect 14188 1241 14197 1275
rect 14197 1241 14231 1275
rect 14231 1241 14240 1275
rect 14188 1232 14240 1241
rect 12072 1164 12124 1216
rect 12348 1207 12400 1216
rect 12348 1173 12357 1207
rect 12357 1173 12391 1207
rect 12391 1173 12400 1207
rect 12348 1164 12400 1173
rect 13084 1207 13136 1216
rect 13084 1173 13093 1207
rect 13093 1173 13127 1207
rect 13127 1173 13136 1207
rect 13084 1164 13136 1173
rect 13452 1207 13504 1216
rect 13452 1173 13461 1207
rect 13461 1173 13495 1207
rect 13495 1173 13504 1207
rect 13452 1164 13504 1173
rect 14004 1164 14056 1216
rect 15108 1368 15160 1420
rect 16120 1504 16172 1556
rect 16120 1368 16172 1420
rect 15200 1300 15252 1352
rect 16304 1300 16356 1352
rect 16580 1300 16632 1352
rect 17040 1368 17092 1420
rect 19156 1504 19208 1556
rect 17592 1436 17644 1488
rect 18696 1436 18748 1488
rect 20720 1504 20772 1556
rect 21640 1504 21692 1556
rect 22192 1504 22244 1556
rect 22008 1436 22060 1488
rect 16948 1232 17000 1284
rect 17224 1232 17276 1284
rect 17776 1300 17828 1352
rect 18052 1232 18104 1284
rect 18604 1300 18656 1352
rect 19340 1275 19392 1284
rect 19340 1241 19349 1275
rect 19349 1241 19383 1275
rect 19383 1241 19392 1275
rect 19340 1232 19392 1241
rect 19432 1232 19484 1284
rect 16396 1164 16448 1216
rect 18512 1164 18564 1216
rect 20812 1164 20864 1216
rect 20996 1232 21048 1284
rect 22284 1343 22336 1352
rect 22284 1309 22293 1343
rect 22293 1309 22327 1343
rect 22327 1309 22336 1343
rect 22284 1300 22336 1309
rect 22560 1343 22612 1352
rect 22560 1309 22569 1343
rect 22569 1309 22603 1343
rect 22603 1309 22612 1343
rect 22560 1300 22612 1309
rect 22744 1300 22796 1352
rect 23020 1300 23072 1352
rect 23388 1343 23440 1352
rect 23388 1309 23397 1343
rect 23397 1309 23431 1343
rect 23431 1309 23440 1343
rect 23388 1300 23440 1309
rect 23756 1436 23808 1488
rect 24032 1436 24084 1488
rect 23756 1343 23808 1352
rect 23756 1309 23765 1343
rect 23765 1309 23799 1343
rect 23799 1309 23808 1343
rect 23756 1300 23808 1309
rect 23940 1300 23992 1352
rect 24216 1343 24268 1352
rect 24216 1309 24225 1343
rect 24225 1309 24259 1343
rect 24259 1309 24268 1343
rect 24216 1300 24268 1309
rect 21456 1207 21508 1216
rect 21456 1173 21465 1207
rect 21465 1173 21499 1207
rect 21499 1173 21508 1207
rect 21456 1164 21508 1173
rect 23112 1207 23164 1216
rect 23112 1173 23121 1207
rect 23121 1173 23155 1207
rect 23155 1173 23164 1207
rect 23112 1164 23164 1173
rect 23480 1164 23532 1216
rect 23940 1207 23992 1216
rect 23940 1173 23949 1207
rect 23949 1173 23983 1207
rect 23983 1173 23992 1207
rect 23940 1164 23992 1173
rect 6884 1062 6936 1114
rect 6948 1062 7000 1114
rect 7012 1062 7064 1114
rect 7076 1062 7128 1114
rect 7140 1062 7192 1114
rect 12818 1062 12870 1114
rect 12882 1062 12934 1114
rect 12946 1062 12998 1114
rect 13010 1062 13062 1114
rect 13074 1062 13126 1114
rect 18752 1062 18804 1114
rect 18816 1062 18868 1114
rect 18880 1062 18932 1114
rect 18944 1062 18996 1114
rect 19008 1062 19060 1114
rect 24686 1062 24738 1114
rect 24750 1062 24802 1114
rect 24814 1062 24866 1114
rect 24878 1062 24930 1114
rect 24942 1062 24994 1114
rect 4988 960 5040 1012
rect 5540 960 5592 1012
rect 6184 960 6236 1012
rect 7380 960 7432 1012
rect 10784 960 10836 1012
rect 11520 960 11572 1012
rect 1768 892 1820 944
rect 3516 892 3568 944
rect 8024 892 8076 944
rect 9772 892 9824 944
rect 12256 892 12308 944
rect 5448 824 5500 876
rect 9404 824 9456 876
rect 9496 824 9548 876
rect 18052 960 18104 1012
rect 18328 960 18380 1012
rect 18512 960 18564 1012
rect 19708 960 19760 1012
rect 20628 960 20680 1012
rect 22560 960 22612 1012
rect 23940 960 23992 1012
rect 21456 892 21508 944
rect 5632 756 5684 808
rect 6644 756 6696 808
rect 14188 756 14240 808
rect 1952 688 2004 740
rect 2688 688 2740 740
rect 3332 688 3384 740
rect 4068 688 4120 740
rect 4528 688 4580 740
rect 5448 688 5500 740
rect 6736 688 6788 740
rect 7380 688 7432 740
rect 7472 688 7524 740
rect 9036 688 9088 740
rect 9680 688 9732 740
rect 1492 620 1544 672
rect 2412 620 2464 672
rect 4712 620 4764 672
rect 5724 620 5776 672
rect 6828 620 6880 672
rect 16856 688 16908 740
rect 12440 620 12492 672
rect 12900 620 12952 672
rect 13268 620 13320 672
rect 13912 620 13964 672
rect 21640 756 21692 808
rect 23020 824 23072 876
rect 23480 756 23532 808
rect 24216 756 24268 808
rect 21088 688 21140 740
rect 22744 688 22796 740
rect 22008 620 22060 672
rect 23756 620 23808 672
rect 2320 552 2372 604
rect 12072 552 12124 604
rect 4252 484 4304 536
rect 11612 484 11664 536
rect 11980 484 12032 536
rect 2596 416 2648 468
rect 6736 416 6788 468
rect 7748 416 7800 468
rect 19248 484 19300 536
rect 20444 484 20496 536
rect 21180 416 21232 468
rect 21640 416 21692 468
rect 7840 280 7892 332
rect 4804 212 4856 264
rect 8944 212 8996 264
rect 15476 212 15528 264
<< metal2 >>
rect 938 9840 994 10000
rect 1044 9846 1256 9874
rect 952 9738 980 9840
rect 1044 9738 1072 9846
rect 952 9710 1072 9738
rect 1228 8634 1256 9846
rect 2134 9840 2190 10000
rect 3330 9840 3386 10000
rect 4526 9840 4582 10000
rect 5722 9840 5778 10000
rect 6918 9840 6974 10000
rect 7024 9846 7328 9874
rect 2148 8634 2176 9840
rect 3344 8634 3372 9840
rect 4540 8634 4568 9840
rect 5736 8634 5764 9840
rect 6932 9738 6960 9840
rect 7024 9738 7052 9846
rect 6932 9710 7052 9738
rect 6884 8732 7192 8741
rect 6884 8730 6890 8732
rect 6946 8730 6970 8732
rect 7026 8730 7050 8732
rect 7106 8730 7130 8732
rect 7186 8730 7192 8732
rect 6946 8678 6948 8730
rect 7128 8678 7130 8730
rect 6884 8676 6890 8678
rect 6946 8676 6970 8678
rect 7026 8676 7050 8678
rect 7106 8676 7130 8678
rect 7186 8676 7192 8678
rect 6884 8667 7192 8676
rect 1216 8628 1268 8634
rect 1216 8570 1268 8576
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 7300 8566 7328 9846
rect 8114 9840 8170 10000
rect 9310 9840 9366 10000
rect 10506 9840 10562 10000
rect 11702 9840 11758 10000
rect 12898 9840 12954 10000
rect 13004 9846 13216 9874
rect 8128 9058 8156 9840
rect 8128 9030 8248 9058
rect 8220 8634 8248 9030
rect 9324 8634 9352 9840
rect 10520 8634 10548 9840
rect 11716 8634 11744 9840
rect 12912 9738 12940 9840
rect 13004 9738 13032 9846
rect 12912 9710 13032 9738
rect 12818 8732 13126 8741
rect 12818 8730 12824 8732
rect 12880 8730 12904 8732
rect 12960 8730 12984 8732
rect 13040 8730 13064 8732
rect 13120 8730 13126 8732
rect 12880 8678 12882 8730
rect 13062 8678 13064 8730
rect 12818 8676 12824 8678
rect 12880 8676 12904 8678
rect 12960 8676 12984 8678
rect 13040 8676 13064 8678
rect 13120 8676 13126 8678
rect 12818 8667 13126 8676
rect 13188 8634 13216 9846
rect 14094 9840 14150 10000
rect 15290 9840 15346 10000
rect 16486 9840 16542 10000
rect 17682 9840 17738 10000
rect 18878 9840 18934 10000
rect 18984 9846 19196 9874
rect 14108 8634 14136 9840
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 14096 8628 14148 8634
rect 15304 8616 15332 9840
rect 15384 8628 15436 8634
rect 15304 8588 15384 8616
rect 14096 8570 14148 8576
rect 15384 8570 15436 8576
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 1504 5574 1532 8434
rect 2240 5778 2268 8434
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 3804 3670 3832 8434
rect 3917 8188 4225 8197
rect 3917 8186 3923 8188
rect 3979 8186 4003 8188
rect 4059 8186 4083 8188
rect 4139 8186 4163 8188
rect 4219 8186 4225 8188
rect 3979 8134 3981 8186
rect 4161 8134 4163 8186
rect 3917 8132 3923 8134
rect 3979 8132 4003 8134
rect 4059 8132 4083 8134
rect 4139 8132 4163 8134
rect 4219 8132 4225 8134
rect 3917 8123 4225 8132
rect 3917 7100 4225 7109
rect 3917 7098 3923 7100
rect 3979 7098 4003 7100
rect 4059 7098 4083 7100
rect 4139 7098 4163 7100
rect 4219 7098 4225 7100
rect 3979 7046 3981 7098
rect 4161 7046 4163 7098
rect 3917 7044 3923 7046
rect 3979 7044 4003 7046
rect 4059 7044 4083 7046
rect 4139 7044 4163 7046
rect 4219 7044 4225 7046
rect 3917 7035 4225 7044
rect 3917 6012 4225 6021
rect 3917 6010 3923 6012
rect 3979 6010 4003 6012
rect 4059 6010 4083 6012
rect 4139 6010 4163 6012
rect 4219 6010 4225 6012
rect 3979 5958 3981 6010
rect 4161 5958 4163 6010
rect 3917 5956 3923 5958
rect 3979 5956 4003 5958
rect 4059 5956 4083 5958
rect 4139 5956 4163 5958
rect 4219 5956 4225 5958
rect 3917 5947 4225 5956
rect 3917 4924 4225 4933
rect 3917 4922 3923 4924
rect 3979 4922 4003 4924
rect 4059 4922 4083 4924
rect 4139 4922 4163 4924
rect 4219 4922 4225 4924
rect 3979 4870 3981 4922
rect 4161 4870 4163 4922
rect 3917 4868 3923 4870
rect 3979 4868 4003 4870
rect 4059 4868 4083 4870
rect 4139 4868 4163 4870
rect 4219 4868 4225 4870
rect 3917 4859 4225 4868
rect 3917 3836 4225 3845
rect 3917 3834 3923 3836
rect 3979 3834 4003 3836
rect 4059 3834 4083 3836
rect 4139 3834 4163 3836
rect 4219 3834 4225 3836
rect 3979 3782 3981 3834
rect 4161 3782 4163 3834
rect 3917 3780 3923 3782
rect 3979 3780 4003 3782
rect 4059 3780 4083 3782
rect 4139 3780 4163 3782
rect 4219 3780 4225 3782
rect 3917 3771 4225 3780
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 4632 3194 4660 8434
rect 6564 8090 6592 8434
rect 7576 8090 7604 8434
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 6288 7546 6316 7822
rect 6884 7644 7192 7653
rect 6884 7642 6890 7644
rect 6946 7642 6970 7644
rect 7026 7642 7050 7644
rect 7106 7642 7130 7644
rect 7186 7642 7192 7644
rect 6946 7590 6948 7642
rect 7128 7590 7130 7642
rect 6884 7588 6890 7590
rect 6946 7588 6970 7590
rect 7026 7588 7050 7590
rect 7106 7588 7130 7590
rect 7186 7588 7192 7590
rect 6884 7579 7192 7588
rect 7484 7546 7512 7822
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 6884 6556 7192 6565
rect 6884 6554 6890 6556
rect 6946 6554 6970 6556
rect 7026 6554 7050 6556
rect 7106 6554 7130 6556
rect 7186 6554 7192 6556
rect 6946 6502 6948 6554
rect 7128 6502 7130 6554
rect 6884 6500 6890 6502
rect 6946 6500 6970 6502
rect 7026 6500 7050 6502
rect 7106 6500 7130 6502
rect 7186 6500 7192 6502
rect 6884 6491 7192 6500
rect 8220 6225 8248 7142
rect 8206 6216 8262 6225
rect 8206 6151 8262 6160
rect 6884 5468 7192 5477
rect 6884 5466 6890 5468
rect 6946 5466 6970 5468
rect 7026 5466 7050 5468
rect 7106 5466 7130 5468
rect 7186 5466 7192 5468
rect 6946 5414 6948 5466
rect 7128 5414 7130 5466
rect 6884 5412 6890 5414
rect 6946 5412 6970 5414
rect 7026 5412 7050 5414
rect 7106 5412 7130 5414
rect 7186 5412 7192 5414
rect 6884 5403 7192 5412
rect 6884 4380 7192 4389
rect 6884 4378 6890 4380
rect 6946 4378 6970 4380
rect 7026 4378 7050 4380
rect 7106 4378 7130 4380
rect 7186 4378 7192 4380
rect 6946 4326 6948 4378
rect 7128 4326 7130 4378
rect 6884 4324 6890 4326
rect 6946 4324 6970 4326
rect 7026 4324 7050 4326
rect 7106 4324 7130 4326
rect 7186 4324 7192 4326
rect 6884 4315 7192 4324
rect 8312 4078 8340 8434
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8864 3738 8892 4082
rect 9508 4010 9536 8434
rect 9851 8188 10159 8197
rect 9851 8186 9857 8188
rect 9913 8186 9937 8188
rect 9993 8186 10017 8188
rect 10073 8186 10097 8188
rect 10153 8186 10159 8188
rect 9913 8134 9915 8186
rect 10095 8134 10097 8186
rect 9851 8132 9857 8134
rect 9913 8132 9937 8134
rect 9993 8132 10017 8134
rect 10073 8132 10097 8134
rect 10153 8132 10159 8134
rect 9851 8123 10159 8132
rect 11164 8090 11192 8434
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11072 7546 11100 7822
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 9851 7100 10159 7109
rect 9851 7098 9857 7100
rect 9913 7098 9937 7100
rect 9993 7098 10017 7100
rect 10073 7098 10097 7100
rect 10153 7098 10159 7100
rect 9913 7046 9915 7098
rect 10095 7046 10097 7098
rect 9851 7044 9857 7046
rect 9913 7044 9937 7046
rect 9993 7044 10017 7046
rect 10073 7044 10097 7046
rect 10153 7044 10159 7046
rect 9851 7035 10159 7044
rect 9851 6012 10159 6021
rect 9851 6010 9857 6012
rect 9913 6010 9937 6012
rect 9993 6010 10017 6012
rect 10073 6010 10097 6012
rect 10153 6010 10159 6012
rect 9913 5958 9915 6010
rect 10095 5958 10097 6010
rect 9851 5956 9857 5958
rect 9913 5956 9937 5958
rect 9993 5956 10017 5958
rect 10073 5956 10097 5958
rect 10153 5956 10159 5958
rect 9851 5947 10159 5956
rect 11808 5370 11836 8434
rect 13556 8090 13584 8434
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 12818 7644 13126 7653
rect 12818 7642 12824 7644
rect 12880 7642 12904 7644
rect 12960 7642 12984 7644
rect 13040 7642 13064 7644
rect 13120 7642 13126 7644
rect 12880 7590 12882 7642
rect 13062 7590 13064 7642
rect 12818 7588 12824 7590
rect 12880 7588 12904 7590
rect 12960 7588 12984 7590
rect 13040 7588 13064 7590
rect 13120 7588 13126 7590
rect 12818 7579 13126 7588
rect 12818 6556 13126 6565
rect 12818 6554 12824 6556
rect 12880 6554 12904 6556
rect 12960 6554 12984 6556
rect 13040 6554 13064 6556
rect 13120 6554 13126 6556
rect 12880 6502 12882 6554
rect 13062 6502 13064 6554
rect 12818 6500 12824 6502
rect 12880 6500 12904 6502
rect 12960 6500 12984 6502
rect 13040 6500 13064 6502
rect 13120 6500 13126 6502
rect 12818 6491 13126 6500
rect 14200 5914 14228 8434
rect 16500 8362 16528 9840
rect 17696 8616 17724 9840
rect 18892 9738 18920 9840
rect 18984 9738 19012 9846
rect 18892 9710 19012 9738
rect 18752 8732 19060 8741
rect 18752 8730 18758 8732
rect 18814 8730 18838 8732
rect 18894 8730 18918 8732
rect 18974 8730 18998 8732
rect 19054 8730 19060 8732
rect 18814 8678 18816 8730
rect 18996 8678 18998 8730
rect 18752 8676 18758 8678
rect 18814 8676 18838 8678
rect 18894 8676 18918 8678
rect 18974 8676 18998 8678
rect 19054 8676 19060 8678
rect 18752 8667 19060 8676
rect 19168 8634 19196 9846
rect 20074 9840 20130 10000
rect 21270 9840 21326 10000
rect 22466 9840 22522 10000
rect 23662 9840 23718 10000
rect 24504 9846 24808 9874
rect 20088 8634 20116 9840
rect 21284 8634 21312 9840
rect 22480 8634 22508 9840
rect 23676 8634 23704 9840
rect 17776 8628 17828 8634
rect 17696 8588 17776 8616
rect 17776 8570 17828 8576
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 15785 8188 16093 8197
rect 15785 8186 15791 8188
rect 15847 8186 15871 8188
rect 15927 8186 15951 8188
rect 16007 8186 16031 8188
rect 16087 8186 16093 8188
rect 15847 8134 15849 8186
rect 16029 8134 16031 8186
rect 15785 8132 15791 8134
rect 15847 8132 15871 8134
rect 15927 8132 15951 8134
rect 16007 8132 16031 8134
rect 16087 8132 16093 8134
rect 15785 8123 16093 8132
rect 17420 8090 17448 8434
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 15785 7100 16093 7109
rect 15785 7098 15791 7100
rect 15847 7098 15871 7100
rect 15927 7098 15951 7100
rect 16007 7098 16031 7100
rect 16087 7098 16093 7100
rect 15847 7046 15849 7098
rect 16029 7046 16031 7098
rect 15785 7044 15791 7046
rect 15847 7044 15871 7046
rect 15927 7044 15951 7046
rect 16007 7044 16031 7046
rect 16087 7044 16093 7046
rect 15785 7035 16093 7044
rect 15785 6012 16093 6021
rect 15785 6010 15791 6012
rect 15847 6010 15871 6012
rect 15927 6010 15951 6012
rect 16007 6010 16031 6012
rect 16087 6010 16093 6012
rect 15847 5958 15849 6010
rect 16029 5958 16031 6010
rect 15785 5956 15791 5958
rect 15847 5956 15871 5958
rect 15927 5956 15951 5958
rect 16007 5956 16031 5958
rect 16087 5956 16093 5958
rect 15785 5947 16093 5956
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 12818 5468 13126 5477
rect 12818 5466 12824 5468
rect 12880 5466 12904 5468
rect 12960 5466 12984 5468
rect 13040 5466 13064 5468
rect 13120 5466 13126 5468
rect 12880 5414 12882 5466
rect 13062 5414 13064 5466
rect 12818 5412 12824 5414
rect 12880 5412 12904 5414
rect 12960 5412 12984 5414
rect 13040 5412 13064 5414
rect 13120 5412 13126 5414
rect 12818 5403 13126 5412
rect 14660 5370 14688 5646
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 9851 4924 10159 4933
rect 9851 4922 9857 4924
rect 9913 4922 9937 4924
rect 9993 4922 10017 4924
rect 10073 4922 10097 4924
rect 10153 4922 10159 4924
rect 9913 4870 9915 4922
rect 10095 4870 10097 4922
rect 9851 4868 9857 4870
rect 9913 4868 9937 4870
rect 9993 4868 10017 4870
rect 10073 4868 10097 4870
rect 10153 4868 10159 4870
rect 9851 4859 10159 4868
rect 12360 4826 12388 5170
rect 15785 4924 16093 4933
rect 15785 4922 15791 4924
rect 15847 4922 15871 4924
rect 15927 4922 15951 4924
rect 16007 4922 16031 4924
rect 16087 4922 16093 4924
rect 15847 4870 15849 4922
rect 16029 4870 16031 4922
rect 15785 4868 15791 4870
rect 15847 4868 15871 4870
rect 15927 4868 15951 4870
rect 16007 4868 16031 4870
rect 16087 4868 16093 4870
rect 15785 4859 16093 4868
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12818 4380 13126 4389
rect 12818 4378 12824 4380
rect 12880 4378 12904 4380
rect 12960 4378 12984 4380
rect 13040 4378 13064 4380
rect 13120 4378 13126 4380
rect 12880 4326 12882 4378
rect 13062 4326 13064 4378
rect 12818 4324 12824 4326
rect 12880 4324 12904 4326
rect 12960 4324 12984 4326
rect 13040 4324 13064 4326
rect 13120 4324 13126 4326
rect 12818 4315 13126 4324
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9692 3738 9720 4082
rect 9851 3836 10159 3845
rect 9851 3834 9857 3836
rect 9913 3834 9937 3836
rect 9993 3834 10017 3836
rect 10073 3834 10097 3836
rect 10153 3834 10159 3836
rect 9913 3782 9915 3834
rect 10095 3782 10097 3834
rect 9851 3780 9857 3782
rect 9913 3780 9937 3782
rect 9993 3780 10017 3782
rect 10073 3780 10097 3782
rect 10153 3780 10159 3782
rect 9851 3771 10159 3780
rect 15785 3836 16093 3845
rect 15785 3834 15791 3836
rect 15847 3834 15871 3836
rect 15927 3834 15951 3836
rect 16007 3834 16031 3836
rect 16087 3834 16093 3836
rect 15847 3782 15849 3834
rect 16029 3782 16031 3834
rect 15785 3780 15791 3782
rect 15847 3780 15871 3782
rect 15927 3780 15951 3782
rect 16007 3780 16031 3782
rect 16087 3780 16093 3782
rect 15785 3771 16093 3780
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 13912 3528 13964 3534
rect 9494 3496 9550 3505
rect 13912 3470 13964 3476
rect 9494 3431 9496 3440
rect 9548 3431 9550 3440
rect 9496 3402 9548 3408
rect 6884 3292 7192 3301
rect 6884 3290 6890 3292
rect 6946 3290 6970 3292
rect 7026 3290 7050 3292
rect 7106 3290 7130 3292
rect 7186 3290 7192 3292
rect 6946 3238 6948 3290
rect 7128 3238 7130 3290
rect 6884 3236 6890 3238
rect 6946 3236 6970 3238
rect 7026 3236 7050 3238
rect 7106 3236 7130 3238
rect 7186 3236 7192 3238
rect 6884 3227 7192 3236
rect 12818 3292 13126 3301
rect 12818 3290 12824 3292
rect 12880 3290 12904 3292
rect 12960 3290 12984 3292
rect 13040 3290 13064 3292
rect 13120 3290 13126 3292
rect 12880 3238 12882 3290
rect 13062 3238 13064 3290
rect 12818 3236 12824 3238
rect 12880 3236 12904 3238
rect 12960 3236 12984 3238
rect 13040 3236 13064 3238
rect 13120 3236 13126 3238
rect 12818 3227 13126 3236
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 756 3120 808 3126
rect 756 3062 808 3068
rect 7378 3088 7434 3097
rect 204 3052 256 3058
rect 204 2994 256 3000
rect 216 160 244 2994
rect 480 2984 532 2990
rect 480 2926 532 2932
rect 492 160 520 2926
rect 768 160 796 3062
rect 2228 3052 2280 3058
rect 7378 3023 7434 3032
rect 2228 2994 2280 3000
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1492 2576 1544 2582
rect 1490 2544 1492 2553
rect 1544 2544 1546 2553
rect 1490 2479 1546 2488
rect 1596 2446 1624 2790
rect 1688 2650 1716 2790
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1032 1828 1084 1834
rect 1032 1770 1084 1776
rect 1044 160 1072 1770
rect 1320 160 1348 2382
rect 1492 2372 1544 2378
rect 1492 2314 1544 2320
rect 1504 1442 1532 2314
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 1688 2106 1716 2246
rect 1676 2100 1728 2106
rect 1676 2042 1728 2048
rect 1584 1964 1636 1970
rect 1636 1924 1900 1952
rect 1584 1906 1636 1912
rect 1504 1414 1624 1442
rect 1492 1352 1544 1358
rect 1492 1294 1544 1300
rect 1504 678 1532 1294
rect 1492 672 1544 678
rect 1492 614 1544 620
rect 1596 160 1624 1414
rect 1676 1216 1728 1222
rect 1676 1158 1728 1164
rect 1768 1216 1820 1222
rect 1768 1158 1820 1164
rect 1688 241 1716 1158
rect 1780 950 1808 1158
rect 1768 944 1820 950
rect 1768 886 1820 892
rect 1674 232 1730 241
rect 1674 167 1730 176
rect 1872 160 1900 1924
rect 2056 1766 2084 2586
rect 2240 2394 2268 2994
rect 3917 2748 4225 2757
rect 3917 2746 3923 2748
rect 3979 2746 4003 2748
rect 4059 2746 4083 2748
rect 4139 2746 4163 2748
rect 4219 2746 4225 2748
rect 3979 2694 3981 2746
rect 4161 2694 4163 2746
rect 3917 2692 3923 2694
rect 3979 2692 4003 2694
rect 4059 2692 4083 2694
rect 4139 2692 4163 2694
rect 4219 2692 4225 2694
rect 3917 2683 4225 2692
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 2148 2366 2268 2394
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 2044 1760 2096 1766
rect 2044 1702 2096 1708
rect 1952 1352 2004 1358
rect 1952 1294 2004 1300
rect 1964 746 1992 1294
rect 1952 740 2004 746
rect 1952 682 2004 688
rect 2148 160 2176 2366
rect 2228 2304 2280 2310
rect 2228 2246 2280 2252
rect 2240 2038 2268 2246
rect 2228 2032 2280 2038
rect 2228 1974 2280 1980
rect 2700 1970 2728 2382
rect 3160 2038 3188 2450
rect 4620 2440 4672 2446
rect 5172 2440 5224 2446
rect 4620 2382 4672 2388
rect 4908 2400 5172 2428
rect 4252 2100 4304 2106
rect 4252 2042 4304 2048
rect 3148 2032 3200 2038
rect 3148 1974 3200 1980
rect 2688 1964 2740 1970
rect 2688 1906 2740 1912
rect 2780 1964 2832 1970
rect 2780 1906 2832 1912
rect 3056 1964 3108 1970
rect 3056 1906 3108 1912
rect 3608 1964 3660 1970
rect 3884 1964 3936 1970
rect 3608 1906 3660 1912
rect 3804 1924 3884 1952
rect 2688 1760 2740 1766
rect 2688 1702 2740 1708
rect 2700 1562 2728 1702
rect 2688 1556 2740 1562
rect 2688 1498 2740 1504
rect 2320 1216 2372 1222
rect 2320 1158 2372 1164
rect 2596 1216 2648 1222
rect 2596 1158 2648 1164
rect 2332 610 2360 1158
rect 2412 672 2464 678
rect 2412 614 2464 620
rect 2320 604 2372 610
rect 2320 546 2372 552
rect 2424 160 2452 614
rect 2608 474 2636 1158
rect 2688 740 2740 746
rect 2688 682 2740 688
rect 2596 468 2648 474
rect 2596 410 2648 416
rect 2700 160 2728 682
rect 202 0 258 160
rect 478 0 534 160
rect 754 0 810 160
rect 1030 0 1086 160
rect 1306 0 1362 160
rect 1582 0 1638 160
rect 1858 0 1914 160
rect 2134 0 2190 160
rect 2410 0 2466 160
rect 2686 0 2742 160
rect 2792 82 2820 1906
rect 2964 1760 3016 1766
rect 2964 1702 3016 1708
rect 2976 1358 3004 1702
rect 2964 1352 3016 1358
rect 2964 1294 3016 1300
rect 2962 82 3018 160
rect 2792 54 3018 82
rect 3068 82 3096 1906
rect 3516 1828 3568 1834
rect 3516 1770 3568 1776
rect 3240 1760 3292 1766
rect 3240 1702 3292 1708
rect 3252 1358 3280 1702
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 3344 746 3372 1294
rect 3528 950 3556 1770
rect 3516 944 3568 950
rect 3516 886 3568 892
rect 3332 740 3384 746
rect 3332 682 3384 688
rect 3238 82 3294 160
rect 3068 54 3294 82
rect 2962 0 3018 54
rect 3238 0 3294 54
rect 3514 82 3570 160
rect 3620 82 3648 1906
rect 3804 160 3832 1924
rect 3884 1906 3936 1912
rect 3917 1660 4225 1669
rect 3917 1658 3923 1660
rect 3979 1658 4003 1660
rect 4059 1658 4083 1660
rect 4139 1658 4163 1660
rect 4219 1658 4225 1660
rect 3979 1606 3981 1658
rect 4161 1606 4163 1658
rect 3917 1604 3923 1606
rect 3979 1604 4003 1606
rect 4059 1604 4083 1606
rect 4139 1604 4163 1606
rect 4219 1604 4225 1606
rect 3917 1595 4225 1604
rect 4158 1456 4214 1465
rect 4158 1391 4214 1400
rect 4172 1222 4200 1391
rect 4160 1216 4212 1222
rect 4160 1158 4212 1164
rect 4068 740 4120 746
rect 4068 682 4120 688
rect 4080 160 4108 682
rect 4264 542 4292 2042
rect 4344 1964 4396 1970
rect 4344 1906 4396 1912
rect 4436 1964 4488 1970
rect 4436 1906 4488 1912
rect 4252 536 4304 542
rect 4252 478 4304 484
rect 4356 160 4384 1906
rect 4448 1562 4476 1906
rect 4436 1556 4488 1562
rect 4436 1498 4488 1504
rect 4528 1556 4580 1562
rect 4528 1498 4580 1504
rect 4540 1442 4568 1498
rect 4448 1414 4568 1442
rect 4448 1290 4476 1414
rect 4528 1352 4580 1358
rect 4528 1294 4580 1300
rect 4436 1284 4488 1290
rect 4436 1226 4488 1232
rect 4540 746 4568 1294
rect 4528 740 4580 746
rect 4528 682 4580 688
rect 4632 160 4660 2382
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4724 2106 4752 2246
rect 4712 2100 4764 2106
rect 4712 2042 4764 2048
rect 4712 1760 4764 1766
rect 4712 1702 4764 1708
rect 4724 678 4752 1702
rect 4816 1426 4844 2246
rect 4804 1420 4856 1426
rect 4804 1362 4856 1368
rect 4804 1216 4856 1222
rect 4804 1158 4856 1164
rect 4712 672 4764 678
rect 4712 614 4764 620
rect 4816 270 4844 1158
rect 4804 264 4856 270
rect 4804 206 4856 212
rect 4908 160 4936 2400
rect 5448 2440 5500 2446
rect 5172 2382 5224 2388
rect 5276 2400 5448 2428
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 5092 1358 5120 2246
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 5080 1352 5132 1358
rect 5080 1294 5132 1300
rect 5000 1018 5028 1294
rect 5276 1204 5304 2400
rect 5448 2382 5500 2388
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6550 2408 6606 2417
rect 5908 1964 5960 1970
rect 5908 1906 5960 1912
rect 5632 1828 5684 1834
rect 5632 1770 5684 1776
rect 5540 1760 5592 1766
rect 5540 1702 5592 1708
rect 5552 1358 5580 1702
rect 5540 1352 5592 1358
rect 5540 1294 5592 1300
rect 5184 1176 5304 1204
rect 5356 1216 5408 1222
rect 4988 1012 5040 1018
rect 4988 954 5040 960
rect 5184 160 5212 1176
rect 5356 1158 5408 1164
rect 5448 1216 5500 1222
rect 5448 1158 5500 1164
rect 5368 921 5396 1158
rect 5354 912 5410 921
rect 5460 882 5488 1158
rect 5540 1012 5592 1018
rect 5540 954 5592 960
rect 5354 847 5410 856
rect 5448 876 5500 882
rect 5448 818 5500 824
rect 5448 740 5500 746
rect 5448 682 5500 688
rect 5460 160 5488 682
rect 5552 490 5580 954
rect 5644 814 5672 1770
rect 5724 1352 5776 1358
rect 5724 1294 5776 1300
rect 5632 808 5684 814
rect 5632 750 5684 756
rect 5736 678 5764 1294
rect 5816 1216 5868 1222
rect 5816 1158 5868 1164
rect 5828 785 5856 1158
rect 5814 776 5870 785
rect 5814 711 5870 720
rect 5724 672 5776 678
rect 5724 614 5776 620
rect 5552 462 5764 490
rect 5736 160 5764 462
rect 3514 54 3648 82
rect 3514 0 3570 54
rect 3790 0 3846 160
rect 4066 0 4122 160
rect 4342 0 4398 160
rect 4618 0 4674 160
rect 4894 0 4950 160
rect 5170 0 5226 160
rect 5446 0 5502 160
rect 5722 0 5778 160
rect 5920 82 5948 1906
rect 6184 1352 6236 1358
rect 6184 1294 6236 1300
rect 6196 1018 6224 1294
rect 6184 1012 6236 1018
rect 6184 954 6236 960
rect 5998 82 6054 160
rect 5920 54 6054 82
rect 5998 0 6054 54
rect 6274 82 6330 160
rect 6380 82 6408 2382
rect 6550 2343 6606 2352
rect 6564 2310 6592 2343
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6460 1964 6512 1970
rect 6460 1906 6512 1912
rect 6274 54 6408 82
rect 6472 82 6500 1906
rect 6656 1873 6684 2042
rect 6642 1864 6698 1873
rect 6642 1799 6698 1808
rect 6748 1562 6776 2246
rect 6884 2204 7192 2213
rect 6884 2202 6890 2204
rect 6946 2202 6970 2204
rect 7026 2202 7050 2204
rect 7106 2202 7130 2204
rect 7186 2202 7192 2204
rect 6946 2150 6948 2202
rect 7128 2150 7130 2202
rect 6884 2148 6890 2150
rect 6946 2148 6970 2150
rect 7026 2148 7050 2150
rect 7106 2148 7130 2150
rect 7186 2148 7192 2150
rect 6884 2139 7192 2148
rect 7392 2106 7420 3023
rect 9404 2916 9456 2922
rect 9404 2858 9456 2864
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 8114 2272 8170 2281
rect 8114 2207 8170 2216
rect 8128 2106 8156 2207
rect 7380 2100 7432 2106
rect 7380 2042 7432 2048
rect 7932 2100 7984 2106
rect 7932 2042 7984 2048
rect 8116 2100 8168 2106
rect 8116 2042 8168 2048
rect 7288 2032 7340 2038
rect 6826 2000 6882 2009
rect 7288 1974 7340 1980
rect 6826 1935 6828 1944
rect 6880 1935 6882 1944
rect 6828 1906 6880 1912
rect 7012 1828 7064 1834
rect 7012 1770 7064 1776
rect 7024 1562 7052 1770
rect 6736 1556 6788 1562
rect 6736 1498 6788 1504
rect 7012 1556 7064 1562
rect 7012 1498 7064 1504
rect 6736 1352 6788 1358
rect 6920 1352 6972 1358
rect 6736 1294 6788 1300
rect 6918 1320 6920 1329
rect 6972 1320 6974 1329
rect 6552 1216 6604 1222
rect 6552 1158 6604 1164
rect 6644 1216 6696 1222
rect 6644 1158 6696 1164
rect 6564 649 6592 1158
rect 6656 814 6684 1158
rect 6644 808 6696 814
rect 6644 750 6696 756
rect 6748 746 6776 1294
rect 6918 1255 6974 1264
rect 6884 1116 7192 1125
rect 6884 1114 6890 1116
rect 6946 1114 6970 1116
rect 7026 1114 7050 1116
rect 7106 1114 7130 1116
rect 7186 1114 7192 1116
rect 6946 1062 6948 1114
rect 7128 1062 7130 1114
rect 6884 1060 6890 1062
rect 6946 1060 6970 1062
rect 7026 1060 7050 1062
rect 7106 1060 7130 1062
rect 7186 1060 7192 1062
rect 6884 1051 7192 1060
rect 6736 740 6788 746
rect 6736 682 6788 688
rect 6828 672 6880 678
rect 6550 640 6606 649
rect 6828 614 6880 620
rect 6550 575 6606 584
rect 6736 468 6788 474
rect 6736 410 6788 416
rect 6748 241 6776 410
rect 6734 232 6790 241
rect 6734 167 6790 176
rect 6840 160 6868 614
rect 6550 82 6606 160
rect 6472 54 6606 82
rect 6274 0 6330 54
rect 6550 0 6606 54
rect 6826 0 6882 160
rect 7102 82 7158 160
rect 7300 82 7328 1974
rect 7484 1970 7696 1986
rect 7472 1964 7696 1970
rect 7524 1958 7696 1964
rect 7472 1906 7524 1912
rect 7564 1896 7616 1902
rect 7564 1838 7616 1844
rect 7576 1562 7604 1838
rect 7564 1556 7616 1562
rect 7564 1498 7616 1504
rect 7472 1488 7524 1494
rect 7472 1430 7524 1436
rect 7380 1216 7432 1222
rect 7380 1158 7432 1164
rect 7392 1018 7420 1158
rect 7380 1012 7432 1018
rect 7380 954 7432 960
rect 7484 746 7512 1430
rect 7562 1184 7618 1193
rect 7562 1119 7618 1128
rect 7380 740 7432 746
rect 7380 682 7432 688
rect 7472 740 7524 746
rect 7472 682 7524 688
rect 7392 160 7420 682
rect 7576 377 7604 1119
rect 7562 368 7618 377
rect 7562 303 7618 312
rect 7668 160 7696 1958
rect 7840 1964 7892 1970
rect 7760 1924 7840 1952
rect 7760 1358 7788 1924
rect 7840 1906 7892 1912
rect 7840 1828 7892 1834
rect 7840 1770 7892 1776
rect 7852 1358 7880 1770
rect 7944 1562 7972 2042
rect 8864 1970 8892 2314
rect 8942 2136 8998 2145
rect 8942 2071 8944 2080
rect 8996 2071 8998 2080
rect 8944 2042 8996 2048
rect 8024 1964 8076 1970
rect 8300 1964 8352 1970
rect 8024 1906 8076 1912
rect 8220 1924 8300 1952
rect 7932 1556 7984 1562
rect 7932 1498 7984 1504
rect 8036 1494 8064 1906
rect 8024 1488 8076 1494
rect 8024 1430 8076 1436
rect 7748 1352 7800 1358
rect 7748 1294 7800 1300
rect 7840 1352 7892 1358
rect 7840 1294 7892 1300
rect 7930 1320 7986 1329
rect 7930 1255 7986 1264
rect 7748 1216 7800 1222
rect 7748 1158 7800 1164
rect 7840 1216 7892 1222
rect 7840 1158 7892 1164
rect 7760 474 7788 1158
rect 7748 468 7800 474
rect 7748 410 7800 416
rect 7852 338 7880 1158
rect 7840 332 7892 338
rect 7840 274 7892 280
rect 7944 160 7972 1255
rect 8024 1216 8076 1222
rect 8024 1158 8076 1164
rect 8036 950 8064 1158
rect 8024 944 8076 950
rect 8024 886 8076 892
rect 8220 160 8248 1924
rect 8300 1906 8352 1912
rect 8576 1964 8628 1970
rect 8852 1964 8904 1970
rect 8628 1924 8800 1952
rect 8576 1906 8628 1912
rect 8668 1760 8720 1766
rect 8668 1702 8720 1708
rect 8680 1358 8708 1702
rect 8668 1352 8720 1358
rect 8668 1294 8720 1300
rect 8300 1284 8352 1290
rect 8300 1226 8352 1232
rect 8312 728 8340 1226
rect 8312 700 8524 728
rect 8496 160 8524 700
rect 8772 160 8800 1924
rect 8852 1906 8904 1912
rect 9048 1737 9076 2586
rect 9324 2582 9352 2790
rect 9312 2576 9364 2582
rect 9312 2518 9364 2524
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9232 2394 9260 2450
rect 9232 2366 9352 2394
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9232 2106 9260 2246
rect 9220 2100 9272 2106
rect 9220 2042 9272 2048
rect 9128 1964 9180 1970
rect 9128 1906 9180 1912
rect 9034 1728 9090 1737
rect 9034 1663 9090 1672
rect 8852 1420 8904 1426
rect 8852 1362 8904 1368
rect 7102 54 7328 82
rect 7102 0 7158 54
rect 7378 0 7434 160
rect 7654 0 7710 160
rect 7930 0 7986 160
rect 8206 0 8262 160
rect 8482 0 8538 160
rect 8758 0 8814 160
rect 8864 82 8892 1362
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 9048 746 9076 1294
rect 9036 740 9088 746
rect 9036 682 9088 688
rect 8942 504 8998 513
rect 8942 439 8998 448
rect 8956 270 8984 439
rect 8944 264 8996 270
rect 8944 206 8996 212
rect 9034 82 9090 160
rect 8864 54 9090 82
rect 9140 82 9168 1906
rect 9324 1426 9352 2366
rect 9416 1970 9444 2858
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 9851 2748 10159 2757
rect 9851 2746 9857 2748
rect 9913 2746 9937 2748
rect 9993 2746 10017 2748
rect 10073 2746 10097 2748
rect 10153 2746 10159 2748
rect 9913 2694 9915 2746
rect 10095 2694 10097 2746
rect 9851 2692 9857 2694
rect 9913 2692 9937 2694
rect 9993 2692 10017 2694
rect 10073 2692 10097 2694
rect 10153 2692 10159 2694
rect 9851 2683 10159 2692
rect 9862 2544 9918 2553
rect 9508 2502 9862 2530
rect 9404 1964 9456 1970
rect 9404 1906 9456 1912
rect 9508 1850 9536 2502
rect 12438 2544 12494 2553
rect 9862 2479 9918 2488
rect 9956 2508 10008 2514
rect 12438 2479 12494 2488
rect 9956 2450 10008 2456
rect 9864 2440 9916 2446
rect 9416 1834 9536 1850
rect 9404 1828 9536 1834
rect 9456 1822 9536 1828
rect 9600 2400 9864 2428
rect 9404 1770 9456 1776
rect 9312 1420 9364 1426
rect 9312 1362 9364 1368
rect 9324 1278 9536 1306
rect 9324 1222 9352 1278
rect 9220 1216 9272 1222
rect 9220 1158 9272 1164
rect 9312 1216 9364 1222
rect 9312 1158 9364 1164
rect 9404 1216 9456 1222
rect 9404 1158 9456 1164
rect 9232 649 9260 1158
rect 9416 882 9444 1158
rect 9508 882 9536 1278
rect 9404 876 9456 882
rect 9404 818 9456 824
rect 9496 876 9548 882
rect 9496 818 9548 824
rect 9218 640 9274 649
rect 9218 575 9274 584
rect 9600 160 9628 2400
rect 9864 2382 9916 2388
rect 9680 2100 9732 2106
rect 9968 2088 9996 2450
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 10324 2372 10376 2378
rect 10324 2314 10376 2320
rect 9732 2060 9996 2088
rect 9680 2042 9732 2048
rect 10336 1970 10364 2314
rect 10980 2145 11008 2382
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 10966 2136 11022 2145
rect 11532 2106 11560 2246
rect 10966 2071 11022 2080
rect 11520 2100 11572 2106
rect 11520 2042 11572 2048
rect 9772 1964 9824 1970
rect 9772 1906 9824 1912
rect 9864 1964 9916 1970
rect 9864 1906 9916 1912
rect 10324 1964 10376 1970
rect 10324 1906 10376 1912
rect 9678 1728 9734 1737
rect 9678 1663 9734 1672
rect 9692 1358 9720 1663
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 9784 950 9812 1906
rect 9876 1766 9904 1906
rect 9864 1760 9916 1766
rect 9864 1702 9916 1708
rect 10508 1760 10560 1766
rect 11060 1760 11112 1766
rect 10508 1702 10560 1708
rect 10980 1720 11060 1748
rect 9851 1660 10159 1669
rect 9851 1658 9857 1660
rect 9913 1658 9937 1660
rect 9993 1658 10017 1660
rect 10073 1658 10097 1660
rect 10153 1658 10159 1660
rect 9913 1606 9915 1658
rect 10095 1606 10097 1658
rect 9851 1604 9857 1606
rect 9913 1604 9937 1606
rect 9993 1604 10017 1606
rect 10073 1604 10097 1606
rect 10153 1604 10159 1606
rect 9851 1595 10159 1604
rect 10048 1216 10100 1222
rect 10048 1158 10100 1164
rect 9772 944 9824 950
rect 9772 886 9824 892
rect 9680 740 9732 746
rect 9732 700 9904 728
rect 9680 682 9732 688
rect 9876 160 9904 700
rect 9310 82 9366 160
rect 9140 54 9366 82
rect 9034 0 9090 54
rect 9310 0 9366 54
rect 9586 0 9642 160
rect 9862 0 9918 160
rect 10060 82 10088 1158
rect 10138 82 10194 160
rect 10060 54 10194 82
rect 10138 0 10194 54
rect 10414 82 10470 160
rect 10520 82 10548 1702
rect 10692 1284 10744 1290
rect 10692 1226 10744 1232
rect 10784 1284 10836 1290
rect 10784 1226 10836 1232
rect 10704 160 10732 1226
rect 10796 1018 10824 1226
rect 10784 1012 10836 1018
rect 10784 954 10836 960
rect 10980 160 11008 1720
rect 11060 1702 11112 1708
rect 11060 1420 11112 1426
rect 11060 1362 11112 1368
rect 10414 54 10548 82
rect 10414 0 10470 54
rect 10690 0 10746 160
rect 10966 0 11022 160
rect 11072 82 11100 1362
rect 11716 1358 11744 2246
rect 11888 1828 11940 1834
rect 11888 1770 11940 1776
rect 11796 1760 11848 1766
rect 11796 1702 11848 1708
rect 11704 1352 11756 1358
rect 11704 1294 11756 1300
rect 11152 1216 11204 1222
rect 11520 1216 11572 1222
rect 11204 1176 11468 1204
rect 11152 1158 11204 1164
rect 11440 626 11468 1176
rect 11520 1158 11572 1164
rect 11612 1216 11664 1222
rect 11612 1158 11664 1164
rect 11532 1018 11560 1158
rect 11520 1012 11572 1018
rect 11520 954 11572 960
rect 11440 598 11560 626
rect 11532 160 11560 598
rect 11624 542 11652 1158
rect 11612 536 11664 542
rect 11612 478 11664 484
rect 11808 160 11836 1702
rect 11242 82 11298 160
rect 11072 54 11298 82
rect 11242 0 11298 54
rect 11518 0 11574 160
rect 11794 0 11850 160
rect 11900 82 11928 1770
rect 11992 542 12020 2382
rect 12346 2272 12402 2281
rect 12346 2207 12402 2216
rect 12256 2100 12308 2106
rect 12256 2042 12308 2048
rect 12072 1216 12124 1222
rect 12072 1158 12124 1164
rect 12084 610 12112 1158
rect 12268 950 12296 2042
rect 12360 1737 12388 2207
rect 12346 1728 12402 1737
rect 12346 1663 12402 1672
rect 12452 1601 12480 2479
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12438 1592 12494 1601
rect 12438 1527 12494 1536
rect 12440 1352 12492 1358
rect 12440 1294 12492 1300
rect 12348 1216 12400 1222
rect 12348 1158 12400 1164
rect 12256 944 12308 950
rect 12256 886 12308 892
rect 12072 604 12124 610
rect 12072 546 12124 552
rect 11980 536 12032 542
rect 11980 478 12032 484
rect 12360 160 12388 1158
rect 12452 678 12480 1294
rect 12544 1193 12572 2382
rect 12636 1970 12664 2790
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13280 2394 13308 2450
rect 13464 2446 13492 2858
rect 13188 2366 13308 2394
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 13728 2372 13780 2378
rect 12818 2204 13126 2213
rect 12818 2202 12824 2204
rect 12880 2202 12904 2204
rect 12960 2202 12984 2204
rect 13040 2202 13064 2204
rect 13120 2202 13126 2204
rect 12880 2150 12882 2202
rect 13062 2150 13064 2202
rect 12818 2148 12824 2150
rect 12880 2148 12904 2150
rect 12960 2148 12984 2150
rect 13040 2148 13064 2150
rect 13120 2148 13126 2150
rect 12818 2139 13126 2148
rect 13188 2106 13216 2366
rect 13728 2314 13780 2320
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 13280 2106 13308 2246
rect 13740 2106 13768 2314
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 13268 2100 13320 2106
rect 13268 2042 13320 2048
rect 13728 2100 13780 2106
rect 13728 2042 13780 2048
rect 13634 2000 13690 2009
rect 12624 1964 12676 1970
rect 12624 1906 12676 1912
rect 12808 1964 12860 1970
rect 13634 1935 13636 1944
rect 12808 1906 12860 1912
rect 13688 1935 13690 1944
rect 13636 1906 13688 1912
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 12530 1184 12586 1193
rect 12530 1119 12586 1128
rect 12440 672 12492 678
rect 12440 614 12492 620
rect 12636 160 12664 1702
rect 12820 1465 12848 1906
rect 13360 1896 13412 1902
rect 13360 1838 13412 1844
rect 13372 1562 13400 1838
rect 13360 1556 13412 1562
rect 13820 1556 13872 1562
rect 13360 1498 13412 1504
rect 13740 1516 13820 1544
rect 12806 1456 12862 1465
rect 12806 1391 12862 1400
rect 12900 1352 12952 1358
rect 12728 1312 12900 1340
rect 12728 241 12756 1312
rect 12900 1294 12952 1300
rect 13268 1352 13320 1358
rect 13268 1294 13320 1300
rect 13084 1216 13136 1222
rect 13136 1176 13216 1204
rect 13084 1158 13136 1164
rect 12818 1116 13126 1125
rect 12818 1114 12824 1116
rect 12880 1114 12904 1116
rect 12960 1114 12984 1116
rect 13040 1114 13064 1116
rect 13120 1114 13126 1116
rect 12880 1062 12882 1114
rect 13062 1062 13064 1114
rect 12818 1060 12824 1062
rect 12880 1060 12904 1062
rect 12960 1060 12984 1062
rect 13040 1060 13064 1062
rect 13120 1060 13126 1062
rect 12818 1051 13126 1060
rect 12900 672 12952 678
rect 12900 614 12952 620
rect 12714 232 12770 241
rect 12714 167 12770 176
rect 12912 160 12940 614
rect 13188 160 13216 1176
rect 13280 678 13308 1294
rect 13452 1216 13504 1222
rect 13452 1158 13504 1164
rect 13268 672 13320 678
rect 13268 614 13320 620
rect 13464 160 13492 1158
rect 13740 160 13768 1516
rect 13820 1498 13872 1504
rect 13924 678 13952 3470
rect 15785 2748 16093 2757
rect 15785 2746 15791 2748
rect 15847 2746 15871 2748
rect 15927 2746 15951 2748
rect 16007 2746 16031 2748
rect 16087 2746 16093 2748
rect 15847 2694 15849 2746
rect 16029 2694 16031 2746
rect 15785 2692 15791 2694
rect 15847 2692 15871 2694
rect 15927 2692 15951 2694
rect 16007 2692 16031 2694
rect 16087 2692 16093 2694
rect 15658 2680 15714 2689
rect 15785 2683 16093 2692
rect 17696 2650 17724 8434
rect 18752 7644 19060 7653
rect 18752 7642 18758 7644
rect 18814 7642 18838 7644
rect 18894 7642 18918 7644
rect 18974 7642 18998 7644
rect 19054 7642 19060 7644
rect 18814 7590 18816 7642
rect 18996 7590 18998 7642
rect 18752 7588 18758 7590
rect 18814 7588 18838 7590
rect 18894 7588 18918 7590
rect 18974 7588 18998 7590
rect 19054 7588 19060 7590
rect 18752 7579 19060 7588
rect 18752 6556 19060 6565
rect 18752 6554 18758 6556
rect 18814 6554 18838 6556
rect 18894 6554 18918 6556
rect 18974 6554 18998 6556
rect 19054 6554 19060 6556
rect 18814 6502 18816 6554
rect 18996 6502 18998 6554
rect 18752 6500 18758 6502
rect 18814 6500 18838 6502
rect 18894 6500 18918 6502
rect 18974 6500 18998 6502
rect 19054 6500 19060 6502
rect 18752 6491 19060 6500
rect 18752 5468 19060 5477
rect 18752 5466 18758 5468
rect 18814 5466 18838 5468
rect 18894 5466 18918 5468
rect 18974 5466 18998 5468
rect 19054 5466 19060 5468
rect 18814 5414 18816 5466
rect 18996 5414 18998 5466
rect 18752 5412 18758 5414
rect 18814 5412 18838 5414
rect 18894 5412 18918 5414
rect 18974 5412 18998 5414
rect 19054 5412 19060 5414
rect 18752 5403 19060 5412
rect 18752 4380 19060 4389
rect 18752 4378 18758 4380
rect 18814 4378 18838 4380
rect 18894 4378 18918 4380
rect 18974 4378 18998 4380
rect 19054 4378 19060 4380
rect 18814 4326 18816 4378
rect 18996 4326 18998 4378
rect 18752 4324 18758 4326
rect 18814 4324 18838 4326
rect 18894 4324 18918 4326
rect 18974 4324 18998 4326
rect 19054 4324 19060 4326
rect 18752 4315 19060 4324
rect 18752 3292 19060 3301
rect 18752 3290 18758 3292
rect 18814 3290 18838 3292
rect 18894 3290 18918 3292
rect 18974 3290 18998 3292
rect 19054 3290 19060 3292
rect 18814 3238 18816 3290
rect 18996 3238 18998 3290
rect 18752 3236 18758 3238
rect 18814 3236 18838 3238
rect 18894 3236 18918 3238
rect 18974 3236 18998 3238
rect 19054 3236 19060 3238
rect 18752 3227 19060 3236
rect 19168 2650 19196 8434
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 21719 8188 22027 8197
rect 21719 8186 21725 8188
rect 21781 8186 21805 8188
rect 21861 8186 21885 8188
rect 21941 8186 21965 8188
rect 22021 8186 22027 8188
rect 21781 8134 21783 8186
rect 21963 8134 21965 8186
rect 21719 8132 21725 8134
rect 21781 8132 21805 8134
rect 21861 8132 21885 8134
rect 21941 8132 21965 8134
rect 22021 8132 22027 8134
rect 21719 8123 22027 8132
rect 21719 7100 22027 7109
rect 21719 7098 21725 7100
rect 21781 7098 21805 7100
rect 21861 7098 21885 7100
rect 21941 7098 21965 7100
rect 22021 7098 22027 7100
rect 21781 7046 21783 7098
rect 21963 7046 21965 7098
rect 21719 7044 21725 7046
rect 21781 7044 21805 7046
rect 21861 7044 21885 7046
rect 21941 7044 21965 7046
rect 22021 7044 22027 7046
rect 21719 7035 22027 7044
rect 21719 6012 22027 6021
rect 21719 6010 21725 6012
rect 21781 6010 21805 6012
rect 21861 6010 21885 6012
rect 21941 6010 21965 6012
rect 22021 6010 22027 6012
rect 21781 5958 21783 6010
rect 21963 5958 21965 6010
rect 21719 5956 21725 5958
rect 21781 5956 21805 5958
rect 21861 5956 21885 5958
rect 21941 5956 21965 5958
rect 22021 5956 22027 5958
rect 21719 5947 22027 5956
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19444 5370 19472 5646
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 19628 4826 19656 5170
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20088 3194 20116 3470
rect 20732 3194 20760 5102
rect 21719 4924 22027 4933
rect 21719 4922 21725 4924
rect 21781 4922 21805 4924
rect 21861 4922 21885 4924
rect 21941 4922 21965 4924
rect 22021 4922 22027 4924
rect 21781 4870 21783 4922
rect 21963 4870 21965 4922
rect 21719 4868 21725 4870
rect 21781 4868 21805 4870
rect 21861 4868 21885 4870
rect 21941 4868 21965 4870
rect 22021 4868 22027 4870
rect 21719 4859 22027 4868
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 15658 2615 15714 2624
rect 17684 2644 17736 2650
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15120 1970 15148 2382
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 15212 2106 15240 2246
rect 15200 2100 15252 2106
rect 15200 2042 15252 2048
rect 14096 1964 14148 1970
rect 14096 1906 14148 1912
rect 15108 1964 15160 1970
rect 15108 1906 15160 1912
rect 14108 1850 14136 1906
rect 14016 1822 14136 1850
rect 15292 1896 15344 1902
rect 15292 1838 15344 1844
rect 14016 1766 14044 1822
rect 14004 1760 14056 1766
rect 14004 1702 14056 1708
rect 14096 1760 14148 1766
rect 14096 1702 14148 1708
rect 14280 1760 14332 1766
rect 14280 1702 14332 1708
rect 14740 1760 14792 1766
rect 14740 1702 14792 1708
rect 15200 1760 15252 1766
rect 15304 1737 15332 1838
rect 15200 1702 15252 1708
rect 15290 1728 15346 1737
rect 14108 1494 14136 1702
rect 14096 1488 14148 1494
rect 14096 1430 14148 1436
rect 14188 1284 14240 1290
rect 14188 1226 14240 1232
rect 14004 1216 14056 1222
rect 14004 1158 14056 1164
rect 13912 672 13964 678
rect 13912 614 13964 620
rect 14016 160 14044 1158
rect 14200 814 14228 1226
rect 14188 808 14240 814
rect 14188 750 14240 756
rect 14292 160 14320 1702
rect 12070 82 12126 160
rect 11900 54 12126 82
rect 12070 0 12126 54
rect 12346 0 12402 160
rect 12622 0 12678 160
rect 12898 0 12954 160
rect 13174 0 13230 160
rect 13450 0 13506 160
rect 13726 0 13782 160
rect 14002 0 14058 160
rect 14278 0 14334 160
rect 14554 82 14610 160
rect 14752 82 14780 1702
rect 15108 1556 15160 1562
rect 14844 1516 15108 1544
rect 14844 160 14872 1516
rect 15108 1498 15160 1504
rect 15108 1420 15160 1426
rect 15108 1362 15160 1368
rect 15120 160 15148 1362
rect 15212 1358 15240 1702
rect 15290 1663 15346 1672
rect 15200 1352 15252 1358
rect 15200 1294 15252 1300
rect 15396 160 15424 2246
rect 15488 270 15516 2450
rect 15672 1970 15700 2615
rect 17684 2586 17736 2592
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 19340 2576 19392 2582
rect 19340 2518 19392 2524
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16580 2304 16632 2310
rect 16580 2246 16632 2252
rect 15660 1964 15712 1970
rect 15660 1906 15712 1912
rect 16212 1964 16264 1970
rect 16212 1906 16264 1912
rect 15660 1760 15712 1766
rect 15660 1702 15712 1708
rect 15476 264 15528 270
rect 15476 206 15528 212
rect 15672 160 15700 1702
rect 15785 1660 16093 1669
rect 15785 1658 15791 1660
rect 15847 1658 15871 1660
rect 15927 1658 15951 1660
rect 16007 1658 16031 1660
rect 16087 1658 16093 1660
rect 15847 1606 15849 1658
rect 16029 1606 16031 1658
rect 15785 1604 15791 1606
rect 15847 1604 15871 1606
rect 15927 1604 15951 1606
rect 16007 1604 16031 1606
rect 16087 1604 16093 1606
rect 15785 1595 16093 1604
rect 16120 1556 16172 1562
rect 15948 1516 16120 1544
rect 15948 160 15976 1516
rect 16120 1498 16172 1504
rect 16120 1420 16172 1426
rect 16120 1362 16172 1368
rect 14554 54 14780 82
rect 14554 0 14610 54
rect 14830 0 14886 160
rect 15106 0 15162 160
rect 15382 0 15438 160
rect 15658 0 15714 160
rect 15934 0 15990 160
rect 16132 82 16160 1362
rect 16224 649 16252 1906
rect 16500 1834 16528 2246
rect 16592 2106 16620 2246
rect 16684 2106 16712 2382
rect 16580 2100 16632 2106
rect 16580 2042 16632 2048
rect 16672 2100 16724 2106
rect 16672 2042 16724 2048
rect 16488 1828 16540 1834
rect 16488 1770 16540 1776
rect 16580 1760 16632 1766
rect 16580 1702 16632 1708
rect 16764 1760 16816 1766
rect 16764 1702 16816 1708
rect 16302 1456 16358 1465
rect 16302 1391 16358 1400
rect 16316 1358 16344 1391
rect 16592 1358 16620 1702
rect 16304 1352 16356 1358
rect 16304 1294 16356 1300
rect 16580 1352 16632 1358
rect 16580 1294 16632 1300
rect 16396 1216 16448 1222
rect 16396 1158 16448 1164
rect 16210 640 16266 649
rect 16210 575 16266 584
rect 16408 218 16436 1158
rect 16408 190 16528 218
rect 16500 160 16528 190
rect 16776 160 16804 1702
rect 16868 746 16896 2382
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 16948 1896 17000 1902
rect 16948 1838 17000 1844
rect 16960 1290 16988 1838
rect 17040 1420 17092 1426
rect 17040 1362 17092 1368
rect 16948 1284 17000 1290
rect 16948 1226 17000 1232
rect 16856 740 16908 746
rect 16856 682 16908 688
rect 17052 160 17080 1362
rect 17144 377 17172 2246
rect 17236 1290 17264 2518
rect 18420 2440 18472 2446
rect 18340 2400 18420 2428
rect 18144 2304 18196 2310
rect 18144 2246 18196 2252
rect 18156 2106 18184 2246
rect 18144 2100 18196 2106
rect 18144 2042 18196 2048
rect 17880 1822 18000 1850
rect 17592 1488 17644 1494
rect 17328 1436 17592 1442
rect 17328 1430 17644 1436
rect 17328 1414 17632 1430
rect 17224 1284 17276 1290
rect 17224 1226 17276 1232
rect 17130 368 17186 377
rect 17130 303 17186 312
rect 17328 160 17356 1414
rect 17776 1352 17828 1358
rect 17604 1312 17776 1340
rect 17604 160 17632 1312
rect 17776 1294 17828 1300
rect 17880 160 17908 1822
rect 17972 1766 18000 1822
rect 17960 1760 18012 1766
rect 17960 1702 18012 1708
rect 18236 1760 18288 1766
rect 18236 1702 18288 1708
rect 17958 1320 18014 1329
rect 17958 1255 18014 1264
rect 18052 1284 18104 1290
rect 17972 785 18000 1255
rect 18052 1226 18104 1232
rect 18064 1018 18092 1226
rect 18052 1012 18104 1018
rect 18052 954 18104 960
rect 18248 898 18276 1702
rect 18340 1018 18368 2400
rect 18420 2382 18472 2388
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 18432 2106 18460 2246
rect 18420 2100 18472 2106
rect 18420 2042 18472 2048
rect 18524 1222 18552 2246
rect 18752 2204 19060 2213
rect 18752 2202 18758 2204
rect 18814 2202 18838 2204
rect 18894 2202 18918 2204
rect 18974 2202 18998 2204
rect 19054 2202 19060 2204
rect 18814 2150 18816 2202
rect 18996 2150 18998 2202
rect 18752 2148 18758 2150
rect 18814 2148 18838 2150
rect 18894 2148 18918 2150
rect 18974 2148 18998 2150
rect 19054 2148 19060 2150
rect 18752 2139 19060 2148
rect 18972 1896 19024 1902
rect 18972 1838 19024 1844
rect 18984 1737 19012 1838
rect 18970 1728 19026 1737
rect 18970 1663 19026 1672
rect 19168 1562 19196 2382
rect 19352 1952 19380 2518
rect 19444 2446 19472 2790
rect 20088 2650 20116 2994
rect 20444 2916 20496 2922
rect 20444 2858 20496 2864
rect 20456 2774 20484 2858
rect 20272 2746 20484 2774
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 19616 2576 19668 2582
rect 19616 2518 19668 2524
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19524 2304 19576 2310
rect 19524 2246 19576 2252
rect 19536 2106 19564 2246
rect 19524 2100 19576 2106
rect 19524 2042 19576 2048
rect 19352 1924 19472 1952
rect 19340 1828 19392 1834
rect 19260 1788 19340 1816
rect 19156 1556 19208 1562
rect 19156 1498 19208 1504
rect 18696 1488 18748 1494
rect 18696 1430 18748 1436
rect 18604 1352 18656 1358
rect 18602 1320 18604 1329
rect 18656 1320 18658 1329
rect 18602 1255 18658 1264
rect 18512 1216 18564 1222
rect 18708 1204 18736 1430
rect 18512 1158 18564 1164
rect 18616 1176 18736 1204
rect 18328 1012 18380 1018
rect 18328 954 18380 960
rect 18512 1012 18564 1018
rect 18512 954 18564 960
rect 18156 870 18276 898
rect 17958 776 18014 785
rect 17958 711 18014 720
rect 18156 160 18184 870
rect 16210 82 16266 160
rect 16132 54 16266 82
rect 16210 0 16266 54
rect 16486 0 16542 160
rect 16762 0 16818 160
rect 17038 0 17094 160
rect 17314 0 17370 160
rect 17590 0 17646 160
rect 17866 0 17922 160
rect 18142 0 18198 160
rect 18418 82 18474 160
rect 18524 82 18552 954
rect 18418 54 18552 82
rect 18616 82 18644 1176
rect 18752 1116 19060 1125
rect 18752 1114 18758 1116
rect 18814 1114 18838 1116
rect 18894 1114 18918 1116
rect 18974 1114 18998 1116
rect 19054 1114 19060 1116
rect 18814 1062 18816 1114
rect 18996 1062 18998 1114
rect 18752 1060 18758 1062
rect 18814 1060 18838 1062
rect 18894 1060 18918 1062
rect 18974 1060 18998 1062
rect 19054 1060 19060 1062
rect 18752 1051 19060 1060
rect 19260 626 19288 1788
rect 19340 1770 19392 1776
rect 19338 1728 19394 1737
rect 19338 1663 19394 1672
rect 19352 1290 19380 1663
rect 19444 1290 19472 1924
rect 19340 1284 19392 1290
rect 19340 1226 19392 1232
rect 19432 1284 19484 1290
rect 19432 1226 19484 1232
rect 19628 1170 19656 2518
rect 19892 2440 19944 2446
rect 19892 2382 19944 2388
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19800 2100 19852 2106
rect 19800 2042 19852 2048
rect 19708 1760 19760 1766
rect 19708 1702 19760 1708
rect 19076 598 19288 626
rect 19536 1142 19656 1170
rect 18694 82 18750 160
rect 18616 54 18750 82
rect 18418 0 18474 54
rect 18694 0 18750 54
rect 18970 82 19026 160
rect 19076 82 19104 598
rect 19248 536 19300 542
rect 19248 478 19300 484
rect 19260 160 19288 478
rect 19536 160 19564 1142
rect 19720 1018 19748 1702
rect 19708 1012 19760 1018
rect 19708 954 19760 960
rect 19812 160 19840 2042
rect 19904 1766 19932 2382
rect 19996 1873 20024 2382
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 20088 1970 20116 2246
rect 20076 1964 20128 1970
rect 20076 1906 20128 1912
rect 19982 1864 20038 1873
rect 19982 1799 20038 1808
rect 19892 1760 19944 1766
rect 19892 1702 19944 1708
rect 18970 54 19104 82
rect 18970 0 19026 54
rect 19246 0 19302 160
rect 19522 0 19578 160
rect 19798 0 19854 160
rect 20074 82 20130 160
rect 20272 82 20300 2746
rect 20626 2544 20682 2553
rect 20626 2479 20628 2488
rect 20680 2479 20682 2488
rect 20628 2450 20680 2456
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 20628 1896 20680 1902
rect 20628 1838 20680 1844
rect 20444 1828 20496 1834
rect 20444 1770 20496 1776
rect 20456 542 20484 1770
rect 20640 1170 20668 1838
rect 20732 1562 20760 2382
rect 20720 1556 20772 1562
rect 20720 1498 20772 1504
rect 21008 1290 21036 4558
rect 21719 3836 22027 3845
rect 21719 3834 21725 3836
rect 21781 3834 21805 3836
rect 21861 3834 21885 3836
rect 21941 3834 21965 3836
rect 22021 3834 22027 3836
rect 21781 3782 21783 3834
rect 21963 3782 21965 3834
rect 21719 3780 21725 3782
rect 21781 3780 21805 3782
rect 21861 3780 21885 3782
rect 21941 3780 21965 3782
rect 22021 3780 22027 3782
rect 21719 3771 22027 3780
rect 21088 3052 21140 3058
rect 21088 2994 21140 3000
rect 21100 2650 21128 2994
rect 21719 2748 22027 2757
rect 21719 2746 21725 2748
rect 21781 2746 21805 2748
rect 21861 2746 21885 2748
rect 21941 2746 21965 2748
rect 22021 2746 22027 2748
rect 21781 2694 21783 2746
rect 21963 2694 21965 2746
rect 21719 2692 21725 2694
rect 21781 2692 21805 2694
rect 21861 2692 21885 2694
rect 21941 2692 21965 2694
rect 22021 2692 22027 2694
rect 21719 2683 22027 2692
rect 22112 2650 22140 8366
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22204 2650 22232 7686
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 22284 2916 22336 2922
rect 22284 2858 22336 2864
rect 21088 2644 21140 2650
rect 21088 2586 21140 2592
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 21640 2508 21692 2514
rect 21640 2450 21692 2456
rect 22020 2502 22232 2530
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 21192 1834 21220 2382
rect 21456 2304 21508 2310
rect 21456 2246 21508 2252
rect 21468 2106 21496 2246
rect 21456 2100 21508 2106
rect 21456 2042 21508 2048
rect 21548 2032 21600 2038
rect 21548 1974 21600 1980
rect 21560 1850 21588 1974
rect 21180 1828 21232 1834
rect 21180 1770 21232 1776
rect 21468 1822 21588 1850
rect 21468 1306 21496 1822
rect 21548 1760 21600 1766
rect 21548 1702 21600 1708
rect 20996 1284 21048 1290
rect 20996 1226 21048 1232
rect 21376 1278 21496 1306
rect 20812 1216 20864 1222
rect 20640 1142 20760 1170
rect 20812 1158 20864 1164
rect 20628 1012 20680 1018
rect 20628 954 20680 960
rect 20444 536 20496 542
rect 20444 478 20496 484
rect 20640 218 20668 954
rect 20548 190 20668 218
rect 20074 54 20300 82
rect 20350 82 20406 160
rect 20548 82 20576 190
rect 20350 54 20576 82
rect 20626 82 20682 160
rect 20732 82 20760 1142
rect 20824 649 20852 1158
rect 21088 740 21140 746
rect 21088 682 21140 688
rect 20810 640 20866 649
rect 20810 575 20866 584
rect 20626 54 20760 82
rect 20902 82 20958 160
rect 21100 82 21128 682
rect 21376 513 21404 1278
rect 21456 1216 21508 1222
rect 21456 1158 21508 1164
rect 21468 950 21496 1158
rect 21456 944 21508 950
rect 21456 886 21508 892
rect 21362 504 21418 513
rect 21180 468 21232 474
rect 21362 439 21418 448
rect 21180 410 21232 416
rect 21192 160 21220 410
rect 20902 54 21128 82
rect 20074 0 20130 54
rect 20350 0 20406 54
rect 20626 0 20682 54
rect 20902 0 20958 54
rect 21178 0 21234 160
rect 21454 82 21510 160
rect 21560 82 21588 1702
rect 21652 1562 21680 2450
rect 21824 2440 21876 2446
rect 21730 2408 21786 2417
rect 21824 2382 21876 2388
rect 21730 2343 21786 2352
rect 21744 1970 21772 2343
rect 21836 2106 21864 2382
rect 22020 2378 22048 2502
rect 22008 2372 22060 2378
rect 22008 2314 22060 2320
rect 21824 2100 21876 2106
rect 21824 2042 21876 2048
rect 21732 1964 21784 1970
rect 21732 1906 21784 1912
rect 21719 1660 22027 1669
rect 21719 1658 21725 1660
rect 21781 1658 21805 1660
rect 21861 1658 21885 1660
rect 21941 1658 21965 1660
rect 22021 1658 22027 1660
rect 21781 1606 21783 1658
rect 21963 1606 21965 1658
rect 21719 1604 21725 1606
rect 21781 1604 21805 1606
rect 21861 1604 21885 1606
rect 21941 1604 21965 1606
rect 22021 1604 22027 1606
rect 21719 1595 22027 1604
rect 22204 1562 22232 2502
rect 22296 1970 22324 2858
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 22388 2106 22416 2382
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 22480 2038 22508 5510
rect 22572 2650 22600 8434
rect 23124 8090 23152 8434
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 22664 2496 22692 3470
rect 22836 3460 22888 3466
rect 22836 3402 22888 3408
rect 22848 2774 22876 3402
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 22572 2468 22692 2496
rect 22756 2746 22876 2774
rect 22468 2032 22520 2038
rect 22468 1974 22520 1980
rect 22284 1964 22336 1970
rect 22284 1906 22336 1912
rect 21640 1556 21692 1562
rect 21640 1498 21692 1504
rect 22192 1556 22244 1562
rect 22192 1498 22244 1504
rect 22008 1488 22060 1494
rect 22572 1442 22600 2468
rect 22756 2394 22784 2746
rect 22836 2576 22888 2582
rect 22834 2544 22836 2553
rect 22888 2544 22890 2553
rect 22834 2479 22890 2488
rect 22008 1430 22060 1436
rect 21640 808 21692 814
rect 22020 762 22048 1430
rect 22388 1414 22600 1442
rect 22664 2366 22784 2394
rect 22836 2440 22888 2446
rect 22836 2382 22888 2388
rect 22284 1352 22336 1358
rect 22284 1294 22336 1300
rect 22296 921 22324 1294
rect 22282 912 22338 921
rect 22282 847 22338 856
rect 22388 796 22416 1414
rect 22560 1352 22612 1358
rect 22560 1294 22612 1300
rect 22572 1018 22600 1294
rect 22560 1012 22612 1018
rect 22560 954 22612 960
rect 22664 898 22692 2366
rect 22744 2304 22796 2310
rect 22744 2246 22796 2252
rect 22756 2106 22784 2246
rect 22744 2100 22796 2106
rect 22744 2042 22796 2048
rect 22744 1352 22796 1358
rect 22744 1294 22796 1300
rect 21640 750 21692 756
rect 21652 474 21680 750
rect 21928 734 22048 762
rect 22296 768 22416 796
rect 22572 870 22692 898
rect 21640 468 21692 474
rect 21640 410 21692 416
rect 21454 54 21588 82
rect 21730 82 21786 160
rect 21928 82 21956 734
rect 22008 672 22060 678
rect 22008 614 22060 620
rect 22020 160 22048 614
rect 22296 160 22324 768
rect 22572 160 22600 870
rect 22756 746 22784 1294
rect 22744 740 22796 746
rect 22744 682 22796 688
rect 22848 160 22876 2382
rect 21730 54 21956 82
rect 21454 0 21510 54
rect 21730 0 21786 54
rect 22006 0 22062 160
rect 22282 0 22338 160
rect 22558 0 22614 160
rect 22834 0 22890 160
rect 22940 82 22968 2994
rect 23032 2938 23060 7346
rect 23112 3596 23164 3602
rect 23112 3538 23164 3544
rect 23124 3058 23152 3538
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23032 2910 23152 2938
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 23032 1970 23060 2790
rect 23020 1964 23072 1970
rect 23020 1906 23072 1912
rect 23124 1834 23152 2910
rect 23216 2854 23244 7346
rect 23400 3738 23428 7482
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 23480 3664 23532 3670
rect 23480 3606 23532 3612
rect 23296 3120 23348 3126
rect 23296 3062 23348 3068
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 23308 2650 23336 3062
rect 23492 3058 23520 3606
rect 23480 3052 23532 3058
rect 23480 2994 23532 3000
rect 23584 2938 23612 8434
rect 23676 8090 23704 8434
rect 24504 8090 24532 9846
rect 24780 9738 24808 9846
rect 24858 9840 24914 10000
rect 24872 9738 24900 9840
rect 24780 9710 24900 9738
rect 24686 8732 24994 8741
rect 24686 8730 24692 8732
rect 24748 8730 24772 8732
rect 24828 8730 24852 8732
rect 24908 8730 24932 8732
rect 24988 8730 24994 8732
rect 24748 8678 24750 8730
rect 24930 8678 24932 8730
rect 24686 8676 24692 8678
rect 24748 8676 24772 8678
rect 24828 8676 24852 8678
rect 24908 8676 24932 8678
rect 24988 8676 24994 8678
rect 24686 8667 24994 8676
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 24492 8084 24544 8090
rect 24492 8026 24544 8032
rect 23848 7948 23900 7954
rect 23848 7890 23900 7896
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23676 7546 23704 7822
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23664 4548 23716 4554
rect 23664 4490 23716 4496
rect 23676 3738 23704 4490
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 23400 2910 23612 2938
rect 23296 2644 23348 2650
rect 23296 2586 23348 2592
rect 23400 2514 23428 2910
rect 23478 2816 23534 2825
rect 23478 2751 23534 2760
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23216 2106 23244 2382
rect 23204 2100 23256 2106
rect 23204 2042 23256 2048
rect 23112 1828 23164 1834
rect 23112 1770 23164 1776
rect 23492 1442 23520 2751
rect 23676 2496 23704 2994
rect 23768 2825 23796 3334
rect 23754 2816 23810 2825
rect 23754 2751 23810 2760
rect 23860 2774 23888 7890
rect 23940 7812 23992 7818
rect 23940 7754 23992 7760
rect 23952 2922 23980 7754
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 24308 4140 24360 4146
rect 24308 4082 24360 4088
rect 24124 3936 24176 3942
rect 24124 3878 24176 3884
rect 23940 2916 23992 2922
rect 23940 2858 23992 2864
rect 24032 2916 24084 2922
rect 24032 2858 24084 2864
rect 23860 2746 23980 2774
rect 23952 2650 23980 2746
rect 23940 2644 23992 2650
rect 23940 2586 23992 2592
rect 23940 2508 23992 2514
rect 23676 2468 23888 2496
rect 23572 2440 23624 2446
rect 23624 2400 23704 2428
rect 23572 2382 23624 2388
rect 23400 1414 23520 1442
rect 23400 1358 23428 1414
rect 23020 1352 23072 1358
rect 23020 1294 23072 1300
rect 23388 1352 23440 1358
rect 23388 1294 23440 1300
rect 23032 882 23060 1294
rect 23112 1216 23164 1222
rect 23110 1184 23112 1193
rect 23480 1216 23532 1222
rect 23164 1184 23166 1193
rect 23480 1158 23532 1164
rect 23110 1119 23166 1128
rect 23492 1057 23520 1158
rect 23478 1048 23534 1057
rect 23478 983 23534 992
rect 23020 876 23072 882
rect 23020 818 23072 824
rect 23480 808 23532 814
rect 23400 768 23480 796
rect 23400 160 23428 768
rect 23480 750 23532 756
rect 23676 160 23704 2400
rect 23756 2372 23808 2378
rect 23756 2314 23808 2320
rect 23768 1494 23796 2314
rect 23756 1488 23808 1494
rect 23756 1430 23808 1436
rect 23756 1352 23808 1358
rect 23756 1294 23808 1300
rect 23768 678 23796 1294
rect 23860 898 23888 2468
rect 23940 2450 23992 2456
rect 23952 1358 23980 2450
rect 24044 2106 24072 2858
rect 24032 2100 24084 2106
rect 24032 2042 24084 2048
rect 24136 1952 24164 3878
rect 24320 3738 24348 4082
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24228 2530 24256 3130
rect 24412 2650 24440 7686
rect 24686 7644 24994 7653
rect 24686 7642 24692 7644
rect 24748 7642 24772 7644
rect 24828 7642 24852 7644
rect 24908 7642 24932 7644
rect 24988 7642 24994 7644
rect 24748 7590 24750 7642
rect 24930 7590 24932 7642
rect 24686 7588 24692 7590
rect 24748 7588 24772 7590
rect 24828 7588 24852 7590
rect 24908 7588 24932 7590
rect 24988 7588 24994 7590
rect 24686 7579 24994 7588
rect 24686 6556 24994 6565
rect 24686 6554 24692 6556
rect 24748 6554 24772 6556
rect 24828 6554 24852 6556
rect 24908 6554 24932 6556
rect 24988 6554 24994 6556
rect 24748 6502 24750 6554
rect 24930 6502 24932 6554
rect 24686 6500 24692 6502
rect 24748 6500 24772 6502
rect 24828 6500 24852 6502
rect 24908 6500 24932 6502
rect 24988 6500 24994 6502
rect 24686 6491 24994 6500
rect 24686 5468 24994 5477
rect 24686 5466 24692 5468
rect 24748 5466 24772 5468
rect 24828 5466 24852 5468
rect 24908 5466 24932 5468
rect 24988 5466 24994 5468
rect 24748 5414 24750 5466
rect 24930 5414 24932 5466
rect 24686 5412 24692 5414
rect 24748 5412 24772 5414
rect 24828 5412 24852 5414
rect 24908 5412 24932 5414
rect 24988 5412 24994 5414
rect 24686 5403 24994 5412
rect 24686 4380 24994 4389
rect 24686 4378 24692 4380
rect 24748 4378 24772 4380
rect 24828 4378 24852 4380
rect 24908 4378 24932 4380
rect 24988 4378 24994 4380
rect 24748 4326 24750 4378
rect 24930 4326 24932 4378
rect 24686 4324 24692 4326
rect 24748 4324 24772 4326
rect 24828 4324 24852 4326
rect 24908 4324 24932 4326
rect 24988 4324 24994 4326
rect 24686 4315 24994 4324
rect 25320 3664 25372 3670
rect 25320 3606 25372 3612
rect 24584 3596 24636 3602
rect 24584 3538 24636 3544
rect 24492 3528 24544 3534
rect 24492 3470 24544 3476
rect 24400 2644 24452 2650
rect 24400 2586 24452 2592
rect 24228 2502 24440 2530
rect 24308 2440 24360 2446
rect 24308 2382 24360 2388
rect 24320 2106 24348 2382
rect 24308 2100 24360 2106
rect 24308 2042 24360 2048
rect 24412 1970 24440 2502
rect 24216 1964 24268 1970
rect 24136 1924 24216 1952
rect 24216 1906 24268 1912
rect 24400 1964 24452 1970
rect 24400 1906 24452 1912
rect 24032 1488 24084 1494
rect 24084 1448 24164 1476
rect 24032 1430 24084 1436
rect 23940 1352 23992 1358
rect 23940 1294 23992 1300
rect 23940 1216 23992 1222
rect 23940 1158 23992 1164
rect 23952 1018 23980 1158
rect 23940 1012 23992 1018
rect 23940 954 23992 960
rect 23860 870 23980 898
rect 23756 672 23808 678
rect 23756 614 23808 620
rect 23952 160 23980 870
rect 24136 660 24164 1448
rect 24216 1352 24268 1358
rect 24216 1294 24268 1300
rect 24228 814 24256 1294
rect 24216 808 24268 814
rect 24216 750 24268 756
rect 24136 632 24256 660
rect 24228 160 24256 632
rect 24504 160 24532 3470
rect 23110 82 23166 160
rect 22940 54 23166 82
rect 23110 0 23166 54
rect 23386 0 23442 160
rect 23662 0 23718 160
rect 23938 0 23994 160
rect 24214 0 24270 160
rect 24490 0 24546 160
rect 24596 82 24624 3538
rect 24686 3292 24994 3301
rect 24686 3290 24692 3292
rect 24748 3290 24772 3292
rect 24828 3290 24852 3292
rect 24908 3290 24932 3292
rect 24988 3290 24994 3292
rect 24748 3238 24750 3290
rect 24930 3238 24932 3290
rect 24686 3236 24692 3238
rect 24748 3236 24772 3238
rect 24828 3236 24852 3238
rect 24908 3236 24932 3238
rect 24988 3236 24994 3238
rect 24686 3227 24994 3236
rect 25044 2304 25096 2310
rect 25044 2246 25096 2252
rect 24686 2204 24994 2213
rect 24686 2202 24692 2204
rect 24748 2202 24772 2204
rect 24828 2202 24852 2204
rect 24908 2202 24932 2204
rect 24988 2202 24994 2204
rect 24748 2150 24750 2202
rect 24930 2150 24932 2202
rect 24686 2148 24692 2150
rect 24748 2148 24772 2150
rect 24828 2148 24852 2150
rect 24908 2148 24932 2150
rect 24988 2148 24994 2150
rect 24686 2139 24994 2148
rect 24686 1116 24994 1125
rect 24686 1114 24692 1116
rect 24748 1114 24772 1116
rect 24828 1114 24852 1116
rect 24908 1114 24932 1116
rect 24988 1114 24994 1116
rect 24748 1062 24750 1114
rect 24930 1062 24932 1114
rect 24686 1060 24692 1062
rect 24748 1060 24772 1062
rect 24828 1060 24852 1062
rect 24908 1060 24932 1062
rect 24988 1060 24994 1062
rect 24686 1051 24994 1060
rect 25056 160 25084 2246
rect 25332 160 25360 3606
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 25608 160 25636 3402
rect 24766 82 24822 160
rect 24596 54 24822 82
rect 24766 0 24822 54
rect 25042 0 25098 160
rect 25318 0 25374 160
rect 25594 0 25650 160
<< via2 >>
rect 6890 8730 6946 8732
rect 6970 8730 7026 8732
rect 7050 8730 7106 8732
rect 7130 8730 7186 8732
rect 6890 8678 6936 8730
rect 6936 8678 6946 8730
rect 6970 8678 7000 8730
rect 7000 8678 7012 8730
rect 7012 8678 7026 8730
rect 7050 8678 7064 8730
rect 7064 8678 7076 8730
rect 7076 8678 7106 8730
rect 7130 8678 7140 8730
rect 7140 8678 7186 8730
rect 6890 8676 6946 8678
rect 6970 8676 7026 8678
rect 7050 8676 7106 8678
rect 7130 8676 7186 8678
rect 12824 8730 12880 8732
rect 12904 8730 12960 8732
rect 12984 8730 13040 8732
rect 13064 8730 13120 8732
rect 12824 8678 12870 8730
rect 12870 8678 12880 8730
rect 12904 8678 12934 8730
rect 12934 8678 12946 8730
rect 12946 8678 12960 8730
rect 12984 8678 12998 8730
rect 12998 8678 13010 8730
rect 13010 8678 13040 8730
rect 13064 8678 13074 8730
rect 13074 8678 13120 8730
rect 12824 8676 12880 8678
rect 12904 8676 12960 8678
rect 12984 8676 13040 8678
rect 13064 8676 13120 8678
rect 3923 8186 3979 8188
rect 4003 8186 4059 8188
rect 4083 8186 4139 8188
rect 4163 8186 4219 8188
rect 3923 8134 3969 8186
rect 3969 8134 3979 8186
rect 4003 8134 4033 8186
rect 4033 8134 4045 8186
rect 4045 8134 4059 8186
rect 4083 8134 4097 8186
rect 4097 8134 4109 8186
rect 4109 8134 4139 8186
rect 4163 8134 4173 8186
rect 4173 8134 4219 8186
rect 3923 8132 3979 8134
rect 4003 8132 4059 8134
rect 4083 8132 4139 8134
rect 4163 8132 4219 8134
rect 3923 7098 3979 7100
rect 4003 7098 4059 7100
rect 4083 7098 4139 7100
rect 4163 7098 4219 7100
rect 3923 7046 3969 7098
rect 3969 7046 3979 7098
rect 4003 7046 4033 7098
rect 4033 7046 4045 7098
rect 4045 7046 4059 7098
rect 4083 7046 4097 7098
rect 4097 7046 4109 7098
rect 4109 7046 4139 7098
rect 4163 7046 4173 7098
rect 4173 7046 4219 7098
rect 3923 7044 3979 7046
rect 4003 7044 4059 7046
rect 4083 7044 4139 7046
rect 4163 7044 4219 7046
rect 3923 6010 3979 6012
rect 4003 6010 4059 6012
rect 4083 6010 4139 6012
rect 4163 6010 4219 6012
rect 3923 5958 3969 6010
rect 3969 5958 3979 6010
rect 4003 5958 4033 6010
rect 4033 5958 4045 6010
rect 4045 5958 4059 6010
rect 4083 5958 4097 6010
rect 4097 5958 4109 6010
rect 4109 5958 4139 6010
rect 4163 5958 4173 6010
rect 4173 5958 4219 6010
rect 3923 5956 3979 5958
rect 4003 5956 4059 5958
rect 4083 5956 4139 5958
rect 4163 5956 4219 5958
rect 3923 4922 3979 4924
rect 4003 4922 4059 4924
rect 4083 4922 4139 4924
rect 4163 4922 4219 4924
rect 3923 4870 3969 4922
rect 3969 4870 3979 4922
rect 4003 4870 4033 4922
rect 4033 4870 4045 4922
rect 4045 4870 4059 4922
rect 4083 4870 4097 4922
rect 4097 4870 4109 4922
rect 4109 4870 4139 4922
rect 4163 4870 4173 4922
rect 4173 4870 4219 4922
rect 3923 4868 3979 4870
rect 4003 4868 4059 4870
rect 4083 4868 4139 4870
rect 4163 4868 4219 4870
rect 3923 3834 3979 3836
rect 4003 3834 4059 3836
rect 4083 3834 4139 3836
rect 4163 3834 4219 3836
rect 3923 3782 3969 3834
rect 3969 3782 3979 3834
rect 4003 3782 4033 3834
rect 4033 3782 4045 3834
rect 4045 3782 4059 3834
rect 4083 3782 4097 3834
rect 4097 3782 4109 3834
rect 4109 3782 4139 3834
rect 4163 3782 4173 3834
rect 4173 3782 4219 3834
rect 3923 3780 3979 3782
rect 4003 3780 4059 3782
rect 4083 3780 4139 3782
rect 4163 3780 4219 3782
rect 6890 7642 6946 7644
rect 6970 7642 7026 7644
rect 7050 7642 7106 7644
rect 7130 7642 7186 7644
rect 6890 7590 6936 7642
rect 6936 7590 6946 7642
rect 6970 7590 7000 7642
rect 7000 7590 7012 7642
rect 7012 7590 7026 7642
rect 7050 7590 7064 7642
rect 7064 7590 7076 7642
rect 7076 7590 7106 7642
rect 7130 7590 7140 7642
rect 7140 7590 7186 7642
rect 6890 7588 6946 7590
rect 6970 7588 7026 7590
rect 7050 7588 7106 7590
rect 7130 7588 7186 7590
rect 6890 6554 6946 6556
rect 6970 6554 7026 6556
rect 7050 6554 7106 6556
rect 7130 6554 7186 6556
rect 6890 6502 6936 6554
rect 6936 6502 6946 6554
rect 6970 6502 7000 6554
rect 7000 6502 7012 6554
rect 7012 6502 7026 6554
rect 7050 6502 7064 6554
rect 7064 6502 7076 6554
rect 7076 6502 7106 6554
rect 7130 6502 7140 6554
rect 7140 6502 7186 6554
rect 6890 6500 6946 6502
rect 6970 6500 7026 6502
rect 7050 6500 7106 6502
rect 7130 6500 7186 6502
rect 8206 6160 8262 6216
rect 6890 5466 6946 5468
rect 6970 5466 7026 5468
rect 7050 5466 7106 5468
rect 7130 5466 7186 5468
rect 6890 5414 6936 5466
rect 6936 5414 6946 5466
rect 6970 5414 7000 5466
rect 7000 5414 7012 5466
rect 7012 5414 7026 5466
rect 7050 5414 7064 5466
rect 7064 5414 7076 5466
rect 7076 5414 7106 5466
rect 7130 5414 7140 5466
rect 7140 5414 7186 5466
rect 6890 5412 6946 5414
rect 6970 5412 7026 5414
rect 7050 5412 7106 5414
rect 7130 5412 7186 5414
rect 6890 4378 6946 4380
rect 6970 4378 7026 4380
rect 7050 4378 7106 4380
rect 7130 4378 7186 4380
rect 6890 4326 6936 4378
rect 6936 4326 6946 4378
rect 6970 4326 7000 4378
rect 7000 4326 7012 4378
rect 7012 4326 7026 4378
rect 7050 4326 7064 4378
rect 7064 4326 7076 4378
rect 7076 4326 7106 4378
rect 7130 4326 7140 4378
rect 7140 4326 7186 4378
rect 6890 4324 6946 4326
rect 6970 4324 7026 4326
rect 7050 4324 7106 4326
rect 7130 4324 7186 4326
rect 9857 8186 9913 8188
rect 9937 8186 9993 8188
rect 10017 8186 10073 8188
rect 10097 8186 10153 8188
rect 9857 8134 9903 8186
rect 9903 8134 9913 8186
rect 9937 8134 9967 8186
rect 9967 8134 9979 8186
rect 9979 8134 9993 8186
rect 10017 8134 10031 8186
rect 10031 8134 10043 8186
rect 10043 8134 10073 8186
rect 10097 8134 10107 8186
rect 10107 8134 10153 8186
rect 9857 8132 9913 8134
rect 9937 8132 9993 8134
rect 10017 8132 10073 8134
rect 10097 8132 10153 8134
rect 9857 7098 9913 7100
rect 9937 7098 9993 7100
rect 10017 7098 10073 7100
rect 10097 7098 10153 7100
rect 9857 7046 9903 7098
rect 9903 7046 9913 7098
rect 9937 7046 9967 7098
rect 9967 7046 9979 7098
rect 9979 7046 9993 7098
rect 10017 7046 10031 7098
rect 10031 7046 10043 7098
rect 10043 7046 10073 7098
rect 10097 7046 10107 7098
rect 10107 7046 10153 7098
rect 9857 7044 9913 7046
rect 9937 7044 9993 7046
rect 10017 7044 10073 7046
rect 10097 7044 10153 7046
rect 9857 6010 9913 6012
rect 9937 6010 9993 6012
rect 10017 6010 10073 6012
rect 10097 6010 10153 6012
rect 9857 5958 9903 6010
rect 9903 5958 9913 6010
rect 9937 5958 9967 6010
rect 9967 5958 9979 6010
rect 9979 5958 9993 6010
rect 10017 5958 10031 6010
rect 10031 5958 10043 6010
rect 10043 5958 10073 6010
rect 10097 5958 10107 6010
rect 10107 5958 10153 6010
rect 9857 5956 9913 5958
rect 9937 5956 9993 5958
rect 10017 5956 10073 5958
rect 10097 5956 10153 5958
rect 12824 7642 12880 7644
rect 12904 7642 12960 7644
rect 12984 7642 13040 7644
rect 13064 7642 13120 7644
rect 12824 7590 12870 7642
rect 12870 7590 12880 7642
rect 12904 7590 12934 7642
rect 12934 7590 12946 7642
rect 12946 7590 12960 7642
rect 12984 7590 12998 7642
rect 12998 7590 13010 7642
rect 13010 7590 13040 7642
rect 13064 7590 13074 7642
rect 13074 7590 13120 7642
rect 12824 7588 12880 7590
rect 12904 7588 12960 7590
rect 12984 7588 13040 7590
rect 13064 7588 13120 7590
rect 12824 6554 12880 6556
rect 12904 6554 12960 6556
rect 12984 6554 13040 6556
rect 13064 6554 13120 6556
rect 12824 6502 12870 6554
rect 12870 6502 12880 6554
rect 12904 6502 12934 6554
rect 12934 6502 12946 6554
rect 12946 6502 12960 6554
rect 12984 6502 12998 6554
rect 12998 6502 13010 6554
rect 13010 6502 13040 6554
rect 13064 6502 13074 6554
rect 13074 6502 13120 6554
rect 12824 6500 12880 6502
rect 12904 6500 12960 6502
rect 12984 6500 13040 6502
rect 13064 6500 13120 6502
rect 18758 8730 18814 8732
rect 18838 8730 18894 8732
rect 18918 8730 18974 8732
rect 18998 8730 19054 8732
rect 18758 8678 18804 8730
rect 18804 8678 18814 8730
rect 18838 8678 18868 8730
rect 18868 8678 18880 8730
rect 18880 8678 18894 8730
rect 18918 8678 18932 8730
rect 18932 8678 18944 8730
rect 18944 8678 18974 8730
rect 18998 8678 19008 8730
rect 19008 8678 19054 8730
rect 18758 8676 18814 8678
rect 18838 8676 18894 8678
rect 18918 8676 18974 8678
rect 18998 8676 19054 8678
rect 15791 8186 15847 8188
rect 15871 8186 15927 8188
rect 15951 8186 16007 8188
rect 16031 8186 16087 8188
rect 15791 8134 15837 8186
rect 15837 8134 15847 8186
rect 15871 8134 15901 8186
rect 15901 8134 15913 8186
rect 15913 8134 15927 8186
rect 15951 8134 15965 8186
rect 15965 8134 15977 8186
rect 15977 8134 16007 8186
rect 16031 8134 16041 8186
rect 16041 8134 16087 8186
rect 15791 8132 15847 8134
rect 15871 8132 15927 8134
rect 15951 8132 16007 8134
rect 16031 8132 16087 8134
rect 15791 7098 15847 7100
rect 15871 7098 15927 7100
rect 15951 7098 16007 7100
rect 16031 7098 16087 7100
rect 15791 7046 15837 7098
rect 15837 7046 15847 7098
rect 15871 7046 15901 7098
rect 15901 7046 15913 7098
rect 15913 7046 15927 7098
rect 15951 7046 15965 7098
rect 15965 7046 15977 7098
rect 15977 7046 16007 7098
rect 16031 7046 16041 7098
rect 16041 7046 16087 7098
rect 15791 7044 15847 7046
rect 15871 7044 15927 7046
rect 15951 7044 16007 7046
rect 16031 7044 16087 7046
rect 15791 6010 15847 6012
rect 15871 6010 15927 6012
rect 15951 6010 16007 6012
rect 16031 6010 16087 6012
rect 15791 5958 15837 6010
rect 15837 5958 15847 6010
rect 15871 5958 15901 6010
rect 15901 5958 15913 6010
rect 15913 5958 15927 6010
rect 15951 5958 15965 6010
rect 15965 5958 15977 6010
rect 15977 5958 16007 6010
rect 16031 5958 16041 6010
rect 16041 5958 16087 6010
rect 15791 5956 15847 5958
rect 15871 5956 15927 5958
rect 15951 5956 16007 5958
rect 16031 5956 16087 5958
rect 12824 5466 12880 5468
rect 12904 5466 12960 5468
rect 12984 5466 13040 5468
rect 13064 5466 13120 5468
rect 12824 5414 12870 5466
rect 12870 5414 12880 5466
rect 12904 5414 12934 5466
rect 12934 5414 12946 5466
rect 12946 5414 12960 5466
rect 12984 5414 12998 5466
rect 12998 5414 13010 5466
rect 13010 5414 13040 5466
rect 13064 5414 13074 5466
rect 13074 5414 13120 5466
rect 12824 5412 12880 5414
rect 12904 5412 12960 5414
rect 12984 5412 13040 5414
rect 13064 5412 13120 5414
rect 9857 4922 9913 4924
rect 9937 4922 9993 4924
rect 10017 4922 10073 4924
rect 10097 4922 10153 4924
rect 9857 4870 9903 4922
rect 9903 4870 9913 4922
rect 9937 4870 9967 4922
rect 9967 4870 9979 4922
rect 9979 4870 9993 4922
rect 10017 4870 10031 4922
rect 10031 4870 10043 4922
rect 10043 4870 10073 4922
rect 10097 4870 10107 4922
rect 10107 4870 10153 4922
rect 9857 4868 9913 4870
rect 9937 4868 9993 4870
rect 10017 4868 10073 4870
rect 10097 4868 10153 4870
rect 15791 4922 15847 4924
rect 15871 4922 15927 4924
rect 15951 4922 16007 4924
rect 16031 4922 16087 4924
rect 15791 4870 15837 4922
rect 15837 4870 15847 4922
rect 15871 4870 15901 4922
rect 15901 4870 15913 4922
rect 15913 4870 15927 4922
rect 15951 4870 15965 4922
rect 15965 4870 15977 4922
rect 15977 4870 16007 4922
rect 16031 4870 16041 4922
rect 16041 4870 16087 4922
rect 15791 4868 15847 4870
rect 15871 4868 15927 4870
rect 15951 4868 16007 4870
rect 16031 4868 16087 4870
rect 12824 4378 12880 4380
rect 12904 4378 12960 4380
rect 12984 4378 13040 4380
rect 13064 4378 13120 4380
rect 12824 4326 12870 4378
rect 12870 4326 12880 4378
rect 12904 4326 12934 4378
rect 12934 4326 12946 4378
rect 12946 4326 12960 4378
rect 12984 4326 12998 4378
rect 12998 4326 13010 4378
rect 13010 4326 13040 4378
rect 13064 4326 13074 4378
rect 13074 4326 13120 4378
rect 12824 4324 12880 4326
rect 12904 4324 12960 4326
rect 12984 4324 13040 4326
rect 13064 4324 13120 4326
rect 9857 3834 9913 3836
rect 9937 3834 9993 3836
rect 10017 3834 10073 3836
rect 10097 3834 10153 3836
rect 9857 3782 9903 3834
rect 9903 3782 9913 3834
rect 9937 3782 9967 3834
rect 9967 3782 9979 3834
rect 9979 3782 9993 3834
rect 10017 3782 10031 3834
rect 10031 3782 10043 3834
rect 10043 3782 10073 3834
rect 10097 3782 10107 3834
rect 10107 3782 10153 3834
rect 9857 3780 9913 3782
rect 9937 3780 9993 3782
rect 10017 3780 10073 3782
rect 10097 3780 10153 3782
rect 15791 3834 15847 3836
rect 15871 3834 15927 3836
rect 15951 3834 16007 3836
rect 16031 3834 16087 3836
rect 15791 3782 15837 3834
rect 15837 3782 15847 3834
rect 15871 3782 15901 3834
rect 15901 3782 15913 3834
rect 15913 3782 15927 3834
rect 15951 3782 15965 3834
rect 15965 3782 15977 3834
rect 15977 3782 16007 3834
rect 16031 3782 16041 3834
rect 16041 3782 16087 3834
rect 15791 3780 15847 3782
rect 15871 3780 15927 3782
rect 15951 3780 16007 3782
rect 16031 3780 16087 3782
rect 9494 3460 9550 3496
rect 9494 3440 9496 3460
rect 9496 3440 9548 3460
rect 9548 3440 9550 3460
rect 6890 3290 6946 3292
rect 6970 3290 7026 3292
rect 7050 3290 7106 3292
rect 7130 3290 7186 3292
rect 6890 3238 6936 3290
rect 6936 3238 6946 3290
rect 6970 3238 7000 3290
rect 7000 3238 7012 3290
rect 7012 3238 7026 3290
rect 7050 3238 7064 3290
rect 7064 3238 7076 3290
rect 7076 3238 7106 3290
rect 7130 3238 7140 3290
rect 7140 3238 7186 3290
rect 6890 3236 6946 3238
rect 6970 3236 7026 3238
rect 7050 3236 7106 3238
rect 7130 3236 7186 3238
rect 12824 3290 12880 3292
rect 12904 3290 12960 3292
rect 12984 3290 13040 3292
rect 13064 3290 13120 3292
rect 12824 3238 12870 3290
rect 12870 3238 12880 3290
rect 12904 3238 12934 3290
rect 12934 3238 12946 3290
rect 12946 3238 12960 3290
rect 12984 3238 12998 3290
rect 12998 3238 13010 3290
rect 13010 3238 13040 3290
rect 13064 3238 13074 3290
rect 13074 3238 13120 3290
rect 12824 3236 12880 3238
rect 12904 3236 12960 3238
rect 12984 3236 13040 3238
rect 13064 3236 13120 3238
rect 7378 3032 7434 3088
rect 1490 2524 1492 2544
rect 1492 2524 1544 2544
rect 1544 2524 1546 2544
rect 1490 2488 1546 2524
rect 1674 176 1730 232
rect 3923 2746 3979 2748
rect 4003 2746 4059 2748
rect 4083 2746 4139 2748
rect 4163 2746 4219 2748
rect 3923 2694 3969 2746
rect 3969 2694 3979 2746
rect 4003 2694 4033 2746
rect 4033 2694 4045 2746
rect 4045 2694 4059 2746
rect 4083 2694 4097 2746
rect 4097 2694 4109 2746
rect 4109 2694 4139 2746
rect 4163 2694 4173 2746
rect 4173 2694 4219 2746
rect 3923 2692 3979 2694
rect 4003 2692 4059 2694
rect 4083 2692 4139 2694
rect 4163 2692 4219 2694
rect 3923 1658 3979 1660
rect 4003 1658 4059 1660
rect 4083 1658 4139 1660
rect 4163 1658 4219 1660
rect 3923 1606 3969 1658
rect 3969 1606 3979 1658
rect 4003 1606 4033 1658
rect 4033 1606 4045 1658
rect 4045 1606 4059 1658
rect 4083 1606 4097 1658
rect 4097 1606 4109 1658
rect 4109 1606 4139 1658
rect 4163 1606 4173 1658
rect 4173 1606 4219 1658
rect 3923 1604 3979 1606
rect 4003 1604 4059 1606
rect 4083 1604 4139 1606
rect 4163 1604 4219 1606
rect 4158 1400 4214 1456
rect 5354 856 5410 912
rect 5814 720 5870 776
rect 6550 2352 6606 2408
rect 6642 1808 6698 1864
rect 6890 2202 6946 2204
rect 6970 2202 7026 2204
rect 7050 2202 7106 2204
rect 7130 2202 7186 2204
rect 6890 2150 6936 2202
rect 6936 2150 6946 2202
rect 6970 2150 7000 2202
rect 7000 2150 7012 2202
rect 7012 2150 7026 2202
rect 7050 2150 7064 2202
rect 7064 2150 7076 2202
rect 7076 2150 7106 2202
rect 7130 2150 7140 2202
rect 7140 2150 7186 2202
rect 6890 2148 6946 2150
rect 6970 2148 7026 2150
rect 7050 2148 7106 2150
rect 7130 2148 7186 2150
rect 8114 2216 8170 2272
rect 6826 1964 6882 2000
rect 6826 1944 6828 1964
rect 6828 1944 6880 1964
rect 6880 1944 6882 1964
rect 6918 1300 6920 1320
rect 6920 1300 6972 1320
rect 6972 1300 6974 1320
rect 6918 1264 6974 1300
rect 6890 1114 6946 1116
rect 6970 1114 7026 1116
rect 7050 1114 7106 1116
rect 7130 1114 7186 1116
rect 6890 1062 6936 1114
rect 6936 1062 6946 1114
rect 6970 1062 7000 1114
rect 7000 1062 7012 1114
rect 7012 1062 7026 1114
rect 7050 1062 7064 1114
rect 7064 1062 7076 1114
rect 7076 1062 7106 1114
rect 7130 1062 7140 1114
rect 7140 1062 7186 1114
rect 6890 1060 6946 1062
rect 6970 1060 7026 1062
rect 7050 1060 7106 1062
rect 7130 1060 7186 1062
rect 6550 584 6606 640
rect 6734 176 6790 232
rect 7562 1128 7618 1184
rect 7562 312 7618 368
rect 8942 2100 8998 2136
rect 8942 2080 8944 2100
rect 8944 2080 8996 2100
rect 8996 2080 8998 2100
rect 7930 1264 7986 1320
rect 9034 1672 9090 1728
rect 8942 448 8998 504
rect 9857 2746 9913 2748
rect 9937 2746 9993 2748
rect 10017 2746 10073 2748
rect 10097 2746 10153 2748
rect 9857 2694 9903 2746
rect 9903 2694 9913 2746
rect 9937 2694 9967 2746
rect 9967 2694 9979 2746
rect 9979 2694 9993 2746
rect 10017 2694 10031 2746
rect 10031 2694 10043 2746
rect 10043 2694 10073 2746
rect 10097 2694 10107 2746
rect 10107 2694 10153 2746
rect 9857 2692 9913 2694
rect 9937 2692 9993 2694
rect 10017 2692 10073 2694
rect 10097 2692 10153 2694
rect 9862 2488 9918 2544
rect 12438 2488 12494 2544
rect 9218 584 9274 640
rect 10966 2080 11022 2136
rect 9678 1672 9734 1728
rect 9857 1658 9913 1660
rect 9937 1658 9993 1660
rect 10017 1658 10073 1660
rect 10097 1658 10153 1660
rect 9857 1606 9903 1658
rect 9903 1606 9913 1658
rect 9937 1606 9967 1658
rect 9967 1606 9979 1658
rect 9979 1606 9993 1658
rect 10017 1606 10031 1658
rect 10031 1606 10043 1658
rect 10043 1606 10073 1658
rect 10097 1606 10107 1658
rect 10107 1606 10153 1658
rect 9857 1604 9913 1606
rect 9937 1604 9993 1606
rect 10017 1604 10073 1606
rect 10097 1604 10153 1606
rect 12346 2216 12402 2272
rect 12346 1672 12402 1728
rect 12438 1536 12494 1592
rect 12824 2202 12880 2204
rect 12904 2202 12960 2204
rect 12984 2202 13040 2204
rect 13064 2202 13120 2204
rect 12824 2150 12870 2202
rect 12870 2150 12880 2202
rect 12904 2150 12934 2202
rect 12934 2150 12946 2202
rect 12946 2150 12960 2202
rect 12984 2150 12998 2202
rect 12998 2150 13010 2202
rect 13010 2150 13040 2202
rect 13064 2150 13074 2202
rect 13074 2150 13120 2202
rect 12824 2148 12880 2150
rect 12904 2148 12960 2150
rect 12984 2148 13040 2150
rect 13064 2148 13120 2150
rect 13634 1964 13690 2000
rect 13634 1944 13636 1964
rect 13636 1944 13688 1964
rect 13688 1944 13690 1964
rect 12530 1128 12586 1184
rect 12806 1400 12862 1456
rect 12824 1114 12880 1116
rect 12904 1114 12960 1116
rect 12984 1114 13040 1116
rect 13064 1114 13120 1116
rect 12824 1062 12870 1114
rect 12870 1062 12880 1114
rect 12904 1062 12934 1114
rect 12934 1062 12946 1114
rect 12946 1062 12960 1114
rect 12984 1062 12998 1114
rect 12998 1062 13010 1114
rect 13010 1062 13040 1114
rect 13064 1062 13074 1114
rect 13074 1062 13120 1114
rect 12824 1060 12880 1062
rect 12904 1060 12960 1062
rect 12984 1060 13040 1062
rect 13064 1060 13120 1062
rect 12714 176 12770 232
rect 15791 2746 15847 2748
rect 15871 2746 15927 2748
rect 15951 2746 16007 2748
rect 16031 2746 16087 2748
rect 15791 2694 15837 2746
rect 15837 2694 15847 2746
rect 15871 2694 15901 2746
rect 15901 2694 15913 2746
rect 15913 2694 15927 2746
rect 15951 2694 15965 2746
rect 15965 2694 15977 2746
rect 15977 2694 16007 2746
rect 16031 2694 16041 2746
rect 16041 2694 16087 2746
rect 15791 2692 15847 2694
rect 15871 2692 15927 2694
rect 15951 2692 16007 2694
rect 16031 2692 16087 2694
rect 15658 2624 15714 2680
rect 18758 7642 18814 7644
rect 18838 7642 18894 7644
rect 18918 7642 18974 7644
rect 18998 7642 19054 7644
rect 18758 7590 18804 7642
rect 18804 7590 18814 7642
rect 18838 7590 18868 7642
rect 18868 7590 18880 7642
rect 18880 7590 18894 7642
rect 18918 7590 18932 7642
rect 18932 7590 18944 7642
rect 18944 7590 18974 7642
rect 18998 7590 19008 7642
rect 19008 7590 19054 7642
rect 18758 7588 18814 7590
rect 18838 7588 18894 7590
rect 18918 7588 18974 7590
rect 18998 7588 19054 7590
rect 18758 6554 18814 6556
rect 18838 6554 18894 6556
rect 18918 6554 18974 6556
rect 18998 6554 19054 6556
rect 18758 6502 18804 6554
rect 18804 6502 18814 6554
rect 18838 6502 18868 6554
rect 18868 6502 18880 6554
rect 18880 6502 18894 6554
rect 18918 6502 18932 6554
rect 18932 6502 18944 6554
rect 18944 6502 18974 6554
rect 18998 6502 19008 6554
rect 19008 6502 19054 6554
rect 18758 6500 18814 6502
rect 18838 6500 18894 6502
rect 18918 6500 18974 6502
rect 18998 6500 19054 6502
rect 18758 5466 18814 5468
rect 18838 5466 18894 5468
rect 18918 5466 18974 5468
rect 18998 5466 19054 5468
rect 18758 5414 18804 5466
rect 18804 5414 18814 5466
rect 18838 5414 18868 5466
rect 18868 5414 18880 5466
rect 18880 5414 18894 5466
rect 18918 5414 18932 5466
rect 18932 5414 18944 5466
rect 18944 5414 18974 5466
rect 18998 5414 19008 5466
rect 19008 5414 19054 5466
rect 18758 5412 18814 5414
rect 18838 5412 18894 5414
rect 18918 5412 18974 5414
rect 18998 5412 19054 5414
rect 18758 4378 18814 4380
rect 18838 4378 18894 4380
rect 18918 4378 18974 4380
rect 18998 4378 19054 4380
rect 18758 4326 18804 4378
rect 18804 4326 18814 4378
rect 18838 4326 18868 4378
rect 18868 4326 18880 4378
rect 18880 4326 18894 4378
rect 18918 4326 18932 4378
rect 18932 4326 18944 4378
rect 18944 4326 18974 4378
rect 18998 4326 19008 4378
rect 19008 4326 19054 4378
rect 18758 4324 18814 4326
rect 18838 4324 18894 4326
rect 18918 4324 18974 4326
rect 18998 4324 19054 4326
rect 18758 3290 18814 3292
rect 18838 3290 18894 3292
rect 18918 3290 18974 3292
rect 18998 3290 19054 3292
rect 18758 3238 18804 3290
rect 18804 3238 18814 3290
rect 18838 3238 18868 3290
rect 18868 3238 18880 3290
rect 18880 3238 18894 3290
rect 18918 3238 18932 3290
rect 18932 3238 18944 3290
rect 18944 3238 18974 3290
rect 18998 3238 19008 3290
rect 19008 3238 19054 3290
rect 18758 3236 18814 3238
rect 18838 3236 18894 3238
rect 18918 3236 18974 3238
rect 18998 3236 19054 3238
rect 21725 8186 21781 8188
rect 21805 8186 21861 8188
rect 21885 8186 21941 8188
rect 21965 8186 22021 8188
rect 21725 8134 21771 8186
rect 21771 8134 21781 8186
rect 21805 8134 21835 8186
rect 21835 8134 21847 8186
rect 21847 8134 21861 8186
rect 21885 8134 21899 8186
rect 21899 8134 21911 8186
rect 21911 8134 21941 8186
rect 21965 8134 21975 8186
rect 21975 8134 22021 8186
rect 21725 8132 21781 8134
rect 21805 8132 21861 8134
rect 21885 8132 21941 8134
rect 21965 8132 22021 8134
rect 21725 7098 21781 7100
rect 21805 7098 21861 7100
rect 21885 7098 21941 7100
rect 21965 7098 22021 7100
rect 21725 7046 21771 7098
rect 21771 7046 21781 7098
rect 21805 7046 21835 7098
rect 21835 7046 21847 7098
rect 21847 7046 21861 7098
rect 21885 7046 21899 7098
rect 21899 7046 21911 7098
rect 21911 7046 21941 7098
rect 21965 7046 21975 7098
rect 21975 7046 22021 7098
rect 21725 7044 21781 7046
rect 21805 7044 21861 7046
rect 21885 7044 21941 7046
rect 21965 7044 22021 7046
rect 21725 6010 21781 6012
rect 21805 6010 21861 6012
rect 21885 6010 21941 6012
rect 21965 6010 22021 6012
rect 21725 5958 21771 6010
rect 21771 5958 21781 6010
rect 21805 5958 21835 6010
rect 21835 5958 21847 6010
rect 21847 5958 21861 6010
rect 21885 5958 21899 6010
rect 21899 5958 21911 6010
rect 21911 5958 21941 6010
rect 21965 5958 21975 6010
rect 21975 5958 22021 6010
rect 21725 5956 21781 5958
rect 21805 5956 21861 5958
rect 21885 5956 21941 5958
rect 21965 5956 22021 5958
rect 21725 4922 21781 4924
rect 21805 4922 21861 4924
rect 21885 4922 21941 4924
rect 21965 4922 22021 4924
rect 21725 4870 21771 4922
rect 21771 4870 21781 4922
rect 21805 4870 21835 4922
rect 21835 4870 21847 4922
rect 21847 4870 21861 4922
rect 21885 4870 21899 4922
rect 21899 4870 21911 4922
rect 21911 4870 21941 4922
rect 21965 4870 21975 4922
rect 21975 4870 22021 4922
rect 21725 4868 21781 4870
rect 21805 4868 21861 4870
rect 21885 4868 21941 4870
rect 21965 4868 22021 4870
rect 15290 1672 15346 1728
rect 15791 1658 15847 1660
rect 15871 1658 15927 1660
rect 15951 1658 16007 1660
rect 16031 1658 16087 1660
rect 15791 1606 15837 1658
rect 15837 1606 15847 1658
rect 15871 1606 15901 1658
rect 15901 1606 15913 1658
rect 15913 1606 15927 1658
rect 15951 1606 15965 1658
rect 15965 1606 15977 1658
rect 15977 1606 16007 1658
rect 16031 1606 16041 1658
rect 16041 1606 16087 1658
rect 15791 1604 15847 1606
rect 15871 1604 15927 1606
rect 15951 1604 16007 1606
rect 16031 1604 16087 1606
rect 16302 1400 16358 1456
rect 16210 584 16266 640
rect 17130 312 17186 368
rect 17958 1264 18014 1320
rect 18758 2202 18814 2204
rect 18838 2202 18894 2204
rect 18918 2202 18974 2204
rect 18998 2202 19054 2204
rect 18758 2150 18804 2202
rect 18804 2150 18814 2202
rect 18838 2150 18868 2202
rect 18868 2150 18880 2202
rect 18880 2150 18894 2202
rect 18918 2150 18932 2202
rect 18932 2150 18944 2202
rect 18944 2150 18974 2202
rect 18998 2150 19008 2202
rect 19008 2150 19054 2202
rect 18758 2148 18814 2150
rect 18838 2148 18894 2150
rect 18918 2148 18974 2150
rect 18998 2148 19054 2150
rect 18970 1672 19026 1728
rect 18602 1300 18604 1320
rect 18604 1300 18656 1320
rect 18656 1300 18658 1320
rect 18602 1264 18658 1300
rect 17958 720 18014 776
rect 18758 1114 18814 1116
rect 18838 1114 18894 1116
rect 18918 1114 18974 1116
rect 18998 1114 19054 1116
rect 18758 1062 18804 1114
rect 18804 1062 18814 1114
rect 18838 1062 18868 1114
rect 18868 1062 18880 1114
rect 18880 1062 18894 1114
rect 18918 1062 18932 1114
rect 18932 1062 18944 1114
rect 18944 1062 18974 1114
rect 18998 1062 19008 1114
rect 19008 1062 19054 1114
rect 18758 1060 18814 1062
rect 18838 1060 18894 1062
rect 18918 1060 18974 1062
rect 18998 1060 19054 1062
rect 19338 1672 19394 1728
rect 19982 1808 20038 1864
rect 20626 2508 20682 2544
rect 20626 2488 20628 2508
rect 20628 2488 20680 2508
rect 20680 2488 20682 2508
rect 21725 3834 21781 3836
rect 21805 3834 21861 3836
rect 21885 3834 21941 3836
rect 21965 3834 22021 3836
rect 21725 3782 21771 3834
rect 21771 3782 21781 3834
rect 21805 3782 21835 3834
rect 21835 3782 21847 3834
rect 21847 3782 21861 3834
rect 21885 3782 21899 3834
rect 21899 3782 21911 3834
rect 21911 3782 21941 3834
rect 21965 3782 21975 3834
rect 21975 3782 22021 3834
rect 21725 3780 21781 3782
rect 21805 3780 21861 3782
rect 21885 3780 21941 3782
rect 21965 3780 22021 3782
rect 21725 2746 21781 2748
rect 21805 2746 21861 2748
rect 21885 2746 21941 2748
rect 21965 2746 22021 2748
rect 21725 2694 21771 2746
rect 21771 2694 21781 2746
rect 21805 2694 21835 2746
rect 21835 2694 21847 2746
rect 21847 2694 21861 2746
rect 21885 2694 21899 2746
rect 21899 2694 21911 2746
rect 21911 2694 21941 2746
rect 21965 2694 21975 2746
rect 21975 2694 22021 2746
rect 21725 2692 21781 2694
rect 21805 2692 21861 2694
rect 21885 2692 21941 2694
rect 21965 2692 22021 2694
rect 20810 584 20866 640
rect 21362 448 21418 504
rect 21730 2352 21786 2408
rect 21725 1658 21781 1660
rect 21805 1658 21861 1660
rect 21885 1658 21941 1660
rect 21965 1658 22021 1660
rect 21725 1606 21771 1658
rect 21771 1606 21781 1658
rect 21805 1606 21835 1658
rect 21835 1606 21847 1658
rect 21847 1606 21861 1658
rect 21885 1606 21899 1658
rect 21899 1606 21911 1658
rect 21911 1606 21941 1658
rect 21965 1606 21975 1658
rect 21975 1606 22021 1658
rect 21725 1604 21781 1606
rect 21805 1604 21861 1606
rect 21885 1604 21941 1606
rect 21965 1604 22021 1606
rect 22834 2524 22836 2544
rect 22836 2524 22888 2544
rect 22888 2524 22890 2544
rect 22834 2488 22890 2524
rect 22282 856 22338 912
rect 24692 8730 24748 8732
rect 24772 8730 24828 8732
rect 24852 8730 24908 8732
rect 24932 8730 24988 8732
rect 24692 8678 24738 8730
rect 24738 8678 24748 8730
rect 24772 8678 24802 8730
rect 24802 8678 24814 8730
rect 24814 8678 24828 8730
rect 24852 8678 24866 8730
rect 24866 8678 24878 8730
rect 24878 8678 24908 8730
rect 24932 8678 24942 8730
rect 24942 8678 24988 8730
rect 24692 8676 24748 8678
rect 24772 8676 24828 8678
rect 24852 8676 24908 8678
rect 24932 8676 24988 8678
rect 23478 2760 23534 2816
rect 23754 2760 23810 2816
rect 23110 1164 23112 1184
rect 23112 1164 23164 1184
rect 23164 1164 23166 1184
rect 23110 1128 23166 1164
rect 23478 992 23534 1048
rect 24692 7642 24748 7644
rect 24772 7642 24828 7644
rect 24852 7642 24908 7644
rect 24932 7642 24988 7644
rect 24692 7590 24738 7642
rect 24738 7590 24748 7642
rect 24772 7590 24802 7642
rect 24802 7590 24814 7642
rect 24814 7590 24828 7642
rect 24852 7590 24866 7642
rect 24866 7590 24878 7642
rect 24878 7590 24908 7642
rect 24932 7590 24942 7642
rect 24942 7590 24988 7642
rect 24692 7588 24748 7590
rect 24772 7588 24828 7590
rect 24852 7588 24908 7590
rect 24932 7588 24988 7590
rect 24692 6554 24748 6556
rect 24772 6554 24828 6556
rect 24852 6554 24908 6556
rect 24932 6554 24988 6556
rect 24692 6502 24738 6554
rect 24738 6502 24748 6554
rect 24772 6502 24802 6554
rect 24802 6502 24814 6554
rect 24814 6502 24828 6554
rect 24852 6502 24866 6554
rect 24866 6502 24878 6554
rect 24878 6502 24908 6554
rect 24932 6502 24942 6554
rect 24942 6502 24988 6554
rect 24692 6500 24748 6502
rect 24772 6500 24828 6502
rect 24852 6500 24908 6502
rect 24932 6500 24988 6502
rect 24692 5466 24748 5468
rect 24772 5466 24828 5468
rect 24852 5466 24908 5468
rect 24932 5466 24988 5468
rect 24692 5414 24738 5466
rect 24738 5414 24748 5466
rect 24772 5414 24802 5466
rect 24802 5414 24814 5466
rect 24814 5414 24828 5466
rect 24852 5414 24866 5466
rect 24866 5414 24878 5466
rect 24878 5414 24908 5466
rect 24932 5414 24942 5466
rect 24942 5414 24988 5466
rect 24692 5412 24748 5414
rect 24772 5412 24828 5414
rect 24852 5412 24908 5414
rect 24932 5412 24988 5414
rect 24692 4378 24748 4380
rect 24772 4378 24828 4380
rect 24852 4378 24908 4380
rect 24932 4378 24988 4380
rect 24692 4326 24738 4378
rect 24738 4326 24748 4378
rect 24772 4326 24802 4378
rect 24802 4326 24814 4378
rect 24814 4326 24828 4378
rect 24852 4326 24866 4378
rect 24866 4326 24878 4378
rect 24878 4326 24908 4378
rect 24932 4326 24942 4378
rect 24942 4326 24988 4378
rect 24692 4324 24748 4326
rect 24772 4324 24828 4326
rect 24852 4324 24908 4326
rect 24932 4324 24988 4326
rect 24692 3290 24748 3292
rect 24772 3290 24828 3292
rect 24852 3290 24908 3292
rect 24932 3290 24988 3292
rect 24692 3238 24738 3290
rect 24738 3238 24748 3290
rect 24772 3238 24802 3290
rect 24802 3238 24814 3290
rect 24814 3238 24828 3290
rect 24852 3238 24866 3290
rect 24866 3238 24878 3290
rect 24878 3238 24908 3290
rect 24932 3238 24942 3290
rect 24942 3238 24988 3290
rect 24692 3236 24748 3238
rect 24772 3236 24828 3238
rect 24852 3236 24908 3238
rect 24932 3236 24988 3238
rect 24692 2202 24748 2204
rect 24772 2202 24828 2204
rect 24852 2202 24908 2204
rect 24932 2202 24988 2204
rect 24692 2150 24738 2202
rect 24738 2150 24748 2202
rect 24772 2150 24802 2202
rect 24802 2150 24814 2202
rect 24814 2150 24828 2202
rect 24852 2150 24866 2202
rect 24866 2150 24878 2202
rect 24878 2150 24908 2202
rect 24932 2150 24942 2202
rect 24942 2150 24988 2202
rect 24692 2148 24748 2150
rect 24772 2148 24828 2150
rect 24852 2148 24908 2150
rect 24932 2148 24988 2150
rect 24692 1114 24748 1116
rect 24772 1114 24828 1116
rect 24852 1114 24908 1116
rect 24932 1114 24988 1116
rect 24692 1062 24738 1114
rect 24738 1062 24748 1114
rect 24772 1062 24802 1114
rect 24802 1062 24814 1114
rect 24814 1062 24828 1114
rect 24852 1062 24866 1114
rect 24866 1062 24878 1114
rect 24878 1062 24908 1114
rect 24932 1062 24942 1114
rect 24942 1062 24988 1114
rect 24692 1060 24748 1062
rect 24772 1060 24828 1062
rect 24852 1060 24908 1062
rect 24932 1060 24988 1062
<< metal3 >>
rect 6880 8736 7196 8737
rect 6880 8672 6886 8736
rect 6950 8672 6966 8736
rect 7030 8672 7046 8736
rect 7110 8672 7126 8736
rect 7190 8672 7196 8736
rect 6880 8671 7196 8672
rect 12814 8736 13130 8737
rect 12814 8672 12820 8736
rect 12884 8672 12900 8736
rect 12964 8672 12980 8736
rect 13044 8672 13060 8736
rect 13124 8672 13130 8736
rect 12814 8671 13130 8672
rect 18748 8736 19064 8737
rect 18748 8672 18754 8736
rect 18818 8672 18834 8736
rect 18898 8672 18914 8736
rect 18978 8672 18994 8736
rect 19058 8672 19064 8736
rect 18748 8671 19064 8672
rect 24682 8736 24998 8737
rect 24682 8672 24688 8736
rect 24752 8672 24768 8736
rect 24832 8672 24848 8736
rect 24912 8672 24928 8736
rect 24992 8672 24998 8736
rect 24682 8671 24998 8672
rect 3913 8192 4229 8193
rect 3913 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4229 8192
rect 3913 8127 4229 8128
rect 9847 8192 10163 8193
rect 9847 8128 9853 8192
rect 9917 8128 9933 8192
rect 9997 8128 10013 8192
rect 10077 8128 10093 8192
rect 10157 8128 10163 8192
rect 9847 8127 10163 8128
rect 15781 8192 16097 8193
rect 15781 8128 15787 8192
rect 15851 8128 15867 8192
rect 15931 8128 15947 8192
rect 16011 8128 16027 8192
rect 16091 8128 16097 8192
rect 15781 8127 16097 8128
rect 21715 8192 22031 8193
rect 21715 8128 21721 8192
rect 21785 8128 21801 8192
rect 21865 8128 21881 8192
rect 21945 8128 21961 8192
rect 22025 8128 22031 8192
rect 21715 8127 22031 8128
rect 6880 7648 7196 7649
rect 6880 7584 6886 7648
rect 6950 7584 6966 7648
rect 7030 7584 7046 7648
rect 7110 7584 7126 7648
rect 7190 7584 7196 7648
rect 6880 7583 7196 7584
rect 12814 7648 13130 7649
rect 12814 7584 12820 7648
rect 12884 7584 12900 7648
rect 12964 7584 12980 7648
rect 13044 7584 13060 7648
rect 13124 7584 13130 7648
rect 12814 7583 13130 7584
rect 18748 7648 19064 7649
rect 18748 7584 18754 7648
rect 18818 7584 18834 7648
rect 18898 7584 18914 7648
rect 18978 7584 18994 7648
rect 19058 7584 19064 7648
rect 18748 7583 19064 7584
rect 24682 7648 24998 7649
rect 24682 7584 24688 7648
rect 24752 7584 24768 7648
rect 24832 7584 24848 7648
rect 24912 7584 24928 7648
rect 24992 7584 24998 7648
rect 24682 7583 24998 7584
rect 3913 7104 4229 7105
rect 3913 7040 3919 7104
rect 3983 7040 3999 7104
rect 4063 7040 4079 7104
rect 4143 7040 4159 7104
rect 4223 7040 4229 7104
rect 3913 7039 4229 7040
rect 9847 7104 10163 7105
rect 9847 7040 9853 7104
rect 9917 7040 9933 7104
rect 9997 7040 10013 7104
rect 10077 7040 10093 7104
rect 10157 7040 10163 7104
rect 9847 7039 10163 7040
rect 15781 7104 16097 7105
rect 15781 7040 15787 7104
rect 15851 7040 15867 7104
rect 15931 7040 15947 7104
rect 16011 7040 16027 7104
rect 16091 7040 16097 7104
rect 15781 7039 16097 7040
rect 21715 7104 22031 7105
rect 21715 7040 21721 7104
rect 21785 7040 21801 7104
rect 21865 7040 21881 7104
rect 21945 7040 21961 7104
rect 22025 7040 22031 7104
rect 21715 7039 22031 7040
rect 6880 6560 7196 6561
rect 6880 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7196 6560
rect 6880 6495 7196 6496
rect 12814 6560 13130 6561
rect 12814 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13130 6560
rect 12814 6495 13130 6496
rect 18748 6560 19064 6561
rect 18748 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19064 6560
rect 18748 6495 19064 6496
rect 24682 6560 24998 6561
rect 24682 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 24998 6560
rect 24682 6495 24998 6496
rect 8201 6218 8267 6221
rect 19742 6218 19748 6220
rect 8201 6216 19748 6218
rect 8201 6160 8206 6216
rect 8262 6160 19748 6216
rect 8201 6158 19748 6160
rect 8201 6155 8267 6158
rect 19742 6156 19748 6158
rect 19812 6156 19818 6220
rect 3913 6016 4229 6017
rect 3913 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4229 6016
rect 3913 5951 4229 5952
rect 9847 6016 10163 6017
rect 9847 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10163 6016
rect 9847 5951 10163 5952
rect 15781 6016 16097 6017
rect 15781 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16097 6016
rect 15781 5951 16097 5952
rect 21715 6016 22031 6017
rect 21715 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22031 6016
rect 21715 5951 22031 5952
rect 6880 5472 7196 5473
rect 6880 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7196 5472
rect 6880 5407 7196 5408
rect 12814 5472 13130 5473
rect 12814 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13130 5472
rect 12814 5407 13130 5408
rect 18748 5472 19064 5473
rect 18748 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19064 5472
rect 18748 5407 19064 5408
rect 24682 5472 24998 5473
rect 24682 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 24998 5472
rect 24682 5407 24998 5408
rect 3913 4928 4229 4929
rect 3913 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4229 4928
rect 3913 4863 4229 4864
rect 9847 4928 10163 4929
rect 9847 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10163 4928
rect 9847 4863 10163 4864
rect 15781 4928 16097 4929
rect 15781 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16097 4928
rect 15781 4863 16097 4864
rect 21715 4928 22031 4929
rect 21715 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22031 4928
rect 21715 4863 22031 4864
rect 6880 4384 7196 4385
rect 6880 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7196 4384
rect 6880 4319 7196 4320
rect 12814 4384 13130 4385
rect 12814 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13130 4384
rect 12814 4319 13130 4320
rect 18748 4384 19064 4385
rect 18748 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19064 4384
rect 18748 4319 19064 4320
rect 24682 4384 24998 4385
rect 24682 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 24998 4384
rect 24682 4319 24998 4320
rect 3913 3840 4229 3841
rect 3913 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4229 3840
rect 3913 3775 4229 3776
rect 9847 3840 10163 3841
rect 9847 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10163 3840
rect 9847 3775 10163 3776
rect 15781 3840 16097 3841
rect 15781 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16097 3840
rect 15781 3775 16097 3776
rect 21715 3840 22031 3841
rect 21715 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22031 3840
rect 21715 3775 22031 3776
rect 9489 3498 9555 3501
rect 19558 3498 19564 3500
rect 9489 3496 19564 3498
rect 9489 3440 9494 3496
rect 9550 3440 19564 3496
rect 9489 3438 19564 3440
rect 9489 3435 9555 3438
rect 19558 3436 19564 3438
rect 19628 3436 19634 3500
rect 6880 3296 7196 3297
rect 6880 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7196 3296
rect 6880 3231 7196 3232
rect 12814 3296 13130 3297
rect 12814 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13130 3296
rect 12814 3231 13130 3232
rect 18748 3296 19064 3297
rect 18748 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19064 3296
rect 18748 3231 19064 3232
rect 24682 3296 24998 3297
rect 24682 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 24998 3296
rect 24682 3231 24998 3232
rect 7373 3090 7439 3093
rect 17902 3090 17908 3092
rect 7373 3088 17908 3090
rect 7373 3032 7378 3088
rect 7434 3032 17908 3088
rect 7373 3030 17908 3032
rect 7373 3027 7439 3030
rect 17902 3028 17908 3030
rect 17972 3028 17978 3092
rect 9630 2894 10426 2954
rect 3913 2752 4229 2753
rect 3913 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4229 2752
rect 3913 2687 4229 2688
rect 1485 2546 1551 2549
rect 9630 2546 9690 2894
rect 9847 2752 10163 2753
rect 9847 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10163 2752
rect 9847 2687 10163 2688
rect 10366 2682 10426 2894
rect 23473 2818 23539 2821
rect 23749 2818 23815 2821
rect 23473 2816 23815 2818
rect 23473 2760 23478 2816
rect 23534 2760 23754 2816
rect 23810 2760 23815 2816
rect 23473 2758 23815 2760
rect 23473 2755 23539 2758
rect 23749 2755 23815 2758
rect 15781 2752 16097 2753
rect 15781 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16097 2752
rect 15781 2687 16097 2688
rect 21715 2752 22031 2753
rect 21715 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22031 2752
rect 21715 2687 22031 2688
rect 15653 2682 15719 2685
rect 10366 2680 15719 2682
rect 10366 2624 15658 2680
rect 15714 2624 15719 2680
rect 10366 2622 15719 2624
rect 15653 2619 15719 2622
rect 1485 2544 9690 2546
rect 1485 2488 1490 2544
rect 1546 2488 9690 2544
rect 1485 2486 9690 2488
rect 9857 2546 9923 2549
rect 12433 2546 12499 2549
rect 20621 2546 20687 2549
rect 22829 2546 22895 2549
rect 9857 2544 12499 2546
rect 9857 2488 9862 2544
rect 9918 2488 12438 2544
rect 12494 2488 12499 2544
rect 9857 2486 12499 2488
rect 1485 2483 1551 2486
rect 9857 2483 9923 2486
rect 12433 2483 12499 2486
rect 12574 2486 15578 2546
rect 6545 2410 6611 2413
rect 12574 2410 12634 2486
rect 6545 2408 12634 2410
rect 6545 2352 6550 2408
rect 6606 2352 12634 2408
rect 6545 2350 12634 2352
rect 15518 2410 15578 2486
rect 20621 2544 22895 2546
rect 20621 2488 20626 2544
rect 20682 2488 22834 2544
rect 22890 2488 22895 2544
rect 20621 2486 22895 2488
rect 20621 2483 20687 2486
rect 22829 2483 22895 2486
rect 21725 2410 21791 2413
rect 15518 2408 21791 2410
rect 15518 2352 21730 2408
rect 21786 2352 21791 2408
rect 15518 2350 21791 2352
rect 6545 2347 6611 2350
rect 21725 2347 21791 2350
rect 8109 2274 8175 2277
rect 12341 2274 12407 2277
rect 8109 2272 12407 2274
rect 8109 2216 8114 2272
rect 8170 2216 12346 2272
rect 12402 2216 12407 2272
rect 8109 2214 12407 2216
rect 8109 2211 8175 2214
rect 12341 2211 12407 2214
rect 6880 2208 7196 2209
rect 6880 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7196 2208
rect 6880 2143 7196 2144
rect 12814 2208 13130 2209
rect 12814 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13130 2208
rect 12814 2143 13130 2144
rect 18748 2208 19064 2209
rect 18748 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19064 2208
rect 18748 2143 19064 2144
rect 24682 2208 24998 2209
rect 24682 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 24998 2208
rect 24682 2143 24998 2144
rect 8937 2138 9003 2141
rect 10961 2138 11027 2141
rect 8937 2136 11027 2138
rect 8937 2080 8942 2136
rect 8998 2080 10966 2136
rect 11022 2080 11027 2136
rect 8937 2078 11027 2080
rect 8937 2075 9003 2078
rect 10961 2075 11027 2078
rect 6821 2002 6887 2005
rect 13629 2002 13695 2005
rect 6821 2000 13695 2002
rect 6821 1944 6826 2000
rect 6882 1944 13634 2000
rect 13690 1944 13695 2000
rect 6821 1942 13695 1944
rect 6821 1939 6887 1942
rect 13629 1939 13695 1942
rect 6637 1866 6703 1869
rect 19977 1866 20043 1869
rect 6637 1864 20043 1866
rect 6637 1808 6642 1864
rect 6698 1808 19982 1864
rect 20038 1808 20043 1864
rect 6637 1806 20043 1808
rect 6637 1803 6703 1806
rect 19977 1803 20043 1806
rect 9029 1730 9095 1733
rect 9673 1730 9739 1733
rect 9029 1728 9739 1730
rect 9029 1672 9034 1728
rect 9090 1672 9678 1728
rect 9734 1672 9739 1728
rect 9029 1670 9739 1672
rect 9029 1667 9095 1670
rect 9673 1667 9739 1670
rect 12341 1730 12407 1733
rect 15285 1730 15351 1733
rect 12341 1728 15351 1730
rect 12341 1672 12346 1728
rect 12402 1672 15290 1728
rect 15346 1672 15351 1728
rect 12341 1670 15351 1672
rect 12341 1667 12407 1670
rect 15285 1667 15351 1670
rect 18965 1730 19031 1733
rect 19333 1730 19399 1733
rect 18965 1728 19399 1730
rect 18965 1672 18970 1728
rect 19026 1672 19338 1728
rect 19394 1672 19399 1728
rect 18965 1670 19399 1672
rect 18965 1667 19031 1670
rect 19333 1667 19399 1670
rect 3913 1664 4229 1665
rect 3913 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4229 1664
rect 3913 1599 4229 1600
rect 9847 1664 10163 1665
rect 9847 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10163 1664
rect 9847 1599 10163 1600
rect 15781 1664 16097 1665
rect 15781 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16097 1664
rect 15781 1599 16097 1600
rect 21715 1664 22031 1665
rect 21715 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22031 1664
rect 21715 1599 22031 1600
rect 12433 1594 12499 1597
rect 12433 1592 13002 1594
rect 12433 1536 12438 1592
rect 12494 1536 13002 1592
rect 12433 1534 13002 1536
rect 12433 1531 12499 1534
rect 4153 1458 4219 1461
rect 12801 1458 12867 1461
rect 4153 1456 12867 1458
rect 4153 1400 4158 1456
rect 4214 1400 12806 1456
rect 12862 1400 12867 1456
rect 4153 1398 12867 1400
rect 12942 1458 13002 1534
rect 16297 1458 16363 1461
rect 12942 1456 16363 1458
rect 12942 1400 16302 1456
rect 16358 1400 16363 1456
rect 12942 1398 16363 1400
rect 4153 1395 4219 1398
rect 12801 1395 12867 1398
rect 16297 1395 16363 1398
rect 6913 1322 6979 1325
rect 7925 1322 7991 1325
rect 6913 1320 7991 1322
rect 6913 1264 6918 1320
rect 6974 1264 7930 1320
rect 7986 1264 7991 1320
rect 6913 1262 7991 1264
rect 6913 1259 6979 1262
rect 7925 1259 7991 1262
rect 17953 1322 18019 1325
rect 18597 1322 18663 1325
rect 17953 1320 18663 1322
rect 17953 1264 17958 1320
rect 18014 1264 18602 1320
rect 18658 1264 18663 1320
rect 17953 1262 18663 1264
rect 17953 1259 18019 1262
rect 18597 1259 18663 1262
rect 7557 1186 7623 1189
rect 12525 1186 12591 1189
rect 7557 1184 12591 1186
rect 7557 1128 7562 1184
rect 7618 1128 12530 1184
rect 12586 1128 12591 1184
rect 7557 1126 12591 1128
rect 7557 1123 7623 1126
rect 12525 1123 12591 1126
rect 19742 1124 19748 1188
rect 19812 1186 19818 1188
rect 23105 1186 23171 1189
rect 19812 1184 23171 1186
rect 19812 1128 23110 1184
rect 23166 1128 23171 1184
rect 19812 1126 23171 1128
rect 19812 1124 19818 1126
rect 23105 1123 23171 1126
rect 6880 1120 7196 1121
rect 6880 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7196 1120
rect 6880 1055 7196 1056
rect 12814 1120 13130 1121
rect 12814 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13130 1120
rect 12814 1055 13130 1056
rect 18748 1120 19064 1121
rect 18748 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19064 1120
rect 18748 1055 19064 1056
rect 24682 1120 24998 1121
rect 24682 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 24998 1120
rect 24682 1055 24998 1056
rect 19558 988 19564 1052
rect 19628 1050 19634 1052
rect 23473 1050 23539 1053
rect 19628 1048 23539 1050
rect 19628 992 23478 1048
rect 23534 992 23539 1048
rect 19628 990 23539 992
rect 19628 988 19634 990
rect 23473 987 23539 990
rect 5349 914 5415 917
rect 22277 914 22343 917
rect 5349 912 22343 914
rect 5349 856 5354 912
rect 5410 856 22282 912
rect 22338 856 22343 912
rect 5349 854 22343 856
rect 5349 851 5415 854
rect 22277 851 22343 854
rect 5809 778 5875 781
rect 17953 778 18019 781
rect 5809 776 18019 778
rect 5809 720 5814 776
rect 5870 720 17958 776
rect 18014 720 18019 776
rect 5809 718 18019 720
rect 5809 715 5875 718
rect 17953 715 18019 718
rect 6545 640 6611 645
rect 6545 584 6550 640
rect 6606 584 6611 640
rect 6545 579 6611 584
rect 9213 642 9279 645
rect 16205 642 16271 645
rect 9213 640 16271 642
rect 9213 584 9218 640
rect 9274 584 16210 640
rect 16266 584 16271 640
rect 9213 582 16271 584
rect 9213 579 9279 582
rect 16205 579 16271 582
rect 17902 580 17908 644
rect 17972 642 17978 644
rect 20805 642 20871 645
rect 17972 640 20871 642
rect 17972 584 20810 640
rect 20866 584 20871 640
rect 17972 582 20871 584
rect 17972 580 17978 582
rect 20805 579 20871 582
rect 6548 506 6608 579
rect 8937 506 9003 509
rect 21357 506 21423 509
rect 6548 446 8172 506
rect 7557 370 7623 373
rect 2730 368 7623 370
rect 2730 312 7562 368
rect 7618 312 7623 368
rect 2730 310 7623 312
rect 8112 370 8172 446
rect 8937 504 21423 506
rect 8937 448 8942 504
rect 8998 448 21362 504
rect 21418 448 21423 504
rect 8937 446 21423 448
rect 8937 443 9003 446
rect 21357 443 21423 446
rect 17125 370 17191 373
rect 8112 368 17191 370
rect 8112 312 17130 368
rect 17186 312 17191 368
rect 8112 310 17191 312
rect 1669 234 1735 237
rect 2730 234 2790 310
rect 7557 307 7623 310
rect 17125 307 17191 310
rect 1669 232 2790 234
rect 1669 176 1674 232
rect 1730 176 2790 232
rect 1669 174 2790 176
rect 6729 234 6795 237
rect 12709 234 12775 237
rect 6729 232 12775 234
rect 6729 176 6734 232
rect 6790 176 12714 232
rect 12770 176 12775 232
rect 6729 174 12775 176
rect 1669 171 1735 174
rect 6729 171 6795 174
rect 12709 171 12775 174
<< via3 >>
rect 6886 8732 6950 8736
rect 6886 8676 6890 8732
rect 6890 8676 6946 8732
rect 6946 8676 6950 8732
rect 6886 8672 6950 8676
rect 6966 8732 7030 8736
rect 6966 8676 6970 8732
rect 6970 8676 7026 8732
rect 7026 8676 7030 8732
rect 6966 8672 7030 8676
rect 7046 8732 7110 8736
rect 7046 8676 7050 8732
rect 7050 8676 7106 8732
rect 7106 8676 7110 8732
rect 7046 8672 7110 8676
rect 7126 8732 7190 8736
rect 7126 8676 7130 8732
rect 7130 8676 7186 8732
rect 7186 8676 7190 8732
rect 7126 8672 7190 8676
rect 12820 8732 12884 8736
rect 12820 8676 12824 8732
rect 12824 8676 12880 8732
rect 12880 8676 12884 8732
rect 12820 8672 12884 8676
rect 12900 8732 12964 8736
rect 12900 8676 12904 8732
rect 12904 8676 12960 8732
rect 12960 8676 12964 8732
rect 12900 8672 12964 8676
rect 12980 8732 13044 8736
rect 12980 8676 12984 8732
rect 12984 8676 13040 8732
rect 13040 8676 13044 8732
rect 12980 8672 13044 8676
rect 13060 8732 13124 8736
rect 13060 8676 13064 8732
rect 13064 8676 13120 8732
rect 13120 8676 13124 8732
rect 13060 8672 13124 8676
rect 18754 8732 18818 8736
rect 18754 8676 18758 8732
rect 18758 8676 18814 8732
rect 18814 8676 18818 8732
rect 18754 8672 18818 8676
rect 18834 8732 18898 8736
rect 18834 8676 18838 8732
rect 18838 8676 18894 8732
rect 18894 8676 18898 8732
rect 18834 8672 18898 8676
rect 18914 8732 18978 8736
rect 18914 8676 18918 8732
rect 18918 8676 18974 8732
rect 18974 8676 18978 8732
rect 18914 8672 18978 8676
rect 18994 8732 19058 8736
rect 18994 8676 18998 8732
rect 18998 8676 19054 8732
rect 19054 8676 19058 8732
rect 18994 8672 19058 8676
rect 24688 8732 24752 8736
rect 24688 8676 24692 8732
rect 24692 8676 24748 8732
rect 24748 8676 24752 8732
rect 24688 8672 24752 8676
rect 24768 8732 24832 8736
rect 24768 8676 24772 8732
rect 24772 8676 24828 8732
rect 24828 8676 24832 8732
rect 24768 8672 24832 8676
rect 24848 8732 24912 8736
rect 24848 8676 24852 8732
rect 24852 8676 24908 8732
rect 24908 8676 24912 8732
rect 24848 8672 24912 8676
rect 24928 8732 24992 8736
rect 24928 8676 24932 8732
rect 24932 8676 24988 8732
rect 24988 8676 24992 8732
rect 24928 8672 24992 8676
rect 3919 8188 3983 8192
rect 3919 8132 3923 8188
rect 3923 8132 3979 8188
rect 3979 8132 3983 8188
rect 3919 8128 3983 8132
rect 3999 8188 4063 8192
rect 3999 8132 4003 8188
rect 4003 8132 4059 8188
rect 4059 8132 4063 8188
rect 3999 8128 4063 8132
rect 4079 8188 4143 8192
rect 4079 8132 4083 8188
rect 4083 8132 4139 8188
rect 4139 8132 4143 8188
rect 4079 8128 4143 8132
rect 4159 8188 4223 8192
rect 4159 8132 4163 8188
rect 4163 8132 4219 8188
rect 4219 8132 4223 8188
rect 4159 8128 4223 8132
rect 9853 8188 9917 8192
rect 9853 8132 9857 8188
rect 9857 8132 9913 8188
rect 9913 8132 9917 8188
rect 9853 8128 9917 8132
rect 9933 8188 9997 8192
rect 9933 8132 9937 8188
rect 9937 8132 9993 8188
rect 9993 8132 9997 8188
rect 9933 8128 9997 8132
rect 10013 8188 10077 8192
rect 10013 8132 10017 8188
rect 10017 8132 10073 8188
rect 10073 8132 10077 8188
rect 10013 8128 10077 8132
rect 10093 8188 10157 8192
rect 10093 8132 10097 8188
rect 10097 8132 10153 8188
rect 10153 8132 10157 8188
rect 10093 8128 10157 8132
rect 15787 8188 15851 8192
rect 15787 8132 15791 8188
rect 15791 8132 15847 8188
rect 15847 8132 15851 8188
rect 15787 8128 15851 8132
rect 15867 8188 15931 8192
rect 15867 8132 15871 8188
rect 15871 8132 15927 8188
rect 15927 8132 15931 8188
rect 15867 8128 15931 8132
rect 15947 8188 16011 8192
rect 15947 8132 15951 8188
rect 15951 8132 16007 8188
rect 16007 8132 16011 8188
rect 15947 8128 16011 8132
rect 16027 8188 16091 8192
rect 16027 8132 16031 8188
rect 16031 8132 16087 8188
rect 16087 8132 16091 8188
rect 16027 8128 16091 8132
rect 21721 8188 21785 8192
rect 21721 8132 21725 8188
rect 21725 8132 21781 8188
rect 21781 8132 21785 8188
rect 21721 8128 21785 8132
rect 21801 8188 21865 8192
rect 21801 8132 21805 8188
rect 21805 8132 21861 8188
rect 21861 8132 21865 8188
rect 21801 8128 21865 8132
rect 21881 8188 21945 8192
rect 21881 8132 21885 8188
rect 21885 8132 21941 8188
rect 21941 8132 21945 8188
rect 21881 8128 21945 8132
rect 21961 8188 22025 8192
rect 21961 8132 21965 8188
rect 21965 8132 22021 8188
rect 22021 8132 22025 8188
rect 21961 8128 22025 8132
rect 6886 7644 6950 7648
rect 6886 7588 6890 7644
rect 6890 7588 6946 7644
rect 6946 7588 6950 7644
rect 6886 7584 6950 7588
rect 6966 7644 7030 7648
rect 6966 7588 6970 7644
rect 6970 7588 7026 7644
rect 7026 7588 7030 7644
rect 6966 7584 7030 7588
rect 7046 7644 7110 7648
rect 7046 7588 7050 7644
rect 7050 7588 7106 7644
rect 7106 7588 7110 7644
rect 7046 7584 7110 7588
rect 7126 7644 7190 7648
rect 7126 7588 7130 7644
rect 7130 7588 7186 7644
rect 7186 7588 7190 7644
rect 7126 7584 7190 7588
rect 12820 7644 12884 7648
rect 12820 7588 12824 7644
rect 12824 7588 12880 7644
rect 12880 7588 12884 7644
rect 12820 7584 12884 7588
rect 12900 7644 12964 7648
rect 12900 7588 12904 7644
rect 12904 7588 12960 7644
rect 12960 7588 12964 7644
rect 12900 7584 12964 7588
rect 12980 7644 13044 7648
rect 12980 7588 12984 7644
rect 12984 7588 13040 7644
rect 13040 7588 13044 7644
rect 12980 7584 13044 7588
rect 13060 7644 13124 7648
rect 13060 7588 13064 7644
rect 13064 7588 13120 7644
rect 13120 7588 13124 7644
rect 13060 7584 13124 7588
rect 18754 7644 18818 7648
rect 18754 7588 18758 7644
rect 18758 7588 18814 7644
rect 18814 7588 18818 7644
rect 18754 7584 18818 7588
rect 18834 7644 18898 7648
rect 18834 7588 18838 7644
rect 18838 7588 18894 7644
rect 18894 7588 18898 7644
rect 18834 7584 18898 7588
rect 18914 7644 18978 7648
rect 18914 7588 18918 7644
rect 18918 7588 18974 7644
rect 18974 7588 18978 7644
rect 18914 7584 18978 7588
rect 18994 7644 19058 7648
rect 18994 7588 18998 7644
rect 18998 7588 19054 7644
rect 19054 7588 19058 7644
rect 18994 7584 19058 7588
rect 24688 7644 24752 7648
rect 24688 7588 24692 7644
rect 24692 7588 24748 7644
rect 24748 7588 24752 7644
rect 24688 7584 24752 7588
rect 24768 7644 24832 7648
rect 24768 7588 24772 7644
rect 24772 7588 24828 7644
rect 24828 7588 24832 7644
rect 24768 7584 24832 7588
rect 24848 7644 24912 7648
rect 24848 7588 24852 7644
rect 24852 7588 24908 7644
rect 24908 7588 24912 7644
rect 24848 7584 24912 7588
rect 24928 7644 24992 7648
rect 24928 7588 24932 7644
rect 24932 7588 24988 7644
rect 24988 7588 24992 7644
rect 24928 7584 24992 7588
rect 3919 7100 3983 7104
rect 3919 7044 3923 7100
rect 3923 7044 3979 7100
rect 3979 7044 3983 7100
rect 3919 7040 3983 7044
rect 3999 7100 4063 7104
rect 3999 7044 4003 7100
rect 4003 7044 4059 7100
rect 4059 7044 4063 7100
rect 3999 7040 4063 7044
rect 4079 7100 4143 7104
rect 4079 7044 4083 7100
rect 4083 7044 4139 7100
rect 4139 7044 4143 7100
rect 4079 7040 4143 7044
rect 4159 7100 4223 7104
rect 4159 7044 4163 7100
rect 4163 7044 4219 7100
rect 4219 7044 4223 7100
rect 4159 7040 4223 7044
rect 9853 7100 9917 7104
rect 9853 7044 9857 7100
rect 9857 7044 9913 7100
rect 9913 7044 9917 7100
rect 9853 7040 9917 7044
rect 9933 7100 9997 7104
rect 9933 7044 9937 7100
rect 9937 7044 9993 7100
rect 9993 7044 9997 7100
rect 9933 7040 9997 7044
rect 10013 7100 10077 7104
rect 10013 7044 10017 7100
rect 10017 7044 10073 7100
rect 10073 7044 10077 7100
rect 10013 7040 10077 7044
rect 10093 7100 10157 7104
rect 10093 7044 10097 7100
rect 10097 7044 10153 7100
rect 10153 7044 10157 7100
rect 10093 7040 10157 7044
rect 15787 7100 15851 7104
rect 15787 7044 15791 7100
rect 15791 7044 15847 7100
rect 15847 7044 15851 7100
rect 15787 7040 15851 7044
rect 15867 7100 15931 7104
rect 15867 7044 15871 7100
rect 15871 7044 15927 7100
rect 15927 7044 15931 7100
rect 15867 7040 15931 7044
rect 15947 7100 16011 7104
rect 15947 7044 15951 7100
rect 15951 7044 16007 7100
rect 16007 7044 16011 7100
rect 15947 7040 16011 7044
rect 16027 7100 16091 7104
rect 16027 7044 16031 7100
rect 16031 7044 16087 7100
rect 16087 7044 16091 7100
rect 16027 7040 16091 7044
rect 21721 7100 21785 7104
rect 21721 7044 21725 7100
rect 21725 7044 21781 7100
rect 21781 7044 21785 7100
rect 21721 7040 21785 7044
rect 21801 7100 21865 7104
rect 21801 7044 21805 7100
rect 21805 7044 21861 7100
rect 21861 7044 21865 7100
rect 21801 7040 21865 7044
rect 21881 7100 21945 7104
rect 21881 7044 21885 7100
rect 21885 7044 21941 7100
rect 21941 7044 21945 7100
rect 21881 7040 21945 7044
rect 21961 7100 22025 7104
rect 21961 7044 21965 7100
rect 21965 7044 22021 7100
rect 22021 7044 22025 7100
rect 21961 7040 22025 7044
rect 6886 6556 6950 6560
rect 6886 6500 6890 6556
rect 6890 6500 6946 6556
rect 6946 6500 6950 6556
rect 6886 6496 6950 6500
rect 6966 6556 7030 6560
rect 6966 6500 6970 6556
rect 6970 6500 7026 6556
rect 7026 6500 7030 6556
rect 6966 6496 7030 6500
rect 7046 6556 7110 6560
rect 7046 6500 7050 6556
rect 7050 6500 7106 6556
rect 7106 6500 7110 6556
rect 7046 6496 7110 6500
rect 7126 6556 7190 6560
rect 7126 6500 7130 6556
rect 7130 6500 7186 6556
rect 7186 6500 7190 6556
rect 7126 6496 7190 6500
rect 12820 6556 12884 6560
rect 12820 6500 12824 6556
rect 12824 6500 12880 6556
rect 12880 6500 12884 6556
rect 12820 6496 12884 6500
rect 12900 6556 12964 6560
rect 12900 6500 12904 6556
rect 12904 6500 12960 6556
rect 12960 6500 12964 6556
rect 12900 6496 12964 6500
rect 12980 6556 13044 6560
rect 12980 6500 12984 6556
rect 12984 6500 13040 6556
rect 13040 6500 13044 6556
rect 12980 6496 13044 6500
rect 13060 6556 13124 6560
rect 13060 6500 13064 6556
rect 13064 6500 13120 6556
rect 13120 6500 13124 6556
rect 13060 6496 13124 6500
rect 18754 6556 18818 6560
rect 18754 6500 18758 6556
rect 18758 6500 18814 6556
rect 18814 6500 18818 6556
rect 18754 6496 18818 6500
rect 18834 6556 18898 6560
rect 18834 6500 18838 6556
rect 18838 6500 18894 6556
rect 18894 6500 18898 6556
rect 18834 6496 18898 6500
rect 18914 6556 18978 6560
rect 18914 6500 18918 6556
rect 18918 6500 18974 6556
rect 18974 6500 18978 6556
rect 18914 6496 18978 6500
rect 18994 6556 19058 6560
rect 18994 6500 18998 6556
rect 18998 6500 19054 6556
rect 19054 6500 19058 6556
rect 18994 6496 19058 6500
rect 24688 6556 24752 6560
rect 24688 6500 24692 6556
rect 24692 6500 24748 6556
rect 24748 6500 24752 6556
rect 24688 6496 24752 6500
rect 24768 6556 24832 6560
rect 24768 6500 24772 6556
rect 24772 6500 24828 6556
rect 24828 6500 24832 6556
rect 24768 6496 24832 6500
rect 24848 6556 24912 6560
rect 24848 6500 24852 6556
rect 24852 6500 24908 6556
rect 24908 6500 24912 6556
rect 24848 6496 24912 6500
rect 24928 6556 24992 6560
rect 24928 6500 24932 6556
rect 24932 6500 24988 6556
rect 24988 6500 24992 6556
rect 24928 6496 24992 6500
rect 19748 6156 19812 6220
rect 3919 6012 3983 6016
rect 3919 5956 3923 6012
rect 3923 5956 3979 6012
rect 3979 5956 3983 6012
rect 3919 5952 3983 5956
rect 3999 6012 4063 6016
rect 3999 5956 4003 6012
rect 4003 5956 4059 6012
rect 4059 5956 4063 6012
rect 3999 5952 4063 5956
rect 4079 6012 4143 6016
rect 4079 5956 4083 6012
rect 4083 5956 4139 6012
rect 4139 5956 4143 6012
rect 4079 5952 4143 5956
rect 4159 6012 4223 6016
rect 4159 5956 4163 6012
rect 4163 5956 4219 6012
rect 4219 5956 4223 6012
rect 4159 5952 4223 5956
rect 9853 6012 9917 6016
rect 9853 5956 9857 6012
rect 9857 5956 9913 6012
rect 9913 5956 9917 6012
rect 9853 5952 9917 5956
rect 9933 6012 9997 6016
rect 9933 5956 9937 6012
rect 9937 5956 9993 6012
rect 9993 5956 9997 6012
rect 9933 5952 9997 5956
rect 10013 6012 10077 6016
rect 10013 5956 10017 6012
rect 10017 5956 10073 6012
rect 10073 5956 10077 6012
rect 10013 5952 10077 5956
rect 10093 6012 10157 6016
rect 10093 5956 10097 6012
rect 10097 5956 10153 6012
rect 10153 5956 10157 6012
rect 10093 5952 10157 5956
rect 15787 6012 15851 6016
rect 15787 5956 15791 6012
rect 15791 5956 15847 6012
rect 15847 5956 15851 6012
rect 15787 5952 15851 5956
rect 15867 6012 15931 6016
rect 15867 5956 15871 6012
rect 15871 5956 15927 6012
rect 15927 5956 15931 6012
rect 15867 5952 15931 5956
rect 15947 6012 16011 6016
rect 15947 5956 15951 6012
rect 15951 5956 16007 6012
rect 16007 5956 16011 6012
rect 15947 5952 16011 5956
rect 16027 6012 16091 6016
rect 16027 5956 16031 6012
rect 16031 5956 16087 6012
rect 16087 5956 16091 6012
rect 16027 5952 16091 5956
rect 21721 6012 21785 6016
rect 21721 5956 21725 6012
rect 21725 5956 21781 6012
rect 21781 5956 21785 6012
rect 21721 5952 21785 5956
rect 21801 6012 21865 6016
rect 21801 5956 21805 6012
rect 21805 5956 21861 6012
rect 21861 5956 21865 6012
rect 21801 5952 21865 5956
rect 21881 6012 21945 6016
rect 21881 5956 21885 6012
rect 21885 5956 21941 6012
rect 21941 5956 21945 6012
rect 21881 5952 21945 5956
rect 21961 6012 22025 6016
rect 21961 5956 21965 6012
rect 21965 5956 22021 6012
rect 22021 5956 22025 6012
rect 21961 5952 22025 5956
rect 6886 5468 6950 5472
rect 6886 5412 6890 5468
rect 6890 5412 6946 5468
rect 6946 5412 6950 5468
rect 6886 5408 6950 5412
rect 6966 5468 7030 5472
rect 6966 5412 6970 5468
rect 6970 5412 7026 5468
rect 7026 5412 7030 5468
rect 6966 5408 7030 5412
rect 7046 5468 7110 5472
rect 7046 5412 7050 5468
rect 7050 5412 7106 5468
rect 7106 5412 7110 5468
rect 7046 5408 7110 5412
rect 7126 5468 7190 5472
rect 7126 5412 7130 5468
rect 7130 5412 7186 5468
rect 7186 5412 7190 5468
rect 7126 5408 7190 5412
rect 12820 5468 12884 5472
rect 12820 5412 12824 5468
rect 12824 5412 12880 5468
rect 12880 5412 12884 5468
rect 12820 5408 12884 5412
rect 12900 5468 12964 5472
rect 12900 5412 12904 5468
rect 12904 5412 12960 5468
rect 12960 5412 12964 5468
rect 12900 5408 12964 5412
rect 12980 5468 13044 5472
rect 12980 5412 12984 5468
rect 12984 5412 13040 5468
rect 13040 5412 13044 5468
rect 12980 5408 13044 5412
rect 13060 5468 13124 5472
rect 13060 5412 13064 5468
rect 13064 5412 13120 5468
rect 13120 5412 13124 5468
rect 13060 5408 13124 5412
rect 18754 5468 18818 5472
rect 18754 5412 18758 5468
rect 18758 5412 18814 5468
rect 18814 5412 18818 5468
rect 18754 5408 18818 5412
rect 18834 5468 18898 5472
rect 18834 5412 18838 5468
rect 18838 5412 18894 5468
rect 18894 5412 18898 5468
rect 18834 5408 18898 5412
rect 18914 5468 18978 5472
rect 18914 5412 18918 5468
rect 18918 5412 18974 5468
rect 18974 5412 18978 5468
rect 18914 5408 18978 5412
rect 18994 5468 19058 5472
rect 18994 5412 18998 5468
rect 18998 5412 19054 5468
rect 19054 5412 19058 5468
rect 18994 5408 19058 5412
rect 24688 5468 24752 5472
rect 24688 5412 24692 5468
rect 24692 5412 24748 5468
rect 24748 5412 24752 5468
rect 24688 5408 24752 5412
rect 24768 5468 24832 5472
rect 24768 5412 24772 5468
rect 24772 5412 24828 5468
rect 24828 5412 24832 5468
rect 24768 5408 24832 5412
rect 24848 5468 24912 5472
rect 24848 5412 24852 5468
rect 24852 5412 24908 5468
rect 24908 5412 24912 5468
rect 24848 5408 24912 5412
rect 24928 5468 24992 5472
rect 24928 5412 24932 5468
rect 24932 5412 24988 5468
rect 24988 5412 24992 5468
rect 24928 5408 24992 5412
rect 3919 4924 3983 4928
rect 3919 4868 3923 4924
rect 3923 4868 3979 4924
rect 3979 4868 3983 4924
rect 3919 4864 3983 4868
rect 3999 4924 4063 4928
rect 3999 4868 4003 4924
rect 4003 4868 4059 4924
rect 4059 4868 4063 4924
rect 3999 4864 4063 4868
rect 4079 4924 4143 4928
rect 4079 4868 4083 4924
rect 4083 4868 4139 4924
rect 4139 4868 4143 4924
rect 4079 4864 4143 4868
rect 4159 4924 4223 4928
rect 4159 4868 4163 4924
rect 4163 4868 4219 4924
rect 4219 4868 4223 4924
rect 4159 4864 4223 4868
rect 9853 4924 9917 4928
rect 9853 4868 9857 4924
rect 9857 4868 9913 4924
rect 9913 4868 9917 4924
rect 9853 4864 9917 4868
rect 9933 4924 9997 4928
rect 9933 4868 9937 4924
rect 9937 4868 9993 4924
rect 9993 4868 9997 4924
rect 9933 4864 9997 4868
rect 10013 4924 10077 4928
rect 10013 4868 10017 4924
rect 10017 4868 10073 4924
rect 10073 4868 10077 4924
rect 10013 4864 10077 4868
rect 10093 4924 10157 4928
rect 10093 4868 10097 4924
rect 10097 4868 10153 4924
rect 10153 4868 10157 4924
rect 10093 4864 10157 4868
rect 15787 4924 15851 4928
rect 15787 4868 15791 4924
rect 15791 4868 15847 4924
rect 15847 4868 15851 4924
rect 15787 4864 15851 4868
rect 15867 4924 15931 4928
rect 15867 4868 15871 4924
rect 15871 4868 15927 4924
rect 15927 4868 15931 4924
rect 15867 4864 15931 4868
rect 15947 4924 16011 4928
rect 15947 4868 15951 4924
rect 15951 4868 16007 4924
rect 16007 4868 16011 4924
rect 15947 4864 16011 4868
rect 16027 4924 16091 4928
rect 16027 4868 16031 4924
rect 16031 4868 16087 4924
rect 16087 4868 16091 4924
rect 16027 4864 16091 4868
rect 21721 4924 21785 4928
rect 21721 4868 21725 4924
rect 21725 4868 21781 4924
rect 21781 4868 21785 4924
rect 21721 4864 21785 4868
rect 21801 4924 21865 4928
rect 21801 4868 21805 4924
rect 21805 4868 21861 4924
rect 21861 4868 21865 4924
rect 21801 4864 21865 4868
rect 21881 4924 21945 4928
rect 21881 4868 21885 4924
rect 21885 4868 21941 4924
rect 21941 4868 21945 4924
rect 21881 4864 21945 4868
rect 21961 4924 22025 4928
rect 21961 4868 21965 4924
rect 21965 4868 22021 4924
rect 22021 4868 22025 4924
rect 21961 4864 22025 4868
rect 6886 4380 6950 4384
rect 6886 4324 6890 4380
rect 6890 4324 6946 4380
rect 6946 4324 6950 4380
rect 6886 4320 6950 4324
rect 6966 4380 7030 4384
rect 6966 4324 6970 4380
rect 6970 4324 7026 4380
rect 7026 4324 7030 4380
rect 6966 4320 7030 4324
rect 7046 4380 7110 4384
rect 7046 4324 7050 4380
rect 7050 4324 7106 4380
rect 7106 4324 7110 4380
rect 7046 4320 7110 4324
rect 7126 4380 7190 4384
rect 7126 4324 7130 4380
rect 7130 4324 7186 4380
rect 7186 4324 7190 4380
rect 7126 4320 7190 4324
rect 12820 4380 12884 4384
rect 12820 4324 12824 4380
rect 12824 4324 12880 4380
rect 12880 4324 12884 4380
rect 12820 4320 12884 4324
rect 12900 4380 12964 4384
rect 12900 4324 12904 4380
rect 12904 4324 12960 4380
rect 12960 4324 12964 4380
rect 12900 4320 12964 4324
rect 12980 4380 13044 4384
rect 12980 4324 12984 4380
rect 12984 4324 13040 4380
rect 13040 4324 13044 4380
rect 12980 4320 13044 4324
rect 13060 4380 13124 4384
rect 13060 4324 13064 4380
rect 13064 4324 13120 4380
rect 13120 4324 13124 4380
rect 13060 4320 13124 4324
rect 18754 4380 18818 4384
rect 18754 4324 18758 4380
rect 18758 4324 18814 4380
rect 18814 4324 18818 4380
rect 18754 4320 18818 4324
rect 18834 4380 18898 4384
rect 18834 4324 18838 4380
rect 18838 4324 18894 4380
rect 18894 4324 18898 4380
rect 18834 4320 18898 4324
rect 18914 4380 18978 4384
rect 18914 4324 18918 4380
rect 18918 4324 18974 4380
rect 18974 4324 18978 4380
rect 18914 4320 18978 4324
rect 18994 4380 19058 4384
rect 18994 4324 18998 4380
rect 18998 4324 19054 4380
rect 19054 4324 19058 4380
rect 18994 4320 19058 4324
rect 24688 4380 24752 4384
rect 24688 4324 24692 4380
rect 24692 4324 24748 4380
rect 24748 4324 24752 4380
rect 24688 4320 24752 4324
rect 24768 4380 24832 4384
rect 24768 4324 24772 4380
rect 24772 4324 24828 4380
rect 24828 4324 24832 4380
rect 24768 4320 24832 4324
rect 24848 4380 24912 4384
rect 24848 4324 24852 4380
rect 24852 4324 24908 4380
rect 24908 4324 24912 4380
rect 24848 4320 24912 4324
rect 24928 4380 24992 4384
rect 24928 4324 24932 4380
rect 24932 4324 24988 4380
rect 24988 4324 24992 4380
rect 24928 4320 24992 4324
rect 3919 3836 3983 3840
rect 3919 3780 3923 3836
rect 3923 3780 3979 3836
rect 3979 3780 3983 3836
rect 3919 3776 3983 3780
rect 3999 3836 4063 3840
rect 3999 3780 4003 3836
rect 4003 3780 4059 3836
rect 4059 3780 4063 3836
rect 3999 3776 4063 3780
rect 4079 3836 4143 3840
rect 4079 3780 4083 3836
rect 4083 3780 4139 3836
rect 4139 3780 4143 3836
rect 4079 3776 4143 3780
rect 4159 3836 4223 3840
rect 4159 3780 4163 3836
rect 4163 3780 4219 3836
rect 4219 3780 4223 3836
rect 4159 3776 4223 3780
rect 9853 3836 9917 3840
rect 9853 3780 9857 3836
rect 9857 3780 9913 3836
rect 9913 3780 9917 3836
rect 9853 3776 9917 3780
rect 9933 3836 9997 3840
rect 9933 3780 9937 3836
rect 9937 3780 9993 3836
rect 9993 3780 9997 3836
rect 9933 3776 9997 3780
rect 10013 3836 10077 3840
rect 10013 3780 10017 3836
rect 10017 3780 10073 3836
rect 10073 3780 10077 3836
rect 10013 3776 10077 3780
rect 10093 3836 10157 3840
rect 10093 3780 10097 3836
rect 10097 3780 10153 3836
rect 10153 3780 10157 3836
rect 10093 3776 10157 3780
rect 15787 3836 15851 3840
rect 15787 3780 15791 3836
rect 15791 3780 15847 3836
rect 15847 3780 15851 3836
rect 15787 3776 15851 3780
rect 15867 3836 15931 3840
rect 15867 3780 15871 3836
rect 15871 3780 15927 3836
rect 15927 3780 15931 3836
rect 15867 3776 15931 3780
rect 15947 3836 16011 3840
rect 15947 3780 15951 3836
rect 15951 3780 16007 3836
rect 16007 3780 16011 3836
rect 15947 3776 16011 3780
rect 16027 3836 16091 3840
rect 16027 3780 16031 3836
rect 16031 3780 16087 3836
rect 16087 3780 16091 3836
rect 16027 3776 16091 3780
rect 21721 3836 21785 3840
rect 21721 3780 21725 3836
rect 21725 3780 21781 3836
rect 21781 3780 21785 3836
rect 21721 3776 21785 3780
rect 21801 3836 21865 3840
rect 21801 3780 21805 3836
rect 21805 3780 21861 3836
rect 21861 3780 21865 3836
rect 21801 3776 21865 3780
rect 21881 3836 21945 3840
rect 21881 3780 21885 3836
rect 21885 3780 21941 3836
rect 21941 3780 21945 3836
rect 21881 3776 21945 3780
rect 21961 3836 22025 3840
rect 21961 3780 21965 3836
rect 21965 3780 22021 3836
rect 22021 3780 22025 3836
rect 21961 3776 22025 3780
rect 19564 3436 19628 3500
rect 6886 3292 6950 3296
rect 6886 3236 6890 3292
rect 6890 3236 6946 3292
rect 6946 3236 6950 3292
rect 6886 3232 6950 3236
rect 6966 3292 7030 3296
rect 6966 3236 6970 3292
rect 6970 3236 7026 3292
rect 7026 3236 7030 3292
rect 6966 3232 7030 3236
rect 7046 3292 7110 3296
rect 7046 3236 7050 3292
rect 7050 3236 7106 3292
rect 7106 3236 7110 3292
rect 7046 3232 7110 3236
rect 7126 3292 7190 3296
rect 7126 3236 7130 3292
rect 7130 3236 7186 3292
rect 7186 3236 7190 3292
rect 7126 3232 7190 3236
rect 12820 3292 12884 3296
rect 12820 3236 12824 3292
rect 12824 3236 12880 3292
rect 12880 3236 12884 3292
rect 12820 3232 12884 3236
rect 12900 3292 12964 3296
rect 12900 3236 12904 3292
rect 12904 3236 12960 3292
rect 12960 3236 12964 3292
rect 12900 3232 12964 3236
rect 12980 3292 13044 3296
rect 12980 3236 12984 3292
rect 12984 3236 13040 3292
rect 13040 3236 13044 3292
rect 12980 3232 13044 3236
rect 13060 3292 13124 3296
rect 13060 3236 13064 3292
rect 13064 3236 13120 3292
rect 13120 3236 13124 3292
rect 13060 3232 13124 3236
rect 18754 3292 18818 3296
rect 18754 3236 18758 3292
rect 18758 3236 18814 3292
rect 18814 3236 18818 3292
rect 18754 3232 18818 3236
rect 18834 3292 18898 3296
rect 18834 3236 18838 3292
rect 18838 3236 18894 3292
rect 18894 3236 18898 3292
rect 18834 3232 18898 3236
rect 18914 3292 18978 3296
rect 18914 3236 18918 3292
rect 18918 3236 18974 3292
rect 18974 3236 18978 3292
rect 18914 3232 18978 3236
rect 18994 3292 19058 3296
rect 18994 3236 18998 3292
rect 18998 3236 19054 3292
rect 19054 3236 19058 3292
rect 18994 3232 19058 3236
rect 24688 3292 24752 3296
rect 24688 3236 24692 3292
rect 24692 3236 24748 3292
rect 24748 3236 24752 3292
rect 24688 3232 24752 3236
rect 24768 3292 24832 3296
rect 24768 3236 24772 3292
rect 24772 3236 24828 3292
rect 24828 3236 24832 3292
rect 24768 3232 24832 3236
rect 24848 3292 24912 3296
rect 24848 3236 24852 3292
rect 24852 3236 24908 3292
rect 24908 3236 24912 3292
rect 24848 3232 24912 3236
rect 24928 3292 24992 3296
rect 24928 3236 24932 3292
rect 24932 3236 24988 3292
rect 24988 3236 24992 3292
rect 24928 3232 24992 3236
rect 17908 3028 17972 3092
rect 3919 2748 3983 2752
rect 3919 2692 3923 2748
rect 3923 2692 3979 2748
rect 3979 2692 3983 2748
rect 3919 2688 3983 2692
rect 3999 2748 4063 2752
rect 3999 2692 4003 2748
rect 4003 2692 4059 2748
rect 4059 2692 4063 2748
rect 3999 2688 4063 2692
rect 4079 2748 4143 2752
rect 4079 2692 4083 2748
rect 4083 2692 4139 2748
rect 4139 2692 4143 2748
rect 4079 2688 4143 2692
rect 4159 2748 4223 2752
rect 4159 2692 4163 2748
rect 4163 2692 4219 2748
rect 4219 2692 4223 2748
rect 4159 2688 4223 2692
rect 9853 2748 9917 2752
rect 9853 2692 9857 2748
rect 9857 2692 9913 2748
rect 9913 2692 9917 2748
rect 9853 2688 9917 2692
rect 9933 2748 9997 2752
rect 9933 2692 9937 2748
rect 9937 2692 9993 2748
rect 9993 2692 9997 2748
rect 9933 2688 9997 2692
rect 10013 2748 10077 2752
rect 10013 2692 10017 2748
rect 10017 2692 10073 2748
rect 10073 2692 10077 2748
rect 10013 2688 10077 2692
rect 10093 2748 10157 2752
rect 10093 2692 10097 2748
rect 10097 2692 10153 2748
rect 10153 2692 10157 2748
rect 10093 2688 10157 2692
rect 15787 2748 15851 2752
rect 15787 2692 15791 2748
rect 15791 2692 15847 2748
rect 15847 2692 15851 2748
rect 15787 2688 15851 2692
rect 15867 2748 15931 2752
rect 15867 2692 15871 2748
rect 15871 2692 15927 2748
rect 15927 2692 15931 2748
rect 15867 2688 15931 2692
rect 15947 2748 16011 2752
rect 15947 2692 15951 2748
rect 15951 2692 16007 2748
rect 16007 2692 16011 2748
rect 15947 2688 16011 2692
rect 16027 2748 16091 2752
rect 16027 2692 16031 2748
rect 16031 2692 16087 2748
rect 16087 2692 16091 2748
rect 16027 2688 16091 2692
rect 21721 2748 21785 2752
rect 21721 2692 21725 2748
rect 21725 2692 21781 2748
rect 21781 2692 21785 2748
rect 21721 2688 21785 2692
rect 21801 2748 21865 2752
rect 21801 2692 21805 2748
rect 21805 2692 21861 2748
rect 21861 2692 21865 2748
rect 21801 2688 21865 2692
rect 21881 2748 21945 2752
rect 21881 2692 21885 2748
rect 21885 2692 21941 2748
rect 21941 2692 21945 2748
rect 21881 2688 21945 2692
rect 21961 2748 22025 2752
rect 21961 2692 21965 2748
rect 21965 2692 22021 2748
rect 22021 2692 22025 2748
rect 21961 2688 22025 2692
rect 6886 2204 6950 2208
rect 6886 2148 6890 2204
rect 6890 2148 6946 2204
rect 6946 2148 6950 2204
rect 6886 2144 6950 2148
rect 6966 2204 7030 2208
rect 6966 2148 6970 2204
rect 6970 2148 7026 2204
rect 7026 2148 7030 2204
rect 6966 2144 7030 2148
rect 7046 2204 7110 2208
rect 7046 2148 7050 2204
rect 7050 2148 7106 2204
rect 7106 2148 7110 2204
rect 7046 2144 7110 2148
rect 7126 2204 7190 2208
rect 7126 2148 7130 2204
rect 7130 2148 7186 2204
rect 7186 2148 7190 2204
rect 7126 2144 7190 2148
rect 12820 2204 12884 2208
rect 12820 2148 12824 2204
rect 12824 2148 12880 2204
rect 12880 2148 12884 2204
rect 12820 2144 12884 2148
rect 12900 2204 12964 2208
rect 12900 2148 12904 2204
rect 12904 2148 12960 2204
rect 12960 2148 12964 2204
rect 12900 2144 12964 2148
rect 12980 2204 13044 2208
rect 12980 2148 12984 2204
rect 12984 2148 13040 2204
rect 13040 2148 13044 2204
rect 12980 2144 13044 2148
rect 13060 2204 13124 2208
rect 13060 2148 13064 2204
rect 13064 2148 13120 2204
rect 13120 2148 13124 2204
rect 13060 2144 13124 2148
rect 18754 2204 18818 2208
rect 18754 2148 18758 2204
rect 18758 2148 18814 2204
rect 18814 2148 18818 2204
rect 18754 2144 18818 2148
rect 18834 2204 18898 2208
rect 18834 2148 18838 2204
rect 18838 2148 18894 2204
rect 18894 2148 18898 2204
rect 18834 2144 18898 2148
rect 18914 2204 18978 2208
rect 18914 2148 18918 2204
rect 18918 2148 18974 2204
rect 18974 2148 18978 2204
rect 18914 2144 18978 2148
rect 18994 2204 19058 2208
rect 18994 2148 18998 2204
rect 18998 2148 19054 2204
rect 19054 2148 19058 2204
rect 18994 2144 19058 2148
rect 24688 2204 24752 2208
rect 24688 2148 24692 2204
rect 24692 2148 24748 2204
rect 24748 2148 24752 2204
rect 24688 2144 24752 2148
rect 24768 2204 24832 2208
rect 24768 2148 24772 2204
rect 24772 2148 24828 2204
rect 24828 2148 24832 2204
rect 24768 2144 24832 2148
rect 24848 2204 24912 2208
rect 24848 2148 24852 2204
rect 24852 2148 24908 2204
rect 24908 2148 24912 2204
rect 24848 2144 24912 2148
rect 24928 2204 24992 2208
rect 24928 2148 24932 2204
rect 24932 2148 24988 2204
rect 24988 2148 24992 2204
rect 24928 2144 24992 2148
rect 3919 1660 3983 1664
rect 3919 1604 3923 1660
rect 3923 1604 3979 1660
rect 3979 1604 3983 1660
rect 3919 1600 3983 1604
rect 3999 1660 4063 1664
rect 3999 1604 4003 1660
rect 4003 1604 4059 1660
rect 4059 1604 4063 1660
rect 3999 1600 4063 1604
rect 4079 1660 4143 1664
rect 4079 1604 4083 1660
rect 4083 1604 4139 1660
rect 4139 1604 4143 1660
rect 4079 1600 4143 1604
rect 4159 1660 4223 1664
rect 4159 1604 4163 1660
rect 4163 1604 4219 1660
rect 4219 1604 4223 1660
rect 4159 1600 4223 1604
rect 9853 1660 9917 1664
rect 9853 1604 9857 1660
rect 9857 1604 9913 1660
rect 9913 1604 9917 1660
rect 9853 1600 9917 1604
rect 9933 1660 9997 1664
rect 9933 1604 9937 1660
rect 9937 1604 9993 1660
rect 9993 1604 9997 1660
rect 9933 1600 9997 1604
rect 10013 1660 10077 1664
rect 10013 1604 10017 1660
rect 10017 1604 10073 1660
rect 10073 1604 10077 1660
rect 10013 1600 10077 1604
rect 10093 1660 10157 1664
rect 10093 1604 10097 1660
rect 10097 1604 10153 1660
rect 10153 1604 10157 1660
rect 10093 1600 10157 1604
rect 15787 1660 15851 1664
rect 15787 1604 15791 1660
rect 15791 1604 15847 1660
rect 15847 1604 15851 1660
rect 15787 1600 15851 1604
rect 15867 1660 15931 1664
rect 15867 1604 15871 1660
rect 15871 1604 15927 1660
rect 15927 1604 15931 1660
rect 15867 1600 15931 1604
rect 15947 1660 16011 1664
rect 15947 1604 15951 1660
rect 15951 1604 16007 1660
rect 16007 1604 16011 1660
rect 15947 1600 16011 1604
rect 16027 1660 16091 1664
rect 16027 1604 16031 1660
rect 16031 1604 16087 1660
rect 16087 1604 16091 1660
rect 16027 1600 16091 1604
rect 21721 1660 21785 1664
rect 21721 1604 21725 1660
rect 21725 1604 21781 1660
rect 21781 1604 21785 1660
rect 21721 1600 21785 1604
rect 21801 1660 21865 1664
rect 21801 1604 21805 1660
rect 21805 1604 21861 1660
rect 21861 1604 21865 1660
rect 21801 1600 21865 1604
rect 21881 1660 21945 1664
rect 21881 1604 21885 1660
rect 21885 1604 21941 1660
rect 21941 1604 21945 1660
rect 21881 1600 21945 1604
rect 21961 1660 22025 1664
rect 21961 1604 21965 1660
rect 21965 1604 22021 1660
rect 22021 1604 22025 1660
rect 21961 1600 22025 1604
rect 19748 1124 19812 1188
rect 6886 1116 6950 1120
rect 6886 1060 6890 1116
rect 6890 1060 6946 1116
rect 6946 1060 6950 1116
rect 6886 1056 6950 1060
rect 6966 1116 7030 1120
rect 6966 1060 6970 1116
rect 6970 1060 7026 1116
rect 7026 1060 7030 1116
rect 6966 1056 7030 1060
rect 7046 1116 7110 1120
rect 7046 1060 7050 1116
rect 7050 1060 7106 1116
rect 7106 1060 7110 1116
rect 7046 1056 7110 1060
rect 7126 1116 7190 1120
rect 7126 1060 7130 1116
rect 7130 1060 7186 1116
rect 7186 1060 7190 1116
rect 7126 1056 7190 1060
rect 12820 1116 12884 1120
rect 12820 1060 12824 1116
rect 12824 1060 12880 1116
rect 12880 1060 12884 1116
rect 12820 1056 12884 1060
rect 12900 1116 12964 1120
rect 12900 1060 12904 1116
rect 12904 1060 12960 1116
rect 12960 1060 12964 1116
rect 12900 1056 12964 1060
rect 12980 1116 13044 1120
rect 12980 1060 12984 1116
rect 12984 1060 13040 1116
rect 13040 1060 13044 1116
rect 12980 1056 13044 1060
rect 13060 1116 13124 1120
rect 13060 1060 13064 1116
rect 13064 1060 13120 1116
rect 13120 1060 13124 1116
rect 13060 1056 13124 1060
rect 18754 1116 18818 1120
rect 18754 1060 18758 1116
rect 18758 1060 18814 1116
rect 18814 1060 18818 1116
rect 18754 1056 18818 1060
rect 18834 1116 18898 1120
rect 18834 1060 18838 1116
rect 18838 1060 18894 1116
rect 18894 1060 18898 1116
rect 18834 1056 18898 1060
rect 18914 1116 18978 1120
rect 18914 1060 18918 1116
rect 18918 1060 18974 1116
rect 18974 1060 18978 1116
rect 18914 1056 18978 1060
rect 18994 1116 19058 1120
rect 18994 1060 18998 1116
rect 18998 1060 19054 1116
rect 19054 1060 19058 1116
rect 18994 1056 19058 1060
rect 24688 1116 24752 1120
rect 24688 1060 24692 1116
rect 24692 1060 24748 1116
rect 24748 1060 24752 1116
rect 24688 1056 24752 1060
rect 24768 1116 24832 1120
rect 24768 1060 24772 1116
rect 24772 1060 24828 1116
rect 24828 1060 24832 1116
rect 24768 1056 24832 1060
rect 24848 1116 24912 1120
rect 24848 1060 24852 1116
rect 24852 1060 24908 1116
rect 24908 1060 24912 1116
rect 24848 1056 24912 1060
rect 24928 1116 24992 1120
rect 24928 1060 24932 1116
rect 24932 1060 24988 1116
rect 24988 1060 24992 1116
rect 24928 1056 24992 1060
rect 19564 988 19628 1052
rect 17908 580 17972 644
<< metal4 >>
rect 3911 8192 4231 8752
rect 3911 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4231 8192
rect 3911 7104 4231 8128
rect 3911 7040 3919 7104
rect 3983 7040 3999 7104
rect 4063 7040 4079 7104
rect 4143 7040 4159 7104
rect 4223 7040 4231 7104
rect 3911 6016 4231 7040
rect 3911 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4231 6016
rect 3911 4928 4231 5952
rect 3911 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4231 4928
rect 3911 3840 4231 4864
rect 3911 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4231 3840
rect 3911 2752 4231 3776
rect 3911 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4231 2752
rect 3911 1664 4231 2688
rect 3911 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4231 1664
rect 3911 1040 4231 1600
rect 6878 8736 7198 8752
rect 6878 8672 6886 8736
rect 6950 8672 6966 8736
rect 7030 8672 7046 8736
rect 7110 8672 7126 8736
rect 7190 8672 7198 8736
rect 6878 7648 7198 8672
rect 6878 7584 6886 7648
rect 6950 7584 6966 7648
rect 7030 7584 7046 7648
rect 7110 7584 7126 7648
rect 7190 7584 7198 7648
rect 6878 6560 7198 7584
rect 6878 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7198 6560
rect 6878 5472 7198 6496
rect 6878 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7198 5472
rect 6878 4384 7198 5408
rect 6878 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7198 4384
rect 6878 3296 7198 4320
rect 6878 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7198 3296
rect 6878 2208 7198 3232
rect 6878 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7198 2208
rect 6878 1120 7198 2144
rect 6878 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7198 1120
rect 6878 1040 7198 1056
rect 9845 8192 10165 8752
rect 9845 8128 9853 8192
rect 9917 8128 9933 8192
rect 9997 8128 10013 8192
rect 10077 8128 10093 8192
rect 10157 8128 10165 8192
rect 9845 7104 10165 8128
rect 9845 7040 9853 7104
rect 9917 7040 9933 7104
rect 9997 7040 10013 7104
rect 10077 7040 10093 7104
rect 10157 7040 10165 7104
rect 9845 6016 10165 7040
rect 9845 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10165 6016
rect 9845 4928 10165 5952
rect 9845 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10165 4928
rect 9845 3840 10165 4864
rect 9845 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10165 3840
rect 9845 2752 10165 3776
rect 9845 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10165 2752
rect 9845 1664 10165 2688
rect 9845 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10165 1664
rect 9845 1040 10165 1600
rect 12812 8736 13132 8752
rect 12812 8672 12820 8736
rect 12884 8672 12900 8736
rect 12964 8672 12980 8736
rect 13044 8672 13060 8736
rect 13124 8672 13132 8736
rect 12812 7648 13132 8672
rect 12812 7584 12820 7648
rect 12884 7584 12900 7648
rect 12964 7584 12980 7648
rect 13044 7584 13060 7648
rect 13124 7584 13132 7648
rect 12812 6560 13132 7584
rect 12812 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13132 6560
rect 12812 5472 13132 6496
rect 12812 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13132 5472
rect 12812 4384 13132 5408
rect 12812 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13132 4384
rect 12812 3296 13132 4320
rect 12812 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13132 3296
rect 12812 2208 13132 3232
rect 12812 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13132 2208
rect 12812 1120 13132 2144
rect 12812 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13132 1120
rect 12812 1040 13132 1056
rect 15779 8192 16099 8752
rect 15779 8128 15787 8192
rect 15851 8128 15867 8192
rect 15931 8128 15947 8192
rect 16011 8128 16027 8192
rect 16091 8128 16099 8192
rect 15779 7104 16099 8128
rect 15779 7040 15787 7104
rect 15851 7040 15867 7104
rect 15931 7040 15947 7104
rect 16011 7040 16027 7104
rect 16091 7040 16099 7104
rect 15779 6016 16099 7040
rect 15779 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16099 6016
rect 15779 4928 16099 5952
rect 15779 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16099 4928
rect 15779 3840 16099 4864
rect 15779 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16099 3840
rect 15779 2752 16099 3776
rect 18746 8736 19066 8752
rect 18746 8672 18754 8736
rect 18818 8672 18834 8736
rect 18898 8672 18914 8736
rect 18978 8672 18994 8736
rect 19058 8672 19066 8736
rect 18746 7648 19066 8672
rect 18746 7584 18754 7648
rect 18818 7584 18834 7648
rect 18898 7584 18914 7648
rect 18978 7584 18994 7648
rect 19058 7584 19066 7648
rect 18746 6560 19066 7584
rect 18746 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19066 6560
rect 18746 5472 19066 6496
rect 21713 8192 22033 8752
rect 21713 8128 21721 8192
rect 21785 8128 21801 8192
rect 21865 8128 21881 8192
rect 21945 8128 21961 8192
rect 22025 8128 22033 8192
rect 21713 7104 22033 8128
rect 21713 7040 21721 7104
rect 21785 7040 21801 7104
rect 21865 7040 21881 7104
rect 21945 7040 21961 7104
rect 22025 7040 22033 7104
rect 19747 6220 19813 6221
rect 19747 6156 19748 6220
rect 19812 6156 19813 6220
rect 19747 6155 19813 6156
rect 18746 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19066 5472
rect 18746 4384 19066 5408
rect 18746 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19066 4384
rect 18746 3296 19066 4320
rect 19563 3500 19629 3501
rect 19563 3436 19564 3500
rect 19628 3436 19629 3500
rect 19563 3435 19629 3436
rect 18746 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19066 3296
rect 17907 3092 17973 3093
rect 17907 3028 17908 3092
rect 17972 3028 17973 3092
rect 17907 3027 17973 3028
rect 15779 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16099 2752
rect 15779 1664 16099 2688
rect 15779 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16099 1664
rect 15779 1040 16099 1600
rect 17910 645 17970 3027
rect 18746 2208 19066 3232
rect 18746 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19066 2208
rect 18746 1120 19066 2144
rect 18746 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19066 1120
rect 18746 1040 19066 1056
rect 19566 1053 19626 3435
rect 19750 1189 19810 6155
rect 21713 6016 22033 7040
rect 21713 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22033 6016
rect 21713 4928 22033 5952
rect 21713 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22033 4928
rect 21713 3840 22033 4864
rect 21713 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22033 3840
rect 21713 2752 22033 3776
rect 21713 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22033 2752
rect 21713 1664 22033 2688
rect 21713 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22033 1664
rect 19747 1188 19813 1189
rect 19747 1124 19748 1188
rect 19812 1124 19813 1188
rect 19747 1123 19813 1124
rect 19563 1052 19629 1053
rect 19563 988 19564 1052
rect 19628 988 19629 1052
rect 21713 1040 22033 1600
rect 24680 8736 25000 8752
rect 24680 8672 24688 8736
rect 24752 8672 24768 8736
rect 24832 8672 24848 8736
rect 24912 8672 24928 8736
rect 24992 8672 25000 8736
rect 24680 7648 25000 8672
rect 24680 7584 24688 7648
rect 24752 7584 24768 7648
rect 24832 7584 24848 7648
rect 24912 7584 24928 7648
rect 24992 7584 25000 7648
rect 24680 6560 25000 7584
rect 24680 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 25000 6560
rect 24680 5472 25000 6496
rect 24680 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 25000 5472
rect 24680 4384 25000 5408
rect 24680 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 25000 4384
rect 24680 3296 25000 4320
rect 24680 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 25000 3296
rect 24680 2208 25000 3232
rect 24680 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 25000 2208
rect 24680 1120 25000 2144
rect 24680 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 25000 1120
rect 24680 1040 25000 1056
rect 19563 987 19629 988
rect 17907 644 17973 645
rect 17907 580 17908 644
rect 17972 580 17973 644
rect 17907 579 17973 580
use sky130_fd_sc_hd__clkbuf_1  _00_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _01_
timestamp 1688980957
transform 1 0 9752 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _02_
timestamp 1688980957
transform 1 0 1840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _03_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _04_
timestamp 1688980957
transform 1 0 2300 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _05_
timestamp 1688980957
transform 1 0 6624 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp 1688980957
transform 1 0 7544 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1688980957
transform 1 0 13800 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1688980957
transform 1 0 14076 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _11_
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1688980957
transform 1 0 7176 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1688980957
transform 1 0 5428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1688980957
transform 1 0 5980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1688980957
transform 1 0 4968 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _17_
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1688980957
transform 1 0 4232 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1688980957
transform 1 0 2576 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1688980957
transform 1 0 16284 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1688980957
transform 1 0 11224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1688980957
transform 1 0 10028 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1688980957
transform 1 0 17112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1688980957
transform 1 0 17664 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1688980957
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1688980957
transform 1 0 18400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1688980957
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1688980957
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1688980957
transform 1 0 22080 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _36_
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _37_
timestamp 1688980957
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _38_
timestamp 1688980957
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1688980957
transform 1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1688980957
transform 1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1688980957
transform 1 0 9476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1688980957
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1688980957
transform 1 0 11868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1688980957
transform 1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1688980957
transform 1 0 14444 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1688980957
transform 1 0 17204 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1688980957
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _51_
timestamp 1688980957
transform 1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1688980957
transform 1 0 22172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1688980957
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1688980957
transform 1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1688980957
transform 1 0 24104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 21068 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_126
timestamp 1688980957
transform 1 0 12696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_136 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13616 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_151
timestamp 1688980957
transform 1 0 14996 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_215
timestamp 1688980957
transform 1 0 20884 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_219
timestamp 1688980957
transform 1 0 21252 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_14
timestamp 1688980957
transform 1 0 2392 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_40
timestamp 1688980957
transform 1 0 4784 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_45
timestamp 1688980957
transform 1 0 5244 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_132
timestamp 1688980957
transform 1 0 13248 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_213
timestamp 1688980957
transform 1 0 20700 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 1688980957
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_48
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_56
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_60 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_72
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_96
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_104
timestamp 1688980957
transform 1 0 10672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_108
timestamp 1688980957
transform 1 0 11040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_119 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_128
timestamp 1688980957
transform 1 0 12880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_135
timestamp 1688980957
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_149
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_156
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_160
timestamp 1688980957
transform 1 0 15824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_194
timestamp 1688980957
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_212
timestamp 1688980957
transform 1 0 20608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 1688980957
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_212
timestamp 1688980957
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_231
timestamp 1688980957
transform 1 0 22356 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_253
timestamp 1688980957
transform 1 0 24380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_88
timestamp 1688980957
transform 1 0 9200 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_92
timestamp 1688980957
transform 1 0 9568 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_100
timestamp 1688980957
transform 1 0 10304 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_112
timestamp 1688980957
transform 1 0 11408 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_124
timestamp 1688980957
transform 1 0 12512 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_136
timestamp 1688980957
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_205
timestamp 1688980957
transform 1 0 19964 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_239
timestamp 1688980957
transform 1 0 23092 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_77
timestamp 1688980957
transform 1 0 8188 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_85
timestamp 1688980957
transform 1 0 8924 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_94
timestamp 1688980957
transform 1 0 9752 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_106
timestamp 1688980957
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_253
timestamp 1688980957
transform 1 0 24380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_117 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_123
timestamp 1688980957
transform 1 0 12420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_135
timestamp 1688980957
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_206
timestamp 1688980957
transform 1 0 20056 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_218
timestamp 1688980957
transform 1 0 21160 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_230
timestamp 1688980957
transform 1 0 22264 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_242
timestamp 1688980957
transform 1 0 23368 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_250
timestamp 1688980957
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_123
timestamp 1688980957
transform 1 0 12420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_135
timestamp 1688980957
transform 1 0 13524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_153
timestamp 1688980957
transform 1 0 15180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1688980957
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_202
timestamp 1688980957
transform 1 0 19688 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_214
timestamp 1688980957
transform 1 0 20792 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 1688980957
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_148
timestamp 1688980957
transform 1 0 14720 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_160
timestamp 1688980957
transform 1 0 15824 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_172
timestamp 1688980957
transform 1 0 16928 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_184
timestamp 1688980957
transform 1 0 18032 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_200
timestamp 1688980957
transform 1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_207
timestamp 1688980957
transform 1 0 20148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_219
timestamp 1688980957
transform 1 0 21252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_231
timestamp 1688980957
transform 1 0 22356 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_243
timestamp 1688980957
transform 1 0 23460 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_60
timestamp 1688980957
transform 1 0 6624 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_64
timestamp 1688980957
transform 1 0 6992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_71
timestamp 1688980957
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_75
timestamp 1688980957
transform 1 0 8004 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_87
timestamp 1688980957
transform 1 0 9108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_99
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_252
timestamp 1688980957
transform 1 0 24288 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_57
timestamp 1688980957
transform 1 0 6348 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_70
timestamp 1688980957
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_105
timestamp 1688980957
transform 1 0 10764 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_112
timestamp 1688980957
transform 1 0 11408 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_124
timestamp 1688980957
transform 1 0 12512 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_132
timestamp 1688980957
transform 1 0 13248 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_171
timestamp 1688980957
transform 1 0 16836 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_178
timestamp 1688980957
transform 1 0 17480 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_190
timestamp 1688980957
transform 1 0 18584 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_241
timestamp 1688980957
transform 1 0 23276 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_16
timestamp 1688980957
transform 1 0 2576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_37
timestamp 1688980957
transform 1 0 4508 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_42
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_50
timestamp 1688980957
transform 1 0 5704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_60
timestamp 1688980957
transform 1 0 6624 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_71
timestamp 1688980957
transform 1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_89
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_94
timestamp 1688980957
transform 1 0 9752 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_102
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1688980957
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_120
timestamp 1688980957
transform 1 0 12144 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_128
timestamp 1688980957
transform 1 0 12880 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_136
timestamp 1688980957
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_146
timestamp 1688980957
transform 1 0 14536 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_152
timestamp 1688980957
transform 1 0 15088 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_159
timestamp 1688980957
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_178
timestamp 1688980957
transform 1 0 17480 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_185
timestamp 1688980957
transform 1 0 18124 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_203
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_211
timestamp 1688980957
transform 1 0 20516 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_219
timestamp 1688980957
transform 1 0 21252 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_240
timestamp 1688980957
transform 1 0 23184 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_250
timestamp 1688980957
transform 1 0 24104 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_253
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 22356 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 22724 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 24012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 23552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 22724 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 23276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 23736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 22356 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 22632 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 22908 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 22908 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 23460 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 23736 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 22448 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 3404 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 3680 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 3128 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 3956 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 4324 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 1564 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 1472 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 1748 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 2576 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 2852 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 4600 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 8372 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 8924 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 5704 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1688980957
transform 1 0 6440 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform 1 0 5704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1688980957
transform 1 0 6716 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 7268 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1688980957
transform 1 0 6900 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 8096 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 22080 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._00_
timestamp 1688980957
transform 1 0 8648 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._01_
timestamp 1688980957
transform 1 0 9200 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._02_
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._03_
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._04_
timestamp 1688980957
transform 1 0 2024 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._05_
timestamp 1688980957
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._06_
timestamp 1688980957
transform 1 0 6992 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._07_
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._08_
timestamp 1688980957
transform 1 0 13248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._09_
timestamp 1688980957
transform 1 0 13432 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._10_
timestamp 1688980957
transform 1 0 12420 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._11_
timestamp 1688980957
transform 1 0 15456 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._12_
timestamp 1688980957
transform 1 0 7820 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._13_
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_RAM_IO_switch_matrix._14_
timestamp 1688980957
transform 1 0 4048 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._15_
timestamp 1688980957
transform 1 0 5428 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._16_
timestamp 1688980957
transform 1 0 4508 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._17_
timestamp 1688980957
transform 1 0 3404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._18_
timestamp 1688980957
transform 1 0 2852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._19_
timestamp 1688980957
transform 1 0 3128 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._20_
timestamp 1688980957
transform 1 0 9292 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._21_
timestamp 1688980957
transform 1 0 9016 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._22_
timestamp 1688980957
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._23_
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._24_
timestamp 1688980957
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._25_
timestamp 1688980957
transform 1 0 21436 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_RAM_IO_switch_matrix._26_
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._27_
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._28_
timestamp 1688980957
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._29_
timestamp 1688980957
transform 1 0 9476 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_RAM_IO_switch_matrix._30_
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._31_
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._32_
timestamp 1688980957
transform 1 0 17388 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._33_
timestamp 1688980957
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._34_
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._35_
timestamp 1688980957
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output58 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1688980957
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output60 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output62
timestamp 1688980957
transform 1 0 17572 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output63
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1688980957
transform 1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1688980957
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1688980957
transform 1 0 22540 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1688980957
transform 1 0 23736 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output68
timestamp 1688980957
transform 1 0 23736 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1688980957
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1688980957
transform 1 0 6808 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1688980957
transform 1 0 10580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1688980957
transform 1 0 11776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1688980957
transform 1 0 12972 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1688980957
transform 1 0 9568 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 10304 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1688980957
transform 1 0 9936 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 10856 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1688980957
transform 1 0 13248 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1688980957
transform 1 0 14628 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1688980957
transform 1 0 14444 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1688980957
transform 1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 10672 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1688980957
transform 1 0 10304 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 11868 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 12144 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 12696 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform 1 0 11776 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 15732 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 19596 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 20332 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output101
timestamp 1688980957
transform 1 0 19044 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 20148 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1688980957
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 20884 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 16836 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 19780 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 17940 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 18492 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 24840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 24840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 24840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 24840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 24840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 24840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 24840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 24840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0._0_
timestamp 1688980957
transform 1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1._0_
timestamp 1688980957
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2._0_
timestamp 1688980957
transform 1 0 21344 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3._0_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4._0_
timestamp 1688980957
transform 1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5._0_
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6._0_
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7._0_
timestamp 1688980957
transform 1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8._0_
timestamp 1688980957
transform 1 0 12144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9._0_
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10._0_
timestamp 1688980957
transform 1 0 14904 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11._0_
timestamp 1688980957
transform 1 0 23000 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12._0_
timestamp 1688980957
transform 1 0 16928 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13._0_
timestamp 1688980957
transform 1 0 24288 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14._0_
timestamp 1688980957
transform 1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15._0_
timestamp 1688980957
transform 1 0 23184 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16._0_
timestamp 1688980957
transform 1 0 23184 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17._0_
timestamp 1688980957
transform 1 0 23736 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18._0_
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19._0_
timestamp 1688980957
transform 1 0 24104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0._0_
timestamp 1688980957
transform 1 0 19412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1._0_
timestamp 1688980957
transform 1 0 20332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_2._0_
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3._0_
timestamp 1688980957
transform 1 0 6072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4._0_
timestamp 1688980957
transform 1 0 7268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5._0_
timestamp 1688980957
transform 1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6._0_
timestamp 1688980957
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7._0_
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8._0_
timestamp 1688980957
transform 1 0 12144 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9._0_
timestamp 1688980957
transform 1 0 13616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10._0_
timestamp 1688980957
transform 1 0 14628 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11._0_
timestamp 1688980957
transform 1 0 22724 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12._0_
timestamp 1688980957
transform 1 0 17204 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13._0_
timestamp 1688980957
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14._0_
timestamp 1688980957
transform 1 0 22448 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15._0_
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16._0_
timestamp 1688980957
transform 1 0 22632 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17._0_
timestamp 1688980957
transform 1 0 23460 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18._0_
timestamp 1688980957
transform 1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19._0_
timestamp 1688980957
transform 1 0 24012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 20350 0 20406 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 23110 0 23166 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 23386 0 23442 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 23662 0 23718 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 23938 0 23994 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 24214 0 24270 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 24490 0 24546 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 24766 0 24822 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 25042 0 25098 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 25318 0 25374 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 25594 0 25650 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 20626 0 20682 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 20902 0 20958 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 21178 0 21234 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 21454 0 21510 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 21730 0 21786 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 22006 0 22062 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 22282 0 22338 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 22558 0 22614 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 22834 0 22890 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 2134 9840 2190 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 14094 9840 14150 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 15290 9840 15346 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 16486 9840 16542 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 17682 9840 17738 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 18878 9840 18934 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 20074 9840 20130 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 21270 9840 21326 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 22466 9840 22522 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 23662 9840 23718 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 24858 9840 24914 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 3330 9840 3386 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 4526 9840 4582 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 5722 9840 5778 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 6918 9840 6974 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 8114 9840 8170 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 9310 9840 9366 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 10506 9840 10562 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 11702 9840 11758 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 12898 9840 12954 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 202 0 258 160 0 FreeSans 224 90 0 0 N1END[0]
port 40 nsew signal input
flabel metal2 s 478 0 534 160 0 FreeSans 224 90 0 0 N1END[1]
port 41 nsew signal input
flabel metal2 s 754 0 810 160 0 FreeSans 224 90 0 0 N1END[2]
port 42 nsew signal input
flabel metal2 s 1030 0 1086 160 0 FreeSans 224 90 0 0 N1END[3]
port 43 nsew signal input
flabel metal2 s 3514 0 3570 160 0 FreeSans 224 90 0 0 N2END[0]
port 44 nsew signal input
flabel metal2 s 3790 0 3846 160 0 FreeSans 224 90 0 0 N2END[1]
port 45 nsew signal input
flabel metal2 s 4066 0 4122 160 0 FreeSans 224 90 0 0 N2END[2]
port 46 nsew signal input
flabel metal2 s 4342 0 4398 160 0 FreeSans 224 90 0 0 N2END[3]
port 47 nsew signal input
flabel metal2 s 4618 0 4674 160 0 FreeSans 224 90 0 0 N2END[4]
port 48 nsew signal input
flabel metal2 s 4894 0 4950 160 0 FreeSans 224 90 0 0 N2END[5]
port 49 nsew signal input
flabel metal2 s 5170 0 5226 160 0 FreeSans 224 90 0 0 N2END[6]
port 50 nsew signal input
flabel metal2 s 5446 0 5502 160 0 FreeSans 224 90 0 0 N2END[7]
port 51 nsew signal input
flabel metal2 s 1306 0 1362 160 0 FreeSans 224 90 0 0 N2MID[0]
port 52 nsew signal input
flabel metal2 s 1582 0 1638 160 0 FreeSans 224 90 0 0 N2MID[1]
port 53 nsew signal input
flabel metal2 s 1858 0 1914 160 0 FreeSans 224 90 0 0 N2MID[2]
port 54 nsew signal input
flabel metal2 s 2134 0 2190 160 0 FreeSans 224 90 0 0 N2MID[3]
port 55 nsew signal input
flabel metal2 s 2410 0 2466 160 0 FreeSans 224 90 0 0 N2MID[4]
port 56 nsew signal input
flabel metal2 s 2686 0 2742 160 0 FreeSans 224 90 0 0 N2MID[5]
port 57 nsew signal input
flabel metal2 s 2962 0 3018 160 0 FreeSans 224 90 0 0 N2MID[6]
port 58 nsew signal input
flabel metal2 s 3238 0 3294 160 0 FreeSans 224 90 0 0 N2MID[7]
port 59 nsew signal input
flabel metal2 s 5722 0 5778 160 0 FreeSans 224 90 0 0 N4END[0]
port 60 nsew signal input
flabel metal2 s 8482 0 8538 160 0 FreeSans 224 90 0 0 N4END[10]
port 61 nsew signal input
flabel metal2 s 8758 0 8814 160 0 FreeSans 224 90 0 0 N4END[11]
port 62 nsew signal input
flabel metal2 s 9034 0 9090 160 0 FreeSans 224 90 0 0 N4END[12]
port 63 nsew signal input
flabel metal2 s 9310 0 9366 160 0 FreeSans 224 90 0 0 N4END[13]
port 64 nsew signal input
flabel metal2 s 9586 0 9642 160 0 FreeSans 224 90 0 0 N4END[14]
port 65 nsew signal input
flabel metal2 s 9862 0 9918 160 0 FreeSans 224 90 0 0 N4END[15]
port 66 nsew signal input
flabel metal2 s 5998 0 6054 160 0 FreeSans 224 90 0 0 N4END[1]
port 67 nsew signal input
flabel metal2 s 6274 0 6330 160 0 FreeSans 224 90 0 0 N4END[2]
port 68 nsew signal input
flabel metal2 s 6550 0 6606 160 0 FreeSans 224 90 0 0 N4END[3]
port 69 nsew signal input
flabel metal2 s 6826 0 6882 160 0 FreeSans 224 90 0 0 N4END[4]
port 70 nsew signal input
flabel metal2 s 7102 0 7158 160 0 FreeSans 224 90 0 0 N4END[5]
port 71 nsew signal input
flabel metal2 s 7378 0 7434 160 0 FreeSans 224 90 0 0 N4END[6]
port 72 nsew signal input
flabel metal2 s 7654 0 7710 160 0 FreeSans 224 90 0 0 N4END[7]
port 73 nsew signal input
flabel metal2 s 7930 0 7986 160 0 FreeSans 224 90 0 0 N4END[8]
port 74 nsew signal input
flabel metal2 s 8206 0 8262 160 0 FreeSans 224 90 0 0 N4END[9]
port 75 nsew signal input
flabel metal2 s 10138 0 10194 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 76 nsew signal tristate
flabel metal2 s 10414 0 10470 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 77 nsew signal tristate
flabel metal2 s 10690 0 10746 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 78 nsew signal tristate
flabel metal2 s 10966 0 11022 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 79 nsew signal tristate
flabel metal2 s 13450 0 13506 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 80 nsew signal tristate
flabel metal2 s 13726 0 13782 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 81 nsew signal tristate
flabel metal2 s 14002 0 14058 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 82 nsew signal tristate
flabel metal2 s 14278 0 14334 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 83 nsew signal tristate
flabel metal2 s 14554 0 14610 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 84 nsew signal tristate
flabel metal2 s 14830 0 14886 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 85 nsew signal tristate
flabel metal2 s 15106 0 15162 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 86 nsew signal tristate
flabel metal2 s 15382 0 15438 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 87 nsew signal tristate
flabel metal2 s 11242 0 11298 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 88 nsew signal tristate
flabel metal2 s 11518 0 11574 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 89 nsew signal tristate
flabel metal2 s 11794 0 11850 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 90 nsew signal tristate
flabel metal2 s 12070 0 12126 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 91 nsew signal tristate
flabel metal2 s 12346 0 12402 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 92 nsew signal tristate
flabel metal2 s 12622 0 12678 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 93 nsew signal tristate
flabel metal2 s 12898 0 12954 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 94 nsew signal tristate
flabel metal2 s 13174 0 13230 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 95 nsew signal tristate
flabel metal2 s 15658 0 15714 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 96 nsew signal tristate
flabel metal2 s 18418 0 18474 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 97 nsew signal tristate
flabel metal2 s 18694 0 18750 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 98 nsew signal tristate
flabel metal2 s 18970 0 19026 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 99 nsew signal tristate
flabel metal2 s 19246 0 19302 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 100 nsew signal tristate
flabel metal2 s 19522 0 19578 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 101 nsew signal tristate
flabel metal2 s 19798 0 19854 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 102 nsew signal tristate
flabel metal2 s 15934 0 15990 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 103 nsew signal tristate
flabel metal2 s 16210 0 16266 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 104 nsew signal tristate
flabel metal2 s 16486 0 16542 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 105 nsew signal tristate
flabel metal2 s 16762 0 16818 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 106 nsew signal tristate
flabel metal2 s 17038 0 17094 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 107 nsew signal tristate
flabel metal2 s 17314 0 17370 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 108 nsew signal tristate
flabel metal2 s 17590 0 17646 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 109 nsew signal tristate
flabel metal2 s 17866 0 17922 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 110 nsew signal tristate
flabel metal2 s 18142 0 18198 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 111 nsew signal tristate
flabel metal2 s 20074 0 20130 160 0 FreeSans 224 90 0 0 UserCLK
port 112 nsew signal input
flabel metal2 s 938 9840 994 10000 0 FreeSans 224 90 0 0 UserCLKo
port 113 nsew signal tristate
flabel metal4 s 6878 1040 7198 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 12812 1040 13132 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 18746 1040 19066 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 24680 1040 25000 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 3911 1040 4231 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 9845 1040 10165 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 15779 1040 16099 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 21713 1040 22033 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
rlabel via1 13052 8704 13052 8704 0 VGND
rlabel metal1 12972 8160 12972 8160 0 VPWR
rlabel metal2 20477 68 20477 68 0 FrameStrobe[0]
rlabel metal2 23039 68 23039 68 0 FrameStrobe[10]
rlabel metal2 23414 432 23414 432 0 FrameStrobe[11]
rlabel metal2 23690 1248 23690 1248 0 FrameStrobe[12]
rlabel metal2 23966 483 23966 483 0 FrameStrobe[13]
rlabel metal2 24242 364 24242 364 0 FrameStrobe[14]
rlabel metal1 24380 3502 24380 3502 0 FrameStrobe[15]
rlabel metal2 24695 68 24695 68 0 FrameStrobe[16]
rlabel metal2 25070 1180 25070 1180 0 FrameStrobe[17]
rlabel metal1 24426 3638 24426 3638 0 FrameStrobe[18]
rlabel metal1 24794 3434 24794 3434 0 FrameStrobe[19]
rlabel metal2 20707 68 20707 68 0 FrameStrobe[1]
rlabel metal2 21029 68 21029 68 0 FrameStrobe[2]
rlabel metal2 21206 262 21206 262 0 FrameStrobe[3]
rlabel metal2 21535 68 21535 68 0 FrameStrobe[4]
rlabel metal2 21857 68 21857 68 0 FrameStrobe[5]
rlabel metal2 22034 364 22034 364 0 FrameStrobe[6]
rlabel metal2 22310 432 22310 432 0 FrameStrobe[7]
rlabel metal2 22586 483 22586 483 0 FrameStrobe[8]
rlabel metal2 22862 1248 22862 1248 0 FrameStrobe[9]
rlabel metal1 2300 8602 2300 8602 0 FrameStrobe_O[0]
rlabel metal1 14260 8602 14260 8602 0 FrameStrobe_O[10]
rlabel metal2 15318 9224 15318 9224 0 FrameStrobe_O[11]
rlabel metal2 16514 9088 16514 9088 0 FrameStrobe_O[12]
rlabel metal2 17710 9224 17710 9224 0 FrameStrobe_O[13]
rlabel metal2 18906 9785 18906 9785 0 FrameStrobe_O[14]
rlabel metal1 20240 8602 20240 8602 0 FrameStrobe_O[15]
rlabel metal1 21436 8602 21436 8602 0 FrameStrobe_O[16]
rlabel metal1 22632 8602 22632 8602 0 FrameStrobe_O[17]
rlabel metal1 23828 8602 23828 8602 0 FrameStrobe_O[18]
rlabel metal1 24334 8058 24334 8058 0 FrameStrobe_O[19]
rlabel metal1 3680 8602 3680 8602 0 FrameStrobe_O[1]
rlabel metal1 4692 8602 4692 8602 0 FrameStrobe_O[2]
rlabel metal1 5888 8602 5888 8602 0 FrameStrobe_O[3]
rlabel metal2 6946 9785 6946 9785 0 FrameStrobe_O[4]
rlabel metal2 8142 9445 8142 9445 0 FrameStrobe_O[5]
rlabel metal1 9476 8602 9476 8602 0 FrameStrobe_O[6]
rlabel metal1 10672 8602 10672 8602 0 FrameStrobe_O[7]
rlabel metal1 11868 8602 11868 8602 0 FrameStrobe_O[8]
rlabel metal2 13202 9231 13202 9231 0 FrameStrobe_O[9]
rlabel metal1 8602 1326 8602 1326 0 Inst_N_term_RAM_IO_switch_matrix.S1BEG0
rlabel metal1 9982 1904 9982 1904 0 Inst_N_term_RAM_IO_switch_matrix.S1BEG1
rlabel metal1 2070 1972 2070 1972 0 Inst_N_term_RAM_IO_switch_matrix.S1BEG2
rlabel metal1 2162 1904 2162 1904 0 Inst_N_term_RAM_IO_switch_matrix.S1BEG3
rlabel metal1 2530 1292 2530 1292 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG0
rlabel metal1 6854 1292 6854 1292 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG1
rlabel metal1 7682 1938 7682 1938 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG2
rlabel metal1 13202 2448 13202 2448 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG3
rlabel metal1 14030 1972 14030 1972 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG4
rlabel metal1 14306 1904 14306 1904 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG5
rlabel metal1 15410 1972 15410 1972 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG6
rlabel metal1 15318 1802 15318 1802 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG7
rlabel metal1 7406 1292 7406 1292 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb0
rlabel metal1 5658 1292 5658 1292 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb1
rlabel metal1 4278 1224 4278 1224 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb2
rlabel metal1 6210 1972 6210 1972 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb3
rlabel metal1 5198 1972 5198 1972 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb4
rlabel metal1 3818 1292 3818 1292 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb5
rlabel metal1 3680 1530 3680 1530 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb6
rlabel metal1 2898 1326 2898 1326 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb7
rlabel metal2 13202 2227 13202 2227 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG0
rlabel metal2 16238 1275 16238 1275 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG1
rlabel metal2 21482 1054 21482 1054 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG10
rlabel metal1 19044 1530 19044 1530 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG11
rlabel metal1 20286 2380 20286 2380 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG12
rlabel metal1 20700 1734 20700 1734 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG13
rlabel metal2 5382 1037 5382 1037 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG14
rlabel metal2 21850 2244 21850 2244 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG15
rlabel metal1 11454 2380 11454 2380 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG2
rlabel metal1 10258 1870 10258 1870 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG3
rlabel metal2 15502 1360 15502 1360 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG4
rlabel metal2 11730 1802 11730 1802 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG5
rlabel metal1 17066 2074 17066 2074 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG6
rlabel metal1 17342 2380 17342 2380 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG7
rlabel metal1 16330 1224 16330 1224 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG8
rlabel metal1 18354 2448 18354 2448 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG9
rlabel metal2 230 1554 230 1554 0 N1END[0]
rlabel metal2 506 1520 506 1520 0 N1END[1]
rlabel metal2 782 1588 782 1588 0 N1END[2]
rlabel metal2 1058 942 1058 942 0 N1END[3]
rlabel metal2 3595 68 3595 68 0 N2END[0]
rlabel metal2 3818 1010 3818 1010 0 N2END[1]
rlabel metal2 4094 398 4094 398 0 N2END[2]
rlabel metal2 4370 1010 4370 1010 0 N2END[3]
rlabel metal2 4646 1248 4646 1248 0 N2END[4]
rlabel metal2 4922 1248 4922 1248 0 N2END[5]
rlabel metal2 5198 636 5198 636 0 N2END[6]
rlabel metal2 5474 398 5474 398 0 N2END[7]
rlabel metal2 1334 1248 1334 1248 0 N2MID[0]
rlabel metal2 1610 755 1610 755 0 N2MID[1]
rlabel metal2 1886 1010 1886 1010 0 N2MID[2]
rlabel metal2 2162 1231 2162 1231 0 N2MID[3]
rlabel metal2 2438 364 2438 364 0 N2MID[4]
rlabel metal2 2714 398 2714 398 0 N2MID[5]
rlabel metal2 2891 68 2891 68 0 N2MID[6]
rlabel metal2 3167 68 3167 68 0 N2MID[7]
rlabel metal2 5750 279 5750 279 0 N4END[0]
rlabel metal2 8510 398 8510 398 0 N4END[10]
rlabel metal2 8786 1010 8786 1010 0 N4END[11]
rlabel metal2 8963 68 8963 68 0 N4END[12]
rlabel metal2 9239 68 9239 68 0 N4END[13]
rlabel metal2 9614 1248 9614 1248 0 N4END[14]
rlabel metal2 9890 398 9890 398 0 N4END[15]
rlabel metal2 5973 68 5973 68 0 N4END[1]
rlabel metal2 6355 68 6355 68 0 N4END[2]
rlabel metal2 6525 68 6525 68 0 N4END[3]
rlabel metal2 6854 364 6854 364 0 N4END[4]
rlabel metal2 7229 68 7229 68 0 N4END[5]
rlabel metal2 7406 398 7406 398 0 N4END[6]
rlabel metal2 7682 1027 7682 1027 0 N4END[7]
rlabel metal2 7958 687 7958 687 0 N4END[8]
rlabel metal2 8234 1010 8234 1010 0 N4END[9]
rlabel metal2 10113 68 10113 68 0 S1BEG[0]
rlabel metal2 10495 68 10495 68 0 S1BEG[1]
rlabel metal2 10718 670 10718 670 0 S1BEG[2]
rlabel metal2 10994 908 10994 908 0 S1BEG[3]
rlabel metal2 13478 636 13478 636 0 S2BEG[0]
rlabel metal2 13754 806 13754 806 0 S2BEG[1]
rlabel metal2 14030 636 14030 636 0 S2BEG[2]
rlabel metal2 14306 908 14306 908 0 S2BEG[3]
rlabel metal2 14681 68 14681 68 0 S2BEG[4]
rlabel metal2 14858 806 14858 806 0 S2BEG[5]
rlabel metal2 15134 738 15134 738 0 S2BEG[6]
rlabel metal2 15410 1180 15410 1180 0 S2BEG[7]
rlabel metal2 11171 68 11171 68 0 S2BEGb[0]
rlabel metal2 11546 347 11546 347 0 S2BEGb[1]
rlabel metal2 11822 908 11822 908 0 S2BEGb[2]
rlabel metal2 11999 68 11999 68 0 S2BEGb[3]
rlabel metal2 12374 636 12374 636 0 S2BEGb[4]
rlabel metal2 12650 908 12650 908 0 S2BEGb[5]
rlabel metal2 12926 364 12926 364 0 S2BEGb[6]
rlabel metal2 13202 636 13202 636 0 S2BEGb[7]
rlabel metal2 15686 908 15686 908 0 S4BEG[0]
rlabel metal2 18499 68 18499 68 0 S4BEG[10]
rlabel metal2 18669 68 18669 68 0 S4BEG[11]
rlabel metal2 19051 68 19051 68 0 S4BEG[12]
rlabel metal2 19274 296 19274 296 0 S4BEG[13]
rlabel metal2 19550 619 19550 619 0 S4BEG[14]
rlabel metal2 19826 1078 19826 1078 0 S4BEG[15]
rlabel metal2 15962 806 15962 806 0 S4BEG[1]
rlabel metal2 16185 68 16185 68 0 S4BEG[2]
rlabel metal2 16514 143 16514 143 0 S4BEG[3]
rlabel metal2 16790 908 16790 908 0 S4BEG[4]
rlabel metal2 17066 738 17066 738 0 S4BEG[5]
rlabel metal2 17342 755 17342 755 0 S4BEG[6]
rlabel metal2 17618 704 17618 704 0 S4BEG[7]
rlabel metal2 17894 959 17894 959 0 S4BEG[8]
rlabel metal2 18170 483 18170 483 0 S4BEG[9]
rlabel metal2 20201 68 20201 68 0 UserCLK
rlabel metal2 966 9785 966 9785 0 UserCLKo
rlabel metal1 21298 1258 21298 1258 0 net1
rlabel metal1 23276 2822 23276 2822 0 net10
rlabel metal1 20470 1224 20470 1224 0 net100
rlabel metal1 19182 1904 19182 1904 0 net101
rlabel metal1 19918 2006 19918 2006 0 net102
rlabel metal1 22034 1530 22034 1530 0 net103
rlabel metal1 21252 2006 21252 2006 0 net104
rlabel metal1 16698 1326 16698 1326 0 net105
rlabel metal1 17296 1258 17296 1258 0 net106
rlabel metal1 17664 1258 17664 1258 0 net107
rlabel metal1 16790 2006 16790 2006 0 net108
rlabel metal1 18078 918 18078 918 0 net109
rlabel metal1 24058 3706 24058 3706 0 net11
rlabel metal2 19366 1479 19366 1479 0 net110
rlabel metal1 19688 1258 19688 1258 0 net111
rlabel metal1 18078 2040 18078 2040 0 net112
rlabel metal1 18400 2006 18400 2006 0 net113
rlabel metal2 1518 7004 1518 7004 0 net114
rlabel metal2 21206 2108 21206 2108 0 net12
rlabel metal2 22034 2431 22034 2431 0 net13
rlabel metal4 19780 3672 19780 3672 0 net14
rlabel metal1 7774 7378 7774 7378 0 net15
rlabel metal4 19596 2244 19596 2244 0 net16
rlabel metal1 15456 646 15456 646 0 net17
rlabel metal2 11086 7684 11086 7684 0 net18
rlabel metal1 12466 4564 12466 4564 0 net19
rlabel metal2 20746 4148 20746 4148 0 net2
rlabel metal1 13570 7786 13570 7786 0 net20
rlabel metal1 1748 2414 1748 2414 0 net21
rlabel metal1 2438 2448 2438 2448 0 net22
rlabel metal1 1978 2856 1978 2856 0 net23
rlabel metal1 2530 2312 2530 2312 0 net24
rlabel metal1 3404 1938 3404 1938 0 net25
rlabel metal1 3174 1326 3174 1326 0 net26
rlabel metal1 3542 1326 3542 1326 0 net27
rlabel metal1 4646 1938 4646 1938 0 net28
rlabel metal1 5474 1938 5474 1938 0 net29
rlabel metal1 24058 1224 24058 1224 0 net3
rlabel metal1 4278 1326 4278 1326 0 net30
rlabel metal2 5106 1802 5106 1802 0 net31
rlabel metal1 4968 1462 4968 1462 0 net32
rlabel via2 1518 2533 1518 2533 0 net33
rlabel metal2 9338 2686 9338 2686 0 net34
rlabel via2 13662 1955 13662 1955 0 net35
rlabel metal1 2438 3060 2438 3060 0 net36
rlabel metal2 1702 697 1702 697 0 net37
rlabel metal2 1794 1054 1794 1054 0 net38
rlabel metal2 3542 1360 3542 1360 0 net39
rlabel metal1 17158 7820 17158 7820 0 net4
rlabel metal1 2254 1360 2254 1360 0 net40
rlabel metal2 21390 884 21390 884 0 net41
rlabel metal1 7636 1190 7636 1190 0 net42
rlabel metal2 7774 1632 7774 1632 0 net43
rlabel metal2 8050 1054 8050 1054 0 net44
rlabel via2 8970 2091 8970 2091 0 net45
rlabel metal1 9246 1360 9246 1360 0 net46
rlabel viali 9522 1324 9522 1324 0 net47
rlabel metal1 5382 1326 5382 1326 0 net48
rlabel metal3 12604 2448 12604 2448 0 net49
rlabel metal2 24334 2516 24334 2516 0 net5
rlabel metal2 20010 2125 20010 2125 0 net50
rlabel metal2 17986 1020 17986 1020 0 net51
rlabel metal1 20976 1190 20976 1190 0 net52
rlabel metal2 17158 1309 17158 1309 0 net53
rlabel metal2 12466 2040 12466 2040 0 net54
rlabel metal2 16882 1564 16882 1564 0 net55
rlabel metal2 8142 2159 8142 2159 0 net56
rlabel metal1 22126 2040 22126 2040 0 net57
rlabel metal2 2254 7106 2254 7106 0 net58
rlabel metal1 14352 5882 14352 5882 0 net59
rlabel metal1 23690 3094 23690 3094 0 net6
rlabel metal1 18722 8364 18722 8364 0 net60
rlabel metal1 16790 8568 16790 8568 0 net61
rlabel metal1 17802 2618 17802 2618 0 net62
rlabel metal1 19228 2618 19228 2618 0 net63
rlabel metal1 20194 8432 20194 8432 0 net64
rlabel metal1 22264 2278 22264 2278 0 net65
rlabel metal1 22816 2618 22816 2618 0 net66
rlabel metal1 23782 8432 23782 8432 0 net67
rlabel metal1 24058 2822 24058 2822 0 net68
rlabel metal2 3818 6052 3818 6052 0 net69
rlabel metal2 23460 1428 23460 1428 0 net7
rlabel metal1 20286 2924 20286 2924 0 net70
rlabel metal1 6118 8466 6118 8466 0 net71
rlabel metal1 6946 8568 6946 8568 0 net72
rlabel metal1 8372 3978 8372 3978 0 net73
rlabel metal2 9522 6222 9522 6222 0 net74
rlabel metal1 10810 8466 10810 8466 0 net75
rlabel metal1 11868 5338 11868 5338 0 net76
rlabel metal1 13202 8466 13202 8466 0 net77
rlabel metal1 9614 1394 9614 1394 0 net78
rlabel metal1 10166 2006 10166 2006 0 net79
rlabel metal1 23230 1938 23230 1938 0 net8
rlabel metal1 1978 1734 1978 1734 0 net80
rlabel metal1 2346 1802 2346 1802 0 net81
rlabel metal1 2346 476 2346 476 0 net82
rlabel metal2 14214 1020 14214 1020 0 net83
rlabel metal1 12558 1326 12558 1326 0 net84
rlabel metal1 14490 2006 14490 2006 0 net85
rlabel metal1 14858 1870 14858 1870 0 net86
rlabel metal1 15180 1258 15180 1258 0 net87
rlabel metal1 15548 1326 15548 1326 0 net88
rlabel metal1 15962 2380 15962 2380 0 net89
rlabel metal1 23966 1972 23966 1972 0 net9
rlabel metal2 10810 1122 10810 1122 0 net90
rlabel metal1 10212 1326 10212 1326 0 net91
rlabel metal1 11776 2006 11776 2006 0 net92
rlabel metal1 11316 1938 11316 1938 0 net93
rlabel metal1 12190 1258 12190 1258 0 net94
rlabel metal2 12834 1683 12834 1683 0 net95
rlabel metal1 11822 1292 11822 1292 0 net96
rlabel metal2 2622 816 2622 816 0 net97
rlabel metal1 15870 2040 15870 2040 0 net98
rlabel metal1 19504 1938 19504 1938 0 net99
rlabel metal1 19734 4794 19734 4794 0 strobe_inbuf_0.X
rlabel metal1 20838 3026 20838 3026 0 strobe_inbuf_1.X
rlabel metal1 14904 5202 14904 5202 0 strobe_inbuf_10.X
rlabel metal1 23000 7854 23000 7854 0 strobe_inbuf_11.X
rlabel metal1 17434 7888 17434 7888 0 strobe_inbuf_12.X
rlabel metal2 24334 2244 24334 2244 0 strobe_inbuf_13.X
rlabel metal1 22678 2992 22678 2992 0 strobe_inbuf_14.X
rlabel metal1 22034 1292 22034 1292 0 strobe_inbuf_15.X
rlabel metal1 22862 1904 22862 1904 0 strobe_inbuf_16.X
rlabel metal1 23736 1938 23736 1938 0 strobe_inbuf_17.X
rlabel metal1 23874 7514 23874 7514 0 strobe_inbuf_18.X
rlabel metal2 24196 1938 24196 1938 0 strobe_inbuf_19.X
rlabel metal1 20562 2380 20562 2380 0 strobe_inbuf_2.X
rlabel metal1 6348 7514 6348 7514 0 strobe_inbuf_3.X
rlabel metal1 7452 7514 7452 7514 0 strobe_inbuf_4.X
rlabel metal1 8924 3706 8924 3706 0 strobe_inbuf_5.X
rlabel metal1 10028 3502 10028 3502 0 strobe_inbuf_6.X
rlabel metal1 11362 7820 11362 7820 0 strobe_inbuf_7.X
rlabel metal1 12282 4794 12282 4794 0 strobe_inbuf_8.X
rlabel metal1 13846 7888 13846 7888 0 strobe_inbuf_9.X
rlabel metal2 19458 5508 19458 5508 0 strobe_outbuf_0.X
rlabel metal1 20240 3162 20240 3162 0 strobe_outbuf_1.X
rlabel metal2 14674 5508 14674 5508 0 strobe_outbuf_10.X
rlabel metal1 22954 8058 22954 8058 0 strobe_outbuf_11.X
rlabel metal1 17342 8058 17342 8058 0 strobe_outbuf_12.X
rlabel via2 20654 2499 20654 2499 0 strobe_outbuf_13.X
rlabel metal2 19458 2618 19458 2618 0 strobe_outbuf_14.X
rlabel metal1 21758 1530 21758 1530 0 strobe_outbuf_15.X
rlabel metal1 22540 2074 22540 2074 0 strobe_outbuf_16.X
rlabel metal1 23368 2074 23368 2074 0 strobe_outbuf_17.X
rlabel metal1 23598 8058 23598 8058 0 strobe_outbuf_18.X
rlabel metal1 24196 2890 24196 2890 0 strobe_outbuf_19.X
rlabel metal1 20240 2618 20240 2618 0 strobe_outbuf_2.X
rlabel metal1 6348 8058 6348 8058 0 strobe_outbuf_3.X
rlabel metal1 7452 8058 7452 8058 0 strobe_outbuf_4.X
rlabel metal1 8648 4114 8648 4114 0 strobe_outbuf_5.X
rlabel metal1 9752 3706 9752 3706 0 strobe_outbuf_6.X
rlabel metal2 11178 8262 11178 8262 0 strobe_outbuf_7.X
rlabel metal1 12144 5202 12144 5202 0 strobe_outbuf_8.X
rlabel metal1 13616 8058 13616 8058 0 strobe_outbuf_9.X
<< properties >>
string FIXED_BBOX 0 0 26000 10000
<< end >>
