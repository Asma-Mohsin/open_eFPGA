// This is the unpowered netlist.
module RegFile (UserCLK,
    UserCLKo,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire AD0;
 wire AD1;
 wire AD2;
 wire AD3;
 wire A_ADR0;
 wire A_ADR1;
 wire A_ADR2;
 wire A_ADR3;
 wire A_ADR4;
 wire BD0;
 wire BD1;
 wire BD2;
 wire BD3;
 wire B_ADR0;
 wire B_ADR1;
 wire B_ADR2;
 wire B_ADR3;
 wire B_ADR4;
 wire \ConfigBits[0] ;
 wire \ConfigBits[100] ;
 wire \ConfigBits[101] ;
 wire \ConfigBits[102] ;
 wire \ConfigBits[103] ;
 wire \ConfigBits[104] ;
 wire \ConfigBits[105] ;
 wire \ConfigBits[106] ;
 wire \ConfigBits[107] ;
 wire \ConfigBits[108] ;
 wire \ConfigBits[109] ;
 wire \ConfigBits[10] ;
 wire \ConfigBits[110] ;
 wire \ConfigBits[111] ;
 wire \ConfigBits[112] ;
 wire \ConfigBits[113] ;
 wire \ConfigBits[114] ;
 wire \ConfigBits[115] ;
 wire \ConfigBits[116] ;
 wire \ConfigBits[117] ;
 wire \ConfigBits[118] ;
 wire \ConfigBits[119] ;
 wire \ConfigBits[11] ;
 wire \ConfigBits[120] ;
 wire \ConfigBits[121] ;
 wire \ConfigBits[122] ;
 wire \ConfigBits[123] ;
 wire \ConfigBits[124] ;
 wire \ConfigBits[125] ;
 wire \ConfigBits[126] ;
 wire \ConfigBits[127] ;
 wire \ConfigBits[128] ;
 wire \ConfigBits[129] ;
 wire \ConfigBits[12] ;
 wire \ConfigBits[130] ;
 wire \ConfigBits[131] ;
 wire \ConfigBits[132] ;
 wire \ConfigBits[133] ;
 wire \ConfigBits[134] ;
 wire \ConfigBits[135] ;
 wire \ConfigBits[136] ;
 wire \ConfigBits[137] ;
 wire \ConfigBits[138] ;
 wire \ConfigBits[139] ;
 wire \ConfigBits[13] ;
 wire \ConfigBits[140] ;
 wire \ConfigBits[141] ;
 wire \ConfigBits[142] ;
 wire \ConfigBits[143] ;
 wire \ConfigBits[144] ;
 wire \ConfigBits[145] ;
 wire \ConfigBits[146] ;
 wire \ConfigBits[147] ;
 wire \ConfigBits[148] ;
 wire \ConfigBits[149] ;
 wire \ConfigBits[14] ;
 wire \ConfigBits[150] ;
 wire \ConfigBits[151] ;
 wire \ConfigBits[152] ;
 wire \ConfigBits[153] ;
 wire \ConfigBits[154] ;
 wire \ConfigBits[155] ;
 wire \ConfigBits[156] ;
 wire \ConfigBits[157] ;
 wire \ConfigBits[158] ;
 wire \ConfigBits[159] ;
 wire \ConfigBits[15] ;
 wire \ConfigBits[160] ;
 wire \ConfigBits[161] ;
 wire \ConfigBits[162] ;
 wire \ConfigBits[163] ;
 wire \ConfigBits[164] ;
 wire \ConfigBits[165] ;
 wire \ConfigBits[166] ;
 wire \ConfigBits[167] ;
 wire \ConfigBits[168] ;
 wire \ConfigBits[169] ;
 wire \ConfigBits[16] ;
 wire \ConfigBits[170] ;
 wire \ConfigBits[171] ;
 wire \ConfigBits[172] ;
 wire \ConfigBits[173] ;
 wire \ConfigBits[174] ;
 wire \ConfigBits[175] ;
 wire \ConfigBits[176] ;
 wire \ConfigBits[177] ;
 wire \ConfigBits[178] ;
 wire \ConfigBits[179] ;
 wire \ConfigBits[17] ;
 wire \ConfigBits[180] ;
 wire \ConfigBits[181] ;
 wire \ConfigBits[182] ;
 wire \ConfigBits[183] ;
 wire \ConfigBits[184] ;
 wire \ConfigBits[185] ;
 wire \ConfigBits[186] ;
 wire \ConfigBits[187] ;
 wire \ConfigBits[188] ;
 wire \ConfigBits[189] ;
 wire \ConfigBits[18] ;
 wire \ConfigBits[190] ;
 wire \ConfigBits[191] ;
 wire \ConfigBits[192] ;
 wire \ConfigBits[193] ;
 wire \ConfigBits[194] ;
 wire \ConfigBits[195] ;
 wire \ConfigBits[196] ;
 wire \ConfigBits[197] ;
 wire \ConfigBits[198] ;
 wire \ConfigBits[199] ;
 wire \ConfigBits[19] ;
 wire \ConfigBits[1] ;
 wire \ConfigBits[200] ;
 wire \ConfigBits[201] ;
 wire \ConfigBits[202] ;
 wire \ConfigBits[203] ;
 wire \ConfigBits[204] ;
 wire \ConfigBits[205] ;
 wire \ConfigBits[206] ;
 wire \ConfigBits[207] ;
 wire \ConfigBits[208] ;
 wire \ConfigBits[209] ;
 wire \ConfigBits[20] ;
 wire \ConfigBits[210] ;
 wire \ConfigBits[211] ;
 wire \ConfigBits[212] ;
 wire \ConfigBits[213] ;
 wire \ConfigBits[214] ;
 wire \ConfigBits[215] ;
 wire \ConfigBits[216] ;
 wire \ConfigBits[217] ;
 wire \ConfigBits[218] ;
 wire \ConfigBits[219] ;
 wire \ConfigBits[21] ;
 wire \ConfigBits[220] ;
 wire \ConfigBits[221] ;
 wire \ConfigBits[222] ;
 wire \ConfigBits[223] ;
 wire \ConfigBits[224] ;
 wire \ConfigBits[225] ;
 wire \ConfigBits[226] ;
 wire \ConfigBits[227] ;
 wire \ConfigBits[228] ;
 wire \ConfigBits[229] ;
 wire \ConfigBits[22] ;
 wire \ConfigBits[230] ;
 wire \ConfigBits[231] ;
 wire \ConfigBits[232] ;
 wire \ConfigBits[233] ;
 wire \ConfigBits[234] ;
 wire \ConfigBits[235] ;
 wire \ConfigBits[236] ;
 wire \ConfigBits[237] ;
 wire \ConfigBits[238] ;
 wire \ConfigBits[239] ;
 wire \ConfigBits[23] ;
 wire \ConfigBits[240] ;
 wire \ConfigBits[241] ;
 wire \ConfigBits[242] ;
 wire \ConfigBits[243] ;
 wire \ConfigBits[244] ;
 wire \ConfigBits[245] ;
 wire \ConfigBits[246] ;
 wire \ConfigBits[247] ;
 wire \ConfigBits[248] ;
 wire \ConfigBits[249] ;
 wire \ConfigBits[24] ;
 wire \ConfigBits[250] ;
 wire \ConfigBits[251] ;
 wire \ConfigBits[252] ;
 wire \ConfigBits[253] ;
 wire \ConfigBits[254] ;
 wire \ConfigBits[255] ;
 wire \ConfigBits[256] ;
 wire \ConfigBits[257] ;
 wire \ConfigBits[258] ;
 wire \ConfigBits[259] ;
 wire \ConfigBits[25] ;
 wire \ConfigBits[260] ;
 wire \ConfigBits[261] ;
 wire \ConfigBits[262] ;
 wire \ConfigBits[263] ;
 wire \ConfigBits[264] ;
 wire \ConfigBits[265] ;
 wire \ConfigBits[266] ;
 wire \ConfigBits[267] ;
 wire \ConfigBits[268] ;
 wire \ConfigBits[269] ;
 wire \ConfigBits[26] ;
 wire \ConfigBits[270] ;
 wire \ConfigBits[271] ;
 wire \ConfigBits[272] ;
 wire \ConfigBits[273] ;
 wire \ConfigBits[274] ;
 wire \ConfigBits[275] ;
 wire \ConfigBits[276] ;
 wire \ConfigBits[277] ;
 wire \ConfigBits[278] ;
 wire \ConfigBits[279] ;
 wire \ConfigBits[27] ;
 wire \ConfigBits[280] ;
 wire \ConfigBits[281] ;
 wire \ConfigBits[282] ;
 wire \ConfigBits[283] ;
 wire \ConfigBits[284] ;
 wire \ConfigBits[285] ;
 wire \ConfigBits[286] ;
 wire \ConfigBits[287] ;
 wire \ConfigBits[288] ;
 wire \ConfigBits[289] ;
 wire \ConfigBits[28] ;
 wire \ConfigBits[290] ;
 wire \ConfigBits[291] ;
 wire \ConfigBits[292] ;
 wire \ConfigBits[293] ;
 wire \ConfigBits[294] ;
 wire \ConfigBits[295] ;
 wire \ConfigBits[296] ;
 wire \ConfigBits[297] ;
 wire \ConfigBits[298] ;
 wire \ConfigBits[299] ;
 wire \ConfigBits[29] ;
 wire \ConfigBits[2] ;
 wire \ConfigBits[300] ;
 wire \ConfigBits[301] ;
 wire \ConfigBits[302] ;
 wire \ConfigBits[303] ;
 wire \ConfigBits[304] ;
 wire \ConfigBits[305] ;
 wire \ConfigBits[306] ;
 wire \ConfigBits[307] ;
 wire \ConfigBits[308] ;
 wire \ConfigBits[309] ;
 wire \ConfigBits[30] ;
 wire \ConfigBits[310] ;
 wire \ConfigBits[311] ;
 wire \ConfigBits[312] ;
 wire \ConfigBits[313] ;
 wire \ConfigBits[314] ;
 wire \ConfigBits[315] ;
 wire \ConfigBits[316] ;
 wire \ConfigBits[317] ;
 wire \ConfigBits[318] ;
 wire \ConfigBits[319] ;
 wire \ConfigBits[31] ;
 wire \ConfigBits[320] ;
 wire \ConfigBits[321] ;
 wire \ConfigBits[322] ;
 wire \ConfigBits[323] ;
 wire \ConfigBits[324] ;
 wire \ConfigBits[325] ;
 wire \ConfigBits[326] ;
 wire \ConfigBits[327] ;
 wire \ConfigBits[328] ;
 wire \ConfigBits[329] ;
 wire \ConfigBits[32] ;
 wire \ConfigBits[330] ;
 wire \ConfigBits[331] ;
 wire \ConfigBits[332] ;
 wire \ConfigBits[333] ;
 wire \ConfigBits[334] ;
 wire \ConfigBits[335] ;
 wire \ConfigBits[336] ;
 wire \ConfigBits[337] ;
 wire \ConfigBits[338] ;
 wire \ConfigBits[339] ;
 wire \ConfigBits[33] ;
 wire \ConfigBits[340] ;
 wire \ConfigBits[341] ;
 wire \ConfigBits[342] ;
 wire \ConfigBits[343] ;
 wire \ConfigBits[344] ;
 wire \ConfigBits[345] ;
 wire \ConfigBits[346] ;
 wire \ConfigBits[347] ;
 wire \ConfigBits[348] ;
 wire \ConfigBits[349] ;
 wire \ConfigBits[34] ;
 wire \ConfigBits[350] ;
 wire \ConfigBits[351] ;
 wire \ConfigBits[352] ;
 wire \ConfigBits[353] ;
 wire \ConfigBits[354] ;
 wire \ConfigBits[355] ;
 wire \ConfigBits[356] ;
 wire \ConfigBits[357] ;
 wire \ConfigBits[358] ;
 wire \ConfigBits[359] ;
 wire \ConfigBits[35] ;
 wire \ConfigBits[360] ;
 wire \ConfigBits[361] ;
 wire \ConfigBits[362] ;
 wire \ConfigBits[363] ;
 wire \ConfigBits[364] ;
 wire \ConfigBits[365] ;
 wire \ConfigBits[366] ;
 wire \ConfigBits[367] ;
 wire \ConfigBits[368] ;
 wire \ConfigBits[369] ;
 wire \ConfigBits[36] ;
 wire \ConfigBits[370] ;
 wire \ConfigBits[371] ;
 wire \ConfigBits[372] ;
 wire \ConfigBits[373] ;
 wire \ConfigBits[374] ;
 wire \ConfigBits[375] ;
 wire \ConfigBits[376] ;
 wire \ConfigBits[377] ;
 wire \ConfigBits[378] ;
 wire \ConfigBits[379] ;
 wire \ConfigBits[37] ;
 wire \ConfigBits[380] ;
 wire \ConfigBits[381] ;
 wire \ConfigBits[382] ;
 wire \ConfigBits[383] ;
 wire \ConfigBits[384] ;
 wire \ConfigBits[385] ;
 wire \ConfigBits[386] ;
 wire \ConfigBits[387] ;
 wire \ConfigBits[388] ;
 wire \ConfigBits[389] ;
 wire \ConfigBits[38] ;
 wire \ConfigBits[390] ;
 wire \ConfigBits[391] ;
 wire \ConfigBits[392] ;
 wire \ConfigBits[393] ;
 wire \ConfigBits[394] ;
 wire \ConfigBits[395] ;
 wire \ConfigBits[396] ;
 wire \ConfigBits[397] ;
 wire \ConfigBits[398] ;
 wire \ConfigBits[399] ;
 wire \ConfigBits[39] ;
 wire \ConfigBits[3] ;
 wire \ConfigBits[400] ;
 wire \ConfigBits[401] ;
 wire \ConfigBits[402] ;
 wire \ConfigBits[403] ;
 wire \ConfigBits[404] ;
 wire \ConfigBits[405] ;
 wire \ConfigBits[406] ;
 wire \ConfigBits[407] ;
 wire \ConfigBits[408] ;
 wire \ConfigBits[409] ;
 wire \ConfigBits[40] ;
 wire \ConfigBits[410] ;
 wire \ConfigBits[411] ;
 wire \ConfigBits[412] ;
 wire \ConfigBits[413] ;
 wire \ConfigBits[41] ;
 wire \ConfigBits[42] ;
 wire \ConfigBits[43] ;
 wire \ConfigBits[44] ;
 wire \ConfigBits[45] ;
 wire \ConfigBits[46] ;
 wire \ConfigBits[47] ;
 wire \ConfigBits[48] ;
 wire \ConfigBits[49] ;
 wire \ConfigBits[4] ;
 wire \ConfigBits[50] ;
 wire \ConfigBits[51] ;
 wire \ConfigBits[52] ;
 wire \ConfigBits[53] ;
 wire \ConfigBits[54] ;
 wire \ConfigBits[55] ;
 wire \ConfigBits[56] ;
 wire \ConfigBits[57] ;
 wire \ConfigBits[58] ;
 wire \ConfigBits[59] ;
 wire \ConfigBits[5] ;
 wire \ConfigBits[60] ;
 wire \ConfigBits[61] ;
 wire \ConfigBits[62] ;
 wire \ConfigBits[63] ;
 wire \ConfigBits[64] ;
 wire \ConfigBits[65] ;
 wire \ConfigBits[66] ;
 wire \ConfigBits[67] ;
 wire \ConfigBits[68] ;
 wire \ConfigBits[69] ;
 wire \ConfigBits[6] ;
 wire \ConfigBits[70] ;
 wire \ConfigBits[71] ;
 wire \ConfigBits[72] ;
 wire \ConfigBits[73] ;
 wire \ConfigBits[74] ;
 wire \ConfigBits[75] ;
 wire \ConfigBits[76] ;
 wire \ConfigBits[77] ;
 wire \ConfigBits[78] ;
 wire \ConfigBits[79] ;
 wire \ConfigBits[7] ;
 wire \ConfigBits[80] ;
 wire \ConfigBits[81] ;
 wire \ConfigBits[82] ;
 wire \ConfigBits[83] ;
 wire \ConfigBits[84] ;
 wire \ConfigBits[85] ;
 wire \ConfigBits[86] ;
 wire \ConfigBits[87] ;
 wire \ConfigBits[88] ;
 wire \ConfigBits[89] ;
 wire \ConfigBits[8] ;
 wire \ConfigBits[90] ;
 wire \ConfigBits[91] ;
 wire \ConfigBits[92] ;
 wire \ConfigBits[93] ;
 wire \ConfigBits[94] ;
 wire \ConfigBits[95] ;
 wire \ConfigBits[96] ;
 wire \ConfigBits[97] ;
 wire \ConfigBits[98] ;
 wire \ConfigBits[99] ;
 wire \ConfigBits[9] ;
 wire \ConfigBits_N[0] ;
 wire \ConfigBits_N[100] ;
 wire \ConfigBits_N[101] ;
 wire \ConfigBits_N[102] ;
 wire \ConfigBits_N[103] ;
 wire \ConfigBits_N[104] ;
 wire \ConfigBits_N[105] ;
 wire \ConfigBits_N[106] ;
 wire \ConfigBits_N[107] ;
 wire \ConfigBits_N[108] ;
 wire \ConfigBits_N[109] ;
 wire \ConfigBits_N[10] ;
 wire \ConfigBits_N[110] ;
 wire \ConfigBits_N[111] ;
 wire \ConfigBits_N[112] ;
 wire \ConfigBits_N[113] ;
 wire \ConfigBits_N[114] ;
 wire \ConfigBits_N[115] ;
 wire \ConfigBits_N[116] ;
 wire \ConfigBits_N[117] ;
 wire \ConfigBits_N[118] ;
 wire \ConfigBits_N[119] ;
 wire \ConfigBits_N[11] ;
 wire \ConfigBits_N[120] ;
 wire \ConfigBits_N[121] ;
 wire \ConfigBits_N[122] ;
 wire \ConfigBits_N[123] ;
 wire \ConfigBits_N[124] ;
 wire \ConfigBits_N[125] ;
 wire \ConfigBits_N[126] ;
 wire \ConfigBits_N[127] ;
 wire \ConfigBits_N[128] ;
 wire \ConfigBits_N[129] ;
 wire \ConfigBits_N[12] ;
 wire \ConfigBits_N[130] ;
 wire \ConfigBits_N[131] ;
 wire \ConfigBits_N[132] ;
 wire \ConfigBits_N[133] ;
 wire \ConfigBits_N[134] ;
 wire \ConfigBits_N[135] ;
 wire \ConfigBits_N[136] ;
 wire \ConfigBits_N[137] ;
 wire \ConfigBits_N[138] ;
 wire \ConfigBits_N[139] ;
 wire \ConfigBits_N[13] ;
 wire \ConfigBits_N[140] ;
 wire \ConfigBits_N[141] ;
 wire \ConfigBits_N[142] ;
 wire \ConfigBits_N[143] ;
 wire \ConfigBits_N[144] ;
 wire \ConfigBits_N[145] ;
 wire \ConfigBits_N[146] ;
 wire \ConfigBits_N[147] ;
 wire \ConfigBits_N[148] ;
 wire \ConfigBits_N[149] ;
 wire \ConfigBits_N[14] ;
 wire \ConfigBits_N[150] ;
 wire \ConfigBits_N[151] ;
 wire \ConfigBits_N[152] ;
 wire \ConfigBits_N[153] ;
 wire \ConfigBits_N[154] ;
 wire \ConfigBits_N[155] ;
 wire \ConfigBits_N[156] ;
 wire \ConfigBits_N[157] ;
 wire \ConfigBits_N[158] ;
 wire \ConfigBits_N[159] ;
 wire \ConfigBits_N[15] ;
 wire \ConfigBits_N[160] ;
 wire \ConfigBits_N[161] ;
 wire \ConfigBits_N[162] ;
 wire \ConfigBits_N[163] ;
 wire \ConfigBits_N[164] ;
 wire \ConfigBits_N[165] ;
 wire \ConfigBits_N[166] ;
 wire \ConfigBits_N[167] ;
 wire \ConfigBits_N[168] ;
 wire \ConfigBits_N[169] ;
 wire \ConfigBits_N[16] ;
 wire \ConfigBits_N[170] ;
 wire \ConfigBits_N[171] ;
 wire \ConfigBits_N[172] ;
 wire \ConfigBits_N[173] ;
 wire \ConfigBits_N[174] ;
 wire \ConfigBits_N[175] ;
 wire \ConfigBits_N[176] ;
 wire \ConfigBits_N[177] ;
 wire \ConfigBits_N[178] ;
 wire \ConfigBits_N[179] ;
 wire \ConfigBits_N[17] ;
 wire \ConfigBits_N[180] ;
 wire \ConfigBits_N[181] ;
 wire \ConfigBits_N[182] ;
 wire \ConfigBits_N[183] ;
 wire \ConfigBits_N[184] ;
 wire \ConfigBits_N[185] ;
 wire \ConfigBits_N[186] ;
 wire \ConfigBits_N[187] ;
 wire \ConfigBits_N[188] ;
 wire \ConfigBits_N[189] ;
 wire \ConfigBits_N[18] ;
 wire \ConfigBits_N[190] ;
 wire \ConfigBits_N[191] ;
 wire \ConfigBits_N[192] ;
 wire \ConfigBits_N[193] ;
 wire \ConfigBits_N[194] ;
 wire \ConfigBits_N[195] ;
 wire \ConfigBits_N[196] ;
 wire \ConfigBits_N[197] ;
 wire \ConfigBits_N[198] ;
 wire \ConfigBits_N[199] ;
 wire \ConfigBits_N[19] ;
 wire \ConfigBits_N[1] ;
 wire \ConfigBits_N[200] ;
 wire \ConfigBits_N[201] ;
 wire \ConfigBits_N[202] ;
 wire \ConfigBits_N[203] ;
 wire \ConfigBits_N[204] ;
 wire \ConfigBits_N[205] ;
 wire \ConfigBits_N[206] ;
 wire \ConfigBits_N[207] ;
 wire \ConfigBits_N[208] ;
 wire \ConfigBits_N[209] ;
 wire \ConfigBits_N[20] ;
 wire \ConfigBits_N[210] ;
 wire \ConfigBits_N[211] ;
 wire \ConfigBits_N[212] ;
 wire \ConfigBits_N[213] ;
 wire \ConfigBits_N[214] ;
 wire \ConfigBits_N[215] ;
 wire \ConfigBits_N[216] ;
 wire \ConfigBits_N[217] ;
 wire \ConfigBits_N[218] ;
 wire \ConfigBits_N[219] ;
 wire \ConfigBits_N[21] ;
 wire \ConfigBits_N[220] ;
 wire \ConfigBits_N[221] ;
 wire \ConfigBits_N[222] ;
 wire \ConfigBits_N[223] ;
 wire \ConfigBits_N[224] ;
 wire \ConfigBits_N[225] ;
 wire \ConfigBits_N[226] ;
 wire \ConfigBits_N[227] ;
 wire \ConfigBits_N[228] ;
 wire \ConfigBits_N[229] ;
 wire \ConfigBits_N[22] ;
 wire \ConfigBits_N[230] ;
 wire \ConfigBits_N[231] ;
 wire \ConfigBits_N[232] ;
 wire \ConfigBits_N[233] ;
 wire \ConfigBits_N[234] ;
 wire \ConfigBits_N[235] ;
 wire \ConfigBits_N[236] ;
 wire \ConfigBits_N[237] ;
 wire \ConfigBits_N[238] ;
 wire \ConfigBits_N[239] ;
 wire \ConfigBits_N[23] ;
 wire \ConfigBits_N[240] ;
 wire \ConfigBits_N[241] ;
 wire \ConfigBits_N[242] ;
 wire \ConfigBits_N[243] ;
 wire \ConfigBits_N[244] ;
 wire \ConfigBits_N[245] ;
 wire \ConfigBits_N[246] ;
 wire \ConfigBits_N[247] ;
 wire \ConfigBits_N[248] ;
 wire \ConfigBits_N[249] ;
 wire \ConfigBits_N[24] ;
 wire \ConfigBits_N[250] ;
 wire \ConfigBits_N[251] ;
 wire \ConfigBits_N[252] ;
 wire \ConfigBits_N[253] ;
 wire \ConfigBits_N[254] ;
 wire \ConfigBits_N[255] ;
 wire \ConfigBits_N[256] ;
 wire \ConfigBits_N[257] ;
 wire \ConfigBits_N[258] ;
 wire \ConfigBits_N[259] ;
 wire \ConfigBits_N[25] ;
 wire \ConfigBits_N[260] ;
 wire \ConfigBits_N[261] ;
 wire \ConfigBits_N[262] ;
 wire \ConfigBits_N[263] ;
 wire \ConfigBits_N[264] ;
 wire \ConfigBits_N[265] ;
 wire \ConfigBits_N[266] ;
 wire \ConfigBits_N[267] ;
 wire \ConfigBits_N[268] ;
 wire \ConfigBits_N[269] ;
 wire \ConfigBits_N[26] ;
 wire \ConfigBits_N[270] ;
 wire \ConfigBits_N[271] ;
 wire \ConfigBits_N[272] ;
 wire \ConfigBits_N[273] ;
 wire \ConfigBits_N[274] ;
 wire \ConfigBits_N[275] ;
 wire \ConfigBits_N[276] ;
 wire \ConfigBits_N[277] ;
 wire \ConfigBits_N[278] ;
 wire \ConfigBits_N[279] ;
 wire \ConfigBits_N[27] ;
 wire \ConfigBits_N[280] ;
 wire \ConfigBits_N[281] ;
 wire \ConfigBits_N[282] ;
 wire \ConfigBits_N[283] ;
 wire \ConfigBits_N[284] ;
 wire \ConfigBits_N[285] ;
 wire \ConfigBits_N[286] ;
 wire \ConfigBits_N[287] ;
 wire \ConfigBits_N[288] ;
 wire \ConfigBits_N[289] ;
 wire \ConfigBits_N[28] ;
 wire \ConfigBits_N[290] ;
 wire \ConfigBits_N[291] ;
 wire \ConfigBits_N[292] ;
 wire \ConfigBits_N[293] ;
 wire \ConfigBits_N[294] ;
 wire \ConfigBits_N[295] ;
 wire \ConfigBits_N[296] ;
 wire \ConfigBits_N[297] ;
 wire \ConfigBits_N[298] ;
 wire \ConfigBits_N[299] ;
 wire \ConfigBits_N[29] ;
 wire \ConfigBits_N[2] ;
 wire \ConfigBits_N[300] ;
 wire \ConfigBits_N[301] ;
 wire \ConfigBits_N[302] ;
 wire \ConfigBits_N[303] ;
 wire \ConfigBits_N[304] ;
 wire \ConfigBits_N[305] ;
 wire \ConfigBits_N[306] ;
 wire \ConfigBits_N[307] ;
 wire \ConfigBits_N[308] ;
 wire \ConfigBits_N[309] ;
 wire \ConfigBits_N[30] ;
 wire \ConfigBits_N[310] ;
 wire \ConfigBits_N[311] ;
 wire \ConfigBits_N[312] ;
 wire \ConfigBits_N[313] ;
 wire \ConfigBits_N[314] ;
 wire \ConfigBits_N[315] ;
 wire \ConfigBits_N[316] ;
 wire \ConfigBits_N[317] ;
 wire \ConfigBits_N[318] ;
 wire \ConfigBits_N[319] ;
 wire \ConfigBits_N[31] ;
 wire \ConfigBits_N[320] ;
 wire \ConfigBits_N[321] ;
 wire \ConfigBits_N[322] ;
 wire \ConfigBits_N[323] ;
 wire \ConfigBits_N[324] ;
 wire \ConfigBits_N[325] ;
 wire \ConfigBits_N[326] ;
 wire \ConfigBits_N[327] ;
 wire \ConfigBits_N[328] ;
 wire \ConfigBits_N[329] ;
 wire \ConfigBits_N[32] ;
 wire \ConfigBits_N[330] ;
 wire \ConfigBits_N[331] ;
 wire \ConfigBits_N[332] ;
 wire \ConfigBits_N[333] ;
 wire \ConfigBits_N[334] ;
 wire \ConfigBits_N[335] ;
 wire \ConfigBits_N[336] ;
 wire \ConfigBits_N[337] ;
 wire \ConfigBits_N[338] ;
 wire \ConfigBits_N[339] ;
 wire \ConfigBits_N[33] ;
 wire \ConfigBits_N[340] ;
 wire \ConfigBits_N[341] ;
 wire \ConfigBits_N[342] ;
 wire \ConfigBits_N[343] ;
 wire \ConfigBits_N[344] ;
 wire \ConfigBits_N[345] ;
 wire \ConfigBits_N[346] ;
 wire \ConfigBits_N[347] ;
 wire \ConfigBits_N[348] ;
 wire \ConfigBits_N[349] ;
 wire \ConfigBits_N[34] ;
 wire \ConfigBits_N[350] ;
 wire \ConfigBits_N[351] ;
 wire \ConfigBits_N[352] ;
 wire \ConfigBits_N[353] ;
 wire \ConfigBits_N[354] ;
 wire \ConfigBits_N[355] ;
 wire \ConfigBits_N[356] ;
 wire \ConfigBits_N[357] ;
 wire \ConfigBits_N[358] ;
 wire \ConfigBits_N[359] ;
 wire \ConfigBits_N[35] ;
 wire \ConfigBits_N[360] ;
 wire \ConfigBits_N[361] ;
 wire \ConfigBits_N[362] ;
 wire \ConfigBits_N[363] ;
 wire \ConfigBits_N[364] ;
 wire \ConfigBits_N[365] ;
 wire \ConfigBits_N[366] ;
 wire \ConfigBits_N[367] ;
 wire \ConfigBits_N[368] ;
 wire \ConfigBits_N[369] ;
 wire \ConfigBits_N[36] ;
 wire \ConfigBits_N[370] ;
 wire \ConfigBits_N[371] ;
 wire \ConfigBits_N[372] ;
 wire \ConfigBits_N[373] ;
 wire \ConfigBits_N[374] ;
 wire \ConfigBits_N[375] ;
 wire \ConfigBits_N[376] ;
 wire \ConfigBits_N[377] ;
 wire \ConfigBits_N[378] ;
 wire \ConfigBits_N[379] ;
 wire \ConfigBits_N[37] ;
 wire \ConfigBits_N[380] ;
 wire \ConfigBits_N[381] ;
 wire \ConfigBits_N[382] ;
 wire \ConfigBits_N[383] ;
 wire \ConfigBits_N[384] ;
 wire \ConfigBits_N[385] ;
 wire \ConfigBits_N[386] ;
 wire \ConfigBits_N[387] ;
 wire \ConfigBits_N[388] ;
 wire \ConfigBits_N[389] ;
 wire \ConfigBits_N[38] ;
 wire \ConfigBits_N[390] ;
 wire \ConfigBits_N[391] ;
 wire \ConfigBits_N[392] ;
 wire \ConfigBits_N[393] ;
 wire \ConfigBits_N[394] ;
 wire \ConfigBits_N[395] ;
 wire \ConfigBits_N[396] ;
 wire \ConfigBits_N[397] ;
 wire \ConfigBits_N[398] ;
 wire \ConfigBits_N[399] ;
 wire \ConfigBits_N[39] ;
 wire \ConfigBits_N[3] ;
 wire \ConfigBits_N[400] ;
 wire \ConfigBits_N[401] ;
 wire \ConfigBits_N[402] ;
 wire \ConfigBits_N[403] ;
 wire \ConfigBits_N[404] ;
 wire \ConfigBits_N[405] ;
 wire \ConfigBits_N[406] ;
 wire \ConfigBits_N[407] ;
 wire \ConfigBits_N[408] ;
 wire \ConfigBits_N[409] ;
 wire \ConfigBits_N[40] ;
 wire \ConfigBits_N[410] ;
 wire \ConfigBits_N[411] ;
 wire \ConfigBits_N[412] ;
 wire \ConfigBits_N[413] ;
 wire \ConfigBits_N[41] ;
 wire \ConfigBits_N[42] ;
 wire \ConfigBits_N[43] ;
 wire \ConfigBits_N[44] ;
 wire \ConfigBits_N[45] ;
 wire \ConfigBits_N[46] ;
 wire \ConfigBits_N[47] ;
 wire \ConfigBits_N[48] ;
 wire \ConfigBits_N[49] ;
 wire \ConfigBits_N[4] ;
 wire \ConfigBits_N[50] ;
 wire \ConfigBits_N[51] ;
 wire \ConfigBits_N[52] ;
 wire \ConfigBits_N[53] ;
 wire \ConfigBits_N[54] ;
 wire \ConfigBits_N[55] ;
 wire \ConfigBits_N[56] ;
 wire \ConfigBits_N[57] ;
 wire \ConfigBits_N[58] ;
 wire \ConfigBits_N[59] ;
 wire \ConfigBits_N[5] ;
 wire \ConfigBits_N[60] ;
 wire \ConfigBits_N[61] ;
 wire \ConfigBits_N[62] ;
 wire \ConfigBits_N[63] ;
 wire \ConfigBits_N[64] ;
 wire \ConfigBits_N[65] ;
 wire \ConfigBits_N[66] ;
 wire \ConfigBits_N[67] ;
 wire \ConfigBits_N[68] ;
 wire \ConfigBits_N[69] ;
 wire \ConfigBits_N[6] ;
 wire \ConfigBits_N[70] ;
 wire \ConfigBits_N[71] ;
 wire \ConfigBits_N[72] ;
 wire \ConfigBits_N[73] ;
 wire \ConfigBits_N[74] ;
 wire \ConfigBits_N[75] ;
 wire \ConfigBits_N[76] ;
 wire \ConfigBits_N[77] ;
 wire \ConfigBits_N[78] ;
 wire \ConfigBits_N[79] ;
 wire \ConfigBits_N[7] ;
 wire \ConfigBits_N[80] ;
 wire \ConfigBits_N[81] ;
 wire \ConfigBits_N[82] ;
 wire \ConfigBits_N[83] ;
 wire \ConfigBits_N[84] ;
 wire \ConfigBits_N[85] ;
 wire \ConfigBits_N[86] ;
 wire \ConfigBits_N[87] ;
 wire \ConfigBits_N[88] ;
 wire \ConfigBits_N[89] ;
 wire \ConfigBits_N[8] ;
 wire \ConfigBits_N[90] ;
 wire \ConfigBits_N[91] ;
 wire \ConfigBits_N[92] ;
 wire \ConfigBits_N[93] ;
 wire \ConfigBits_N[94] ;
 wire \ConfigBits_N[95] ;
 wire \ConfigBits_N[96] ;
 wire \ConfigBits_N[97] ;
 wire \ConfigBits_N[98] ;
 wire \ConfigBits_N[99] ;
 wire \ConfigBits_N[9] ;
 wire D0;
 wire D1;
 wire D2;
 wire D3;
 wire \E6BEG_i[0] ;
 wire \E6BEG_i[1] ;
 wire \E6BEG_i[2] ;
 wire \E6BEG_i[3] ;
 wire \E6BEG_i[4] ;
 wire \E6BEG_i[5] ;
 wire \E6BEG_i[6] ;
 wire \E6BEG_i[7] ;
 wire \E6BEG_i[8] ;
 wire \E6BEG_i[9] ;
 wire \EE4BEG_i[0] ;
 wire \EE4BEG_i[10] ;
 wire \EE4BEG_i[11] ;
 wire \EE4BEG_i[1] ;
 wire \EE4BEG_i[2] ;
 wire \EE4BEG_i[3] ;
 wire \EE4BEG_i[4] ;
 wire \EE4BEG_i[5] ;
 wire \EE4BEG_i[6] ;
 wire \EE4BEG_i[7] ;
 wire \EE4BEG_i[8] ;
 wire \EE4BEG_i[9] ;
 wire \FrameData_O_i[0] ;
 wire \FrameData_O_i[10] ;
 wire \FrameData_O_i[11] ;
 wire \FrameData_O_i[12] ;
 wire \FrameData_O_i[13] ;
 wire \FrameData_O_i[14] ;
 wire \FrameData_O_i[15] ;
 wire \FrameData_O_i[16] ;
 wire \FrameData_O_i[17] ;
 wire \FrameData_O_i[18] ;
 wire \FrameData_O_i[19] ;
 wire \FrameData_O_i[1] ;
 wire \FrameData_O_i[20] ;
 wire \FrameData_O_i[21] ;
 wire \FrameData_O_i[22] ;
 wire \FrameData_O_i[23] ;
 wire \FrameData_O_i[24] ;
 wire \FrameData_O_i[25] ;
 wire \FrameData_O_i[26] ;
 wire \FrameData_O_i[27] ;
 wire \FrameData_O_i[28] ;
 wire \FrameData_O_i[29] ;
 wire \FrameData_O_i[2] ;
 wire \FrameData_O_i[30] ;
 wire \FrameData_O_i[31] ;
 wire \FrameData_O_i[3] ;
 wire \FrameData_O_i[4] ;
 wire \FrameData_O_i[5] ;
 wire \FrameData_O_i[6] ;
 wire \FrameData_O_i[7] ;
 wire \FrameData_O_i[8] ;
 wire \FrameData_O_i[9] ;
 wire \FrameStrobe_O_i[0] ;
 wire \FrameStrobe_O_i[10] ;
 wire \FrameStrobe_O_i[11] ;
 wire \FrameStrobe_O_i[12] ;
 wire \FrameStrobe_O_i[13] ;
 wire \FrameStrobe_O_i[14] ;
 wire \FrameStrobe_O_i[15] ;
 wire \FrameStrobe_O_i[16] ;
 wire \FrameStrobe_O_i[17] ;
 wire \FrameStrobe_O_i[18] ;
 wire \FrameStrobe_O_i[19] ;
 wire \FrameStrobe_O_i[1] ;
 wire \FrameStrobe_O_i[2] ;
 wire \FrameStrobe_O_i[3] ;
 wire \FrameStrobe_O_i[4] ;
 wire \FrameStrobe_O_i[5] ;
 wire \FrameStrobe_O_i[6] ;
 wire \FrameStrobe_O_i[7] ;
 wire \FrameStrobe_O_i[8] ;
 wire \FrameStrobe_O_i[9] ;
 wire \Inst_RegFile_32x4/AD_comb[0] ;
 wire \Inst_RegFile_32x4/AD_comb[1] ;
 wire \Inst_RegFile_32x4/AD_comb[2] ;
 wire \Inst_RegFile_32x4/AD_comb[3] ;
 wire \Inst_RegFile_32x4/AD_reg[0] ;
 wire \Inst_RegFile_32x4/AD_reg[1] ;
 wire \Inst_RegFile_32x4/AD_reg[2] ;
 wire \Inst_RegFile_32x4/AD_reg[3] ;
 wire \Inst_RegFile_32x4/BD_comb[0] ;
 wire \Inst_RegFile_32x4/BD_comb[1] ;
 wire \Inst_RegFile_32x4/BD_comb[2] ;
 wire \Inst_RegFile_32x4/BD_comb[3] ;
 wire \Inst_RegFile_32x4/BD_reg[0] ;
 wire \Inst_RegFile_32x4/BD_reg[1] ;
 wire \Inst_RegFile_32x4/BD_reg[2] ;
 wire \Inst_RegFile_32x4/BD_reg[3] ;
 wire \Inst_RegFile_32x4/_0000_ ;
 wire \Inst_RegFile_32x4/_0001_ ;
 wire \Inst_RegFile_32x4/_0002_ ;
 wire \Inst_RegFile_32x4/_0003_ ;
 wire \Inst_RegFile_32x4/_0004_ ;
 wire \Inst_RegFile_32x4/_0005_ ;
 wire \Inst_RegFile_32x4/_0006_ ;
 wire \Inst_RegFile_32x4/_0007_ ;
 wire \Inst_RegFile_32x4/_0008_ ;
 wire \Inst_RegFile_32x4/_0009_ ;
 wire \Inst_RegFile_32x4/_0010_ ;
 wire \Inst_RegFile_32x4/_0011_ ;
 wire \Inst_RegFile_32x4/_0012_ ;
 wire \Inst_RegFile_32x4/_0013_ ;
 wire \Inst_RegFile_32x4/_0014_ ;
 wire \Inst_RegFile_32x4/_0015_ ;
 wire \Inst_RegFile_32x4/_0016_ ;
 wire \Inst_RegFile_32x4/_0017_ ;
 wire \Inst_RegFile_32x4/_0018_ ;
 wire \Inst_RegFile_32x4/_0019_ ;
 wire \Inst_RegFile_32x4/_0020_ ;
 wire \Inst_RegFile_32x4/_0021_ ;
 wire \Inst_RegFile_32x4/_0022_ ;
 wire \Inst_RegFile_32x4/_0023_ ;
 wire \Inst_RegFile_32x4/_0024_ ;
 wire \Inst_RegFile_32x4/_0025_ ;
 wire \Inst_RegFile_32x4/_0026_ ;
 wire \Inst_RegFile_32x4/_0027_ ;
 wire \Inst_RegFile_32x4/_0028_ ;
 wire \Inst_RegFile_32x4/_0029_ ;
 wire \Inst_RegFile_32x4/_0030_ ;
 wire \Inst_RegFile_32x4/_0031_ ;
 wire \Inst_RegFile_32x4/_0032_ ;
 wire \Inst_RegFile_32x4/_0033_ ;
 wire \Inst_RegFile_32x4/_0034_ ;
 wire \Inst_RegFile_32x4/_0035_ ;
 wire \Inst_RegFile_32x4/_0036_ ;
 wire \Inst_RegFile_32x4/_0037_ ;
 wire \Inst_RegFile_32x4/_0038_ ;
 wire \Inst_RegFile_32x4/_0039_ ;
 wire \Inst_RegFile_32x4/_0040_ ;
 wire \Inst_RegFile_32x4/_0041_ ;
 wire \Inst_RegFile_32x4/_0042_ ;
 wire \Inst_RegFile_32x4/_0043_ ;
 wire \Inst_RegFile_32x4/_0044_ ;
 wire \Inst_RegFile_32x4/_0045_ ;
 wire \Inst_RegFile_32x4/_0046_ ;
 wire \Inst_RegFile_32x4/_0047_ ;
 wire \Inst_RegFile_32x4/_0048_ ;
 wire \Inst_RegFile_32x4/_0049_ ;
 wire \Inst_RegFile_32x4/_0050_ ;
 wire \Inst_RegFile_32x4/_0051_ ;
 wire \Inst_RegFile_32x4/_0052_ ;
 wire \Inst_RegFile_32x4/_0053_ ;
 wire \Inst_RegFile_32x4/_0054_ ;
 wire \Inst_RegFile_32x4/_0055_ ;
 wire \Inst_RegFile_32x4/_0056_ ;
 wire \Inst_RegFile_32x4/_0057_ ;
 wire \Inst_RegFile_32x4/_0058_ ;
 wire \Inst_RegFile_32x4/_0059_ ;
 wire \Inst_RegFile_32x4/_0060_ ;
 wire \Inst_RegFile_32x4/_0061_ ;
 wire \Inst_RegFile_32x4/_0062_ ;
 wire \Inst_RegFile_32x4/_0063_ ;
 wire \Inst_RegFile_32x4/_0064_ ;
 wire \Inst_RegFile_32x4/_0065_ ;
 wire \Inst_RegFile_32x4/_0066_ ;
 wire \Inst_RegFile_32x4/_0067_ ;
 wire \Inst_RegFile_32x4/_0068_ ;
 wire \Inst_RegFile_32x4/_0069_ ;
 wire \Inst_RegFile_32x4/_0070_ ;
 wire \Inst_RegFile_32x4/_0071_ ;
 wire \Inst_RegFile_32x4/_0072_ ;
 wire \Inst_RegFile_32x4/_0073_ ;
 wire \Inst_RegFile_32x4/_0074_ ;
 wire \Inst_RegFile_32x4/_0075_ ;
 wire \Inst_RegFile_32x4/_0076_ ;
 wire \Inst_RegFile_32x4/_0077_ ;
 wire \Inst_RegFile_32x4/_0078_ ;
 wire \Inst_RegFile_32x4/_0079_ ;
 wire \Inst_RegFile_32x4/_0080_ ;
 wire \Inst_RegFile_32x4/_0081_ ;
 wire \Inst_RegFile_32x4/_0082_ ;
 wire \Inst_RegFile_32x4/_0083_ ;
 wire \Inst_RegFile_32x4/_0084_ ;
 wire \Inst_RegFile_32x4/_0085_ ;
 wire \Inst_RegFile_32x4/_0086_ ;
 wire \Inst_RegFile_32x4/_0087_ ;
 wire \Inst_RegFile_32x4/_0088_ ;
 wire \Inst_RegFile_32x4/_0089_ ;
 wire \Inst_RegFile_32x4/_0090_ ;
 wire \Inst_RegFile_32x4/_0091_ ;
 wire \Inst_RegFile_32x4/_0092_ ;
 wire \Inst_RegFile_32x4/_0093_ ;
 wire \Inst_RegFile_32x4/_0094_ ;
 wire \Inst_RegFile_32x4/_0095_ ;
 wire \Inst_RegFile_32x4/_0096_ ;
 wire \Inst_RegFile_32x4/_0097_ ;
 wire \Inst_RegFile_32x4/_0098_ ;
 wire \Inst_RegFile_32x4/_0099_ ;
 wire \Inst_RegFile_32x4/_0100_ ;
 wire \Inst_RegFile_32x4/_0101_ ;
 wire \Inst_RegFile_32x4/_0102_ ;
 wire \Inst_RegFile_32x4/_0103_ ;
 wire \Inst_RegFile_32x4/_0104_ ;
 wire \Inst_RegFile_32x4/_0105_ ;
 wire \Inst_RegFile_32x4/_0106_ ;
 wire \Inst_RegFile_32x4/_0107_ ;
 wire \Inst_RegFile_32x4/_0108_ ;
 wire \Inst_RegFile_32x4/_0109_ ;
 wire \Inst_RegFile_32x4/_0110_ ;
 wire \Inst_RegFile_32x4/_0111_ ;
 wire \Inst_RegFile_32x4/_0112_ ;
 wire \Inst_RegFile_32x4/_0113_ ;
 wire \Inst_RegFile_32x4/_0114_ ;
 wire \Inst_RegFile_32x4/_0115_ ;
 wire \Inst_RegFile_32x4/_0116_ ;
 wire \Inst_RegFile_32x4/_0117_ ;
 wire \Inst_RegFile_32x4/_0118_ ;
 wire \Inst_RegFile_32x4/_0119_ ;
 wire \Inst_RegFile_32x4/_0120_ ;
 wire \Inst_RegFile_32x4/_0121_ ;
 wire \Inst_RegFile_32x4/_0122_ ;
 wire \Inst_RegFile_32x4/_0123_ ;
 wire \Inst_RegFile_32x4/_0124_ ;
 wire \Inst_RegFile_32x4/_0125_ ;
 wire \Inst_RegFile_32x4/_0126_ ;
 wire \Inst_RegFile_32x4/_0127_ ;
 wire \Inst_RegFile_32x4/_0128_ ;
 wire \Inst_RegFile_32x4/_0129_ ;
 wire \Inst_RegFile_32x4/_0130_ ;
 wire \Inst_RegFile_32x4/_0131_ ;
 wire \Inst_RegFile_32x4/_0132_ ;
 wire \Inst_RegFile_32x4/_0133_ ;
 wire \Inst_RegFile_32x4/_0134_ ;
 wire \Inst_RegFile_32x4/_0135_ ;
 wire \Inst_RegFile_32x4/_0136_ ;
 wire \Inst_RegFile_32x4/_0137_ ;
 wire \Inst_RegFile_32x4/_0138_ ;
 wire \Inst_RegFile_32x4/_0139_ ;
 wire \Inst_RegFile_32x4/_0140_ ;
 wire \Inst_RegFile_32x4/_0141_ ;
 wire \Inst_RegFile_32x4/_0142_ ;
 wire \Inst_RegFile_32x4/_0143_ ;
 wire \Inst_RegFile_32x4/_0144_ ;
 wire \Inst_RegFile_32x4/_0145_ ;
 wire \Inst_RegFile_32x4/_0146_ ;
 wire \Inst_RegFile_32x4/_0147_ ;
 wire \Inst_RegFile_32x4/_0148_ ;
 wire \Inst_RegFile_32x4/_0149_ ;
 wire \Inst_RegFile_32x4/_0150_ ;
 wire \Inst_RegFile_32x4/_0151_ ;
 wire \Inst_RegFile_32x4/_0152_ ;
 wire \Inst_RegFile_32x4/_0153_ ;
 wire \Inst_RegFile_32x4/_0154_ ;
 wire \Inst_RegFile_32x4/_0155_ ;
 wire \Inst_RegFile_32x4/_0156_ ;
 wire \Inst_RegFile_32x4/_0157_ ;
 wire \Inst_RegFile_32x4/_0158_ ;
 wire \Inst_RegFile_32x4/_0159_ ;
 wire \Inst_RegFile_32x4/_0160_ ;
 wire \Inst_RegFile_32x4/_0161_ ;
 wire \Inst_RegFile_32x4/_0162_ ;
 wire \Inst_RegFile_32x4/_0163_ ;
 wire \Inst_RegFile_32x4/_0164_ ;
 wire \Inst_RegFile_32x4/_0165_ ;
 wire \Inst_RegFile_32x4/_0166_ ;
 wire \Inst_RegFile_32x4/_0167_ ;
 wire \Inst_RegFile_32x4/_0168_ ;
 wire \Inst_RegFile_32x4/_0169_ ;
 wire \Inst_RegFile_32x4/_0170_ ;
 wire \Inst_RegFile_32x4/_0171_ ;
 wire \Inst_RegFile_32x4/_0172_ ;
 wire \Inst_RegFile_32x4/_0173_ ;
 wire \Inst_RegFile_32x4/_0174_ ;
 wire \Inst_RegFile_32x4/_0175_ ;
 wire \Inst_RegFile_32x4/_0176_ ;
 wire \Inst_RegFile_32x4/_0177_ ;
 wire \Inst_RegFile_32x4/_0178_ ;
 wire \Inst_RegFile_32x4/_0179_ ;
 wire \Inst_RegFile_32x4/_0180_ ;
 wire \Inst_RegFile_32x4/_0181_ ;
 wire \Inst_RegFile_32x4/_0182_ ;
 wire \Inst_RegFile_32x4/_0183_ ;
 wire \Inst_RegFile_32x4/_0184_ ;
 wire \Inst_RegFile_32x4/_0185_ ;
 wire \Inst_RegFile_32x4/_0186_ ;
 wire \Inst_RegFile_32x4/_0187_ ;
 wire \Inst_RegFile_32x4/_0188_ ;
 wire \Inst_RegFile_32x4/_0189_ ;
 wire \Inst_RegFile_32x4/_0190_ ;
 wire \Inst_RegFile_32x4/_0191_ ;
 wire \Inst_RegFile_32x4/_0192_ ;
 wire \Inst_RegFile_32x4/_0193_ ;
 wire \Inst_RegFile_32x4/_0194_ ;
 wire \Inst_RegFile_32x4/_0195_ ;
 wire \Inst_RegFile_32x4/_0196_ ;
 wire \Inst_RegFile_32x4/_0197_ ;
 wire \Inst_RegFile_32x4/_0198_ ;
 wire \Inst_RegFile_32x4/_0199_ ;
 wire \Inst_RegFile_32x4/_0200_ ;
 wire \Inst_RegFile_32x4/_0201_ ;
 wire \Inst_RegFile_32x4/_0202_ ;
 wire \Inst_RegFile_32x4/_0203_ ;
 wire \Inst_RegFile_32x4/_0204_ ;
 wire \Inst_RegFile_32x4/_0205_ ;
 wire \Inst_RegFile_32x4/_0206_ ;
 wire \Inst_RegFile_32x4/_0207_ ;
 wire \Inst_RegFile_32x4/_0208_ ;
 wire \Inst_RegFile_32x4/_0209_ ;
 wire \Inst_RegFile_32x4/_0210_ ;
 wire \Inst_RegFile_32x4/_0211_ ;
 wire \Inst_RegFile_32x4/_0212_ ;
 wire \Inst_RegFile_32x4/_0213_ ;
 wire \Inst_RegFile_32x4/_0214_ ;
 wire \Inst_RegFile_32x4/_0215_ ;
 wire \Inst_RegFile_32x4/_0216_ ;
 wire \Inst_RegFile_32x4/_0217_ ;
 wire \Inst_RegFile_32x4/_0218_ ;
 wire \Inst_RegFile_32x4/_0219_ ;
 wire \Inst_RegFile_32x4/_0220_ ;
 wire \Inst_RegFile_32x4/_0221_ ;
 wire \Inst_RegFile_32x4/_0222_ ;
 wire \Inst_RegFile_32x4/_0223_ ;
 wire \Inst_RegFile_32x4/_0224_ ;
 wire \Inst_RegFile_32x4/_0225_ ;
 wire \Inst_RegFile_32x4/_0226_ ;
 wire \Inst_RegFile_32x4/_0227_ ;
 wire \Inst_RegFile_32x4/_0228_ ;
 wire \Inst_RegFile_32x4/_0229_ ;
 wire \Inst_RegFile_32x4/_0230_ ;
 wire \Inst_RegFile_32x4/_0231_ ;
 wire \Inst_RegFile_32x4/_0232_ ;
 wire \Inst_RegFile_32x4/_0233_ ;
 wire \Inst_RegFile_32x4/_0234_ ;
 wire \Inst_RegFile_32x4/_0235_ ;
 wire \Inst_RegFile_32x4/_0236_ ;
 wire \Inst_RegFile_32x4/_0237_ ;
 wire \Inst_RegFile_32x4/_0238_ ;
 wire \Inst_RegFile_32x4/_0239_ ;
 wire \Inst_RegFile_32x4/_0240_ ;
 wire \Inst_RegFile_32x4/_0241_ ;
 wire \Inst_RegFile_32x4/_0242_ ;
 wire \Inst_RegFile_32x4/_0243_ ;
 wire \Inst_RegFile_32x4/_0244_ ;
 wire \Inst_RegFile_32x4/_0245_ ;
 wire \Inst_RegFile_32x4/_0246_ ;
 wire \Inst_RegFile_32x4/_0247_ ;
 wire \Inst_RegFile_32x4/_0248_ ;
 wire \Inst_RegFile_32x4/_0249_ ;
 wire \Inst_RegFile_32x4/_0250_ ;
 wire \Inst_RegFile_32x4/_0251_ ;
 wire \Inst_RegFile_32x4/_0252_ ;
 wire \Inst_RegFile_32x4/_0253_ ;
 wire \Inst_RegFile_32x4/_0254_ ;
 wire \Inst_RegFile_32x4/_0255_ ;
 wire \Inst_RegFile_32x4/_0256_ ;
 wire \Inst_RegFile_32x4/_0257_ ;
 wire \Inst_RegFile_32x4/_0258_ ;
 wire \Inst_RegFile_32x4/_0259_ ;
 wire \Inst_RegFile_32x4/_0260_ ;
 wire \Inst_RegFile_32x4/_0261_ ;
 wire \Inst_RegFile_32x4/_0262_ ;
 wire \Inst_RegFile_32x4/_0263_ ;
 wire \Inst_RegFile_32x4/_0264_ ;
 wire \Inst_RegFile_32x4/_0265_ ;
 wire \Inst_RegFile_32x4/_0266_ ;
 wire \Inst_RegFile_32x4/_0267_ ;
 wire \Inst_RegFile_32x4/_0268_ ;
 wire \Inst_RegFile_32x4/_0269_ ;
 wire \Inst_RegFile_32x4/_0270_ ;
 wire \Inst_RegFile_32x4/_0271_ ;
 wire \Inst_RegFile_32x4/_0272_ ;
 wire \Inst_RegFile_32x4/_0273_ ;
 wire \Inst_RegFile_32x4/_0274_ ;
 wire \Inst_RegFile_32x4/_0275_ ;
 wire \Inst_RegFile_32x4/_0276_ ;
 wire \Inst_RegFile_32x4/_0277_ ;
 wire \Inst_RegFile_32x4/_0278_ ;
 wire \Inst_RegFile_32x4/_0279_ ;
 wire \Inst_RegFile_32x4/_0280_ ;
 wire \Inst_RegFile_32x4/_0281_ ;
 wire \Inst_RegFile_32x4/_0282_ ;
 wire \Inst_RegFile_32x4/_0283_ ;
 wire \Inst_RegFile_32x4/_0284_ ;
 wire \Inst_RegFile_32x4/_0285_ ;
 wire \Inst_RegFile_32x4/_0286_ ;
 wire \Inst_RegFile_32x4/_0287_ ;
 wire \Inst_RegFile_32x4/_0288_ ;
 wire \Inst_RegFile_32x4/_0289_ ;
 wire \Inst_RegFile_32x4/_0290_ ;
 wire \Inst_RegFile_32x4/_0291_ ;
 wire \Inst_RegFile_32x4/_0292_ ;
 wire \Inst_RegFile_32x4/_0293_ ;
 wire \Inst_RegFile_32x4/_0294_ ;
 wire \Inst_RegFile_32x4/_0295_ ;
 wire \Inst_RegFile_32x4/_0296_ ;
 wire \Inst_RegFile_32x4/_0297_ ;
 wire \Inst_RegFile_32x4/_0298_ ;
 wire \Inst_RegFile_32x4/_0299_ ;
 wire \Inst_RegFile_32x4/_0300_ ;
 wire \Inst_RegFile_32x4/_0301_ ;
 wire \Inst_RegFile_32x4/_0302_ ;
 wire \Inst_RegFile_32x4/_0303_ ;
 wire \Inst_RegFile_32x4/_0304_ ;
 wire \Inst_RegFile_32x4/_0305_ ;
 wire \Inst_RegFile_32x4/_0306_ ;
 wire \Inst_RegFile_32x4/_0307_ ;
 wire \Inst_RegFile_32x4/_0308_ ;
 wire \Inst_RegFile_32x4/_0309_ ;
 wire \Inst_RegFile_32x4/_0310_ ;
 wire \Inst_RegFile_32x4/_0311_ ;
 wire \Inst_RegFile_32x4/_0312_ ;
 wire \Inst_RegFile_32x4/_0313_ ;
 wire \Inst_RegFile_32x4/_0314_ ;
 wire \Inst_RegFile_32x4/_0315_ ;
 wire \Inst_RegFile_32x4/_0316_ ;
 wire \Inst_RegFile_32x4/_0317_ ;
 wire \Inst_RegFile_32x4/_0318_ ;
 wire \Inst_RegFile_32x4/_0319_ ;
 wire \Inst_RegFile_32x4/_0320_ ;
 wire \Inst_RegFile_32x4/_0321_ ;
 wire \Inst_RegFile_32x4/_0322_ ;
 wire \Inst_RegFile_32x4/_0323_ ;
 wire \Inst_RegFile_32x4/_0324_ ;
 wire \Inst_RegFile_32x4/_0325_ ;
 wire \Inst_RegFile_32x4/_0326_ ;
 wire \Inst_RegFile_32x4/_0327_ ;
 wire \Inst_RegFile_32x4/_0328_ ;
 wire \Inst_RegFile_32x4/_0329_ ;
 wire \Inst_RegFile_32x4/_0330_ ;
 wire \Inst_RegFile_32x4/_0331_ ;
 wire \Inst_RegFile_32x4/_0332_ ;
 wire \Inst_RegFile_32x4/_0333_ ;
 wire \Inst_RegFile_32x4/_0334_ ;
 wire \Inst_RegFile_32x4/_0335_ ;
 wire \Inst_RegFile_32x4/_0336_ ;
 wire \Inst_RegFile_32x4/_0337_ ;
 wire \Inst_RegFile_32x4/_0338_ ;
 wire \Inst_RegFile_32x4/_0339_ ;
 wire \Inst_RegFile_32x4/_0340_ ;
 wire \Inst_RegFile_32x4/_0341_ ;
 wire \Inst_RegFile_32x4/_0342_ ;
 wire \Inst_RegFile_32x4/_0343_ ;
 wire \Inst_RegFile_32x4/_0344_ ;
 wire \Inst_RegFile_32x4/_0345_ ;
 wire \Inst_RegFile_32x4/_0346_ ;
 wire \Inst_RegFile_32x4/_0347_ ;
 wire \Inst_RegFile_32x4/_0348_ ;
 wire \Inst_RegFile_32x4/_0349_ ;
 wire \Inst_RegFile_32x4/_0350_ ;
 wire \Inst_RegFile_32x4/_0351_ ;
 wire \Inst_RegFile_32x4/_0352_ ;
 wire \Inst_RegFile_32x4/_0353_ ;
 wire \Inst_RegFile_32x4/_0354_ ;
 wire \Inst_RegFile_32x4/_0355_ ;
 wire \Inst_RegFile_32x4/_0356_ ;
 wire \Inst_RegFile_32x4/_0357_ ;
 wire \Inst_RegFile_32x4/_0358_ ;
 wire \Inst_RegFile_32x4/_0359_ ;
 wire \Inst_RegFile_32x4/_0360_ ;
 wire \Inst_RegFile_32x4/_0361_ ;
 wire \Inst_RegFile_32x4/_0362_ ;
 wire \Inst_RegFile_32x4/_0363_ ;
 wire \Inst_RegFile_32x4/_0364_ ;
 wire \Inst_RegFile_32x4/_0365_ ;
 wire \Inst_RegFile_32x4/_0366_ ;
 wire \Inst_RegFile_32x4/_0367_ ;
 wire \Inst_RegFile_32x4/_0368_ ;
 wire \Inst_RegFile_32x4/_0369_ ;
 wire \Inst_RegFile_32x4/_0370_ ;
 wire \Inst_RegFile_32x4/_0371_ ;
 wire \Inst_RegFile_32x4/_0372_ ;
 wire \Inst_RegFile_32x4/_0373_ ;
 wire \Inst_RegFile_32x4/_0374_ ;
 wire \Inst_RegFile_32x4/_0375_ ;
 wire \Inst_RegFile_32x4/_0376_ ;
 wire \Inst_RegFile_32x4/_0377_ ;
 wire \Inst_RegFile_32x4/_0378_ ;
 wire \Inst_RegFile_32x4/_0379_ ;
 wire \Inst_RegFile_32x4/_0380_ ;
 wire \Inst_RegFile_32x4/_0381_ ;
 wire \Inst_RegFile_32x4/_0382_ ;
 wire \Inst_RegFile_32x4/_0383_ ;
 wire \Inst_RegFile_32x4/_0384_ ;
 wire \Inst_RegFile_32x4/_0385_ ;
 wire \Inst_RegFile_32x4/_0386_ ;
 wire \Inst_RegFile_32x4/_0387_ ;
 wire \Inst_RegFile_32x4/_0388_ ;
 wire \Inst_RegFile_32x4/_0389_ ;
 wire \Inst_RegFile_32x4/_0390_ ;
 wire \Inst_RegFile_32x4/_0391_ ;
 wire \Inst_RegFile_32x4/_0392_ ;
 wire \Inst_RegFile_32x4/_0393_ ;
 wire \Inst_RegFile_32x4/_0394_ ;
 wire \Inst_RegFile_32x4/_0395_ ;
 wire \Inst_RegFile_32x4/_0396_ ;
 wire \Inst_RegFile_32x4/_0397_ ;
 wire \Inst_RegFile_32x4/_0398_ ;
 wire \Inst_RegFile_32x4/_0399_ ;
 wire \Inst_RegFile_32x4/_0400_ ;
 wire \Inst_RegFile_32x4/_0401_ ;
 wire \Inst_RegFile_32x4/_0402_ ;
 wire \Inst_RegFile_32x4/_0403_ ;
 wire \Inst_RegFile_32x4/_0404_ ;
 wire \Inst_RegFile_32x4/_0405_ ;
 wire \Inst_RegFile_32x4/_0406_ ;
 wire \Inst_RegFile_32x4/_0407_ ;
 wire \Inst_RegFile_32x4/_0408_ ;
 wire \Inst_RegFile_32x4/_0409_ ;
 wire \Inst_RegFile_32x4/_0410_ ;
 wire \Inst_RegFile_32x4/_0411_ ;
 wire \Inst_RegFile_32x4/_0412_ ;
 wire \Inst_RegFile_32x4/_0413_ ;
 wire \Inst_RegFile_32x4/_0414_ ;
 wire \Inst_RegFile_32x4/_0415_ ;
 wire \Inst_RegFile_32x4/_0416_ ;
 wire \Inst_RegFile_32x4/_0417_ ;
 wire \Inst_RegFile_32x4/_0418_ ;
 wire \Inst_RegFile_32x4/_0419_ ;
 wire \Inst_RegFile_32x4/_0420_ ;
 wire \Inst_RegFile_32x4/_0421_ ;
 wire \Inst_RegFile_32x4/_0422_ ;
 wire \Inst_RegFile_32x4/_0423_ ;
 wire \Inst_RegFile_32x4/_0424_ ;
 wire \Inst_RegFile_32x4/_0425_ ;
 wire \Inst_RegFile_32x4/_0426_ ;
 wire \Inst_RegFile_32x4/_0427_ ;
 wire \Inst_RegFile_32x4/_0428_ ;
 wire \Inst_RegFile_32x4/_0429_ ;
 wire \Inst_RegFile_32x4/_0430_ ;
 wire \Inst_RegFile_32x4/_0431_ ;
 wire \Inst_RegFile_32x4/_0432_ ;
 wire \Inst_RegFile_32x4/_0433_ ;
 wire \Inst_RegFile_32x4/_0434_ ;
 wire \Inst_RegFile_32x4/_0435_ ;
 wire \Inst_RegFile_32x4/_0436_ ;
 wire \Inst_RegFile_32x4/_0437_ ;
 wire \Inst_RegFile_32x4/_0438_ ;
 wire \Inst_RegFile_32x4/_0439_ ;
 wire \Inst_RegFile_32x4/_0440_ ;
 wire \Inst_RegFile_32x4/_0441_ ;
 wire \Inst_RegFile_32x4/_0442_ ;
 wire \Inst_RegFile_32x4/_0443_ ;
 wire \Inst_RegFile_32x4/_0444_ ;
 wire \Inst_RegFile_32x4/_0445_ ;
 wire \Inst_RegFile_32x4/_0446_ ;
 wire \Inst_RegFile_32x4/_0447_ ;
 wire \Inst_RegFile_32x4/_0448_ ;
 wire \Inst_RegFile_32x4/_0449_ ;
 wire \Inst_RegFile_32x4/_0450_ ;
 wire \Inst_RegFile_32x4/_0451_ ;
 wire \Inst_RegFile_32x4/_0452_ ;
 wire \Inst_RegFile_32x4/_0453_ ;
 wire \Inst_RegFile_32x4/_0454_ ;
 wire \Inst_RegFile_32x4/_0455_ ;
 wire \Inst_RegFile_32x4/_0456_ ;
 wire \Inst_RegFile_32x4/_0457_ ;
 wire \Inst_RegFile_32x4/_0458_ ;
 wire \Inst_RegFile_32x4/_0459_ ;
 wire \Inst_RegFile_32x4/_0460_ ;
 wire \Inst_RegFile_32x4/_0461_ ;
 wire \Inst_RegFile_32x4/_0462_ ;
 wire \Inst_RegFile_32x4/_0463_ ;
 wire \Inst_RegFile_32x4/_0464_ ;
 wire \Inst_RegFile_32x4/_0465_ ;
 wire \Inst_RegFile_32x4/_0466_ ;
 wire \Inst_RegFile_32x4/_0467_ ;
 wire \Inst_RegFile_32x4/_0468_ ;
 wire \Inst_RegFile_32x4/_0469_ ;
 wire \Inst_RegFile_32x4/_0470_ ;
 wire \Inst_RegFile_32x4/_0471_ ;
 wire \Inst_RegFile_32x4/_0472_ ;
 wire \Inst_RegFile_32x4/_0473_ ;
 wire \Inst_RegFile_32x4/_0474_ ;
 wire \Inst_RegFile_32x4/_0475_ ;
 wire \Inst_RegFile_32x4/_0476_ ;
 wire \Inst_RegFile_32x4/_0477_ ;
 wire \Inst_RegFile_32x4/_0478_ ;
 wire \Inst_RegFile_32x4/_0479_ ;
 wire \Inst_RegFile_32x4/_0480_ ;
 wire \Inst_RegFile_32x4/_0481_ ;
 wire \Inst_RegFile_32x4/_0482_ ;
 wire \Inst_RegFile_32x4/_0483_ ;
 wire \Inst_RegFile_32x4/_0484_ ;
 wire \Inst_RegFile_32x4/_0485_ ;
 wire \Inst_RegFile_32x4/_0486_ ;
 wire \Inst_RegFile_32x4/_0487_ ;
 wire \Inst_RegFile_32x4/_0488_ ;
 wire \Inst_RegFile_32x4/_0489_ ;
 wire \Inst_RegFile_32x4/_0490_ ;
 wire \Inst_RegFile_32x4/_0491_ ;
 wire \Inst_RegFile_32x4/_0492_ ;
 wire \Inst_RegFile_32x4/_0493_ ;
 wire \Inst_RegFile_32x4/_0494_ ;
 wire \Inst_RegFile_32x4/_0495_ ;
 wire \Inst_RegFile_32x4/_0496_ ;
 wire \Inst_RegFile_32x4/_0497_ ;
 wire \Inst_RegFile_32x4/_0498_ ;
 wire \Inst_RegFile_32x4/_0499_ ;
 wire \Inst_RegFile_32x4/_0500_ ;
 wire \Inst_RegFile_32x4/_0501_ ;
 wire \Inst_RegFile_32x4/_0502_ ;
 wire \Inst_RegFile_32x4/_0503_ ;
 wire \Inst_RegFile_32x4/_0504_ ;
 wire \Inst_RegFile_32x4/_0505_ ;
 wire \Inst_RegFile_32x4/_0506_ ;
 wire \Inst_RegFile_32x4/_0507_ ;
 wire \Inst_RegFile_32x4/_0508_ ;
 wire \Inst_RegFile_32x4/_0509_ ;
 wire \Inst_RegFile_32x4/_0510_ ;
 wire \Inst_RegFile_32x4/_0511_ ;
 wire \Inst_RegFile_32x4/_0512_ ;
 wire \Inst_RegFile_32x4/_0513_ ;
 wire \Inst_RegFile_32x4/_0514_ ;
 wire \Inst_RegFile_32x4/_0515_ ;
 wire \Inst_RegFile_32x4/_0516_ ;
 wire \Inst_RegFile_32x4/_0517_ ;
 wire \Inst_RegFile_32x4/_0518_ ;
 wire \Inst_RegFile_32x4/_0519_ ;
 wire \Inst_RegFile_32x4/_0520_ ;
 wire \Inst_RegFile_32x4/_0521_ ;
 wire \Inst_RegFile_32x4/_0522_ ;
 wire \Inst_RegFile_32x4/_0523_ ;
 wire \Inst_RegFile_32x4/_0524_ ;
 wire \Inst_RegFile_32x4/_0525_ ;
 wire \Inst_RegFile_32x4/_0526_ ;
 wire \Inst_RegFile_32x4/_0527_ ;
 wire \Inst_RegFile_32x4/_0528_ ;
 wire \Inst_RegFile_32x4/_0529_ ;
 wire \Inst_RegFile_32x4/_0530_ ;
 wire \Inst_RegFile_32x4/_0531_ ;
 wire \Inst_RegFile_32x4/_0532_ ;
 wire \Inst_RegFile_32x4/_0533_ ;
 wire \Inst_RegFile_32x4/_0534_ ;
 wire \Inst_RegFile_32x4/_0535_ ;
 wire \Inst_RegFile_32x4/_0536_ ;
 wire \Inst_RegFile_32x4/_0537_ ;
 wire \Inst_RegFile_32x4/_0538_ ;
 wire \Inst_RegFile_32x4/_0539_ ;
 wire \Inst_RegFile_32x4/_0540_ ;
 wire \Inst_RegFile_32x4/_0541_ ;
 wire \Inst_RegFile_32x4/_0542_ ;
 wire \Inst_RegFile_32x4/_0543_ ;
 wire \Inst_RegFile_32x4/_0544_ ;
 wire \Inst_RegFile_32x4/_0545_ ;
 wire \Inst_RegFile_32x4/_0546_ ;
 wire \Inst_RegFile_32x4/_0547_ ;
 wire \Inst_RegFile_32x4/_0548_ ;
 wire \Inst_RegFile_32x4/_0549_ ;
 wire \Inst_RegFile_32x4/_0550_ ;
 wire \Inst_RegFile_32x4/_0551_ ;
 wire \Inst_RegFile_32x4/_0552_ ;
 wire \Inst_RegFile_32x4/_0553_ ;
 wire \Inst_RegFile_32x4/_0554_ ;
 wire \Inst_RegFile_32x4/_0555_ ;
 wire \Inst_RegFile_32x4/_0556_ ;
 wire \Inst_RegFile_32x4/_0557_ ;
 wire \Inst_RegFile_32x4/_0558_ ;
 wire \Inst_RegFile_32x4/_0559_ ;
 wire \Inst_RegFile_32x4/_0560_ ;
 wire \Inst_RegFile_32x4/_0561_ ;
 wire \Inst_RegFile_32x4/_0562_ ;
 wire \Inst_RegFile_32x4/_0563_ ;
 wire \Inst_RegFile_32x4/_0564_ ;
 wire \Inst_RegFile_32x4/_0565_ ;
 wire \Inst_RegFile_32x4/_0566_ ;
 wire \Inst_RegFile_32x4/_0567_ ;
 wire \Inst_RegFile_32x4/_0568_ ;
 wire \Inst_RegFile_32x4/_0569_ ;
 wire \Inst_RegFile_32x4/_0570_ ;
 wire \Inst_RegFile_32x4/_0571_ ;
 wire \Inst_RegFile_32x4/_0572_ ;
 wire \Inst_RegFile_32x4/_0573_ ;
 wire \Inst_RegFile_32x4/_0574_ ;
 wire \Inst_RegFile_32x4/_0575_ ;
 wire \Inst_RegFile_32x4/_0576_ ;
 wire \Inst_RegFile_32x4/_0577_ ;
 wire \Inst_RegFile_32x4/_0578_ ;
 wire \Inst_RegFile_32x4/_0579_ ;
 wire \Inst_RegFile_32x4/_0580_ ;
 wire \Inst_RegFile_32x4/_0581_ ;
 wire \Inst_RegFile_32x4/_0582_ ;
 wire \Inst_RegFile_32x4/_0583_ ;
 wire \Inst_RegFile_32x4/_0584_ ;
 wire \Inst_RegFile_32x4/_0585_ ;
 wire \Inst_RegFile_32x4/_0586_ ;
 wire \Inst_RegFile_32x4/_0587_ ;
 wire \Inst_RegFile_32x4/_0588_ ;
 wire \Inst_RegFile_32x4/_0589_ ;
 wire \Inst_RegFile_32x4/_0590_ ;
 wire \Inst_RegFile_32x4/_0591_ ;
 wire \Inst_RegFile_32x4/_0592_ ;
 wire \Inst_RegFile_32x4/_0593_ ;
 wire \Inst_RegFile_32x4/_0594_ ;
 wire \Inst_RegFile_32x4/_0595_ ;
 wire \Inst_RegFile_32x4/_0596_ ;
 wire \Inst_RegFile_32x4/_0597_ ;
 wire \Inst_RegFile_32x4/_0598_ ;
 wire \Inst_RegFile_32x4/_0599_ ;
 wire \Inst_RegFile_32x4/_0600_ ;
 wire \Inst_RegFile_32x4/_0601_ ;
 wire \Inst_RegFile_32x4/_0602_ ;
 wire \Inst_RegFile_32x4/_0603_ ;
 wire \Inst_RegFile_32x4/_0604_ ;
 wire \Inst_RegFile_32x4/_0605_ ;
 wire \Inst_RegFile_32x4/_0606_ ;
 wire \Inst_RegFile_32x4/_0607_ ;
 wire \Inst_RegFile_32x4/_0608_ ;
 wire \Inst_RegFile_32x4/_0609_ ;
 wire \Inst_RegFile_32x4/_0610_ ;
 wire \Inst_RegFile_32x4/_0611_ ;
 wire \Inst_RegFile_32x4/_0612_ ;
 wire \Inst_RegFile_32x4/_0613_ ;
 wire \Inst_RegFile_32x4/_0614_ ;
 wire \Inst_RegFile_32x4/_0615_ ;
 wire \Inst_RegFile_32x4/_0616_ ;
 wire \Inst_RegFile_32x4/_0617_ ;
 wire \Inst_RegFile_32x4/_0618_ ;
 wire \Inst_RegFile_32x4/_0619_ ;
 wire \Inst_RegFile_32x4/_0620_ ;
 wire \Inst_RegFile_32x4/_0621_ ;
 wire \Inst_RegFile_32x4/_0622_ ;
 wire \Inst_RegFile_32x4/_0623_ ;
 wire \Inst_RegFile_32x4/_0624_ ;
 wire \Inst_RegFile_32x4/_0625_ ;
 wire \Inst_RegFile_32x4/_0626_ ;
 wire \Inst_RegFile_32x4/_0627_ ;
 wire \Inst_RegFile_32x4/_0628_ ;
 wire \Inst_RegFile_32x4/_0629_ ;
 wire \Inst_RegFile_32x4/_0630_ ;
 wire \Inst_RegFile_32x4/_0631_ ;
 wire \Inst_RegFile_32x4/_0632_ ;
 wire \Inst_RegFile_32x4/_0633_ ;
 wire \Inst_RegFile_32x4/_0634_ ;
 wire \Inst_RegFile_32x4/_0635_ ;
 wire \Inst_RegFile_32x4/_0636_ ;
 wire \Inst_RegFile_32x4/_0637_ ;
 wire \Inst_RegFile_32x4/_0638_ ;
 wire \Inst_RegFile_32x4/_0639_ ;
 wire \Inst_RegFile_32x4/_0640_ ;
 wire \Inst_RegFile_32x4/_0641_ ;
 wire \Inst_RegFile_32x4/_0642_ ;
 wire \Inst_RegFile_32x4/_0643_ ;
 wire \Inst_RegFile_32x4/_0644_ ;
 wire \Inst_RegFile_32x4/_0645_ ;
 wire \Inst_RegFile_32x4/_0646_ ;
 wire \Inst_RegFile_32x4/_0647_ ;
 wire \Inst_RegFile_32x4/_0648_ ;
 wire \Inst_RegFile_32x4/_0649_ ;
 wire \Inst_RegFile_32x4/_0650_ ;
 wire \Inst_RegFile_32x4/_0651_ ;
 wire \Inst_RegFile_32x4/_0652_ ;
 wire \Inst_RegFile_32x4/_0653_ ;
 wire \Inst_RegFile_32x4/_0654_ ;
 wire \Inst_RegFile_32x4/_0655_ ;
 wire \Inst_RegFile_32x4/_0656_ ;
 wire \Inst_RegFile_32x4/_0657_ ;
 wire \Inst_RegFile_32x4/_0658_ ;
 wire \Inst_RegFile_32x4/_0659_ ;
 wire \Inst_RegFile_32x4/_0660_ ;
 wire \Inst_RegFile_32x4/_0661_ ;
 wire \Inst_RegFile_32x4/mem[0][0] ;
 wire \Inst_RegFile_32x4/mem[0][1] ;
 wire \Inst_RegFile_32x4/mem[0][2] ;
 wire \Inst_RegFile_32x4/mem[0][3] ;
 wire \Inst_RegFile_32x4/mem[10][0] ;
 wire \Inst_RegFile_32x4/mem[10][1] ;
 wire \Inst_RegFile_32x4/mem[10][2] ;
 wire \Inst_RegFile_32x4/mem[10][3] ;
 wire \Inst_RegFile_32x4/mem[11][0] ;
 wire \Inst_RegFile_32x4/mem[11][1] ;
 wire \Inst_RegFile_32x4/mem[11][2] ;
 wire \Inst_RegFile_32x4/mem[11][3] ;
 wire \Inst_RegFile_32x4/mem[12][0] ;
 wire \Inst_RegFile_32x4/mem[12][1] ;
 wire \Inst_RegFile_32x4/mem[12][2] ;
 wire \Inst_RegFile_32x4/mem[12][3] ;
 wire \Inst_RegFile_32x4/mem[13][0] ;
 wire \Inst_RegFile_32x4/mem[13][1] ;
 wire \Inst_RegFile_32x4/mem[13][2] ;
 wire \Inst_RegFile_32x4/mem[13][3] ;
 wire \Inst_RegFile_32x4/mem[14][0] ;
 wire \Inst_RegFile_32x4/mem[14][1] ;
 wire \Inst_RegFile_32x4/mem[14][2] ;
 wire \Inst_RegFile_32x4/mem[14][3] ;
 wire \Inst_RegFile_32x4/mem[15][0] ;
 wire \Inst_RegFile_32x4/mem[15][1] ;
 wire \Inst_RegFile_32x4/mem[15][2] ;
 wire \Inst_RegFile_32x4/mem[15][3] ;
 wire \Inst_RegFile_32x4/mem[16][0] ;
 wire \Inst_RegFile_32x4/mem[16][1] ;
 wire \Inst_RegFile_32x4/mem[16][2] ;
 wire \Inst_RegFile_32x4/mem[16][3] ;
 wire \Inst_RegFile_32x4/mem[17][0] ;
 wire \Inst_RegFile_32x4/mem[17][1] ;
 wire \Inst_RegFile_32x4/mem[17][2] ;
 wire \Inst_RegFile_32x4/mem[17][3] ;
 wire \Inst_RegFile_32x4/mem[18][0] ;
 wire \Inst_RegFile_32x4/mem[18][1] ;
 wire \Inst_RegFile_32x4/mem[18][2] ;
 wire \Inst_RegFile_32x4/mem[18][3] ;
 wire \Inst_RegFile_32x4/mem[19][0] ;
 wire \Inst_RegFile_32x4/mem[19][1] ;
 wire \Inst_RegFile_32x4/mem[19][2] ;
 wire \Inst_RegFile_32x4/mem[19][3] ;
 wire \Inst_RegFile_32x4/mem[1][0] ;
 wire \Inst_RegFile_32x4/mem[1][1] ;
 wire \Inst_RegFile_32x4/mem[1][2] ;
 wire \Inst_RegFile_32x4/mem[1][3] ;
 wire \Inst_RegFile_32x4/mem[20][0] ;
 wire \Inst_RegFile_32x4/mem[20][1] ;
 wire \Inst_RegFile_32x4/mem[20][2] ;
 wire \Inst_RegFile_32x4/mem[20][3] ;
 wire \Inst_RegFile_32x4/mem[21][0] ;
 wire \Inst_RegFile_32x4/mem[21][1] ;
 wire \Inst_RegFile_32x4/mem[21][2] ;
 wire \Inst_RegFile_32x4/mem[21][3] ;
 wire \Inst_RegFile_32x4/mem[22][0] ;
 wire \Inst_RegFile_32x4/mem[22][1] ;
 wire \Inst_RegFile_32x4/mem[22][2] ;
 wire \Inst_RegFile_32x4/mem[22][3] ;
 wire \Inst_RegFile_32x4/mem[23][0] ;
 wire \Inst_RegFile_32x4/mem[23][1] ;
 wire \Inst_RegFile_32x4/mem[23][2] ;
 wire \Inst_RegFile_32x4/mem[23][3] ;
 wire \Inst_RegFile_32x4/mem[24][0] ;
 wire \Inst_RegFile_32x4/mem[24][1] ;
 wire \Inst_RegFile_32x4/mem[24][2] ;
 wire \Inst_RegFile_32x4/mem[24][3] ;
 wire \Inst_RegFile_32x4/mem[25][0] ;
 wire \Inst_RegFile_32x4/mem[25][1] ;
 wire \Inst_RegFile_32x4/mem[25][2] ;
 wire \Inst_RegFile_32x4/mem[25][3] ;
 wire \Inst_RegFile_32x4/mem[26][0] ;
 wire \Inst_RegFile_32x4/mem[26][1] ;
 wire \Inst_RegFile_32x4/mem[26][2] ;
 wire \Inst_RegFile_32x4/mem[26][3] ;
 wire \Inst_RegFile_32x4/mem[27][0] ;
 wire \Inst_RegFile_32x4/mem[27][1] ;
 wire \Inst_RegFile_32x4/mem[27][2] ;
 wire \Inst_RegFile_32x4/mem[27][3] ;
 wire \Inst_RegFile_32x4/mem[28][0] ;
 wire \Inst_RegFile_32x4/mem[28][1] ;
 wire \Inst_RegFile_32x4/mem[28][2] ;
 wire \Inst_RegFile_32x4/mem[28][3] ;
 wire \Inst_RegFile_32x4/mem[29][0] ;
 wire \Inst_RegFile_32x4/mem[29][1] ;
 wire \Inst_RegFile_32x4/mem[29][2] ;
 wire \Inst_RegFile_32x4/mem[29][3] ;
 wire \Inst_RegFile_32x4/mem[2][0] ;
 wire \Inst_RegFile_32x4/mem[2][1] ;
 wire \Inst_RegFile_32x4/mem[2][2] ;
 wire \Inst_RegFile_32x4/mem[2][3] ;
 wire \Inst_RegFile_32x4/mem[30][0] ;
 wire \Inst_RegFile_32x4/mem[30][1] ;
 wire \Inst_RegFile_32x4/mem[30][2] ;
 wire \Inst_RegFile_32x4/mem[30][3] ;
 wire \Inst_RegFile_32x4/mem[31][0] ;
 wire \Inst_RegFile_32x4/mem[31][1] ;
 wire \Inst_RegFile_32x4/mem[31][2] ;
 wire \Inst_RegFile_32x4/mem[31][3] ;
 wire \Inst_RegFile_32x4/mem[3][0] ;
 wire \Inst_RegFile_32x4/mem[3][1] ;
 wire \Inst_RegFile_32x4/mem[3][2] ;
 wire \Inst_RegFile_32x4/mem[3][3] ;
 wire \Inst_RegFile_32x4/mem[4][0] ;
 wire \Inst_RegFile_32x4/mem[4][1] ;
 wire \Inst_RegFile_32x4/mem[4][2] ;
 wire \Inst_RegFile_32x4/mem[4][3] ;
 wire \Inst_RegFile_32x4/mem[5][0] ;
 wire \Inst_RegFile_32x4/mem[5][1] ;
 wire \Inst_RegFile_32x4/mem[5][2] ;
 wire \Inst_RegFile_32x4/mem[5][3] ;
 wire \Inst_RegFile_32x4/mem[6][0] ;
 wire \Inst_RegFile_32x4/mem[6][1] ;
 wire \Inst_RegFile_32x4/mem[6][2] ;
 wire \Inst_RegFile_32x4/mem[6][3] ;
 wire \Inst_RegFile_32x4/mem[7][0] ;
 wire \Inst_RegFile_32x4/mem[7][1] ;
 wire \Inst_RegFile_32x4/mem[7][2] ;
 wire \Inst_RegFile_32x4/mem[7][3] ;
 wire \Inst_RegFile_32x4/mem[8][0] ;
 wire \Inst_RegFile_32x4/mem[8][1] ;
 wire \Inst_RegFile_32x4/mem[8][2] ;
 wire \Inst_RegFile_32x4/mem[8][3] ;
 wire \Inst_RegFile_32x4/mem[9][0] ;
 wire \Inst_RegFile_32x4/mem[9][1] ;
 wire \Inst_RegFile_32x4/mem[9][2] ;
 wire \Inst_RegFile_32x4/mem[9][3] ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/my_mux2_inst/_0_ ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/cus_mux41_buf_out0 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/cus_mux41_buf_out1 ;
 wire \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/my_mux2_inst/_0_ ;
 wire \J2END_AB_BEG[0] ;
 wire \J2END_AB_BEG[1] ;
 wire \J2END_AB_BEG[2] ;
 wire \J2END_AB_BEG[3] ;
 wire \J2END_CD_BEG[0] ;
 wire \J2END_CD_BEG[1] ;
 wire \J2END_CD_BEG[2] ;
 wire \J2END_CD_BEG[3] ;
 wire \J2END_EF_BEG[0] ;
 wire \J2END_EF_BEG[1] ;
 wire \J2END_EF_BEG[2] ;
 wire \J2END_EF_BEG[3] ;
 wire \J2END_GH_BEG[0] ;
 wire \J2END_GH_BEG[1] ;
 wire \J2END_GH_BEG[2] ;
 wire \J2END_GH_BEG[3] ;
 wire \J2MID_ABa_BEG[0] ;
 wire \J2MID_ABa_BEG[1] ;
 wire \J2MID_ABa_BEG[2] ;
 wire \J2MID_ABa_BEG[3] ;
 wire \J2MID_ABb_BEG[0] ;
 wire \J2MID_ABb_BEG[1] ;
 wire \J2MID_ABb_BEG[2] ;
 wire \J2MID_ABb_BEG[3] ;
 wire \J2MID_CDa_BEG[0] ;
 wire \J2MID_CDa_BEG[1] ;
 wire \J2MID_CDa_BEG[2] ;
 wire \J2MID_CDa_BEG[3] ;
 wire \J2MID_CDb_BEG[0] ;
 wire \J2MID_CDb_BEG[1] ;
 wire \J2MID_CDb_BEG[2] ;
 wire \J2MID_CDb_BEG[3] ;
 wire \J2MID_EFa_BEG[0] ;
 wire \J2MID_EFa_BEG[1] ;
 wire \J2MID_EFa_BEG[2] ;
 wire \J2MID_EFa_BEG[3] ;
 wire \J2MID_EFb_BEG[0] ;
 wire \J2MID_EFb_BEG[1] ;
 wire \J2MID_EFb_BEG[2] ;
 wire \J2MID_EFb_BEG[3] ;
 wire \J2MID_GHa_BEG[0] ;
 wire \J2MID_GHa_BEG[1] ;
 wire \J2MID_GHa_BEG[2] ;
 wire \J2MID_GHa_BEG[3] ;
 wire \J2MID_GHb_BEG[0] ;
 wire \J2MID_GHb_BEG[1] ;
 wire \J2MID_GHb_BEG[2] ;
 wire \J2MID_GHb_BEG[3] ;
 wire \JE2BEG[0] ;
 wire \JE2BEG[1] ;
 wire \JE2BEG[2] ;
 wire \JE2BEG[3] ;
 wire \JE2BEG[4] ;
 wire \JE2BEG[5] ;
 wire \JE2BEG[6] ;
 wire \JE2BEG[7] ;
 wire \JN2BEG[0] ;
 wire \JN2BEG[1] ;
 wire \JN2BEG[2] ;
 wire \JN2BEG[3] ;
 wire \JN2BEG[4] ;
 wire \JN2BEG[5] ;
 wire \JN2BEG[6] ;
 wire \JN2BEG[7] ;
 wire \JS2BEG[0] ;
 wire \JS2BEG[1] ;
 wire \JS2BEG[2] ;
 wire \JS2BEG[3] ;
 wire \JS2BEG[4] ;
 wire \JS2BEG[5] ;
 wire \JS2BEG[6] ;
 wire \JS2BEG[7] ;
 wire \JW2BEG[0] ;
 wire \JW2BEG[1] ;
 wire \JW2BEG[2] ;
 wire \JW2BEG[3] ;
 wire \JW2BEG[4] ;
 wire \JW2BEG[5] ;
 wire \JW2BEG[6] ;
 wire \JW2BEG[7] ;
 wire \J_l_AB_BEG[0] ;
 wire \J_l_AB_BEG[1] ;
 wire \J_l_AB_BEG[2] ;
 wire \J_l_AB_BEG[3] ;
 wire \J_l_CD_BEG[0] ;
 wire \J_l_CD_BEG[1] ;
 wire \J_l_CD_BEG[2] ;
 wire \J_l_CD_BEG[3] ;
 wire \J_l_EF_BEG[0] ;
 wire \J_l_EF_BEG[1] ;
 wire \J_l_EF_BEG[2] ;
 wire \J_l_EF_BEG[3] ;
 wire \J_l_GH_BEG[0] ;
 wire \J_l_GH_BEG[1] ;
 wire \J_l_GH_BEG[2] ;
 wire \J_l_GH_BEG[3] ;
 wire \N4BEG_i[0] ;
 wire \N4BEG_i[10] ;
 wire \N4BEG_i[11] ;
 wire \N4BEG_i[1] ;
 wire \N4BEG_i[2] ;
 wire \N4BEG_i[3] ;
 wire \N4BEG_i[4] ;
 wire \N4BEG_i[5] ;
 wire \N4BEG_i[6] ;
 wire \N4BEG_i[7] ;
 wire \N4BEG_i[8] ;
 wire \N4BEG_i[9] ;
 wire \NN4BEG_i[0] ;
 wire \NN4BEG_i[10] ;
 wire \NN4BEG_i[11] ;
 wire \NN4BEG_i[1] ;
 wire \NN4BEG_i[2] ;
 wire \NN4BEG_i[3] ;
 wire \NN4BEG_i[4] ;
 wire \NN4BEG_i[5] ;
 wire \NN4BEG_i[6] ;
 wire \NN4BEG_i[7] ;
 wire \NN4BEG_i[8] ;
 wire \NN4BEG_i[9] ;
 wire \S4BEG_i[0] ;
 wire \S4BEG_i[10] ;
 wire \S4BEG_i[11] ;
 wire \S4BEG_i[1] ;
 wire \S4BEG_i[2] ;
 wire \S4BEG_i[3] ;
 wire \S4BEG_i[4] ;
 wire \S4BEG_i[5] ;
 wire \S4BEG_i[6] ;
 wire \S4BEG_i[7] ;
 wire \S4BEG_i[8] ;
 wire \S4BEG_i[9] ;
 wire \SS4BEG_i[0] ;
 wire \SS4BEG_i[10] ;
 wire \SS4BEG_i[11] ;
 wire \SS4BEG_i[1] ;
 wire \SS4BEG_i[2] ;
 wire \SS4BEG_i[3] ;
 wire \SS4BEG_i[4] ;
 wire \SS4BEG_i[5] ;
 wire \SS4BEG_i[6] ;
 wire \SS4BEG_i[7] ;
 wire \SS4BEG_i[8] ;
 wire \SS4BEG_i[9] ;
 wire \W6BEG_i[0] ;
 wire \W6BEG_i[1] ;
 wire \W6BEG_i[2] ;
 wire \W6BEG_i[3] ;
 wire \W6BEG_i[4] ;
 wire \W6BEG_i[5] ;
 wire \W6BEG_i[6] ;
 wire \W6BEG_i[7] ;
 wire \W6BEG_i[8] ;
 wire \W6BEG_i[9] ;
 wire \WW4BEG_i[0] ;
 wire \WW4BEG_i[10] ;
 wire \WW4BEG_i[11] ;
 wire \WW4BEG_i[1] ;
 wire \WW4BEG_i[2] ;
 wire \WW4BEG_i[3] ;
 wire \WW4BEG_i[4] ;
 wire \WW4BEG_i[5] ;
 wire \WW4BEG_i[6] ;
 wire \WW4BEG_i[7] ;
 wire \WW4BEG_i[8] ;
 wire \WW4BEG_i[9] ;
 wire W_ADR0;
 wire W_ADR1;
 wire W_ADR2;
 wire W_ADR3;
 wire W_ADR4;
 wire W_en;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\E6BEG_i[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\J2MID_EFb_BEG[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\J2MID_EFb_BEG[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\J2MID_EFb_BEG[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\JN2BEG[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\JS2BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\JW2BEG[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\JW2BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\JW2BEG[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\JW2BEG[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\E6BEG_i[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\JW2BEG[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\J_l_AB_BEG[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\J_l_EF_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\J_l_EF_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\N4BEG_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\N4BEG_i[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\N4BEG_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\NN4BEG_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\NN4BEG_i[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\S4BEG_i[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\E6BEG_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\SS4BEG_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\SS4BEG_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\W6BEG_i[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\E6BEG_i[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\J2END_GH_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\J2MID_ABb_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\J2END_GH_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(\J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(\J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(\JS2BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(\J_l_GH_BEG[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(\J_l_GH_BEG[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(\N4BEG_i[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\J2MID_ABa_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(\S4BEG_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(\J2MID_ABb_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(\J_l_GH_BEG[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(\J_l_GH_BEG[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\J2MID_CDa_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\J2MID_CDa_BEG[2] ));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_0/_0_  (.A(\E6BEG_i[0] ),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_1/_0_  (.A(\E6BEG_i[1] ),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_2/_0_  (.A(\E6BEG_i[2] ),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_3/_0_  (.A(\E6BEG_i[3] ),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_4/_0_  (.A(\E6BEG_i[4] ),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_5/_0_  (.A(\E6BEG_i[5] ),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_6/_0_  (.A(\E6BEG_i[6] ),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_7/_0_  (.A(\E6BEG_i[7] ),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_8/_0_  (.A(\E6BEG_i[8] ),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_9/_0_  (.A(\E6BEG_i[9] ),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_0/_0_  (.A(net25),
    .X(\E6BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_1/_0_  (.A(net26),
    .X(\E6BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_2/_0_  (.A(net27),
    .X(\E6BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_3/_0_  (.A(net28),
    .X(\E6BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_4/_0_  (.A(net29),
    .X(\E6BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_5/_0_  (.A(net30),
    .X(\E6BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_6/_0_  (.A(net31),
    .X(\E6BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_7/_0_  (.A(net32),
    .X(\E6BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_8/_0_  (.A(net22),
    .X(\E6BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_9/_0_  (.A(net23),
    .X(\E6BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_0/_0_  (.A(\EE4BEG_i[0] ),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_1/_0_  (.A(\EE4BEG_i[1] ),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_10/_0_  (.A(\EE4BEG_i[10] ),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_11/_0_  (.A(\EE4BEG_i[11] ),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_2/_0_  (.A(\EE4BEG_i[2] ),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_3/_0_  (.A(\EE4BEG_i[3] ),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_4/_0_  (.A(\EE4BEG_i[4] ),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_5/_0_  (.A(\EE4BEG_i[5] ),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_6/_0_  (.A(\EE4BEG_i[6] ),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_7/_0_  (.A(\EE4BEG_i[7] ),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_8/_0_  (.A(\EE4BEG_i[8] ),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_9/_0_  (.A(\EE4BEG_i[9] ),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_0/_0_  (.A(net43),
    .X(\EE4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_1/_0_  (.A(net44),
    .X(\EE4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_10/_0_  (.A(net38),
    .X(\EE4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_11/_0_  (.A(net39),
    .X(\EE4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_2/_0_  (.A(net45),
    .X(\EE4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_3/_0_  (.A(net46),
    .X(\EE4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_4/_0_  (.A(net47),
    .X(\EE4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_5/_0_  (.A(net48),
    .X(\EE4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_6/_0_  (.A(net34),
    .X(\EE4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_7/_0_  (.A(net35),
    .X(\EE4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_8/_0_  (.A(net36),
    .X(\EE4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_9/_0_  (.A(net37),
    .X(\EE4BEG_i[9] ));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_77 ();
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_0662_  (.A(A_ADR1),
    .X(\Inst_RegFile_32x4/_0128_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RegFile_32x4/_0663_  (.A(\Inst_RegFile_32x4/_0128_ ),
    .X(\Inst_RegFile_32x4/_0129_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0664_  (.A(A_ADR0),
    .X(\Inst_RegFile_32x4/_0130_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0665_  (.A(\Inst_RegFile_32x4/_0130_ ),
    .X(\Inst_RegFile_32x4/_0131_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0666_  (.A0(\Inst_RegFile_32x4/mem[0][0] ),
    .A1(\Inst_RegFile_32x4/mem[1][0] ),
    .S(\Inst_RegFile_32x4/_0131_ ),
    .X(\Inst_RegFile_32x4/_0132_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0667_  (.A_N(\Inst_RegFile_32x4/_0129_ ),
    .B(\Inst_RegFile_32x4/_0132_ ),
    .X(\Inst_RegFile_32x4/_0133_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0668_  (.A(A_ADR1),
    .X(\Inst_RegFile_32x4/_0134_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0669_  (.A(\Inst_RegFile_32x4/_0134_ ),
    .X(\Inst_RegFile_32x4/_0135_ ));
 sky130_fd_sc_hd__buf_2 \Inst_RegFile_32x4/_0670_  (.A(A_ADR0),
    .X(\Inst_RegFile_32x4/_0136_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0671_  (.A(\Inst_RegFile_32x4/_0136_ ),
    .X(\Inst_RegFile_32x4/_0137_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0672_  (.A0(\Inst_RegFile_32x4/mem[2][0] ),
    .A1(\Inst_RegFile_32x4/mem[3][0] ),
    .S(\Inst_RegFile_32x4/_0137_ ),
    .X(\Inst_RegFile_32x4/_0138_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0673_  (.A(A_ADR2),
    .X(\Inst_RegFile_32x4/_0139_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0674_  (.A1(\Inst_RegFile_32x4/_0135_ ),
    .A2(\Inst_RegFile_32x4/_0138_ ),
    .B1(\Inst_RegFile_32x4/_0139_ ),
    .X(\Inst_RegFile_32x4/_0140_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0675_  (.A(\Inst_RegFile_32x4/_0128_ ),
    .X(\Inst_RegFile_32x4/_0141_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0676_  (.A(\Inst_RegFile_32x4/_0130_ ),
    .X(\Inst_RegFile_32x4/_0142_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0677_  (.A0(\Inst_RegFile_32x4/mem[4][0] ),
    .A1(\Inst_RegFile_32x4/mem[5][0] ),
    .S(\Inst_RegFile_32x4/_0142_ ),
    .X(\Inst_RegFile_32x4/_0143_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0678_  (.A_N(\Inst_RegFile_32x4/_0141_ ),
    .B(\Inst_RegFile_32x4/_0143_ ),
    .X(\Inst_RegFile_32x4/_0144_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0679_  (.A(\Inst_RegFile_32x4/_0134_ ),
    .X(\Inst_RegFile_32x4/_0145_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0680_  (.A(\Inst_RegFile_32x4/_0136_ ),
    .X(\Inst_RegFile_32x4/_0146_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0681_  (.A0(\Inst_RegFile_32x4/mem[6][0] ),
    .A1(\Inst_RegFile_32x4/mem[7][0] ),
    .S(\Inst_RegFile_32x4/_0146_ ),
    .X(\Inst_RegFile_32x4/_0147_ ));
 sky130_fd_sc_hd__inv_2 \Inst_RegFile_32x4/_0682_  (.A(A_ADR2),
    .Y(\Inst_RegFile_32x4/_0148_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0683_  (.A(\Inst_RegFile_32x4/_0148_ ),
    .X(\Inst_RegFile_32x4/_0149_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0684_  (.A1(\Inst_RegFile_32x4/_0145_ ),
    .A2(\Inst_RegFile_32x4/_0147_ ),
    .B1(\Inst_RegFile_32x4/_0149_ ),
    .X(\Inst_RegFile_32x4/_0150_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0685_  (.A1(\Inst_RegFile_32x4/_0133_ ),
    .A2(\Inst_RegFile_32x4/_0140_ ),
    .B1(\Inst_RegFile_32x4/_0144_ ),
    .B2(\Inst_RegFile_32x4/_0150_ ),
    .X(\Inst_RegFile_32x4/_0151_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RegFile_32x4/_0686_  (.A(\Inst_RegFile_32x4/_0128_ ),
    .X(\Inst_RegFile_32x4/_0152_ ));
 sky130_fd_sc_hd__buf_2 \Inst_RegFile_32x4/_0687_  (.A(A_ADR0),
    .X(\Inst_RegFile_32x4/_0153_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0688_  (.A0(\Inst_RegFile_32x4/mem[8][0] ),
    .A1(\Inst_RegFile_32x4/mem[9][0] ),
    .S(\Inst_RegFile_32x4/_0153_ ),
    .X(\Inst_RegFile_32x4/_0154_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0689_  (.A_N(\Inst_RegFile_32x4/_0152_ ),
    .B(\Inst_RegFile_32x4/_0154_ ),
    .X(\Inst_RegFile_32x4/_0155_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0690_  (.A(\Inst_RegFile_32x4/_0130_ ),
    .X(\Inst_RegFile_32x4/_0156_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0691_  (.A0(\Inst_RegFile_32x4/mem[10][0] ),
    .A1(\Inst_RegFile_32x4/mem[11][0] ),
    .S(\Inst_RegFile_32x4/_0156_ ),
    .X(\Inst_RegFile_32x4/_0157_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0692_  (.A(A_ADR2),
    .X(\Inst_RegFile_32x4/_0158_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0693_  (.A1(\Inst_RegFile_32x4/_0141_ ),
    .A2(\Inst_RegFile_32x4/_0157_ ),
    .B1(\Inst_RegFile_32x4/_0158_ ),
    .X(\Inst_RegFile_32x4/_0159_ ));
 sky130_fd_sc_hd__buf_2 \Inst_RegFile_32x4/_0694_  (.A(\Inst_RegFile_32x4/_0136_ ),
    .X(\Inst_RegFile_32x4/_0160_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0695_  (.A(A_ADR1),
    .X(\Inst_RegFile_32x4/_0161_ ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_32x4/_0696_  (.A0(\Inst_RegFile_32x4/mem[12][0] ),
    .A1(\Inst_RegFile_32x4/mem[13][0] ),
    .A2(\Inst_RegFile_32x4/mem[14][0] ),
    .A3(\Inst_RegFile_32x4/mem[15][0] ),
    .S0(\Inst_RegFile_32x4/_0160_ ),
    .S1(\Inst_RegFile_32x4/_0161_ ),
    .X(\Inst_RegFile_32x4/_0162_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0697_  (.A(\Inst_RegFile_32x4/_0148_ ),
    .X(\Inst_RegFile_32x4/_0163_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0698_  (.A1(\Inst_RegFile_32x4/_0155_ ),
    .A2(\Inst_RegFile_32x4/_0159_ ),
    .B1(\Inst_RegFile_32x4/_0162_ ),
    .B2(\Inst_RegFile_32x4/_0163_ ),
    .X(\Inst_RegFile_32x4/_0164_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0699_  (.A(A_ADR0),
    .X(\Inst_RegFile_32x4/_0165_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0700_  (.A0(\Inst_RegFile_32x4/mem[16][0] ),
    .A1(\Inst_RegFile_32x4/mem[17][0] ),
    .S(\Inst_RegFile_32x4/_0165_ ),
    .X(\Inst_RegFile_32x4/_0166_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0701_  (.A_N(\Inst_RegFile_32x4/_0152_ ),
    .B(\Inst_RegFile_32x4/_0166_ ),
    .X(\Inst_RegFile_32x4/_0167_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0702_  (.A(\Inst_RegFile_32x4/_0134_ ),
    .X(\Inst_RegFile_32x4/_0168_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0703_  (.A(\Inst_RegFile_32x4/_0130_ ),
    .X(\Inst_RegFile_32x4/_0169_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0704_  (.A0(\Inst_RegFile_32x4/mem[18][0] ),
    .A1(\Inst_RegFile_32x4/mem[19][0] ),
    .S(\Inst_RegFile_32x4/_0169_ ),
    .X(\Inst_RegFile_32x4/_0170_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0705_  (.A(A_ADR2),
    .X(\Inst_RegFile_32x4/_0171_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0706_  (.A1(\Inst_RegFile_32x4/_0168_ ),
    .A2(\Inst_RegFile_32x4/_0170_ ),
    .B1(\Inst_RegFile_32x4/_0171_ ),
    .X(\Inst_RegFile_32x4/_0172_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RegFile_32x4/_0707_  (.A(\Inst_RegFile_32x4/_0128_ ),
    .X(\Inst_RegFile_32x4/_0173_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0708_  (.A(\Inst_RegFile_32x4/_0130_ ),
    .X(\Inst_RegFile_32x4/_0174_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0709_  (.A0(\Inst_RegFile_32x4/mem[20][0] ),
    .A1(\Inst_RegFile_32x4/mem[21][0] ),
    .S(\Inst_RegFile_32x4/_0174_ ),
    .X(\Inst_RegFile_32x4/_0175_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0710_  (.A_N(\Inst_RegFile_32x4/_0173_ ),
    .B(\Inst_RegFile_32x4/_0175_ ),
    .X(\Inst_RegFile_32x4/_0176_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0711_  (.A(\Inst_RegFile_32x4/_0136_ ),
    .X(\Inst_RegFile_32x4/_0177_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0712_  (.A0(\Inst_RegFile_32x4/mem[22][0] ),
    .A1(\Inst_RegFile_32x4/mem[23][0] ),
    .S(\Inst_RegFile_32x4/_0177_ ),
    .X(\Inst_RegFile_32x4/_0178_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0713_  (.A(\Inst_RegFile_32x4/_0148_ ),
    .X(\Inst_RegFile_32x4/_0179_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0714_  (.A1(\Inst_RegFile_32x4/_0145_ ),
    .A2(\Inst_RegFile_32x4/_0178_ ),
    .B1(\Inst_RegFile_32x4/_0179_ ),
    .X(\Inst_RegFile_32x4/_0180_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0715_  (.A1(\Inst_RegFile_32x4/_0167_ ),
    .A2(\Inst_RegFile_32x4/_0172_ ),
    .B1(\Inst_RegFile_32x4/_0176_ ),
    .B2(\Inst_RegFile_32x4/_0180_ ),
    .X(\Inst_RegFile_32x4/_0181_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_0716_  (.A(\Inst_RegFile_32x4/_0128_ ),
    .X(\Inst_RegFile_32x4/_0182_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0717_  (.A0(\Inst_RegFile_32x4/mem[24][0] ),
    .A1(\Inst_RegFile_32x4/mem[25][0] ),
    .S(\Inst_RegFile_32x4/_0131_ ),
    .X(\Inst_RegFile_32x4/_0183_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0718_  (.A_N(\Inst_RegFile_32x4/_0182_ ),
    .B(\Inst_RegFile_32x4/_0183_ ),
    .X(\Inst_RegFile_32x4/_0184_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0719_  (.A(\Inst_RegFile_32x4/_0134_ ),
    .X(\Inst_RegFile_32x4/_0185_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0720_  (.A0(\Inst_RegFile_32x4/mem[26][0] ),
    .A1(\Inst_RegFile_32x4/mem[27][0] ),
    .S(\Inst_RegFile_32x4/_0169_ ),
    .X(\Inst_RegFile_32x4/_0186_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0721_  (.A1(\Inst_RegFile_32x4/_0185_ ),
    .A2(\Inst_RegFile_32x4/_0186_ ),
    .B1(\Inst_RegFile_32x4/_0139_ ),
    .X(\Inst_RegFile_32x4/_0187_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_0722_  (.A(A_ADR1),
    .X(\Inst_RegFile_32x4/_0188_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0723_  (.A0(\Inst_RegFile_32x4/mem[28][0] ),
    .A1(\Inst_RegFile_32x4/mem[29][0] ),
    .A2(\Inst_RegFile_32x4/mem[30][0] ),
    .A3(\Inst_RegFile_32x4/mem[31][0] ),
    .S0(\Inst_RegFile_32x4/_0160_ ),
    .S1(\Inst_RegFile_32x4/_0188_ ),
    .X(\Inst_RegFile_32x4/_0189_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0724_  (.A1(\Inst_RegFile_32x4/_0184_ ),
    .A2(\Inst_RegFile_32x4/_0187_ ),
    .B1(\Inst_RegFile_32x4/_0189_ ),
    .B2(\Inst_RegFile_32x4/_0163_ ),
    .X(\Inst_RegFile_32x4/_0190_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0725_  (.A0(\Inst_RegFile_32x4/_0151_ ),
    .A1(\Inst_RegFile_32x4/_0164_ ),
    .A2(\Inst_RegFile_32x4/_0181_ ),
    .A3(\Inst_RegFile_32x4/_0190_ ),
    .S0(A_ADR3),
    .S1(A_ADR4),
    .X(\Inst_RegFile_32x4/_0191_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_0726_  (.A(\Inst_RegFile_32x4/_0191_ ),
    .X(\Inst_RegFile_32x4/AD_comb[0] ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0727_  (.A0(\Inst_RegFile_32x4/mem[0][1] ),
    .A1(\Inst_RegFile_32x4/mem[1][1] ),
    .S(\Inst_RegFile_32x4/_0131_ ),
    .X(\Inst_RegFile_32x4/_0192_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0728_  (.A_N(\Inst_RegFile_32x4/_0129_ ),
    .B(\Inst_RegFile_32x4/_0192_ ),
    .X(\Inst_RegFile_32x4/_0193_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0729_  (.A0(\Inst_RegFile_32x4/mem[2][1] ),
    .A1(\Inst_RegFile_32x4/mem[3][1] ),
    .S(\Inst_RegFile_32x4/_0137_ ),
    .X(\Inst_RegFile_32x4/_0194_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0730_  (.A1(\Inst_RegFile_32x4/_0135_ ),
    .A2(\Inst_RegFile_32x4/_0194_ ),
    .B1(\Inst_RegFile_32x4/_0139_ ),
    .X(\Inst_RegFile_32x4/_0195_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0731_  (.A0(\Inst_RegFile_32x4/mem[4][1] ),
    .A1(\Inst_RegFile_32x4/mem[5][1] ),
    .S(\Inst_RegFile_32x4/_0142_ ),
    .X(\Inst_RegFile_32x4/_0196_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0732_  (.A_N(\Inst_RegFile_32x4/_0173_ ),
    .B(\Inst_RegFile_32x4/_0196_ ),
    .X(\Inst_RegFile_32x4/_0197_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0733_  (.A0(\Inst_RegFile_32x4/mem[6][1] ),
    .A1(\Inst_RegFile_32x4/mem[7][1] ),
    .S(\Inst_RegFile_32x4/_0146_ ),
    .X(\Inst_RegFile_32x4/_0198_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0734_  (.A1(\Inst_RegFile_32x4/_0145_ ),
    .A2(\Inst_RegFile_32x4/_0198_ ),
    .B1(\Inst_RegFile_32x4/_0149_ ),
    .X(\Inst_RegFile_32x4/_0199_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0735_  (.A1(\Inst_RegFile_32x4/_0193_ ),
    .A2(\Inst_RegFile_32x4/_0195_ ),
    .B1(\Inst_RegFile_32x4/_0197_ ),
    .B2(\Inst_RegFile_32x4/_0199_ ),
    .X(\Inst_RegFile_32x4/_0200_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0736_  (.A0(\Inst_RegFile_32x4/mem[8][1] ),
    .A1(\Inst_RegFile_32x4/mem[9][1] ),
    .S(\Inst_RegFile_32x4/_0153_ ),
    .X(\Inst_RegFile_32x4/_0201_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0737_  (.A_N(\Inst_RegFile_32x4/_0188_ ),
    .B(\Inst_RegFile_32x4/_0201_ ),
    .X(\Inst_RegFile_32x4/_0202_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0738_  (.A0(\Inst_RegFile_32x4/mem[10][1] ),
    .A1(\Inst_RegFile_32x4/mem[11][1] ),
    .S(\Inst_RegFile_32x4/_0156_ ),
    .X(\Inst_RegFile_32x4/_0203_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0739_  (.A1(\Inst_RegFile_32x4/_0141_ ),
    .A2(\Inst_RegFile_32x4/_0203_ ),
    .B1(\Inst_RegFile_32x4/_0158_ ),
    .X(\Inst_RegFile_32x4/_0204_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0740_  (.A0(\Inst_RegFile_32x4/mem[12][1] ),
    .A1(\Inst_RegFile_32x4/mem[13][1] ),
    .A2(\Inst_RegFile_32x4/mem[14][1] ),
    .A3(\Inst_RegFile_32x4/mem[15][1] ),
    .S0(\Inst_RegFile_32x4/_0146_ ),
    .S1(\Inst_RegFile_32x4/_0161_ ),
    .X(\Inst_RegFile_32x4/_0205_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0741_  (.A1(\Inst_RegFile_32x4/_0202_ ),
    .A2(\Inst_RegFile_32x4/_0204_ ),
    .B1(\Inst_RegFile_32x4/_0205_ ),
    .B2(\Inst_RegFile_32x4/_0149_ ),
    .X(\Inst_RegFile_32x4/_0206_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0742_  (.A0(\Inst_RegFile_32x4/mem[16][1] ),
    .A1(\Inst_RegFile_32x4/mem[17][1] ),
    .S(\Inst_RegFile_32x4/_0165_ ),
    .X(\Inst_RegFile_32x4/_0207_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0743_  (.A_N(\Inst_RegFile_32x4/_0152_ ),
    .B(\Inst_RegFile_32x4/_0207_ ),
    .X(\Inst_RegFile_32x4/_0208_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0744_  (.A0(\Inst_RegFile_32x4/mem[18][1] ),
    .A1(\Inst_RegFile_32x4/mem[19][1] ),
    .S(\Inst_RegFile_32x4/_0156_ ),
    .X(\Inst_RegFile_32x4/_0209_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0745_  (.A1(\Inst_RegFile_32x4/_0168_ ),
    .A2(\Inst_RegFile_32x4/_0209_ ),
    .B1(\Inst_RegFile_32x4/_0171_ ),
    .X(\Inst_RegFile_32x4/_0210_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0746_  (.A0(\Inst_RegFile_32x4/mem[20][1] ),
    .A1(\Inst_RegFile_32x4/mem[21][1] ),
    .S(\Inst_RegFile_32x4/_0174_ ),
    .X(\Inst_RegFile_32x4/_0211_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0747_  (.A_N(\Inst_RegFile_32x4/_0173_ ),
    .B(\Inst_RegFile_32x4/_0211_ ),
    .X(\Inst_RegFile_32x4/_0212_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0748_  (.A0(\Inst_RegFile_32x4/mem[22][1] ),
    .A1(\Inst_RegFile_32x4/mem[23][1] ),
    .S(\Inst_RegFile_32x4/_0177_ ),
    .X(\Inst_RegFile_32x4/_0213_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0749_  (.A1(\Inst_RegFile_32x4/_0135_ ),
    .A2(\Inst_RegFile_32x4/_0213_ ),
    .B1(\Inst_RegFile_32x4/_0179_ ),
    .X(\Inst_RegFile_32x4/_0214_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0750_  (.A1(\Inst_RegFile_32x4/_0208_ ),
    .A2(\Inst_RegFile_32x4/_0210_ ),
    .B1(\Inst_RegFile_32x4/_0212_ ),
    .B2(\Inst_RegFile_32x4/_0214_ ),
    .X(\Inst_RegFile_32x4/_0215_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0751_  (.A0(\Inst_RegFile_32x4/mem[24][1] ),
    .A1(\Inst_RegFile_32x4/mem[25][1] ),
    .S(\Inst_RegFile_32x4/_0165_ ),
    .X(\Inst_RegFile_32x4/_0216_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0752_  (.A_N(\Inst_RegFile_32x4/_0182_ ),
    .B(\Inst_RegFile_32x4/_0216_ ),
    .X(\Inst_RegFile_32x4/_0217_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0753_  (.A0(\Inst_RegFile_32x4/mem[26][1] ),
    .A1(\Inst_RegFile_32x4/mem[27][1] ),
    .S(\Inst_RegFile_32x4/_0169_ ),
    .X(\Inst_RegFile_32x4/_0218_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0754_  (.A1(\Inst_RegFile_32x4/_0185_ ),
    .A2(\Inst_RegFile_32x4/_0218_ ),
    .B1(\Inst_RegFile_32x4/_0171_ ),
    .X(\Inst_RegFile_32x4/_0219_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0755_  (.A0(\Inst_RegFile_32x4/mem[28][1] ),
    .A1(\Inst_RegFile_32x4/mem[29][1] ),
    .A2(\Inst_RegFile_32x4/mem[30][1] ),
    .A3(\Inst_RegFile_32x4/mem[31][1] ),
    .S0(\Inst_RegFile_32x4/_0160_ ),
    .S1(\Inst_RegFile_32x4/_0188_ ),
    .X(\Inst_RegFile_32x4/_0220_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0756_  (.A1(\Inst_RegFile_32x4/_0217_ ),
    .A2(\Inst_RegFile_32x4/_0219_ ),
    .B1(\Inst_RegFile_32x4/_0220_ ),
    .B2(\Inst_RegFile_32x4/_0163_ ),
    .X(\Inst_RegFile_32x4/_0221_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0757_  (.A0(\Inst_RegFile_32x4/_0200_ ),
    .A1(\Inst_RegFile_32x4/_0206_ ),
    .A2(\Inst_RegFile_32x4/_0215_ ),
    .A3(\Inst_RegFile_32x4/_0221_ ),
    .S0(A_ADR3),
    .S1(A_ADR4),
    .X(\Inst_RegFile_32x4/_0222_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_0758_  (.A(\Inst_RegFile_32x4/_0222_ ),
    .X(\Inst_RegFile_32x4/AD_comb[1] ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0759_  (.A0(\Inst_RegFile_32x4/mem[0][2] ),
    .A1(\Inst_RegFile_32x4/mem[1][2] ),
    .S(\Inst_RegFile_32x4/_0131_ ),
    .X(\Inst_RegFile_32x4/_0223_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0760_  (.A_N(\Inst_RegFile_32x4/_0129_ ),
    .B(\Inst_RegFile_32x4/_0223_ ),
    .X(\Inst_RegFile_32x4/_0224_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0761_  (.A0(\Inst_RegFile_32x4/mem[2][2] ),
    .A1(\Inst_RegFile_32x4/mem[3][2] ),
    .S(\Inst_RegFile_32x4/_0137_ ),
    .X(\Inst_RegFile_32x4/_0225_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0762_  (.A1(\Inst_RegFile_32x4/_0185_ ),
    .A2(\Inst_RegFile_32x4/_0225_ ),
    .B1(\Inst_RegFile_32x4/_0139_ ),
    .X(\Inst_RegFile_32x4/_0226_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0763_  (.A0(\Inst_RegFile_32x4/mem[4][2] ),
    .A1(\Inst_RegFile_32x4/mem[5][2] ),
    .S(\Inst_RegFile_32x4/_0142_ ),
    .X(\Inst_RegFile_32x4/_0227_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0764_  (.A_N(\Inst_RegFile_32x4/_0173_ ),
    .B(\Inst_RegFile_32x4/_0227_ ),
    .X(\Inst_RegFile_32x4/_0228_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0765_  (.A0(\Inst_RegFile_32x4/mem[6][2] ),
    .A1(\Inst_RegFile_32x4/mem[7][2] ),
    .S(\Inst_RegFile_32x4/_0177_ ),
    .X(\Inst_RegFile_32x4/_0229_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0766_  (.A1(\Inst_RegFile_32x4/_0145_ ),
    .A2(\Inst_RegFile_32x4/_0229_ ),
    .B1(\Inst_RegFile_32x4/_0179_ ),
    .X(\Inst_RegFile_32x4/_0230_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0767_  (.A1(\Inst_RegFile_32x4/_0224_ ),
    .A2(\Inst_RegFile_32x4/_0226_ ),
    .B1(\Inst_RegFile_32x4/_0228_ ),
    .B2(\Inst_RegFile_32x4/_0230_ ),
    .X(\Inst_RegFile_32x4/_0231_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0768_  (.A0(\Inst_RegFile_32x4/mem[8][2] ),
    .A1(\Inst_RegFile_32x4/mem[9][2] ),
    .S(\Inst_RegFile_32x4/_0153_ ),
    .X(\Inst_RegFile_32x4/_0232_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0769_  (.A_N(\Inst_RegFile_32x4/_0188_ ),
    .B(\Inst_RegFile_32x4/_0232_ ),
    .X(\Inst_RegFile_32x4/_0233_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0770_  (.A0(\Inst_RegFile_32x4/mem[10][2] ),
    .A1(\Inst_RegFile_32x4/mem[11][2] ),
    .S(\Inst_RegFile_32x4/_0142_ ),
    .X(\Inst_RegFile_32x4/_0234_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0771_  (.A1(\Inst_RegFile_32x4/_0141_ ),
    .A2(\Inst_RegFile_32x4/_0234_ ),
    .B1(\Inst_RegFile_32x4/_0158_ ),
    .X(\Inst_RegFile_32x4/_0235_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0772_  (.A0(\Inst_RegFile_32x4/mem[12][2] ),
    .A1(\Inst_RegFile_32x4/mem[13][2] ),
    .A2(\Inst_RegFile_32x4/mem[14][2] ),
    .A3(\Inst_RegFile_32x4/mem[15][2] ),
    .S0(\Inst_RegFile_32x4/_0146_ ),
    .S1(\Inst_RegFile_32x4/_0161_ ),
    .X(\Inst_RegFile_32x4/_0236_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0773_  (.A1(\Inst_RegFile_32x4/_0233_ ),
    .A2(\Inst_RegFile_32x4/_0235_ ),
    .B1(\Inst_RegFile_32x4/_0236_ ),
    .B2(\Inst_RegFile_32x4/_0149_ ),
    .X(\Inst_RegFile_32x4/_0237_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0774_  (.A0(\Inst_RegFile_32x4/mem[16][2] ),
    .A1(\Inst_RegFile_32x4/mem[17][2] ),
    .S(\Inst_RegFile_32x4/_0153_ ),
    .X(\Inst_RegFile_32x4/_0238_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0775_  (.A_N(\Inst_RegFile_32x4/_0152_ ),
    .B(\Inst_RegFile_32x4/_0238_ ),
    .X(\Inst_RegFile_32x4/_0239_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0776_  (.A0(\Inst_RegFile_32x4/mem[18][2] ),
    .A1(\Inst_RegFile_32x4/mem[19][2] ),
    .S(\Inst_RegFile_32x4/_0156_ ),
    .X(\Inst_RegFile_32x4/_0240_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0777_  (.A1(\Inst_RegFile_32x4/_0168_ ),
    .A2(\Inst_RegFile_32x4/_0240_ ),
    .B1(\Inst_RegFile_32x4/_0158_ ),
    .X(\Inst_RegFile_32x4/_0241_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0778_  (.A0(\Inst_RegFile_32x4/mem[20][2] ),
    .A1(\Inst_RegFile_32x4/mem[21][2] ),
    .S(\Inst_RegFile_32x4/_0174_ ),
    .X(\Inst_RegFile_32x4/_0242_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0779_  (.A_N(\Inst_RegFile_32x4/_0129_ ),
    .B(\Inst_RegFile_32x4/_0242_ ),
    .X(\Inst_RegFile_32x4/_0243_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0780_  (.A0(\Inst_RegFile_32x4/mem[22][2] ),
    .A1(\Inst_RegFile_32x4/mem[23][2] ),
    .S(\Inst_RegFile_32x4/_0177_ ),
    .X(\Inst_RegFile_32x4/_0244_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0781_  (.A1(\Inst_RegFile_32x4/_0135_ ),
    .A2(\Inst_RegFile_32x4/_0244_ ),
    .B1(\Inst_RegFile_32x4/_0179_ ),
    .X(\Inst_RegFile_32x4/_0245_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0782_  (.A1(\Inst_RegFile_32x4/_0239_ ),
    .A2(\Inst_RegFile_32x4/_0241_ ),
    .B1(\Inst_RegFile_32x4/_0243_ ),
    .B2(\Inst_RegFile_32x4/_0245_ ),
    .X(\Inst_RegFile_32x4/_0246_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0783_  (.A0(\Inst_RegFile_32x4/mem[24][2] ),
    .A1(\Inst_RegFile_32x4/mem[25][2] ),
    .S(\Inst_RegFile_32x4/_0165_ ),
    .X(\Inst_RegFile_32x4/_0247_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0784_  (.A_N(\Inst_RegFile_32x4/_0182_ ),
    .B(\Inst_RegFile_32x4/_0247_ ),
    .X(\Inst_RegFile_32x4/_0248_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0785_  (.A0(\Inst_RegFile_32x4/mem[26][2] ),
    .A1(\Inst_RegFile_32x4/mem[27][2] ),
    .S(\Inst_RegFile_32x4/_0169_ ),
    .X(\Inst_RegFile_32x4/_0249_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0786_  (.A1(\Inst_RegFile_32x4/_0185_ ),
    .A2(\Inst_RegFile_32x4/_0249_ ),
    .B1(\Inst_RegFile_32x4/_0171_ ),
    .X(\Inst_RegFile_32x4/_0250_ ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_32x4/_0787_  (.A0(\Inst_RegFile_32x4/mem[28][2] ),
    .A1(\Inst_RegFile_32x4/mem[29][2] ),
    .A2(\Inst_RegFile_32x4/mem[30][2] ),
    .A3(\Inst_RegFile_32x4/mem[31][2] ),
    .S0(\Inst_RegFile_32x4/_0160_ ),
    .S1(\Inst_RegFile_32x4/_0161_ ),
    .X(\Inst_RegFile_32x4/_0251_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0788_  (.A1(\Inst_RegFile_32x4/_0248_ ),
    .A2(\Inst_RegFile_32x4/_0250_ ),
    .B1(\Inst_RegFile_32x4/_0251_ ),
    .B2(\Inst_RegFile_32x4/_0163_ ),
    .X(\Inst_RegFile_32x4/_0252_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0789_  (.A0(\Inst_RegFile_32x4/_0231_ ),
    .A1(\Inst_RegFile_32x4/_0237_ ),
    .A2(\Inst_RegFile_32x4/_0246_ ),
    .A3(\Inst_RegFile_32x4/_0252_ ),
    .S0(A_ADR3),
    .S1(A_ADR4),
    .X(\Inst_RegFile_32x4/_0253_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_0790_  (.A(\Inst_RegFile_32x4/_0253_ ),
    .X(\Inst_RegFile_32x4/AD_comb[2] ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0791_  (.A0(\Inst_RegFile_32x4/mem[0][3] ),
    .A1(\Inst_RegFile_32x4/mem[1][3] ),
    .S(\Inst_RegFile_32x4/_0131_ ),
    .X(\Inst_RegFile_32x4/_0254_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0792_  (.A_N(\Inst_RegFile_32x4/_0182_ ),
    .B(\Inst_RegFile_32x4/_0254_ ),
    .X(\Inst_RegFile_32x4/_0255_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0793_  (.A0(\Inst_RegFile_32x4/mem[2][3] ),
    .A1(\Inst_RegFile_32x4/mem[3][3] ),
    .S(\Inst_RegFile_32x4/_0137_ ),
    .X(\Inst_RegFile_32x4/_0256_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0794_  (.A1(\Inst_RegFile_32x4/_0185_ ),
    .A2(\Inst_RegFile_32x4/_0256_ ),
    .B1(\Inst_RegFile_32x4/_0139_ ),
    .X(\Inst_RegFile_32x4/_0257_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0795_  (.A0(\Inst_RegFile_32x4/mem[4][3] ),
    .A1(\Inst_RegFile_32x4/mem[5][3] ),
    .S(\Inst_RegFile_32x4/_0174_ ),
    .X(\Inst_RegFile_32x4/_0258_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0796_  (.A_N(\Inst_RegFile_32x4/_0173_ ),
    .B(\Inst_RegFile_32x4/_0258_ ),
    .X(\Inst_RegFile_32x4/_0259_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0797_  (.A0(\Inst_RegFile_32x4/mem[6][3] ),
    .A1(\Inst_RegFile_32x4/mem[7][3] ),
    .S(\Inst_RegFile_32x4/_0177_ ),
    .X(\Inst_RegFile_32x4/_0260_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0798_  (.A1(\Inst_RegFile_32x4/_0145_ ),
    .A2(\Inst_RegFile_32x4/_0260_ ),
    .B1(\Inst_RegFile_32x4/_0179_ ),
    .X(\Inst_RegFile_32x4/_0261_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0799_  (.A1(\Inst_RegFile_32x4/_0255_ ),
    .A2(\Inst_RegFile_32x4/_0257_ ),
    .B1(\Inst_RegFile_32x4/_0259_ ),
    .B2(\Inst_RegFile_32x4/_0261_ ),
    .X(\Inst_RegFile_32x4/_0262_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0800_  (.A0(\Inst_RegFile_32x4/mem[8][3] ),
    .A1(\Inst_RegFile_32x4/mem[9][3] ),
    .S(\Inst_RegFile_32x4/_0136_ ),
    .X(\Inst_RegFile_32x4/_0263_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0801_  (.A_N(\Inst_RegFile_32x4/_0188_ ),
    .B(\Inst_RegFile_32x4/_0263_ ),
    .X(\Inst_RegFile_32x4/_0264_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0802_  (.A0(\Inst_RegFile_32x4/mem[10][3] ),
    .A1(\Inst_RegFile_32x4/mem[11][3] ),
    .S(\Inst_RegFile_32x4/_0142_ ),
    .X(\Inst_RegFile_32x4/_0265_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0803_  (.A1(\Inst_RegFile_32x4/_0141_ ),
    .A2(\Inst_RegFile_32x4/_0265_ ),
    .B1(A_ADR2),
    .X(\Inst_RegFile_32x4/_0266_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0804_  (.A0(\Inst_RegFile_32x4/mem[12][3] ),
    .A1(\Inst_RegFile_32x4/mem[13][3] ),
    .A2(\Inst_RegFile_32x4/mem[14][3] ),
    .A3(\Inst_RegFile_32x4/mem[15][3] ),
    .S0(\Inst_RegFile_32x4/_0146_ ),
    .S1(\Inst_RegFile_32x4/_0134_ ),
    .X(\Inst_RegFile_32x4/_0267_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0805_  (.A1(\Inst_RegFile_32x4/_0264_ ),
    .A2(\Inst_RegFile_32x4/_0266_ ),
    .B1(\Inst_RegFile_32x4/_0267_ ),
    .B2(\Inst_RegFile_32x4/_0149_ ),
    .X(\Inst_RegFile_32x4/_0268_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0806_  (.A0(\Inst_RegFile_32x4/mem[16][3] ),
    .A1(\Inst_RegFile_32x4/mem[17][3] ),
    .S(\Inst_RegFile_32x4/_0153_ ),
    .X(\Inst_RegFile_32x4/_0269_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0807_  (.A_N(\Inst_RegFile_32x4/_0152_ ),
    .B(\Inst_RegFile_32x4/_0269_ ),
    .X(\Inst_RegFile_32x4/_0270_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0808_  (.A0(\Inst_RegFile_32x4/mem[18][3] ),
    .A1(\Inst_RegFile_32x4/mem[19][3] ),
    .S(\Inst_RegFile_32x4/_0156_ ),
    .X(\Inst_RegFile_32x4/_0271_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0809_  (.A1(\Inst_RegFile_32x4/_0168_ ),
    .A2(\Inst_RegFile_32x4/_0271_ ),
    .B1(\Inst_RegFile_32x4/_0158_ ),
    .X(\Inst_RegFile_32x4/_0272_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0810_  (.A0(\Inst_RegFile_32x4/mem[20][3] ),
    .A1(\Inst_RegFile_32x4/mem[21][3] ),
    .S(\Inst_RegFile_32x4/_0174_ ),
    .X(\Inst_RegFile_32x4/_0273_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0811_  (.A_N(\Inst_RegFile_32x4/_0129_ ),
    .B(\Inst_RegFile_32x4/_0273_ ),
    .X(\Inst_RegFile_32x4/_0274_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0812_  (.A0(\Inst_RegFile_32x4/mem[22][3] ),
    .A1(\Inst_RegFile_32x4/mem[23][3] ),
    .S(\Inst_RegFile_32x4/_0137_ ),
    .X(\Inst_RegFile_32x4/_0275_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0813_  (.A1(\Inst_RegFile_32x4/_0135_ ),
    .A2(\Inst_RegFile_32x4/_0275_ ),
    .B1(\Inst_RegFile_32x4/_0148_ ),
    .X(\Inst_RegFile_32x4/_0276_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0814_  (.A1(\Inst_RegFile_32x4/_0270_ ),
    .A2(\Inst_RegFile_32x4/_0272_ ),
    .B1(\Inst_RegFile_32x4/_0274_ ),
    .B2(\Inst_RegFile_32x4/_0276_ ),
    .X(\Inst_RegFile_32x4/_0277_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0815_  (.A0(\Inst_RegFile_32x4/mem[24][3] ),
    .A1(\Inst_RegFile_32x4/mem[25][3] ),
    .S(\Inst_RegFile_32x4/_0165_ ),
    .X(\Inst_RegFile_32x4/_0278_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0816_  (.A_N(\Inst_RegFile_32x4/_0182_ ),
    .B(\Inst_RegFile_32x4/_0278_ ),
    .X(\Inst_RegFile_32x4/_0279_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0817_  (.A0(\Inst_RegFile_32x4/mem[26][3] ),
    .A1(\Inst_RegFile_32x4/mem[27][3] ),
    .S(\Inst_RegFile_32x4/_0169_ ),
    .X(\Inst_RegFile_32x4/_0280_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0818_  (.A1(\Inst_RegFile_32x4/_0168_ ),
    .A2(\Inst_RegFile_32x4/_0280_ ),
    .B1(\Inst_RegFile_32x4/_0171_ ),
    .X(\Inst_RegFile_32x4/_0281_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0819_  (.A0(\Inst_RegFile_32x4/mem[28][3] ),
    .A1(\Inst_RegFile_32x4/mem[29][3] ),
    .A2(\Inst_RegFile_32x4/mem[30][3] ),
    .A3(\Inst_RegFile_32x4/mem[31][3] ),
    .S0(\Inst_RegFile_32x4/_0160_ ),
    .S1(\Inst_RegFile_32x4/_0161_ ),
    .X(\Inst_RegFile_32x4/_0282_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0820_  (.A1(\Inst_RegFile_32x4/_0279_ ),
    .A2(\Inst_RegFile_32x4/_0281_ ),
    .B1(\Inst_RegFile_32x4/_0282_ ),
    .B2(\Inst_RegFile_32x4/_0163_ ),
    .X(\Inst_RegFile_32x4/_0283_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0821_  (.A0(\Inst_RegFile_32x4/_0262_ ),
    .A1(\Inst_RegFile_32x4/_0268_ ),
    .A2(\Inst_RegFile_32x4/_0277_ ),
    .A3(\Inst_RegFile_32x4/_0283_ ),
    .S0(A_ADR3),
    .S1(A_ADR4),
    .X(\Inst_RegFile_32x4/_0284_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_0822_  (.A(\Inst_RegFile_32x4/_0284_ ),
    .X(\Inst_RegFile_32x4/AD_comb[3] ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0823_  (.A0(\Inst_RegFile_32x4/AD_comb[0] ),
    .A1(\Inst_RegFile_32x4/AD_reg[0] ),
    .S(\ConfigBits[0] ),
    .X(\Inst_RegFile_32x4/_0285_ ));
 sky130_fd_sc_hd__buf_12 \Inst_RegFile_32x4/_0824_  (.A(\Inst_RegFile_32x4/_0285_ ),
    .X(AD0));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0825_  (.A0(\Inst_RegFile_32x4/AD_comb[1] ),
    .A1(\Inst_RegFile_32x4/AD_reg[1] ),
    .S(\ConfigBits[0] ),
    .X(\Inst_RegFile_32x4/_0286_ ));
 sky130_fd_sc_hd__clkbuf_16 \Inst_RegFile_32x4/_0826_  (.A(\Inst_RegFile_32x4/_0286_ ),
    .X(AD1));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0827_  (.A0(\Inst_RegFile_32x4/AD_comb[2] ),
    .A1(\Inst_RegFile_32x4/AD_reg[2] ),
    .S(\ConfigBits[0] ),
    .X(\Inst_RegFile_32x4/_0287_ ));
 sky130_fd_sc_hd__buf_12 \Inst_RegFile_32x4/_0828_  (.A(\Inst_RegFile_32x4/_0287_ ),
    .X(AD2));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0829_  (.A0(\Inst_RegFile_32x4/AD_comb[3] ),
    .A1(\Inst_RegFile_32x4/AD_reg[3] ),
    .S(\ConfigBits[0] ),
    .X(\Inst_RegFile_32x4/_0288_ ));
 sky130_fd_sc_hd__buf_12 \Inst_RegFile_32x4/_0830_  (.A(\Inst_RegFile_32x4/_0288_ ),
    .X(AD3));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_0831_  (.A(B_ADR1),
    .X(\Inst_RegFile_32x4/_0289_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_0832_  (.A(\Inst_RegFile_32x4/_0289_ ),
    .X(\Inst_RegFile_32x4/_0290_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RegFile_32x4/_0833_  (.A(B_ADR0),
    .X(\Inst_RegFile_32x4/_0291_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0834_  (.A(\Inst_RegFile_32x4/_0291_ ),
    .X(\Inst_RegFile_32x4/_0292_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0835_  (.A0(\Inst_RegFile_32x4/mem[0][0] ),
    .A1(\Inst_RegFile_32x4/mem[1][0] ),
    .S(\Inst_RegFile_32x4/_0292_ ),
    .X(\Inst_RegFile_32x4/_0293_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0836_  (.A_N(\Inst_RegFile_32x4/_0290_ ),
    .B(\Inst_RegFile_32x4/_0293_ ),
    .X(\Inst_RegFile_32x4/_0294_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0837_  (.A(B_ADR1),
    .X(\Inst_RegFile_32x4/_0295_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0838_  (.A(\Inst_RegFile_32x4/_0295_ ),
    .X(\Inst_RegFile_32x4/_0296_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0839_  (.A(B_ADR0),
    .X(\Inst_RegFile_32x4/_0297_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0840_  (.A(\Inst_RegFile_32x4/_0297_ ),
    .X(\Inst_RegFile_32x4/_0298_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0841_  (.A0(\Inst_RegFile_32x4/mem[2][0] ),
    .A1(\Inst_RegFile_32x4/mem[3][0] ),
    .S(\Inst_RegFile_32x4/_0298_ ),
    .X(\Inst_RegFile_32x4/_0299_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0842_  (.A(B_ADR2),
    .X(\Inst_RegFile_32x4/_0300_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0843_  (.A1(\Inst_RegFile_32x4/_0296_ ),
    .A2(\Inst_RegFile_32x4/_0299_ ),
    .B1(\Inst_RegFile_32x4/_0300_ ),
    .X(\Inst_RegFile_32x4/_0301_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RegFile_32x4/_0844_  (.A(\Inst_RegFile_32x4/_0289_ ),
    .X(\Inst_RegFile_32x4/_0302_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0845_  (.A(\Inst_RegFile_32x4/_0291_ ),
    .X(\Inst_RegFile_32x4/_0303_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0846_  (.A0(\Inst_RegFile_32x4/mem[4][0] ),
    .A1(\Inst_RegFile_32x4/mem[5][0] ),
    .S(\Inst_RegFile_32x4/_0303_ ),
    .X(\Inst_RegFile_32x4/_0304_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0847_  (.A_N(\Inst_RegFile_32x4/_0302_ ),
    .B(\Inst_RegFile_32x4/_0304_ ),
    .X(\Inst_RegFile_32x4/_0305_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0848_  (.A(\Inst_RegFile_32x4/_0295_ ),
    .X(\Inst_RegFile_32x4/_0306_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0849_  (.A(\Inst_RegFile_32x4/_0297_ ),
    .X(\Inst_RegFile_32x4/_0307_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0850_  (.A0(\Inst_RegFile_32x4/mem[6][0] ),
    .A1(\Inst_RegFile_32x4/mem[7][0] ),
    .S(\Inst_RegFile_32x4/_0307_ ),
    .X(\Inst_RegFile_32x4/_0308_ ));
 sky130_fd_sc_hd__inv_2 \Inst_RegFile_32x4/_0851_  (.A(B_ADR2),
    .Y(\Inst_RegFile_32x4/_0309_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RegFile_32x4/_0852_  (.A(\Inst_RegFile_32x4/_0309_ ),
    .X(\Inst_RegFile_32x4/_0310_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0853_  (.A1(\Inst_RegFile_32x4/_0306_ ),
    .A2(\Inst_RegFile_32x4/_0308_ ),
    .B1(\Inst_RegFile_32x4/_0310_ ),
    .X(\Inst_RegFile_32x4/_0311_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0854_  (.A1(\Inst_RegFile_32x4/_0294_ ),
    .A2(\Inst_RegFile_32x4/_0301_ ),
    .B1(\Inst_RegFile_32x4/_0305_ ),
    .B2(\Inst_RegFile_32x4/_0311_ ),
    .X(\Inst_RegFile_32x4/_0312_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RegFile_32x4/_0855_  (.A(\Inst_RegFile_32x4/_0289_ ),
    .X(\Inst_RegFile_32x4/_0313_ ));
 sky130_fd_sc_hd__buf_2 \Inst_RegFile_32x4/_0856_  (.A(B_ADR0),
    .X(\Inst_RegFile_32x4/_0314_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0857_  (.A0(\Inst_RegFile_32x4/mem[8][0] ),
    .A1(\Inst_RegFile_32x4/mem[9][0] ),
    .S(\Inst_RegFile_32x4/_0314_ ),
    .X(\Inst_RegFile_32x4/_0315_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0858_  (.A_N(\Inst_RegFile_32x4/_0313_ ),
    .B(\Inst_RegFile_32x4/_0315_ ),
    .X(\Inst_RegFile_32x4/_0316_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0859_  (.A(\Inst_RegFile_32x4/_0291_ ),
    .X(\Inst_RegFile_32x4/_0317_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0860_  (.A0(\Inst_RegFile_32x4/mem[10][0] ),
    .A1(\Inst_RegFile_32x4/mem[11][0] ),
    .S(\Inst_RegFile_32x4/_0317_ ),
    .X(\Inst_RegFile_32x4/_0318_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0861_  (.A(B_ADR2),
    .X(\Inst_RegFile_32x4/_0319_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0862_  (.A1(\Inst_RegFile_32x4/_0302_ ),
    .A2(\Inst_RegFile_32x4/_0318_ ),
    .B1(\Inst_RegFile_32x4/_0319_ ),
    .X(\Inst_RegFile_32x4/_0320_ ));
 sky130_fd_sc_hd__buf_2 \Inst_RegFile_32x4/_0863_  (.A(\Inst_RegFile_32x4/_0297_ ),
    .X(\Inst_RegFile_32x4/_0321_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0864_  (.A(B_ADR1),
    .X(\Inst_RegFile_32x4/_0322_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0865_  (.A0(\Inst_RegFile_32x4/mem[12][0] ),
    .A1(\Inst_RegFile_32x4/mem[13][0] ),
    .A2(\Inst_RegFile_32x4/mem[14][0] ),
    .A3(\Inst_RegFile_32x4/mem[15][0] ),
    .S0(\Inst_RegFile_32x4/_0321_ ),
    .S1(\Inst_RegFile_32x4/_0322_ ),
    .X(\Inst_RegFile_32x4/_0323_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0866_  (.A(\Inst_RegFile_32x4/_0309_ ),
    .X(\Inst_RegFile_32x4/_0324_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0867_  (.A1(\Inst_RegFile_32x4/_0316_ ),
    .A2(\Inst_RegFile_32x4/_0320_ ),
    .B1(\Inst_RegFile_32x4/_0323_ ),
    .B2(\Inst_RegFile_32x4/_0324_ ),
    .X(\Inst_RegFile_32x4/_0325_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0868_  (.A(B_ADR0),
    .X(\Inst_RegFile_32x4/_0326_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0869_  (.A0(\Inst_RegFile_32x4/mem[16][0] ),
    .A1(\Inst_RegFile_32x4/mem[17][0] ),
    .S(\Inst_RegFile_32x4/_0326_ ),
    .X(\Inst_RegFile_32x4/_0327_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0870_  (.A_N(\Inst_RegFile_32x4/_0313_ ),
    .B(\Inst_RegFile_32x4/_0327_ ),
    .X(\Inst_RegFile_32x4/_0328_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0871_  (.A(\Inst_RegFile_32x4/_0295_ ),
    .X(\Inst_RegFile_32x4/_0329_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0872_  (.A(\Inst_RegFile_32x4/_0291_ ),
    .X(\Inst_RegFile_32x4/_0330_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0873_  (.A0(\Inst_RegFile_32x4/mem[18][0] ),
    .A1(\Inst_RegFile_32x4/mem[19][0] ),
    .S(\Inst_RegFile_32x4/_0330_ ),
    .X(\Inst_RegFile_32x4/_0331_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0874_  (.A(B_ADR2),
    .X(\Inst_RegFile_32x4/_0332_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0875_  (.A1(\Inst_RegFile_32x4/_0329_ ),
    .A2(\Inst_RegFile_32x4/_0331_ ),
    .B1(\Inst_RegFile_32x4/_0332_ ),
    .X(\Inst_RegFile_32x4/_0333_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RegFile_32x4/_0876_  (.A(\Inst_RegFile_32x4/_0289_ ),
    .X(\Inst_RegFile_32x4/_0334_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0877_  (.A(\Inst_RegFile_32x4/_0291_ ),
    .X(\Inst_RegFile_32x4/_0335_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0878_  (.A0(\Inst_RegFile_32x4/mem[20][0] ),
    .A1(\Inst_RegFile_32x4/mem[21][0] ),
    .S(\Inst_RegFile_32x4/_0335_ ),
    .X(\Inst_RegFile_32x4/_0336_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0879_  (.A_N(\Inst_RegFile_32x4/_0334_ ),
    .B(\Inst_RegFile_32x4/_0336_ ),
    .X(\Inst_RegFile_32x4/_0337_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0880_  (.A(\Inst_RegFile_32x4/_0297_ ),
    .X(\Inst_RegFile_32x4/_0338_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0881_  (.A0(\Inst_RegFile_32x4/mem[22][0] ),
    .A1(\Inst_RegFile_32x4/mem[23][0] ),
    .S(\Inst_RegFile_32x4/_0338_ ),
    .X(\Inst_RegFile_32x4/_0339_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0882_  (.A(\Inst_RegFile_32x4/_0309_ ),
    .X(\Inst_RegFile_32x4/_0340_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0883_  (.A1(\Inst_RegFile_32x4/_0306_ ),
    .A2(\Inst_RegFile_32x4/_0339_ ),
    .B1(\Inst_RegFile_32x4/_0340_ ),
    .X(\Inst_RegFile_32x4/_0341_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0884_  (.A1(\Inst_RegFile_32x4/_0328_ ),
    .A2(\Inst_RegFile_32x4/_0333_ ),
    .B1(\Inst_RegFile_32x4/_0337_ ),
    .B2(\Inst_RegFile_32x4/_0341_ ),
    .X(\Inst_RegFile_32x4/_0342_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_0885_  (.A(\Inst_RegFile_32x4/_0289_ ),
    .X(\Inst_RegFile_32x4/_0343_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0886_  (.A0(\Inst_RegFile_32x4/mem[24][0] ),
    .A1(\Inst_RegFile_32x4/mem[25][0] ),
    .S(\Inst_RegFile_32x4/_0292_ ),
    .X(\Inst_RegFile_32x4/_0344_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0887_  (.A_N(\Inst_RegFile_32x4/_0343_ ),
    .B(\Inst_RegFile_32x4/_0344_ ),
    .X(\Inst_RegFile_32x4/_0345_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_0888_  (.A(\Inst_RegFile_32x4/_0295_ ),
    .X(\Inst_RegFile_32x4/_0346_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0889_  (.A0(\Inst_RegFile_32x4/mem[26][0] ),
    .A1(\Inst_RegFile_32x4/mem[27][0] ),
    .S(\Inst_RegFile_32x4/_0330_ ),
    .X(\Inst_RegFile_32x4/_0347_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0890_  (.A1(\Inst_RegFile_32x4/_0346_ ),
    .A2(\Inst_RegFile_32x4/_0347_ ),
    .B1(\Inst_RegFile_32x4/_0300_ ),
    .X(\Inst_RegFile_32x4/_0348_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_0891_  (.A(B_ADR1),
    .X(\Inst_RegFile_32x4/_0349_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0892_  (.A0(\Inst_RegFile_32x4/mem[28][0] ),
    .A1(\Inst_RegFile_32x4/mem[29][0] ),
    .A2(\Inst_RegFile_32x4/mem[30][0] ),
    .A3(\Inst_RegFile_32x4/mem[31][0] ),
    .S0(\Inst_RegFile_32x4/_0321_ ),
    .S1(\Inst_RegFile_32x4/_0349_ ),
    .X(\Inst_RegFile_32x4/_0350_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0893_  (.A1(\Inst_RegFile_32x4/_0345_ ),
    .A2(\Inst_RegFile_32x4/_0348_ ),
    .B1(\Inst_RegFile_32x4/_0350_ ),
    .B2(\Inst_RegFile_32x4/_0324_ ),
    .X(\Inst_RegFile_32x4/_0351_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0894_  (.A0(\Inst_RegFile_32x4/_0312_ ),
    .A1(\Inst_RegFile_32x4/_0325_ ),
    .A2(\Inst_RegFile_32x4/_0342_ ),
    .A3(\Inst_RegFile_32x4/_0351_ ),
    .S0(B_ADR3),
    .S1(B_ADR4),
    .X(\Inst_RegFile_32x4/_0352_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_0895_  (.A(\Inst_RegFile_32x4/_0352_ ),
    .X(\Inst_RegFile_32x4/BD_comb[0] ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0896_  (.A0(\Inst_RegFile_32x4/BD_comb[0] ),
    .A1(\Inst_RegFile_32x4/BD_reg[0] ),
    .S(\ConfigBits[1] ),
    .X(\Inst_RegFile_32x4/_0353_ ));
 sky130_fd_sc_hd__buf_12 \Inst_RegFile_32x4/_0897_  (.A(\Inst_RegFile_32x4/_0353_ ),
    .X(BD0));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0898_  (.A0(\Inst_RegFile_32x4/mem[0][1] ),
    .A1(\Inst_RegFile_32x4/mem[1][1] ),
    .S(\Inst_RegFile_32x4/_0292_ ),
    .X(\Inst_RegFile_32x4/_0354_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0899_  (.A_N(\Inst_RegFile_32x4/_0290_ ),
    .B(\Inst_RegFile_32x4/_0354_ ),
    .X(\Inst_RegFile_32x4/_0355_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0900_  (.A0(\Inst_RegFile_32x4/mem[2][1] ),
    .A1(\Inst_RegFile_32x4/mem[3][1] ),
    .S(\Inst_RegFile_32x4/_0298_ ),
    .X(\Inst_RegFile_32x4/_0356_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0901_  (.A1(\Inst_RegFile_32x4/_0296_ ),
    .A2(\Inst_RegFile_32x4/_0356_ ),
    .B1(\Inst_RegFile_32x4/_0300_ ),
    .X(\Inst_RegFile_32x4/_0357_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0902_  (.A0(\Inst_RegFile_32x4/mem[4][1] ),
    .A1(\Inst_RegFile_32x4/mem[5][1] ),
    .S(\Inst_RegFile_32x4/_0303_ ),
    .X(\Inst_RegFile_32x4/_0358_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0903_  (.A_N(\Inst_RegFile_32x4/_0334_ ),
    .B(\Inst_RegFile_32x4/_0358_ ),
    .X(\Inst_RegFile_32x4/_0359_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0904_  (.A0(\Inst_RegFile_32x4/mem[6][1] ),
    .A1(\Inst_RegFile_32x4/mem[7][1] ),
    .S(\Inst_RegFile_32x4/_0307_ ),
    .X(\Inst_RegFile_32x4/_0360_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0905_  (.A1(\Inst_RegFile_32x4/_0306_ ),
    .A2(\Inst_RegFile_32x4/_0360_ ),
    .B1(\Inst_RegFile_32x4/_0310_ ),
    .X(\Inst_RegFile_32x4/_0361_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0906_  (.A1(\Inst_RegFile_32x4/_0355_ ),
    .A2(\Inst_RegFile_32x4/_0357_ ),
    .B1(\Inst_RegFile_32x4/_0359_ ),
    .B2(\Inst_RegFile_32x4/_0361_ ),
    .X(\Inst_RegFile_32x4/_0362_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0907_  (.A0(\Inst_RegFile_32x4/mem[8][1] ),
    .A1(\Inst_RegFile_32x4/mem[9][1] ),
    .S(\Inst_RegFile_32x4/_0314_ ),
    .X(\Inst_RegFile_32x4/_0363_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0908_  (.A_N(\Inst_RegFile_32x4/_0349_ ),
    .B(\Inst_RegFile_32x4/_0363_ ),
    .X(\Inst_RegFile_32x4/_0364_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0909_  (.A0(\Inst_RegFile_32x4/mem[10][1] ),
    .A1(\Inst_RegFile_32x4/mem[11][1] ),
    .S(\Inst_RegFile_32x4/_0317_ ),
    .X(\Inst_RegFile_32x4/_0365_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0910_  (.A1(\Inst_RegFile_32x4/_0302_ ),
    .A2(\Inst_RegFile_32x4/_0365_ ),
    .B1(\Inst_RegFile_32x4/_0319_ ),
    .X(\Inst_RegFile_32x4/_0366_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0911_  (.A0(\Inst_RegFile_32x4/mem[12][1] ),
    .A1(\Inst_RegFile_32x4/mem[13][1] ),
    .A2(\Inst_RegFile_32x4/mem[14][1] ),
    .A3(\Inst_RegFile_32x4/mem[15][1] ),
    .S0(\Inst_RegFile_32x4/_0307_ ),
    .S1(\Inst_RegFile_32x4/_0322_ ),
    .X(\Inst_RegFile_32x4/_0367_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0912_  (.A1(\Inst_RegFile_32x4/_0364_ ),
    .A2(\Inst_RegFile_32x4/_0366_ ),
    .B1(\Inst_RegFile_32x4/_0367_ ),
    .B2(\Inst_RegFile_32x4/_0310_ ),
    .X(\Inst_RegFile_32x4/_0368_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0913_  (.A0(\Inst_RegFile_32x4/mem[16][1] ),
    .A1(\Inst_RegFile_32x4/mem[17][1] ),
    .S(\Inst_RegFile_32x4/_0326_ ),
    .X(\Inst_RegFile_32x4/_0369_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0914_  (.A_N(\Inst_RegFile_32x4/_0313_ ),
    .B(\Inst_RegFile_32x4/_0369_ ),
    .X(\Inst_RegFile_32x4/_0370_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0915_  (.A0(\Inst_RegFile_32x4/mem[18][1] ),
    .A1(\Inst_RegFile_32x4/mem[19][1] ),
    .S(\Inst_RegFile_32x4/_0317_ ),
    .X(\Inst_RegFile_32x4/_0371_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0916_  (.A1(\Inst_RegFile_32x4/_0329_ ),
    .A2(\Inst_RegFile_32x4/_0371_ ),
    .B1(\Inst_RegFile_32x4/_0332_ ),
    .X(\Inst_RegFile_32x4/_0372_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0917_  (.A0(\Inst_RegFile_32x4/mem[20][1] ),
    .A1(\Inst_RegFile_32x4/mem[21][1] ),
    .S(\Inst_RegFile_32x4/_0335_ ),
    .X(\Inst_RegFile_32x4/_0373_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0918_  (.A_N(\Inst_RegFile_32x4/_0334_ ),
    .B(\Inst_RegFile_32x4/_0373_ ),
    .X(\Inst_RegFile_32x4/_0374_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0919_  (.A0(\Inst_RegFile_32x4/mem[22][1] ),
    .A1(\Inst_RegFile_32x4/mem[23][1] ),
    .S(\Inst_RegFile_32x4/_0338_ ),
    .X(\Inst_RegFile_32x4/_0375_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0920_  (.A1(\Inst_RegFile_32x4/_0296_ ),
    .A2(\Inst_RegFile_32x4/_0375_ ),
    .B1(\Inst_RegFile_32x4/_0340_ ),
    .X(\Inst_RegFile_32x4/_0376_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0921_  (.A1(\Inst_RegFile_32x4/_0370_ ),
    .A2(\Inst_RegFile_32x4/_0372_ ),
    .B1(\Inst_RegFile_32x4/_0374_ ),
    .B2(\Inst_RegFile_32x4/_0376_ ),
    .X(\Inst_RegFile_32x4/_0377_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0922_  (.A0(\Inst_RegFile_32x4/mem[24][1] ),
    .A1(\Inst_RegFile_32x4/mem[25][1] ),
    .S(\Inst_RegFile_32x4/_0326_ ),
    .X(\Inst_RegFile_32x4/_0378_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0923_  (.A_N(\Inst_RegFile_32x4/_0343_ ),
    .B(\Inst_RegFile_32x4/_0378_ ),
    .X(\Inst_RegFile_32x4/_0379_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0924_  (.A0(\Inst_RegFile_32x4/mem[26][1] ),
    .A1(\Inst_RegFile_32x4/mem[27][1] ),
    .S(\Inst_RegFile_32x4/_0330_ ),
    .X(\Inst_RegFile_32x4/_0380_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0925_  (.A1(\Inst_RegFile_32x4/_0346_ ),
    .A2(\Inst_RegFile_32x4/_0380_ ),
    .B1(\Inst_RegFile_32x4/_0332_ ),
    .X(\Inst_RegFile_32x4/_0381_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0926_  (.A0(\Inst_RegFile_32x4/mem[28][1] ),
    .A1(\Inst_RegFile_32x4/mem[29][1] ),
    .A2(\Inst_RegFile_32x4/mem[30][1] ),
    .A3(\Inst_RegFile_32x4/mem[31][1] ),
    .S0(\Inst_RegFile_32x4/_0321_ ),
    .S1(\Inst_RegFile_32x4/_0349_ ),
    .X(\Inst_RegFile_32x4/_0382_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0927_  (.A1(\Inst_RegFile_32x4/_0379_ ),
    .A2(\Inst_RegFile_32x4/_0381_ ),
    .B1(\Inst_RegFile_32x4/_0382_ ),
    .B2(\Inst_RegFile_32x4/_0324_ ),
    .X(\Inst_RegFile_32x4/_0383_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0928_  (.A0(\Inst_RegFile_32x4/_0362_ ),
    .A1(\Inst_RegFile_32x4/_0368_ ),
    .A2(\Inst_RegFile_32x4/_0377_ ),
    .A3(\Inst_RegFile_32x4/_0383_ ),
    .S0(B_ADR3),
    .S1(B_ADR4),
    .X(\Inst_RegFile_32x4/_0384_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_0929_  (.A(\Inst_RegFile_32x4/_0384_ ),
    .X(\Inst_RegFile_32x4/BD_comb[1] ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0930_  (.A0(\Inst_RegFile_32x4/BD_comb[1] ),
    .A1(\Inst_RegFile_32x4/BD_reg[1] ),
    .S(\ConfigBits[1] ),
    .X(\Inst_RegFile_32x4/_0385_ ));
 sky130_fd_sc_hd__buf_12 \Inst_RegFile_32x4/_0931_  (.A(\Inst_RegFile_32x4/_0385_ ),
    .X(BD1));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0932_  (.A0(\Inst_RegFile_32x4/mem[0][2] ),
    .A1(\Inst_RegFile_32x4/mem[1][2] ),
    .S(\Inst_RegFile_32x4/_0292_ ),
    .X(\Inst_RegFile_32x4/_0386_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0933_  (.A_N(\Inst_RegFile_32x4/_0290_ ),
    .B(\Inst_RegFile_32x4/_0386_ ),
    .X(\Inst_RegFile_32x4/_0387_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0934_  (.A0(\Inst_RegFile_32x4/mem[2][2] ),
    .A1(\Inst_RegFile_32x4/mem[3][2] ),
    .S(\Inst_RegFile_32x4/_0298_ ),
    .X(\Inst_RegFile_32x4/_0388_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0935_  (.A1(\Inst_RegFile_32x4/_0346_ ),
    .A2(\Inst_RegFile_32x4/_0388_ ),
    .B1(\Inst_RegFile_32x4/_0300_ ),
    .X(\Inst_RegFile_32x4/_0389_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0936_  (.A0(\Inst_RegFile_32x4/mem[4][2] ),
    .A1(\Inst_RegFile_32x4/mem[5][2] ),
    .S(\Inst_RegFile_32x4/_0303_ ),
    .X(\Inst_RegFile_32x4/_0390_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0937_  (.A_N(\Inst_RegFile_32x4/_0334_ ),
    .B(\Inst_RegFile_32x4/_0390_ ),
    .X(\Inst_RegFile_32x4/_0391_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0938_  (.A0(\Inst_RegFile_32x4/mem[6][2] ),
    .A1(\Inst_RegFile_32x4/mem[7][2] ),
    .S(\Inst_RegFile_32x4/_0338_ ),
    .X(\Inst_RegFile_32x4/_0392_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0939_  (.A1(\Inst_RegFile_32x4/_0306_ ),
    .A2(\Inst_RegFile_32x4/_0392_ ),
    .B1(\Inst_RegFile_32x4/_0340_ ),
    .X(\Inst_RegFile_32x4/_0393_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0940_  (.A1(\Inst_RegFile_32x4/_0387_ ),
    .A2(\Inst_RegFile_32x4/_0389_ ),
    .B1(\Inst_RegFile_32x4/_0391_ ),
    .B2(\Inst_RegFile_32x4/_0393_ ),
    .X(\Inst_RegFile_32x4/_0394_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0941_  (.A0(\Inst_RegFile_32x4/mem[8][2] ),
    .A1(\Inst_RegFile_32x4/mem[9][2] ),
    .S(\Inst_RegFile_32x4/_0314_ ),
    .X(\Inst_RegFile_32x4/_0395_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0942_  (.A_N(\Inst_RegFile_32x4/_0349_ ),
    .B(\Inst_RegFile_32x4/_0395_ ),
    .X(\Inst_RegFile_32x4/_0396_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0943_  (.A0(\Inst_RegFile_32x4/mem[10][2] ),
    .A1(\Inst_RegFile_32x4/mem[11][2] ),
    .S(\Inst_RegFile_32x4/_0303_ ),
    .X(\Inst_RegFile_32x4/_0397_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0944_  (.A1(\Inst_RegFile_32x4/_0302_ ),
    .A2(\Inst_RegFile_32x4/_0397_ ),
    .B1(\Inst_RegFile_32x4/_0319_ ),
    .X(\Inst_RegFile_32x4/_0398_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0945_  (.A0(\Inst_RegFile_32x4/mem[12][2] ),
    .A1(\Inst_RegFile_32x4/mem[13][2] ),
    .A2(\Inst_RegFile_32x4/mem[14][2] ),
    .A3(\Inst_RegFile_32x4/mem[15][2] ),
    .S0(\Inst_RegFile_32x4/_0307_ ),
    .S1(\Inst_RegFile_32x4/_0322_ ),
    .X(\Inst_RegFile_32x4/_0399_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0946_  (.A1(\Inst_RegFile_32x4/_0396_ ),
    .A2(\Inst_RegFile_32x4/_0398_ ),
    .B1(\Inst_RegFile_32x4/_0399_ ),
    .B2(\Inst_RegFile_32x4/_0310_ ),
    .X(\Inst_RegFile_32x4/_0400_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0947_  (.A0(\Inst_RegFile_32x4/mem[16][2] ),
    .A1(\Inst_RegFile_32x4/mem[17][2] ),
    .S(\Inst_RegFile_32x4/_0314_ ),
    .X(\Inst_RegFile_32x4/_0401_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0948_  (.A_N(\Inst_RegFile_32x4/_0313_ ),
    .B(\Inst_RegFile_32x4/_0401_ ),
    .X(\Inst_RegFile_32x4/_0402_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0949_  (.A0(\Inst_RegFile_32x4/mem[18][2] ),
    .A1(\Inst_RegFile_32x4/mem[19][2] ),
    .S(\Inst_RegFile_32x4/_0317_ ),
    .X(\Inst_RegFile_32x4/_0403_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0950_  (.A1(\Inst_RegFile_32x4/_0329_ ),
    .A2(\Inst_RegFile_32x4/_0403_ ),
    .B1(\Inst_RegFile_32x4/_0319_ ),
    .X(\Inst_RegFile_32x4/_0404_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0951_  (.A0(\Inst_RegFile_32x4/mem[20][2] ),
    .A1(\Inst_RegFile_32x4/mem[21][2] ),
    .S(\Inst_RegFile_32x4/_0335_ ),
    .X(\Inst_RegFile_32x4/_0405_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0952_  (.A_N(\Inst_RegFile_32x4/_0290_ ),
    .B(\Inst_RegFile_32x4/_0405_ ),
    .X(\Inst_RegFile_32x4/_0406_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0953_  (.A0(\Inst_RegFile_32x4/mem[22][2] ),
    .A1(\Inst_RegFile_32x4/mem[23][2] ),
    .S(\Inst_RegFile_32x4/_0338_ ),
    .X(\Inst_RegFile_32x4/_0407_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0954_  (.A1(\Inst_RegFile_32x4/_0296_ ),
    .A2(\Inst_RegFile_32x4/_0407_ ),
    .B1(\Inst_RegFile_32x4/_0340_ ),
    .X(\Inst_RegFile_32x4/_0408_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0955_  (.A1(\Inst_RegFile_32x4/_0402_ ),
    .A2(\Inst_RegFile_32x4/_0404_ ),
    .B1(\Inst_RegFile_32x4/_0406_ ),
    .B2(\Inst_RegFile_32x4/_0408_ ),
    .X(\Inst_RegFile_32x4/_0409_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0956_  (.A0(\Inst_RegFile_32x4/mem[24][2] ),
    .A1(\Inst_RegFile_32x4/mem[25][2] ),
    .S(\Inst_RegFile_32x4/_0326_ ),
    .X(\Inst_RegFile_32x4/_0410_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0957_  (.A_N(\Inst_RegFile_32x4/_0343_ ),
    .B(\Inst_RegFile_32x4/_0410_ ),
    .X(\Inst_RegFile_32x4/_0411_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0958_  (.A0(\Inst_RegFile_32x4/mem[26][2] ),
    .A1(\Inst_RegFile_32x4/mem[27][2] ),
    .S(\Inst_RegFile_32x4/_0330_ ),
    .X(\Inst_RegFile_32x4/_0412_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0959_  (.A1(\Inst_RegFile_32x4/_0346_ ),
    .A2(\Inst_RegFile_32x4/_0412_ ),
    .B1(\Inst_RegFile_32x4/_0332_ ),
    .X(\Inst_RegFile_32x4/_0413_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0960_  (.A0(\Inst_RegFile_32x4/mem[28][2] ),
    .A1(\Inst_RegFile_32x4/mem[29][2] ),
    .A2(\Inst_RegFile_32x4/mem[30][2] ),
    .A3(\Inst_RegFile_32x4/mem[31][2] ),
    .S0(\Inst_RegFile_32x4/_0321_ ),
    .S1(\Inst_RegFile_32x4/_0322_ ),
    .X(\Inst_RegFile_32x4/_0414_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0961_  (.A1(\Inst_RegFile_32x4/_0411_ ),
    .A2(\Inst_RegFile_32x4/_0413_ ),
    .B1(\Inst_RegFile_32x4/_0414_ ),
    .B2(\Inst_RegFile_32x4/_0324_ ),
    .X(\Inst_RegFile_32x4/_0415_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0962_  (.A0(\Inst_RegFile_32x4/_0394_ ),
    .A1(\Inst_RegFile_32x4/_0400_ ),
    .A2(\Inst_RegFile_32x4/_0409_ ),
    .A3(\Inst_RegFile_32x4/_0415_ ),
    .S0(B_ADR3),
    .S1(B_ADR4),
    .X(\Inst_RegFile_32x4/_0416_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_0963_  (.A(\Inst_RegFile_32x4/_0416_ ),
    .X(\Inst_RegFile_32x4/BD_comb[2] ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0964_  (.A0(\Inst_RegFile_32x4/BD_comb[2] ),
    .A1(\Inst_RegFile_32x4/BD_reg[2] ),
    .S(\ConfigBits[1] ),
    .X(\Inst_RegFile_32x4/_0417_ ));
 sky130_fd_sc_hd__buf_12 \Inst_RegFile_32x4/_0965_  (.A(\Inst_RegFile_32x4/_0417_ ),
    .X(BD2));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0966_  (.A0(\Inst_RegFile_32x4/mem[0][3] ),
    .A1(\Inst_RegFile_32x4/mem[1][3] ),
    .S(\Inst_RegFile_32x4/_0292_ ),
    .X(\Inst_RegFile_32x4/_0418_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0967_  (.A_N(\Inst_RegFile_32x4/_0343_ ),
    .B(\Inst_RegFile_32x4/_0418_ ),
    .X(\Inst_RegFile_32x4/_0419_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0968_  (.A0(\Inst_RegFile_32x4/mem[2][3] ),
    .A1(\Inst_RegFile_32x4/mem[3][3] ),
    .S(\Inst_RegFile_32x4/_0298_ ),
    .X(\Inst_RegFile_32x4/_0420_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0969_  (.A1(\Inst_RegFile_32x4/_0346_ ),
    .A2(\Inst_RegFile_32x4/_0420_ ),
    .B1(\Inst_RegFile_32x4/_0300_ ),
    .X(\Inst_RegFile_32x4/_0421_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0970_  (.A0(\Inst_RegFile_32x4/mem[4][3] ),
    .A1(\Inst_RegFile_32x4/mem[5][3] ),
    .S(\Inst_RegFile_32x4/_0335_ ),
    .X(\Inst_RegFile_32x4/_0422_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0971_  (.A_N(\Inst_RegFile_32x4/_0334_ ),
    .B(\Inst_RegFile_32x4/_0422_ ),
    .X(\Inst_RegFile_32x4/_0423_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0972_  (.A0(\Inst_RegFile_32x4/mem[6][3] ),
    .A1(\Inst_RegFile_32x4/mem[7][3] ),
    .S(\Inst_RegFile_32x4/_0338_ ),
    .X(\Inst_RegFile_32x4/_0424_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0973_  (.A1(\Inst_RegFile_32x4/_0306_ ),
    .A2(\Inst_RegFile_32x4/_0424_ ),
    .B1(\Inst_RegFile_32x4/_0340_ ),
    .X(\Inst_RegFile_32x4/_0425_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0974_  (.A1(\Inst_RegFile_32x4/_0419_ ),
    .A2(\Inst_RegFile_32x4/_0421_ ),
    .B1(\Inst_RegFile_32x4/_0423_ ),
    .B2(\Inst_RegFile_32x4/_0425_ ),
    .X(\Inst_RegFile_32x4/_0426_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0975_  (.A0(\Inst_RegFile_32x4/mem[8][3] ),
    .A1(\Inst_RegFile_32x4/mem[9][3] ),
    .S(\Inst_RegFile_32x4/_0297_ ),
    .X(\Inst_RegFile_32x4/_0427_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0976_  (.A_N(\Inst_RegFile_32x4/_0349_ ),
    .B(\Inst_RegFile_32x4/_0427_ ),
    .X(\Inst_RegFile_32x4/_0428_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0977_  (.A0(\Inst_RegFile_32x4/mem[10][3] ),
    .A1(\Inst_RegFile_32x4/mem[11][3] ),
    .S(\Inst_RegFile_32x4/_0303_ ),
    .X(\Inst_RegFile_32x4/_0429_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0978_  (.A1(\Inst_RegFile_32x4/_0302_ ),
    .A2(\Inst_RegFile_32x4/_0429_ ),
    .B1(B_ADR2),
    .X(\Inst_RegFile_32x4/_0430_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0979_  (.A0(\Inst_RegFile_32x4/mem[12][3] ),
    .A1(\Inst_RegFile_32x4/mem[13][3] ),
    .A2(\Inst_RegFile_32x4/mem[14][3] ),
    .A3(\Inst_RegFile_32x4/mem[15][3] ),
    .S0(\Inst_RegFile_32x4/_0307_ ),
    .S1(\Inst_RegFile_32x4/_0295_ ),
    .X(\Inst_RegFile_32x4/_0431_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0980_  (.A1(\Inst_RegFile_32x4/_0428_ ),
    .A2(\Inst_RegFile_32x4/_0430_ ),
    .B1(\Inst_RegFile_32x4/_0431_ ),
    .B2(\Inst_RegFile_32x4/_0310_ ),
    .X(\Inst_RegFile_32x4/_0432_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0981_  (.A0(\Inst_RegFile_32x4/mem[16][3] ),
    .A1(\Inst_RegFile_32x4/mem[17][3] ),
    .S(\Inst_RegFile_32x4/_0314_ ),
    .X(\Inst_RegFile_32x4/_0433_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0982_  (.A_N(\Inst_RegFile_32x4/_0313_ ),
    .B(\Inst_RegFile_32x4/_0433_ ),
    .X(\Inst_RegFile_32x4/_0434_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0983_  (.A0(\Inst_RegFile_32x4/mem[18][3] ),
    .A1(\Inst_RegFile_32x4/mem[19][3] ),
    .S(\Inst_RegFile_32x4/_0317_ ),
    .X(\Inst_RegFile_32x4/_0435_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0984_  (.A1(\Inst_RegFile_32x4/_0329_ ),
    .A2(\Inst_RegFile_32x4/_0435_ ),
    .B1(\Inst_RegFile_32x4/_0319_ ),
    .X(\Inst_RegFile_32x4/_0436_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0985_  (.A0(\Inst_RegFile_32x4/mem[20][3] ),
    .A1(\Inst_RegFile_32x4/mem[21][3] ),
    .S(\Inst_RegFile_32x4/_0335_ ),
    .X(\Inst_RegFile_32x4/_0437_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0986_  (.A_N(\Inst_RegFile_32x4/_0290_ ),
    .B(\Inst_RegFile_32x4/_0437_ ),
    .X(\Inst_RegFile_32x4/_0438_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0987_  (.A0(\Inst_RegFile_32x4/mem[22][3] ),
    .A1(\Inst_RegFile_32x4/mem[23][3] ),
    .S(\Inst_RegFile_32x4/_0298_ ),
    .X(\Inst_RegFile_32x4/_0439_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0988_  (.A1(\Inst_RegFile_32x4/_0296_ ),
    .A2(\Inst_RegFile_32x4/_0439_ ),
    .B1(\Inst_RegFile_32x4/_0309_ ),
    .X(\Inst_RegFile_32x4/_0440_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0989_  (.A1(\Inst_RegFile_32x4/_0434_ ),
    .A2(\Inst_RegFile_32x4/_0436_ ),
    .B1(\Inst_RegFile_32x4/_0438_ ),
    .B2(\Inst_RegFile_32x4/_0440_ ),
    .X(\Inst_RegFile_32x4/_0441_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0990_  (.A0(\Inst_RegFile_32x4/mem[24][3] ),
    .A1(\Inst_RegFile_32x4/mem[25][3] ),
    .S(\Inst_RegFile_32x4/_0326_ ),
    .X(\Inst_RegFile_32x4/_0442_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_RegFile_32x4/_0991_  (.A_N(\Inst_RegFile_32x4/_0343_ ),
    .B(\Inst_RegFile_32x4/_0442_ ),
    .X(\Inst_RegFile_32x4/_0443_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0992_  (.A0(\Inst_RegFile_32x4/mem[26][3] ),
    .A1(\Inst_RegFile_32x4/mem[27][3] ),
    .S(\Inst_RegFile_32x4/_0330_ ),
    .X(\Inst_RegFile_32x4/_0444_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_RegFile_32x4/_0993_  (.A1(\Inst_RegFile_32x4/_0329_ ),
    .A2(\Inst_RegFile_32x4/_0444_ ),
    .B1(\Inst_RegFile_32x4/_0332_ ),
    .X(\Inst_RegFile_32x4/_0445_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0994_  (.A0(\Inst_RegFile_32x4/mem[28][3] ),
    .A1(\Inst_RegFile_32x4/mem[29][3] ),
    .A2(\Inst_RegFile_32x4/mem[30][3] ),
    .A3(\Inst_RegFile_32x4/mem[31][3] ),
    .S0(\Inst_RegFile_32x4/_0321_ ),
    .S1(\Inst_RegFile_32x4/_0322_ ),
    .X(\Inst_RegFile_32x4/_0446_ ));
 sky130_fd_sc_hd__o22a_1 \Inst_RegFile_32x4/_0995_  (.A1(\Inst_RegFile_32x4/_0443_ ),
    .A2(\Inst_RegFile_32x4/_0445_ ),
    .B1(\Inst_RegFile_32x4/_0446_ ),
    .B2(\Inst_RegFile_32x4/_0324_ ),
    .X(\Inst_RegFile_32x4/_0447_ ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_32x4/_0996_  (.A0(\Inst_RegFile_32x4/_0426_ ),
    .A1(\Inst_RegFile_32x4/_0432_ ),
    .A2(\Inst_RegFile_32x4/_0441_ ),
    .A3(\Inst_RegFile_32x4/_0447_ ),
    .S0(B_ADR3),
    .S1(B_ADR4),
    .X(\Inst_RegFile_32x4/_0448_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_0997_  (.A(\Inst_RegFile_32x4/_0448_ ),
    .X(\Inst_RegFile_32x4/BD_comb[3] ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_0998_  (.A0(\Inst_RegFile_32x4/BD_comb[3] ),
    .A1(\Inst_RegFile_32x4/BD_reg[3] ),
    .S(\ConfigBits[1] ),
    .X(\Inst_RegFile_32x4/_0449_ ));
 sky130_fd_sc_hd__buf_12 \Inst_RegFile_32x4/_0999_  (.A(\Inst_RegFile_32x4/_0449_ ),
    .X(BD3));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1000_  (.A(D0),
    .X(\Inst_RegFile_32x4/_0450_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1001_  (.A(\Inst_RegFile_32x4/_0450_ ),
    .X(\Inst_RegFile_32x4/_0451_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_1002_  (.A(W_ADR4),
    .X(\Inst_RegFile_32x4/_0452_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_1003_  (.A(W_ADR3),
    .X(\Inst_RegFile_32x4/_0453_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_1004_  (.A(W_ADR2),
    .X(\Inst_RegFile_32x4/_0454_ ));
 sky130_fd_sc_hd__and3_2 \Inst_RegFile_32x4/_1005_  (.A(\Inst_RegFile_32x4/_0452_ ),
    .B(\Inst_RegFile_32x4/_0453_ ),
    .C(\Inst_RegFile_32x4/_0454_ ),
    .X(\Inst_RegFile_32x4/_0455_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1006_  (.A(W_ADR1),
    .X(\Inst_RegFile_32x4/_0456_ ));
 sky130_fd_sc_hd__buf_2 \Inst_RegFile_32x4/_1007_  (.A(W_en),
    .X(\Inst_RegFile_32x4/_0457_ ));
 sky130_fd_sc_hd__and3b_4 \Inst_RegFile_32x4/_1008_  (.A_N(\Inst_RegFile_32x4/_0456_ ),
    .B(W_ADR0),
    .C(\Inst_RegFile_32x4/_0457_ ),
    .X(\Inst_RegFile_32x4/_0458_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1009_  (.A(\Inst_RegFile_32x4/_0455_ ),
    .B(\Inst_RegFile_32x4/_0458_ ),
    .Y(\Inst_RegFile_32x4/_0459_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1010_  (.A0(\Inst_RegFile_32x4/_0451_ ),
    .A1(\Inst_RegFile_32x4/mem[29][0] ),
    .S(\Inst_RegFile_32x4/_0459_ ),
    .X(\Inst_RegFile_32x4/_0460_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1011_  (.A(\Inst_RegFile_32x4/_0460_ ),
    .X(\Inst_RegFile_32x4/_0000_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RegFile_32x4/_1012_  (.A(D1),
    .X(\Inst_RegFile_32x4/_0461_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1013_  (.A(\Inst_RegFile_32x4/_0461_ ),
    .X(\Inst_RegFile_32x4/_0462_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1014_  (.A0(\Inst_RegFile_32x4/_0462_ ),
    .A1(\Inst_RegFile_32x4/mem[29][1] ),
    .S(\Inst_RegFile_32x4/_0459_ ),
    .X(\Inst_RegFile_32x4/_0463_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1015_  (.A(\Inst_RegFile_32x4/_0463_ ),
    .X(\Inst_RegFile_32x4/_0001_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_1016_  (.A(D2),
    .X(\Inst_RegFile_32x4/_0464_ ));
 sky130_fd_sc_hd__buf_2 \Inst_RegFile_32x4/_1017_  (.A(\Inst_RegFile_32x4/_0464_ ),
    .X(\Inst_RegFile_32x4/_0465_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1018_  (.A0(\Inst_RegFile_32x4/_0465_ ),
    .A1(\Inst_RegFile_32x4/mem[29][2] ),
    .S(\Inst_RegFile_32x4/_0459_ ),
    .X(\Inst_RegFile_32x4/_0466_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1019_  (.A(\Inst_RegFile_32x4/_0466_ ),
    .X(\Inst_RegFile_32x4/_0002_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RegFile_32x4/_1020_  (.A(D3),
    .X(\Inst_RegFile_32x4/_0467_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1021_  (.A(\Inst_RegFile_32x4/_0467_ ),
    .X(\Inst_RegFile_32x4/_0468_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1022_  (.A0(\Inst_RegFile_32x4/_0468_ ),
    .A1(\Inst_RegFile_32x4/mem[29][3] ),
    .S(\Inst_RegFile_32x4/_0459_ ),
    .X(\Inst_RegFile_32x4/_0469_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1023_  (.A(\Inst_RegFile_32x4/_0469_ ),
    .X(\Inst_RegFile_32x4/_0003_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RegFile_32x4/_1024_  (.A(D0),
    .X(\Inst_RegFile_32x4/_0470_ ));
 sky130_fd_sc_hd__and3b_2 \Inst_RegFile_32x4/_1025_  (.A_N(W_ADR4),
    .B(W_ADR3),
    .C(W_ADR2),
    .X(\Inst_RegFile_32x4/_0471_ ));
 sky130_fd_sc_hd__or3b_1 \Inst_RegFile_32x4/_1026_  (.A(W_ADR1),
    .B(W_ADR0),
    .C_N(W_en),
    .X(\Inst_RegFile_32x4/_0472_ ));
 sky130_fd_sc_hd__clkbuf_4 \Inst_RegFile_32x4/_1027_  (.A(\Inst_RegFile_32x4/_0472_ ),
    .X(\Inst_RegFile_32x4/_0473_ ));
 sky130_fd_sc_hd__inv_2 \Inst_RegFile_32x4/_1028_  (.A(\Inst_RegFile_32x4/_0473_ ),
    .Y(\Inst_RegFile_32x4/_0474_ ));
 sky130_fd_sc_hd__and2_2 \Inst_RegFile_32x4/_1029_  (.A(\Inst_RegFile_32x4/_0471_ ),
    .B(\Inst_RegFile_32x4/_0474_ ),
    .X(\Inst_RegFile_32x4/_0475_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1030_  (.A0(\Inst_RegFile_32x4/mem[12][0] ),
    .A1(\Inst_RegFile_32x4/_0470_ ),
    .S(\Inst_RegFile_32x4/_0475_ ),
    .X(\Inst_RegFile_32x4/_0476_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1031_  (.A(\Inst_RegFile_32x4/_0476_ ),
    .X(\Inst_RegFile_32x4/_0004_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1032_  (.A(D1),
    .X(\Inst_RegFile_32x4/_0477_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1033_  (.A0(\Inst_RegFile_32x4/mem[12][1] ),
    .A1(\Inst_RegFile_32x4/_0477_ ),
    .S(\Inst_RegFile_32x4/_0475_ ),
    .X(\Inst_RegFile_32x4/_0478_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1034_  (.A(\Inst_RegFile_32x4/_0478_ ),
    .X(\Inst_RegFile_32x4/_0005_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1035_  (.A(D2),
    .X(\Inst_RegFile_32x4/_0479_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1036_  (.A0(\Inst_RegFile_32x4/mem[12][2] ),
    .A1(\Inst_RegFile_32x4/_0479_ ),
    .S(\Inst_RegFile_32x4/_0475_ ),
    .X(\Inst_RegFile_32x4/_0480_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1037_  (.A(\Inst_RegFile_32x4/_0480_ ),
    .X(\Inst_RegFile_32x4/_0006_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_1038_  (.A(D3),
    .X(\Inst_RegFile_32x4/_0481_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1039_  (.A0(\Inst_RegFile_32x4/mem[12][3] ),
    .A1(\Inst_RegFile_32x4/_0481_ ),
    .S(\Inst_RegFile_32x4/_0475_ ),
    .X(\Inst_RegFile_32x4/_0482_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1040_  (.A(\Inst_RegFile_32x4/_0482_ ),
    .X(\Inst_RegFile_32x4/_0007_ ));
 sky130_fd_sc_hd__or3b_4 \Inst_RegFile_32x4/_1041_  (.A(\Inst_RegFile_32x4/_0452_ ),
    .B(\Inst_RegFile_32x4/_0454_ ),
    .C_N(\Inst_RegFile_32x4/_0453_ ),
    .X(\Inst_RegFile_32x4/_0483_ ));
 sky130_fd_sc_hd__buf_2 \Inst_RegFile_32x4/_1042_  (.A(W_ADR0),
    .X(\Inst_RegFile_32x4/_0484_ ));
 sky130_fd_sc_hd__nand3_4 \Inst_RegFile_32x4/_1043_  (.A(\Inst_RegFile_32x4/_0456_ ),
    .B(\Inst_RegFile_32x4/_0484_ ),
    .C(\Inst_RegFile_32x4/_0457_ ),
    .Y(\Inst_RegFile_32x4/_0485_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1044_  (.A(\Inst_RegFile_32x4/_0483_ ),
    .B(\Inst_RegFile_32x4/_0485_ ),
    .Y(\Inst_RegFile_32x4/_0486_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1045_  (.A0(\Inst_RegFile_32x4/mem[11][0] ),
    .A1(\Inst_RegFile_32x4/_0470_ ),
    .S(\Inst_RegFile_32x4/_0486_ ),
    .X(\Inst_RegFile_32x4/_0487_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1046_  (.A(\Inst_RegFile_32x4/_0487_ ),
    .X(\Inst_RegFile_32x4/_0008_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1047_  (.A0(\Inst_RegFile_32x4/mem[11][1] ),
    .A1(\Inst_RegFile_32x4/_0477_ ),
    .S(\Inst_RegFile_32x4/_0486_ ),
    .X(\Inst_RegFile_32x4/_0488_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1048_  (.A(\Inst_RegFile_32x4/_0488_ ),
    .X(\Inst_RegFile_32x4/_0009_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1049_  (.A0(\Inst_RegFile_32x4/mem[11][2] ),
    .A1(\Inst_RegFile_32x4/_0479_ ),
    .S(\Inst_RegFile_32x4/_0486_ ),
    .X(\Inst_RegFile_32x4/_0489_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1050_  (.A(\Inst_RegFile_32x4/_0489_ ),
    .X(\Inst_RegFile_32x4/_0010_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1051_  (.A0(\Inst_RegFile_32x4/mem[11][3] ),
    .A1(\Inst_RegFile_32x4/_0481_ ),
    .S(\Inst_RegFile_32x4/_0486_ ),
    .X(\Inst_RegFile_32x4/_0490_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1052_  (.A(\Inst_RegFile_32x4/_0490_ ),
    .X(\Inst_RegFile_32x4/_0011_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1053_  (.A(\Inst_RegFile_32x4/_0450_ ),
    .X(\Inst_RegFile_32x4/_0491_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RegFile_32x4/_1054_  (.A(\Inst_RegFile_32x4/_0456_ ),
    .B(\Inst_RegFile_32x4/_0457_ ),
    .Y(\Inst_RegFile_32x4/_0492_ ));
 sky130_fd_sc_hd__or2_4 \Inst_RegFile_32x4/_1055_  (.A(\Inst_RegFile_32x4/_0484_ ),
    .B(\Inst_RegFile_32x4/_0492_ ),
    .X(\Inst_RegFile_32x4/_0493_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1056_  (.A(\Inst_RegFile_32x4/_0483_ ),
    .B(\Inst_RegFile_32x4/_0493_ ),
    .Y(\Inst_RegFile_32x4/_0494_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1057_  (.A0(\Inst_RegFile_32x4/mem[10][0] ),
    .A1(\Inst_RegFile_32x4/_0491_ ),
    .S(\Inst_RegFile_32x4/_0494_ ),
    .X(\Inst_RegFile_32x4/_0495_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1058_  (.A(\Inst_RegFile_32x4/_0495_ ),
    .X(\Inst_RegFile_32x4/_0012_ ));
 sky130_fd_sc_hd__buf_2 \Inst_RegFile_32x4/_1059_  (.A(\Inst_RegFile_32x4/_0461_ ),
    .X(\Inst_RegFile_32x4/_0496_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1060_  (.A0(\Inst_RegFile_32x4/mem[10][1] ),
    .A1(\Inst_RegFile_32x4/_0496_ ),
    .S(\Inst_RegFile_32x4/_0494_ ),
    .X(\Inst_RegFile_32x4/_0497_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1061_  (.A(\Inst_RegFile_32x4/_0497_ ),
    .X(\Inst_RegFile_32x4/_0013_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1062_  (.A(\Inst_RegFile_32x4/_0464_ ),
    .X(\Inst_RegFile_32x4/_0498_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1063_  (.A0(\Inst_RegFile_32x4/mem[10][2] ),
    .A1(\Inst_RegFile_32x4/_0498_ ),
    .S(\Inst_RegFile_32x4/_0494_ ),
    .X(\Inst_RegFile_32x4/_0499_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1064_  (.A(\Inst_RegFile_32x4/_0499_ ),
    .X(\Inst_RegFile_32x4/_0014_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1065_  (.A(\Inst_RegFile_32x4/_0467_ ),
    .X(\Inst_RegFile_32x4/_0500_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1066_  (.A0(\Inst_RegFile_32x4/mem[10][3] ),
    .A1(\Inst_RegFile_32x4/_0500_ ),
    .S(\Inst_RegFile_32x4/_0494_ ),
    .X(\Inst_RegFile_32x4/_0501_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1067_  (.A(\Inst_RegFile_32x4/_0501_ ),
    .X(\Inst_RegFile_32x4/_0015_ ));
 sky130_fd_sc_hd__or3_4 \Inst_RegFile_32x4/_1068_  (.A(\Inst_RegFile_32x4/_0452_ ),
    .B(\Inst_RegFile_32x4/_0453_ ),
    .C(\Inst_RegFile_32x4/_0454_ ),
    .X(\Inst_RegFile_32x4/_0502_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1069_  (.A(\Inst_RegFile_32x4/_0473_ ),
    .B(\Inst_RegFile_32x4/_0502_ ),
    .Y(\Inst_RegFile_32x4/_0503_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1070_  (.A0(\Inst_RegFile_32x4/mem[0][0] ),
    .A1(\Inst_RegFile_32x4/_0491_ ),
    .S(\Inst_RegFile_32x4/_0503_ ),
    .X(\Inst_RegFile_32x4/_0504_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1071_  (.A(\Inst_RegFile_32x4/_0504_ ),
    .X(\Inst_RegFile_32x4/_0016_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1072_  (.A0(\Inst_RegFile_32x4/mem[0][1] ),
    .A1(\Inst_RegFile_32x4/_0496_ ),
    .S(\Inst_RegFile_32x4/_0503_ ),
    .X(\Inst_RegFile_32x4/_0505_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1073_  (.A(\Inst_RegFile_32x4/_0505_ ),
    .X(\Inst_RegFile_32x4/_0017_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1074_  (.A0(\Inst_RegFile_32x4/mem[0][2] ),
    .A1(\Inst_RegFile_32x4/_0498_ ),
    .S(\Inst_RegFile_32x4/_0503_ ),
    .X(\Inst_RegFile_32x4/_0506_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1075_  (.A(\Inst_RegFile_32x4/_0506_ ),
    .X(\Inst_RegFile_32x4/_0018_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1076_  (.A0(\Inst_RegFile_32x4/mem[0][3] ),
    .A1(\Inst_RegFile_32x4/_0500_ ),
    .S(\Inst_RegFile_32x4/_0503_ ),
    .X(\Inst_RegFile_32x4/_0507_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1077_  (.A(\Inst_RegFile_32x4/_0507_ ),
    .X(\Inst_RegFile_32x4/_0019_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1078_  (.A(\Inst_RegFile_32x4/_0473_ ),
    .B(\Inst_RegFile_32x4/_0483_ ),
    .Y(\Inst_RegFile_32x4/_0508_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1079_  (.A0(\Inst_RegFile_32x4/mem[8][0] ),
    .A1(\Inst_RegFile_32x4/_0491_ ),
    .S(\Inst_RegFile_32x4/_0508_ ),
    .X(\Inst_RegFile_32x4/_0509_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1080_  (.A(\Inst_RegFile_32x4/_0509_ ),
    .X(\Inst_RegFile_32x4/_0020_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1081_  (.A0(\Inst_RegFile_32x4/mem[8][1] ),
    .A1(\Inst_RegFile_32x4/_0496_ ),
    .S(\Inst_RegFile_32x4/_0508_ ),
    .X(\Inst_RegFile_32x4/_0510_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1082_  (.A(\Inst_RegFile_32x4/_0510_ ),
    .X(\Inst_RegFile_32x4/_0021_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1083_  (.A0(\Inst_RegFile_32x4/mem[8][2] ),
    .A1(\Inst_RegFile_32x4/_0498_ ),
    .S(\Inst_RegFile_32x4/_0508_ ),
    .X(\Inst_RegFile_32x4/_0511_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1084_  (.A(\Inst_RegFile_32x4/_0511_ ),
    .X(\Inst_RegFile_32x4/_0022_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1085_  (.A0(\Inst_RegFile_32x4/mem[8][3] ),
    .A1(\Inst_RegFile_32x4/_0500_ ),
    .S(\Inst_RegFile_32x4/_0508_ ),
    .X(\Inst_RegFile_32x4/_0512_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1086_  (.A(\Inst_RegFile_32x4/_0512_ ),
    .X(\Inst_RegFile_32x4/_0023_ ));
 sky130_fd_sc_hd__or3b_4 \Inst_RegFile_32x4/_1087_  (.A(\Inst_RegFile_32x4/_0452_ ),
    .B(\Inst_RegFile_32x4/_0453_ ),
    .C_N(\Inst_RegFile_32x4/_0454_ ),
    .X(\Inst_RegFile_32x4/_0513_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1088_  (.A(\Inst_RegFile_32x4/_0485_ ),
    .B(\Inst_RegFile_32x4/_0513_ ),
    .Y(\Inst_RegFile_32x4/_0514_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1089_  (.A0(\Inst_RegFile_32x4/mem[7][0] ),
    .A1(\Inst_RegFile_32x4/_0491_ ),
    .S(\Inst_RegFile_32x4/_0514_ ),
    .X(\Inst_RegFile_32x4/_0515_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1090_  (.A(\Inst_RegFile_32x4/_0515_ ),
    .X(\Inst_RegFile_32x4/_0024_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1091_  (.A0(\Inst_RegFile_32x4/mem[7][1] ),
    .A1(\Inst_RegFile_32x4/_0496_ ),
    .S(\Inst_RegFile_32x4/_0514_ ),
    .X(\Inst_RegFile_32x4/_0516_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1092_  (.A(\Inst_RegFile_32x4/_0516_ ),
    .X(\Inst_RegFile_32x4/_0025_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1093_  (.A0(\Inst_RegFile_32x4/mem[7][2] ),
    .A1(\Inst_RegFile_32x4/_0498_ ),
    .S(\Inst_RegFile_32x4/_0514_ ),
    .X(\Inst_RegFile_32x4/_0517_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1094_  (.A(\Inst_RegFile_32x4/_0517_ ),
    .X(\Inst_RegFile_32x4/_0026_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1095_  (.A0(\Inst_RegFile_32x4/mem[7][3] ),
    .A1(\Inst_RegFile_32x4/_0500_ ),
    .S(\Inst_RegFile_32x4/_0514_ ),
    .X(\Inst_RegFile_32x4/_0518_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1096_  (.A(\Inst_RegFile_32x4/_0518_ ),
    .X(\Inst_RegFile_32x4/_0027_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1097_  (.A(\Inst_RegFile_32x4/_0493_ ),
    .B(\Inst_RegFile_32x4/_0513_ ),
    .Y(\Inst_RegFile_32x4/_0519_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1098_  (.A0(\Inst_RegFile_32x4/mem[6][0] ),
    .A1(\Inst_RegFile_32x4/_0491_ ),
    .S(\Inst_RegFile_32x4/_0519_ ),
    .X(\Inst_RegFile_32x4/_0520_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1099_  (.A(\Inst_RegFile_32x4/_0520_ ),
    .X(\Inst_RegFile_32x4/_0028_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1100_  (.A0(\Inst_RegFile_32x4/mem[6][1] ),
    .A1(\Inst_RegFile_32x4/_0496_ ),
    .S(\Inst_RegFile_32x4/_0519_ ),
    .X(\Inst_RegFile_32x4/_0521_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1101_  (.A(\Inst_RegFile_32x4/_0521_ ),
    .X(\Inst_RegFile_32x4/_0029_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1102_  (.A0(\Inst_RegFile_32x4/mem[6][2] ),
    .A1(\Inst_RegFile_32x4/_0498_ ),
    .S(\Inst_RegFile_32x4/_0519_ ),
    .X(\Inst_RegFile_32x4/_0522_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1103_  (.A(\Inst_RegFile_32x4/_0522_ ),
    .X(\Inst_RegFile_32x4/_0030_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1104_  (.A0(\Inst_RegFile_32x4/mem[6][3] ),
    .A1(\Inst_RegFile_32x4/_0500_ ),
    .S(\Inst_RegFile_32x4/_0519_ ),
    .X(\Inst_RegFile_32x4/_0523_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1105_  (.A(\Inst_RegFile_32x4/_0523_ ),
    .X(\Inst_RegFile_32x4/_0031_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RegFile_32x4/_1106_  (.A(D0),
    .X(\Inst_RegFile_32x4/_0524_ ));
 sky130_fd_sc_hd__nand3b_4 \Inst_RegFile_32x4/_1107_  (.A_N(\Inst_RegFile_32x4/_0456_ ),
    .B(\Inst_RegFile_32x4/_0484_ ),
    .C(\Inst_RegFile_32x4/_0457_ ),
    .Y(\Inst_RegFile_32x4/_0525_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1108_  (.A(\Inst_RegFile_32x4/_0525_ ),
    .B(\Inst_RegFile_32x4/_0513_ ),
    .Y(\Inst_RegFile_32x4/_0526_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1109_  (.A0(\Inst_RegFile_32x4/mem[5][0] ),
    .A1(\Inst_RegFile_32x4/_0524_ ),
    .S(\Inst_RegFile_32x4/_0526_ ),
    .X(\Inst_RegFile_32x4/_0527_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1110_  (.A(\Inst_RegFile_32x4/_0527_ ),
    .X(\Inst_RegFile_32x4/_0032_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1111_  (.A(D1),
    .X(\Inst_RegFile_32x4/_0528_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1112_  (.A0(\Inst_RegFile_32x4/mem[5][1] ),
    .A1(\Inst_RegFile_32x4/_0528_ ),
    .S(\Inst_RegFile_32x4/_0526_ ),
    .X(\Inst_RegFile_32x4/_0529_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1113_  (.A(\Inst_RegFile_32x4/_0529_ ),
    .X(\Inst_RegFile_32x4/_0033_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1114_  (.A(D2),
    .X(\Inst_RegFile_32x4/_0530_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1115_  (.A0(\Inst_RegFile_32x4/mem[5][2] ),
    .A1(\Inst_RegFile_32x4/_0530_ ),
    .S(\Inst_RegFile_32x4/_0526_ ),
    .X(\Inst_RegFile_32x4/_0531_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1116_  (.A(\Inst_RegFile_32x4/_0531_ ),
    .X(\Inst_RegFile_32x4/_0034_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1117_  (.A(D3),
    .X(\Inst_RegFile_32x4/_0532_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1118_  (.A0(\Inst_RegFile_32x4/mem[5][3] ),
    .A1(\Inst_RegFile_32x4/_0532_ ),
    .S(\Inst_RegFile_32x4/_0526_ ),
    .X(\Inst_RegFile_32x4/_0533_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1119_  (.A(\Inst_RegFile_32x4/_0533_ ),
    .X(\Inst_RegFile_32x4/_0035_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1120_  (.A(\Inst_RegFile_32x4/_0473_ ),
    .B(\Inst_RegFile_32x4/_0513_ ),
    .Y(\Inst_RegFile_32x4/_0534_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1121_  (.A0(\Inst_RegFile_32x4/mem[4][0] ),
    .A1(\Inst_RegFile_32x4/_0524_ ),
    .S(\Inst_RegFile_32x4/_0534_ ),
    .X(\Inst_RegFile_32x4/_0535_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1122_  (.A(\Inst_RegFile_32x4/_0535_ ),
    .X(\Inst_RegFile_32x4/_0036_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1123_  (.A0(\Inst_RegFile_32x4/mem[4][1] ),
    .A1(\Inst_RegFile_32x4/_0528_ ),
    .S(\Inst_RegFile_32x4/_0534_ ),
    .X(\Inst_RegFile_32x4/_0536_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1124_  (.A(\Inst_RegFile_32x4/_0536_ ),
    .X(\Inst_RegFile_32x4/_0037_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1125_  (.A0(\Inst_RegFile_32x4/mem[4][2] ),
    .A1(\Inst_RegFile_32x4/_0530_ ),
    .S(\Inst_RegFile_32x4/_0534_ ),
    .X(\Inst_RegFile_32x4/_0537_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1126_  (.A(\Inst_RegFile_32x4/_0537_ ),
    .X(\Inst_RegFile_32x4/_0038_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1127_  (.A0(\Inst_RegFile_32x4/mem[4][3] ),
    .A1(\Inst_RegFile_32x4/_0532_ ),
    .S(\Inst_RegFile_32x4/_0534_ ),
    .X(\Inst_RegFile_32x4/_0538_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1128_  (.A(\Inst_RegFile_32x4/_0538_ ),
    .X(\Inst_RegFile_32x4/_0039_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1129_  (.A(\Inst_RegFile_32x4/_0485_ ),
    .B(\Inst_RegFile_32x4/_0502_ ),
    .Y(\Inst_RegFile_32x4/_0539_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1130_  (.A0(\Inst_RegFile_32x4/mem[3][0] ),
    .A1(\Inst_RegFile_32x4/_0524_ ),
    .S(\Inst_RegFile_32x4/_0539_ ),
    .X(\Inst_RegFile_32x4/_0540_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1131_  (.A(\Inst_RegFile_32x4/_0540_ ),
    .X(\Inst_RegFile_32x4/_0040_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1132_  (.A0(\Inst_RegFile_32x4/mem[3][1] ),
    .A1(\Inst_RegFile_32x4/_0528_ ),
    .S(\Inst_RegFile_32x4/_0539_ ),
    .X(\Inst_RegFile_32x4/_0541_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1133_  (.A(\Inst_RegFile_32x4/_0541_ ),
    .X(\Inst_RegFile_32x4/_0041_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1134_  (.A0(\Inst_RegFile_32x4/mem[3][2] ),
    .A1(\Inst_RegFile_32x4/_0530_ ),
    .S(\Inst_RegFile_32x4/_0539_ ),
    .X(\Inst_RegFile_32x4/_0542_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1135_  (.A(\Inst_RegFile_32x4/_0542_ ),
    .X(\Inst_RegFile_32x4/_0042_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1136_  (.A0(\Inst_RegFile_32x4/mem[3][3] ),
    .A1(\Inst_RegFile_32x4/_0532_ ),
    .S(\Inst_RegFile_32x4/_0539_ ),
    .X(\Inst_RegFile_32x4/_0543_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1137_  (.A(\Inst_RegFile_32x4/_0543_ ),
    .X(\Inst_RegFile_32x4/_0043_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1138_  (.A(\Inst_RegFile_32x4/_0458_ ),
    .B(\Inst_RegFile_32x4/_0471_ ),
    .Y(\Inst_RegFile_32x4/_0544_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1139_  (.A0(\Inst_RegFile_32x4/_0451_ ),
    .A1(\Inst_RegFile_32x4/mem[13][0] ),
    .S(\Inst_RegFile_32x4/_0544_ ),
    .X(\Inst_RegFile_32x4/_0545_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1140_  (.A(\Inst_RegFile_32x4/_0545_ ),
    .X(\Inst_RegFile_32x4/_0044_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1141_  (.A0(\Inst_RegFile_32x4/_0462_ ),
    .A1(\Inst_RegFile_32x4/mem[13][1] ),
    .S(\Inst_RegFile_32x4/_0544_ ),
    .X(\Inst_RegFile_32x4/_0546_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1142_  (.A(\Inst_RegFile_32x4/_0546_ ),
    .X(\Inst_RegFile_32x4/_0045_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1143_  (.A0(\Inst_RegFile_32x4/_0465_ ),
    .A1(\Inst_RegFile_32x4/mem[13][2] ),
    .S(\Inst_RegFile_32x4/_0544_ ),
    .X(\Inst_RegFile_32x4/_0547_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1144_  (.A(\Inst_RegFile_32x4/_0547_ ),
    .X(\Inst_RegFile_32x4/_0046_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1145_  (.A0(\Inst_RegFile_32x4/_0468_ ),
    .A1(\Inst_RegFile_32x4/mem[13][3] ),
    .S(\Inst_RegFile_32x4/_0544_ ),
    .X(\Inst_RegFile_32x4/_0548_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1146_  (.A(\Inst_RegFile_32x4/_0548_ ),
    .X(\Inst_RegFile_32x4/_0047_ ));
 sky130_fd_sc_hd__nor2_1 \Inst_RegFile_32x4/_1147_  (.A(\Inst_RegFile_32x4/_0525_ ),
    .B(\Inst_RegFile_32x4/_0483_ ),
    .Y(\Inst_RegFile_32x4/_0549_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1148_  (.A0(\Inst_RegFile_32x4/mem[9][0] ),
    .A1(\Inst_RegFile_32x4/_0524_ ),
    .S(\Inst_RegFile_32x4/_0549_ ),
    .X(\Inst_RegFile_32x4/_0550_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1149_  (.A(\Inst_RegFile_32x4/_0550_ ),
    .X(\Inst_RegFile_32x4/_0048_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1150_  (.A0(\Inst_RegFile_32x4/mem[9][1] ),
    .A1(\Inst_RegFile_32x4/_0528_ ),
    .S(\Inst_RegFile_32x4/_0549_ ),
    .X(\Inst_RegFile_32x4/_0551_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1151_  (.A(\Inst_RegFile_32x4/_0551_ ),
    .X(\Inst_RegFile_32x4/_0049_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1152_  (.A0(\Inst_RegFile_32x4/mem[9][2] ),
    .A1(\Inst_RegFile_32x4/_0530_ ),
    .S(\Inst_RegFile_32x4/_0549_ ),
    .X(\Inst_RegFile_32x4/_0552_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1153_  (.A(\Inst_RegFile_32x4/_0552_ ),
    .X(\Inst_RegFile_32x4/_0050_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1154_  (.A0(\Inst_RegFile_32x4/mem[9][3] ),
    .A1(\Inst_RegFile_32x4/_0532_ ),
    .S(\Inst_RegFile_32x4/_0549_ ),
    .X(\Inst_RegFile_32x4/_0553_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1155_  (.A(\Inst_RegFile_32x4/_0553_ ),
    .X(\Inst_RegFile_32x4/_0051_ ));
 sky130_fd_sc_hd__nor2_4 \Inst_RegFile_32x4/_1156_  (.A(\Inst_RegFile_32x4/_0484_ ),
    .B(\Inst_RegFile_32x4/_0492_ ),
    .Y(\Inst_RegFile_32x4/_0554_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1157_  (.A(\Inst_RegFile_32x4/_0455_ ),
    .B(\Inst_RegFile_32x4/_0554_ ),
    .Y(\Inst_RegFile_32x4/_0555_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1158_  (.A0(\Inst_RegFile_32x4/_0451_ ),
    .A1(\Inst_RegFile_32x4/mem[30][0] ),
    .S(\Inst_RegFile_32x4/_0555_ ),
    .X(\Inst_RegFile_32x4/_0556_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1159_  (.A(\Inst_RegFile_32x4/_0556_ ),
    .X(\Inst_RegFile_32x4/_0052_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1160_  (.A0(\Inst_RegFile_32x4/_0462_ ),
    .A1(\Inst_RegFile_32x4/mem[30][1] ),
    .S(\Inst_RegFile_32x4/_0555_ ),
    .X(\Inst_RegFile_32x4/_0557_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1161_  (.A(\Inst_RegFile_32x4/_0557_ ),
    .X(\Inst_RegFile_32x4/_0053_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1162_  (.A0(\Inst_RegFile_32x4/_0465_ ),
    .A1(\Inst_RegFile_32x4/mem[30][2] ),
    .S(\Inst_RegFile_32x4/_0555_ ),
    .X(\Inst_RegFile_32x4/_0558_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1163_  (.A(\Inst_RegFile_32x4/_0558_ ),
    .X(\Inst_RegFile_32x4/_0054_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1164_  (.A0(\Inst_RegFile_32x4/_0468_ ),
    .A1(\Inst_RegFile_32x4/mem[30][3] ),
    .S(\Inst_RegFile_32x4/_0555_ ),
    .X(\Inst_RegFile_32x4/_0559_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1165_  (.A(\Inst_RegFile_32x4/_0559_ ),
    .X(\Inst_RegFile_32x4/_0055_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1166_  (.A(\Inst_RegFile_32x4/_0493_ ),
    .B(\Inst_RegFile_32x4/_0502_ ),
    .Y(\Inst_RegFile_32x4/_0560_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1167_  (.A0(\Inst_RegFile_32x4/mem[2][0] ),
    .A1(\Inst_RegFile_32x4/_0524_ ),
    .S(\Inst_RegFile_32x4/_0560_ ),
    .X(\Inst_RegFile_32x4/_0561_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1168_  (.A(\Inst_RegFile_32x4/_0561_ ),
    .X(\Inst_RegFile_32x4/_0056_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1169_  (.A0(\Inst_RegFile_32x4/mem[2][1] ),
    .A1(\Inst_RegFile_32x4/_0528_ ),
    .S(\Inst_RegFile_32x4/_0560_ ),
    .X(\Inst_RegFile_32x4/_0562_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1170_  (.A(\Inst_RegFile_32x4/_0562_ ),
    .X(\Inst_RegFile_32x4/_0057_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1171_  (.A0(\Inst_RegFile_32x4/mem[2][2] ),
    .A1(\Inst_RegFile_32x4/_0530_ ),
    .S(\Inst_RegFile_32x4/_0560_ ),
    .X(\Inst_RegFile_32x4/_0563_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1172_  (.A(\Inst_RegFile_32x4/_0563_ ),
    .X(\Inst_RegFile_32x4/_0058_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1173_  (.A0(\Inst_RegFile_32x4/mem[2][3] ),
    .A1(\Inst_RegFile_32x4/_0532_ ),
    .S(\Inst_RegFile_32x4/_0560_ ),
    .X(\Inst_RegFile_32x4/_0564_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1174_  (.A(\Inst_RegFile_32x4/_0564_ ),
    .X(\Inst_RegFile_32x4/_0059_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1175_  (.A(\Inst_RegFile_32x4/_0455_ ),
    .B(\Inst_RegFile_32x4/_0474_ ),
    .Y(\Inst_RegFile_32x4/_0565_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1176_  (.A0(\Inst_RegFile_32x4/_0451_ ),
    .A1(\Inst_RegFile_32x4/mem[28][0] ),
    .S(\Inst_RegFile_32x4/_0565_ ),
    .X(\Inst_RegFile_32x4/_0566_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1177_  (.A(\Inst_RegFile_32x4/_0566_ ),
    .X(\Inst_RegFile_32x4/_0060_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1178_  (.A0(\Inst_RegFile_32x4/_0462_ ),
    .A1(\Inst_RegFile_32x4/mem[28][1] ),
    .S(\Inst_RegFile_32x4/_0565_ ),
    .X(\Inst_RegFile_32x4/_0567_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1179_  (.A(\Inst_RegFile_32x4/_0567_ ),
    .X(\Inst_RegFile_32x4/_0061_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1180_  (.A0(\Inst_RegFile_32x4/_0465_ ),
    .A1(\Inst_RegFile_32x4/mem[28][2] ),
    .S(\Inst_RegFile_32x4/_0565_ ),
    .X(\Inst_RegFile_32x4/_0568_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1181_  (.A(\Inst_RegFile_32x4/_0568_ ),
    .X(\Inst_RegFile_32x4/_0062_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1182_  (.A0(\Inst_RegFile_32x4/_0468_ ),
    .A1(\Inst_RegFile_32x4/mem[28][3] ),
    .S(\Inst_RegFile_32x4/_0565_ ),
    .X(\Inst_RegFile_32x4/_0569_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1183_  (.A(\Inst_RegFile_32x4/_0569_ ),
    .X(\Inst_RegFile_32x4/_0063_ ));
 sky130_fd_sc_hd__and3_2 \Inst_RegFile_32x4/_1184_  (.A(\Inst_RegFile_32x4/_0456_ ),
    .B(\Inst_RegFile_32x4/_0484_ ),
    .C(\Inst_RegFile_32x4/_0457_ ),
    .X(\Inst_RegFile_32x4/_0570_ ));
 sky130_fd_sc_hd__and3b_2 \Inst_RegFile_32x4/_1185_  (.A_N(W_ADR2),
    .B(W_ADR3),
    .C(W_ADR4),
    .X(\Inst_RegFile_32x4/_0571_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1186_  (.A(\Inst_RegFile_32x4/_0570_ ),
    .B(\Inst_RegFile_32x4/_0571_ ),
    .Y(\Inst_RegFile_32x4/_0572_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1187_  (.A0(\Inst_RegFile_32x4/_0451_ ),
    .A1(\Inst_RegFile_32x4/mem[27][0] ),
    .S(\Inst_RegFile_32x4/_0572_ ),
    .X(\Inst_RegFile_32x4/_0573_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1188_  (.A(\Inst_RegFile_32x4/_0573_ ),
    .X(\Inst_RegFile_32x4/_0064_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1189_  (.A0(\Inst_RegFile_32x4/_0462_ ),
    .A1(\Inst_RegFile_32x4/mem[27][1] ),
    .S(\Inst_RegFile_32x4/_0572_ ),
    .X(\Inst_RegFile_32x4/_0574_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1190_  (.A(\Inst_RegFile_32x4/_0574_ ),
    .X(\Inst_RegFile_32x4/_0065_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1191_  (.A0(\Inst_RegFile_32x4/_0465_ ),
    .A1(\Inst_RegFile_32x4/mem[27][2] ),
    .S(\Inst_RegFile_32x4/_0572_ ),
    .X(\Inst_RegFile_32x4/_0575_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1192_  (.A(\Inst_RegFile_32x4/_0575_ ),
    .X(\Inst_RegFile_32x4/_0066_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1193_  (.A0(\Inst_RegFile_32x4/_0468_ ),
    .A1(\Inst_RegFile_32x4/mem[27][3] ),
    .S(\Inst_RegFile_32x4/_0572_ ),
    .X(\Inst_RegFile_32x4/_0576_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1194_  (.A(\Inst_RegFile_32x4/_0576_ ),
    .X(\Inst_RegFile_32x4/_0067_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_32x4/_1195_  (.A(\Inst_RegFile_32x4/_0450_ ),
    .X(\Inst_RegFile_32x4/_0577_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1196_  (.A(\Inst_RegFile_32x4/_0554_ ),
    .B(\Inst_RegFile_32x4/_0571_ ),
    .Y(\Inst_RegFile_32x4/_0578_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1197_  (.A0(\Inst_RegFile_32x4/_0577_ ),
    .A1(\Inst_RegFile_32x4/mem[26][0] ),
    .S(\Inst_RegFile_32x4/_0578_ ),
    .X(\Inst_RegFile_32x4/_0579_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1198_  (.A(\Inst_RegFile_32x4/_0579_ ),
    .X(\Inst_RegFile_32x4/_0068_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1199_  (.A(\Inst_RegFile_32x4/_0461_ ),
    .X(\Inst_RegFile_32x4/_0580_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1200_  (.A0(\Inst_RegFile_32x4/_0580_ ),
    .A1(\Inst_RegFile_32x4/mem[26][1] ),
    .S(\Inst_RegFile_32x4/_0578_ ),
    .X(\Inst_RegFile_32x4/_0581_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1201_  (.A(\Inst_RegFile_32x4/_0581_ ),
    .X(\Inst_RegFile_32x4/_0069_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1202_  (.A(\Inst_RegFile_32x4/_0464_ ),
    .X(\Inst_RegFile_32x4/_0582_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1203_  (.A0(\Inst_RegFile_32x4/_0582_ ),
    .A1(\Inst_RegFile_32x4/mem[26][2] ),
    .S(\Inst_RegFile_32x4/_0578_ ),
    .X(\Inst_RegFile_32x4/_0583_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1204_  (.A(\Inst_RegFile_32x4/_0583_ ),
    .X(\Inst_RegFile_32x4/_0070_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1205_  (.A(\Inst_RegFile_32x4/_0467_ ),
    .X(\Inst_RegFile_32x4/_0584_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1206_  (.A0(\Inst_RegFile_32x4/_0584_ ),
    .A1(\Inst_RegFile_32x4/mem[26][3] ),
    .S(\Inst_RegFile_32x4/_0578_ ),
    .X(\Inst_RegFile_32x4/_0585_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1207_  (.A(\Inst_RegFile_32x4/_0585_ ),
    .X(\Inst_RegFile_32x4/_0071_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1208_  (.A(\Inst_RegFile_32x4/_0458_ ),
    .B(\Inst_RegFile_32x4/_0571_ ),
    .Y(\Inst_RegFile_32x4/_0586_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1209_  (.A0(\Inst_RegFile_32x4/_0577_ ),
    .A1(\Inst_RegFile_32x4/mem[25][0] ),
    .S(\Inst_RegFile_32x4/_0586_ ),
    .X(\Inst_RegFile_32x4/_0587_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1210_  (.A(\Inst_RegFile_32x4/_0587_ ),
    .X(\Inst_RegFile_32x4/_0072_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1211_  (.A0(\Inst_RegFile_32x4/_0580_ ),
    .A1(\Inst_RegFile_32x4/mem[25][1] ),
    .S(\Inst_RegFile_32x4/_0586_ ),
    .X(\Inst_RegFile_32x4/_0588_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1212_  (.A(\Inst_RegFile_32x4/_0588_ ),
    .X(\Inst_RegFile_32x4/_0073_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1213_  (.A0(\Inst_RegFile_32x4/_0582_ ),
    .A1(\Inst_RegFile_32x4/mem[25][2] ),
    .S(\Inst_RegFile_32x4/_0586_ ),
    .X(\Inst_RegFile_32x4/_0589_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1214_  (.A(\Inst_RegFile_32x4/_0589_ ),
    .X(\Inst_RegFile_32x4/_0074_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1215_  (.A0(\Inst_RegFile_32x4/_0584_ ),
    .A1(\Inst_RegFile_32x4/mem[25][3] ),
    .S(\Inst_RegFile_32x4/_0586_ ),
    .X(\Inst_RegFile_32x4/_0590_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1216_  (.A(\Inst_RegFile_32x4/_0590_ ),
    .X(\Inst_RegFile_32x4/_0075_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1217_  (.A(D0),
    .X(\Inst_RegFile_32x4/_0591_ ));
 sky130_fd_sc_hd__and2_1 \Inst_RegFile_32x4/_1218_  (.A(\Inst_RegFile_32x4/_0474_ ),
    .B(\Inst_RegFile_32x4/_0571_ ),
    .X(\Inst_RegFile_32x4/_0592_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1219_  (.A0(\Inst_RegFile_32x4/mem[24][0] ),
    .A1(\Inst_RegFile_32x4/_0591_ ),
    .S(\Inst_RegFile_32x4/_0592_ ),
    .X(\Inst_RegFile_32x4/_0593_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1220_  (.A(\Inst_RegFile_32x4/_0593_ ),
    .X(\Inst_RegFile_32x4/_0076_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1221_  (.A(D1),
    .X(\Inst_RegFile_32x4/_0594_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1222_  (.A0(\Inst_RegFile_32x4/mem[24][1] ),
    .A1(\Inst_RegFile_32x4/_0594_ ),
    .S(\Inst_RegFile_32x4/_0592_ ),
    .X(\Inst_RegFile_32x4/_0595_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1223_  (.A(\Inst_RegFile_32x4/_0595_ ),
    .X(\Inst_RegFile_32x4/_0077_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1224_  (.A(D2),
    .X(\Inst_RegFile_32x4/_0596_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1225_  (.A0(\Inst_RegFile_32x4/mem[24][2] ),
    .A1(\Inst_RegFile_32x4/_0596_ ),
    .S(\Inst_RegFile_32x4/_0592_ ),
    .X(\Inst_RegFile_32x4/_0597_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1226_  (.A(\Inst_RegFile_32x4/_0597_ ),
    .X(\Inst_RegFile_32x4/_0078_ ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_32x4/_1227_  (.A(D3),
    .X(\Inst_RegFile_32x4/_0598_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1228_  (.A0(\Inst_RegFile_32x4/mem[24][3] ),
    .A1(\Inst_RegFile_32x4/_0598_ ),
    .S(\Inst_RegFile_32x4/_0592_ ),
    .X(\Inst_RegFile_32x4/_0599_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1229_  (.A(\Inst_RegFile_32x4/_0599_ ),
    .X(\Inst_RegFile_32x4/_0079_ ));
 sky130_fd_sc_hd__and3b_2 \Inst_RegFile_32x4/_1230_  (.A_N(W_ADR3),
    .B(W_ADR2),
    .C(W_ADR4),
    .X(\Inst_RegFile_32x4/_0600_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1231_  (.A(\Inst_RegFile_32x4/_0570_ ),
    .B(\Inst_RegFile_32x4/_0600_ ),
    .Y(\Inst_RegFile_32x4/_0601_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1232_  (.A0(\Inst_RegFile_32x4/_0577_ ),
    .A1(\Inst_RegFile_32x4/mem[23][0] ),
    .S(\Inst_RegFile_32x4/_0601_ ),
    .X(\Inst_RegFile_32x4/_0602_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1233_  (.A(\Inst_RegFile_32x4/_0602_ ),
    .X(\Inst_RegFile_32x4/_0080_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1234_  (.A0(\Inst_RegFile_32x4/_0580_ ),
    .A1(\Inst_RegFile_32x4/mem[23][1] ),
    .S(\Inst_RegFile_32x4/_0601_ ),
    .X(\Inst_RegFile_32x4/_0603_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1235_  (.A(\Inst_RegFile_32x4/_0603_ ),
    .X(\Inst_RegFile_32x4/_0081_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1236_  (.A0(\Inst_RegFile_32x4/_0582_ ),
    .A1(\Inst_RegFile_32x4/mem[23][2] ),
    .S(\Inst_RegFile_32x4/_0601_ ),
    .X(\Inst_RegFile_32x4/_0604_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1237_  (.A(\Inst_RegFile_32x4/_0604_ ),
    .X(\Inst_RegFile_32x4/_0082_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1238_  (.A0(\Inst_RegFile_32x4/_0584_ ),
    .A1(\Inst_RegFile_32x4/mem[23][3] ),
    .S(\Inst_RegFile_32x4/_0601_ ),
    .X(\Inst_RegFile_32x4/_0605_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1239_  (.A(\Inst_RegFile_32x4/_0605_ ),
    .X(\Inst_RegFile_32x4/_0083_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1240_  (.A(\Inst_RegFile_32x4/_0554_ ),
    .B(\Inst_RegFile_32x4/_0600_ ),
    .Y(\Inst_RegFile_32x4/_0606_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1241_  (.A0(\Inst_RegFile_32x4/_0577_ ),
    .A1(\Inst_RegFile_32x4/mem[22][0] ),
    .S(\Inst_RegFile_32x4/_0606_ ),
    .X(\Inst_RegFile_32x4/_0607_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1242_  (.A(\Inst_RegFile_32x4/_0607_ ),
    .X(\Inst_RegFile_32x4/_0084_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1243_  (.A0(\Inst_RegFile_32x4/_0580_ ),
    .A1(\Inst_RegFile_32x4/mem[22][1] ),
    .S(\Inst_RegFile_32x4/_0606_ ),
    .X(\Inst_RegFile_32x4/_0608_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1244_  (.A(\Inst_RegFile_32x4/_0608_ ),
    .X(\Inst_RegFile_32x4/_0085_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1245_  (.A0(\Inst_RegFile_32x4/_0582_ ),
    .A1(\Inst_RegFile_32x4/mem[22][2] ),
    .S(\Inst_RegFile_32x4/_0606_ ),
    .X(\Inst_RegFile_32x4/_0609_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1246_  (.A(\Inst_RegFile_32x4/_0609_ ),
    .X(\Inst_RegFile_32x4/_0086_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1247_  (.A0(\Inst_RegFile_32x4/_0584_ ),
    .A1(\Inst_RegFile_32x4/mem[22][3] ),
    .S(\Inst_RegFile_32x4/_0606_ ),
    .X(\Inst_RegFile_32x4/_0610_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1248_  (.A(\Inst_RegFile_32x4/_0610_ ),
    .X(\Inst_RegFile_32x4/_0087_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1249_  (.A(\Inst_RegFile_32x4/_0458_ ),
    .B(\Inst_RegFile_32x4/_0600_ ),
    .Y(\Inst_RegFile_32x4/_0611_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1250_  (.A0(\Inst_RegFile_32x4/_0577_ ),
    .A1(\Inst_RegFile_32x4/mem[21][0] ),
    .S(\Inst_RegFile_32x4/_0611_ ),
    .X(\Inst_RegFile_32x4/_0612_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1251_  (.A(\Inst_RegFile_32x4/_0612_ ),
    .X(\Inst_RegFile_32x4/_0088_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1252_  (.A0(\Inst_RegFile_32x4/_0580_ ),
    .A1(\Inst_RegFile_32x4/mem[21][1] ),
    .S(\Inst_RegFile_32x4/_0611_ ),
    .X(\Inst_RegFile_32x4/_0613_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1253_  (.A(\Inst_RegFile_32x4/_0613_ ),
    .X(\Inst_RegFile_32x4/_0089_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1254_  (.A0(\Inst_RegFile_32x4/_0582_ ),
    .A1(\Inst_RegFile_32x4/mem[21][2] ),
    .S(\Inst_RegFile_32x4/_0611_ ),
    .X(\Inst_RegFile_32x4/_0614_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1255_  (.A(\Inst_RegFile_32x4/_0614_ ),
    .X(\Inst_RegFile_32x4/_0090_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1256_  (.A0(\Inst_RegFile_32x4/_0584_ ),
    .A1(\Inst_RegFile_32x4/mem[21][3] ),
    .S(\Inst_RegFile_32x4/_0611_ ),
    .X(\Inst_RegFile_32x4/_0615_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1257_  (.A(\Inst_RegFile_32x4/_0615_ ),
    .X(\Inst_RegFile_32x4/_0091_ ));
 sky130_fd_sc_hd__and2_2 \Inst_RegFile_32x4/_1258_  (.A(\Inst_RegFile_32x4/_0474_ ),
    .B(\Inst_RegFile_32x4/_0600_ ),
    .X(\Inst_RegFile_32x4/_0616_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1259_  (.A0(\Inst_RegFile_32x4/mem[20][0] ),
    .A1(\Inst_RegFile_32x4/_0591_ ),
    .S(\Inst_RegFile_32x4/_0616_ ),
    .X(\Inst_RegFile_32x4/_0617_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1260_  (.A(\Inst_RegFile_32x4/_0617_ ),
    .X(\Inst_RegFile_32x4/_0092_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1261_  (.A0(\Inst_RegFile_32x4/mem[20][1] ),
    .A1(\Inst_RegFile_32x4/_0594_ ),
    .S(\Inst_RegFile_32x4/_0616_ ),
    .X(\Inst_RegFile_32x4/_0618_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1262_  (.A(\Inst_RegFile_32x4/_0618_ ),
    .X(\Inst_RegFile_32x4/_0093_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1263_  (.A0(\Inst_RegFile_32x4/mem[20][2] ),
    .A1(\Inst_RegFile_32x4/_0596_ ),
    .S(\Inst_RegFile_32x4/_0616_ ),
    .X(\Inst_RegFile_32x4/_0619_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1264_  (.A(\Inst_RegFile_32x4/_0619_ ),
    .X(\Inst_RegFile_32x4/_0094_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1265_  (.A0(\Inst_RegFile_32x4/mem[20][3] ),
    .A1(\Inst_RegFile_32x4/_0598_ ),
    .S(\Inst_RegFile_32x4/_0616_ ),
    .X(\Inst_RegFile_32x4/_0620_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1266_  (.A(\Inst_RegFile_32x4/_0620_ ),
    .X(\Inst_RegFile_32x4/_0095_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1267_  (.A(\Inst_RegFile_32x4/_0525_ ),
    .B(\Inst_RegFile_32x4/_0502_ ),
    .Y(\Inst_RegFile_32x4/_0621_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1268_  (.A0(\Inst_RegFile_32x4/mem[1][0] ),
    .A1(\Inst_RegFile_32x4/_0591_ ),
    .S(\Inst_RegFile_32x4/_0621_ ),
    .X(\Inst_RegFile_32x4/_0622_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1269_  (.A(\Inst_RegFile_32x4/_0622_ ),
    .X(\Inst_RegFile_32x4/_0096_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1270_  (.A0(\Inst_RegFile_32x4/mem[1][1] ),
    .A1(\Inst_RegFile_32x4/_0594_ ),
    .S(\Inst_RegFile_32x4/_0621_ ),
    .X(\Inst_RegFile_32x4/_0623_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1271_  (.A(\Inst_RegFile_32x4/_0623_ ),
    .X(\Inst_RegFile_32x4/_0097_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1272_  (.A0(\Inst_RegFile_32x4/mem[1][2] ),
    .A1(\Inst_RegFile_32x4/_0596_ ),
    .S(\Inst_RegFile_32x4/_0621_ ),
    .X(\Inst_RegFile_32x4/_0624_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1273_  (.A(\Inst_RegFile_32x4/_0624_ ),
    .X(\Inst_RegFile_32x4/_0098_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1274_  (.A0(\Inst_RegFile_32x4/mem[1][3] ),
    .A1(\Inst_RegFile_32x4/_0598_ ),
    .S(\Inst_RegFile_32x4/_0621_ ),
    .X(\Inst_RegFile_32x4/_0625_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1275_  (.A(\Inst_RegFile_32x4/_0625_ ),
    .X(\Inst_RegFile_32x4/_0099_ ));
 sky130_fd_sc_hd__or3b_4 \Inst_RegFile_32x4/_1276_  (.A(\Inst_RegFile_32x4/_0453_ ),
    .B(\Inst_RegFile_32x4/_0454_ ),
    .C_N(\Inst_RegFile_32x4/_0452_ ),
    .X(\Inst_RegFile_32x4/_0626_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1277_  (.A(\Inst_RegFile_32x4/_0493_ ),
    .B(\Inst_RegFile_32x4/_0626_ ),
    .Y(\Inst_RegFile_32x4/_0627_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1278_  (.A0(\Inst_RegFile_32x4/mem[18][0] ),
    .A1(\Inst_RegFile_32x4/_0591_ ),
    .S(\Inst_RegFile_32x4/_0627_ ),
    .X(\Inst_RegFile_32x4/_0628_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1279_  (.A(\Inst_RegFile_32x4/_0628_ ),
    .X(\Inst_RegFile_32x4/_0100_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1280_  (.A0(\Inst_RegFile_32x4/mem[18][1] ),
    .A1(\Inst_RegFile_32x4/_0594_ ),
    .S(\Inst_RegFile_32x4/_0627_ ),
    .X(\Inst_RegFile_32x4/_0629_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1281_  (.A(\Inst_RegFile_32x4/_0629_ ),
    .X(\Inst_RegFile_32x4/_0101_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1282_  (.A0(\Inst_RegFile_32x4/mem[18][2] ),
    .A1(\Inst_RegFile_32x4/_0596_ ),
    .S(\Inst_RegFile_32x4/_0627_ ),
    .X(\Inst_RegFile_32x4/_0630_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1283_  (.A(\Inst_RegFile_32x4/_0630_ ),
    .X(\Inst_RegFile_32x4/_0102_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1284_  (.A0(\Inst_RegFile_32x4/mem[18][3] ),
    .A1(\Inst_RegFile_32x4/_0598_ ),
    .S(\Inst_RegFile_32x4/_0627_ ),
    .X(\Inst_RegFile_32x4/_0631_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1285_  (.A(\Inst_RegFile_32x4/_0631_ ),
    .X(\Inst_RegFile_32x4/_0103_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1286_  (.A(\Inst_RegFile_32x4/_0525_ ),
    .B(\Inst_RegFile_32x4/_0626_ ),
    .Y(\Inst_RegFile_32x4/_0632_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1287_  (.A0(\Inst_RegFile_32x4/mem[17][0] ),
    .A1(\Inst_RegFile_32x4/_0591_ ),
    .S(\Inst_RegFile_32x4/_0632_ ),
    .X(\Inst_RegFile_32x4/_0633_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1288_  (.A(\Inst_RegFile_32x4/_0633_ ),
    .X(\Inst_RegFile_32x4/_0104_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1289_  (.A0(\Inst_RegFile_32x4/mem[17][1] ),
    .A1(\Inst_RegFile_32x4/_0594_ ),
    .S(\Inst_RegFile_32x4/_0632_ ),
    .X(\Inst_RegFile_32x4/_0634_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1290_  (.A(\Inst_RegFile_32x4/_0634_ ),
    .X(\Inst_RegFile_32x4/_0105_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1291_  (.A0(\Inst_RegFile_32x4/mem[17][2] ),
    .A1(\Inst_RegFile_32x4/_0596_ ),
    .S(\Inst_RegFile_32x4/_0632_ ),
    .X(\Inst_RegFile_32x4/_0635_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1292_  (.A(\Inst_RegFile_32x4/_0635_ ),
    .X(\Inst_RegFile_32x4/_0106_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1293_  (.A0(\Inst_RegFile_32x4/mem[17][3] ),
    .A1(\Inst_RegFile_32x4/_0598_ ),
    .S(\Inst_RegFile_32x4/_0632_ ),
    .X(\Inst_RegFile_32x4/_0636_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1294_  (.A(\Inst_RegFile_32x4/_0636_ ),
    .X(\Inst_RegFile_32x4/_0107_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1295_  (.A(\Inst_RegFile_32x4/_0473_ ),
    .B(\Inst_RegFile_32x4/_0626_ ),
    .Y(\Inst_RegFile_32x4/_0637_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1296_  (.A0(\Inst_RegFile_32x4/mem[16][0] ),
    .A1(\Inst_RegFile_32x4/_0450_ ),
    .S(\Inst_RegFile_32x4/_0637_ ),
    .X(\Inst_RegFile_32x4/_0638_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1297_  (.A(\Inst_RegFile_32x4/_0638_ ),
    .X(\Inst_RegFile_32x4/_0108_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1298_  (.A0(\Inst_RegFile_32x4/mem[16][1] ),
    .A1(\Inst_RegFile_32x4/_0461_ ),
    .S(\Inst_RegFile_32x4/_0637_ ),
    .X(\Inst_RegFile_32x4/_0639_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1299_  (.A(\Inst_RegFile_32x4/_0639_ ),
    .X(\Inst_RegFile_32x4/_0109_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1300_  (.A0(\Inst_RegFile_32x4/mem[16][2] ),
    .A1(\Inst_RegFile_32x4/_0464_ ),
    .S(\Inst_RegFile_32x4/_0637_ ),
    .X(\Inst_RegFile_32x4/_0640_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1301_  (.A(\Inst_RegFile_32x4/_0640_ ),
    .X(\Inst_RegFile_32x4/_0110_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1302_  (.A0(\Inst_RegFile_32x4/mem[16][3] ),
    .A1(\Inst_RegFile_32x4/_0467_ ),
    .S(\Inst_RegFile_32x4/_0637_ ),
    .X(\Inst_RegFile_32x4/_0641_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1303_  (.A(\Inst_RegFile_32x4/_0641_ ),
    .X(\Inst_RegFile_32x4/_0111_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1304_  (.A(\Inst_RegFile_32x4/_0471_ ),
    .B(\Inst_RegFile_32x4/_0570_ ),
    .Y(\Inst_RegFile_32x4/_0642_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1305_  (.A0(\Inst_RegFile_32x4/_0470_ ),
    .A1(\Inst_RegFile_32x4/mem[15][0] ),
    .S(\Inst_RegFile_32x4/_0642_ ),
    .X(\Inst_RegFile_32x4/_0643_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1306_  (.A(\Inst_RegFile_32x4/_0643_ ),
    .X(\Inst_RegFile_32x4/_0112_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1307_  (.A0(\Inst_RegFile_32x4/_0477_ ),
    .A1(\Inst_RegFile_32x4/mem[15][1] ),
    .S(\Inst_RegFile_32x4/_0642_ ),
    .X(\Inst_RegFile_32x4/_0644_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1308_  (.A(\Inst_RegFile_32x4/_0644_ ),
    .X(\Inst_RegFile_32x4/_0113_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1309_  (.A0(\Inst_RegFile_32x4/_0479_ ),
    .A1(\Inst_RegFile_32x4/mem[15][2] ),
    .S(\Inst_RegFile_32x4/_0642_ ),
    .X(\Inst_RegFile_32x4/_0645_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1310_  (.A(\Inst_RegFile_32x4/_0645_ ),
    .X(\Inst_RegFile_32x4/_0114_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1311_  (.A0(\Inst_RegFile_32x4/_0481_ ),
    .A1(\Inst_RegFile_32x4/mem[15][3] ),
    .S(\Inst_RegFile_32x4/_0642_ ),
    .X(\Inst_RegFile_32x4/_0646_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1312_  (.A(\Inst_RegFile_32x4/_0646_ ),
    .X(\Inst_RegFile_32x4/_0115_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1313_  (.A(\Inst_RegFile_32x4/_0471_ ),
    .B(\Inst_RegFile_32x4/_0554_ ),
    .Y(\Inst_RegFile_32x4/_0647_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1314_  (.A0(\Inst_RegFile_32x4/_0470_ ),
    .A1(\Inst_RegFile_32x4/mem[14][0] ),
    .S(\Inst_RegFile_32x4/_0647_ ),
    .X(\Inst_RegFile_32x4/_0648_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1315_  (.A(\Inst_RegFile_32x4/_0648_ ),
    .X(\Inst_RegFile_32x4/_0116_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1316_  (.A0(\Inst_RegFile_32x4/_0477_ ),
    .A1(\Inst_RegFile_32x4/mem[14][1] ),
    .S(\Inst_RegFile_32x4/_0647_ ),
    .X(\Inst_RegFile_32x4/_0649_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1317_  (.A(\Inst_RegFile_32x4/_0649_ ),
    .X(\Inst_RegFile_32x4/_0117_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1318_  (.A0(\Inst_RegFile_32x4/_0479_ ),
    .A1(\Inst_RegFile_32x4/mem[14][2] ),
    .S(\Inst_RegFile_32x4/_0647_ ),
    .X(\Inst_RegFile_32x4/_0650_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1319_  (.A(\Inst_RegFile_32x4/_0650_ ),
    .X(\Inst_RegFile_32x4/_0118_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1320_  (.A0(\Inst_RegFile_32x4/_0481_ ),
    .A1(\Inst_RegFile_32x4/mem[14][3] ),
    .S(\Inst_RegFile_32x4/_0647_ ),
    .X(\Inst_RegFile_32x4/_0651_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1321_  (.A(\Inst_RegFile_32x4/_0651_ ),
    .X(\Inst_RegFile_32x4/_0119_ ));
 sky130_fd_sc_hd__nand2_2 \Inst_RegFile_32x4/_1322_  (.A(\Inst_RegFile_32x4/_0455_ ),
    .B(\Inst_RegFile_32x4/_0570_ ),
    .Y(\Inst_RegFile_32x4/_0652_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1323_  (.A0(\Inst_RegFile_32x4/_0470_ ),
    .A1(\Inst_RegFile_32x4/mem[31][0] ),
    .S(\Inst_RegFile_32x4/_0652_ ),
    .X(\Inst_RegFile_32x4/_0653_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1324_  (.A(\Inst_RegFile_32x4/_0653_ ),
    .X(\Inst_RegFile_32x4/_0120_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1325_  (.A0(\Inst_RegFile_32x4/_0477_ ),
    .A1(\Inst_RegFile_32x4/mem[31][1] ),
    .S(\Inst_RegFile_32x4/_0652_ ),
    .X(\Inst_RegFile_32x4/_0654_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1326_  (.A(\Inst_RegFile_32x4/_0654_ ),
    .X(\Inst_RegFile_32x4/_0121_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1327_  (.A0(\Inst_RegFile_32x4/_0479_ ),
    .A1(\Inst_RegFile_32x4/mem[31][2] ),
    .S(\Inst_RegFile_32x4/_0652_ ),
    .X(\Inst_RegFile_32x4/_0655_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1328_  (.A(\Inst_RegFile_32x4/_0655_ ),
    .X(\Inst_RegFile_32x4/_0122_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1329_  (.A0(\Inst_RegFile_32x4/_0481_ ),
    .A1(\Inst_RegFile_32x4/mem[31][3] ),
    .S(\Inst_RegFile_32x4/_0652_ ),
    .X(\Inst_RegFile_32x4/_0656_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1330_  (.A(\Inst_RegFile_32x4/_0656_ ),
    .X(\Inst_RegFile_32x4/_0123_ ));
 sky130_fd_sc_hd__nor2_2 \Inst_RegFile_32x4/_1331_  (.A(\Inst_RegFile_32x4/_0485_ ),
    .B(\Inst_RegFile_32x4/_0626_ ),
    .Y(\Inst_RegFile_32x4/_0657_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1332_  (.A0(\Inst_RegFile_32x4/mem[19][0] ),
    .A1(\Inst_RegFile_32x4/_0450_ ),
    .S(\Inst_RegFile_32x4/_0657_ ),
    .X(\Inst_RegFile_32x4/_0658_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1333_  (.A(\Inst_RegFile_32x4/_0658_ ),
    .X(\Inst_RegFile_32x4/_0124_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1334_  (.A0(\Inst_RegFile_32x4/mem[19][1] ),
    .A1(\Inst_RegFile_32x4/_0461_ ),
    .S(\Inst_RegFile_32x4/_0657_ ),
    .X(\Inst_RegFile_32x4/_0659_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1335_  (.A(\Inst_RegFile_32x4/_0659_ ),
    .X(\Inst_RegFile_32x4/_0125_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1336_  (.A0(\Inst_RegFile_32x4/mem[19][2] ),
    .A1(\Inst_RegFile_32x4/_0464_ ),
    .S(\Inst_RegFile_32x4/_0657_ ),
    .X(\Inst_RegFile_32x4/_0660_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1337_  (.A(\Inst_RegFile_32x4/_0660_ ),
    .X(\Inst_RegFile_32x4/_0126_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_32x4/_1338_  (.A0(\Inst_RegFile_32x4/mem[19][3] ),
    .A1(\Inst_RegFile_32x4/_0467_ ),
    .S(\Inst_RegFile_32x4/_0657_ ),
    .X(\Inst_RegFile_32x4/_0661_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_32x4/_1339_  (.A(\Inst_RegFile_32x4/_0661_ ),
    .X(\Inst_RegFile_32x4/_0127_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1340_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0000_ ),
    .Q(\Inst_RegFile_32x4/mem[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1341_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0001_ ),
    .Q(\Inst_RegFile_32x4/mem[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1342_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0002_ ),
    .Q(\Inst_RegFile_32x4/mem[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1343_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0003_ ),
    .Q(\Inst_RegFile_32x4/mem[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1344_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0004_ ),
    .Q(\Inst_RegFile_32x4/mem[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1345_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0005_ ),
    .Q(\Inst_RegFile_32x4/mem[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1346_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0006_ ),
    .Q(\Inst_RegFile_32x4/mem[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1347_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0007_ ),
    .Q(\Inst_RegFile_32x4/mem[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1348_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0008_ ),
    .Q(\Inst_RegFile_32x4/mem[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1349_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0009_ ),
    .Q(\Inst_RegFile_32x4/mem[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1350_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0010_ ),
    .Q(\Inst_RegFile_32x4/mem[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1351_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0011_ ),
    .Q(\Inst_RegFile_32x4/mem[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1352_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0012_ ),
    .Q(\Inst_RegFile_32x4/mem[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1353_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0013_ ),
    .Q(\Inst_RegFile_32x4/mem[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1354_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0014_ ),
    .Q(\Inst_RegFile_32x4/mem[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1355_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0015_ ),
    .Q(\Inst_RegFile_32x4/mem[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1356_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0016_ ),
    .Q(\Inst_RegFile_32x4/mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1357_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0017_ ),
    .Q(\Inst_RegFile_32x4/mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1358_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0018_ ),
    .Q(\Inst_RegFile_32x4/mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1359_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0019_ ),
    .Q(\Inst_RegFile_32x4/mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1360_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0020_ ),
    .Q(\Inst_RegFile_32x4/mem[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1361_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0021_ ),
    .Q(\Inst_RegFile_32x4/mem[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1362_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0022_ ),
    .Q(\Inst_RegFile_32x4/mem[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1363_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0023_ ),
    .Q(\Inst_RegFile_32x4/mem[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1364_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0024_ ),
    .Q(\Inst_RegFile_32x4/mem[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1365_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0025_ ),
    .Q(\Inst_RegFile_32x4/mem[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1366_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0026_ ),
    .Q(\Inst_RegFile_32x4/mem[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1367_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0027_ ),
    .Q(\Inst_RegFile_32x4/mem[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1368_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0028_ ),
    .Q(\Inst_RegFile_32x4/mem[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1369_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0029_ ),
    .Q(\Inst_RegFile_32x4/mem[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1370_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0030_ ),
    .Q(\Inst_RegFile_32x4/mem[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1371_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0031_ ),
    .Q(\Inst_RegFile_32x4/mem[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1372_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0032_ ),
    .Q(\Inst_RegFile_32x4/mem[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1373_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0033_ ),
    .Q(\Inst_RegFile_32x4/mem[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1374_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0034_ ),
    .Q(\Inst_RegFile_32x4/mem[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1375_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0035_ ),
    .Q(\Inst_RegFile_32x4/mem[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1376_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0036_ ),
    .Q(\Inst_RegFile_32x4/mem[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1377_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0037_ ),
    .Q(\Inst_RegFile_32x4/mem[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1378_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0038_ ),
    .Q(\Inst_RegFile_32x4/mem[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1379_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0039_ ),
    .Q(\Inst_RegFile_32x4/mem[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1380_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0040_ ),
    .Q(\Inst_RegFile_32x4/mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1381_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0041_ ),
    .Q(\Inst_RegFile_32x4/mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1382_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0042_ ),
    .Q(\Inst_RegFile_32x4/mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1383_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0043_ ),
    .Q(\Inst_RegFile_32x4/mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1384_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/AD_comb[0] ),
    .Q(\Inst_RegFile_32x4/AD_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1385_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/AD_comb[1] ),
    .Q(\Inst_RegFile_32x4/AD_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1386_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/AD_comb[2] ),
    .Q(\Inst_RegFile_32x4/AD_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1387_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/AD_comb[3] ),
    .Q(\Inst_RegFile_32x4/AD_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1388_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/BD_comb[0] ),
    .Q(\Inst_RegFile_32x4/BD_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1389_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/BD_comb[1] ),
    .Q(\Inst_RegFile_32x4/BD_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1390_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/BD_comb[2] ),
    .Q(\Inst_RegFile_32x4/BD_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1391_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/BD_comb[3] ),
    .Q(\Inst_RegFile_32x4/BD_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1392_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0044_ ),
    .Q(\Inst_RegFile_32x4/mem[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1393_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0045_ ),
    .Q(\Inst_RegFile_32x4/mem[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1394_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0046_ ),
    .Q(\Inst_RegFile_32x4/mem[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1395_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0047_ ),
    .Q(\Inst_RegFile_32x4/mem[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1396_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0048_ ),
    .Q(\Inst_RegFile_32x4/mem[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1397_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0049_ ),
    .Q(\Inst_RegFile_32x4/mem[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1398_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0050_ ),
    .Q(\Inst_RegFile_32x4/mem[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1399_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0051_ ),
    .Q(\Inst_RegFile_32x4/mem[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1400_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0052_ ),
    .Q(\Inst_RegFile_32x4/mem[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1401_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0053_ ),
    .Q(\Inst_RegFile_32x4/mem[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1402_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0054_ ),
    .Q(\Inst_RegFile_32x4/mem[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1403_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0055_ ),
    .Q(\Inst_RegFile_32x4/mem[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1404_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0056_ ),
    .Q(\Inst_RegFile_32x4/mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1405_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0057_ ),
    .Q(\Inst_RegFile_32x4/mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1406_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0058_ ),
    .Q(\Inst_RegFile_32x4/mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1407_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0059_ ),
    .Q(\Inst_RegFile_32x4/mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1408_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0060_ ),
    .Q(\Inst_RegFile_32x4/mem[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1409_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0061_ ),
    .Q(\Inst_RegFile_32x4/mem[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1410_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0062_ ),
    .Q(\Inst_RegFile_32x4/mem[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1411_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0063_ ),
    .Q(\Inst_RegFile_32x4/mem[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1412_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0064_ ),
    .Q(\Inst_RegFile_32x4/mem[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1413_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0065_ ),
    .Q(\Inst_RegFile_32x4/mem[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1414_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0066_ ),
    .Q(\Inst_RegFile_32x4/mem[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1415_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0067_ ),
    .Q(\Inst_RegFile_32x4/mem[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1416_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0068_ ),
    .Q(\Inst_RegFile_32x4/mem[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1417_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0069_ ),
    .Q(\Inst_RegFile_32x4/mem[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1418_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0070_ ),
    .Q(\Inst_RegFile_32x4/mem[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1419_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0071_ ),
    .Q(\Inst_RegFile_32x4/mem[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1420_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0072_ ),
    .Q(\Inst_RegFile_32x4/mem[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1421_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0073_ ),
    .Q(\Inst_RegFile_32x4/mem[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1422_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0074_ ),
    .Q(\Inst_RegFile_32x4/mem[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1423_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0075_ ),
    .Q(\Inst_RegFile_32x4/mem[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1424_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0076_ ),
    .Q(\Inst_RegFile_32x4/mem[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1425_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0077_ ),
    .Q(\Inst_RegFile_32x4/mem[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1426_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0078_ ),
    .Q(\Inst_RegFile_32x4/mem[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1427_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0079_ ),
    .Q(\Inst_RegFile_32x4/mem[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1428_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0080_ ),
    .Q(\Inst_RegFile_32x4/mem[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1429_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0081_ ),
    .Q(\Inst_RegFile_32x4/mem[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1430_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0082_ ),
    .Q(\Inst_RegFile_32x4/mem[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1431_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0083_ ),
    .Q(\Inst_RegFile_32x4/mem[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1432_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0084_ ),
    .Q(\Inst_RegFile_32x4/mem[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1433_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0085_ ),
    .Q(\Inst_RegFile_32x4/mem[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1434_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0086_ ),
    .Q(\Inst_RegFile_32x4/mem[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1435_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0087_ ),
    .Q(\Inst_RegFile_32x4/mem[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1436_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0088_ ),
    .Q(\Inst_RegFile_32x4/mem[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1437_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0089_ ),
    .Q(\Inst_RegFile_32x4/mem[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1438_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0090_ ),
    .Q(\Inst_RegFile_32x4/mem[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1439_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0091_ ),
    .Q(\Inst_RegFile_32x4/mem[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1440_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0092_ ),
    .Q(\Inst_RegFile_32x4/mem[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1441_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0093_ ),
    .Q(\Inst_RegFile_32x4/mem[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1442_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0094_ ),
    .Q(\Inst_RegFile_32x4/mem[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1443_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0095_ ),
    .Q(\Inst_RegFile_32x4/mem[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1444_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0096_ ),
    .Q(\Inst_RegFile_32x4/mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1445_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0097_ ),
    .Q(\Inst_RegFile_32x4/mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1446_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0098_ ),
    .Q(\Inst_RegFile_32x4/mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1447_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0099_ ),
    .Q(\Inst_RegFile_32x4/mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1448_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0100_ ),
    .Q(\Inst_RegFile_32x4/mem[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1449_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0101_ ),
    .Q(\Inst_RegFile_32x4/mem[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1450_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0102_ ),
    .Q(\Inst_RegFile_32x4/mem[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1451_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0103_ ),
    .Q(\Inst_RegFile_32x4/mem[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1452_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0104_ ),
    .Q(\Inst_RegFile_32x4/mem[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1453_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0105_ ),
    .Q(\Inst_RegFile_32x4/mem[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1454_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0106_ ),
    .Q(\Inst_RegFile_32x4/mem[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1455_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0107_ ),
    .Q(\Inst_RegFile_32x4/mem[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1456_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0108_ ),
    .Q(\Inst_RegFile_32x4/mem[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1457_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0109_ ),
    .Q(\Inst_RegFile_32x4/mem[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1458_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0110_ ),
    .Q(\Inst_RegFile_32x4/mem[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1459_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0111_ ),
    .Q(\Inst_RegFile_32x4/mem[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1460_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0112_ ),
    .Q(\Inst_RegFile_32x4/mem[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1461_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0113_ ),
    .Q(\Inst_RegFile_32x4/mem[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1462_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0114_ ),
    .Q(\Inst_RegFile_32x4/mem[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1463_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0115_ ),
    .Q(\Inst_RegFile_32x4/mem[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1464_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0116_ ),
    .Q(\Inst_RegFile_32x4/mem[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1465_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0117_ ),
    .Q(\Inst_RegFile_32x4/mem[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1466_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0118_ ),
    .Q(\Inst_RegFile_32x4/mem[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1467_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0119_ ),
    .Q(\Inst_RegFile_32x4/mem[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1468_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0120_ ),
    .Q(\Inst_RegFile_32x4/mem[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1469_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0121_ ),
    .Q(\Inst_RegFile_32x4/mem[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1470_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0122_ ),
    .Q(\Inst_RegFile_32x4/mem[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1471_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0123_ ),
    .Q(\Inst_RegFile_32x4/mem[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1472_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0124_ ),
    .Q(\Inst_RegFile_32x4/mem[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1473_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0125_ ),
    .Q(\Inst_RegFile_32x4/mem[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1474_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0126_ ),
    .Q(\Inst_RegFile_32x4/mem[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RegFile_32x4/_1475_  (.CLK(net205),
    .D(\Inst_RegFile_32x4/_0127_ ),
    .Q(\Inst_RegFile_32x4/mem[19][3] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit0  (.D(net49),
    .GATE(net81),
    .Q(\ConfigBits[382] ),
    .Q_N(\ConfigBits_N[382] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit1  (.D(net60),
    .GATE(net81),
    .Q(\ConfigBits[383] ),
    .Q_N(\ConfigBits_N[383] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit10  (.D(net50),
    .GATE(net81),
    .Q(\ConfigBits[392] ),
    .Q_N(\ConfigBits_N[392] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit11  (.D(net51),
    .GATE(net81),
    .Q(\ConfigBits[393] ),
    .Q_N(\ConfigBits_N[393] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit12  (.D(net52),
    .GATE(net81),
    .Q(\ConfigBits[394] ),
    .Q_N(\ConfigBits_N[394] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit13  (.D(net53),
    .GATE(net81),
    .Q(\ConfigBits[395] ),
    .Q_N(\ConfigBits_N[395] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit14  (.D(net54),
    .GATE(net81),
    .Q(\ConfigBits[396] ),
    .Q_N(\ConfigBits_N[396] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit15  (.D(net55),
    .GATE(net81),
    .Q(\ConfigBits[397] ),
    .Q_N(\ConfigBits_N[397] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit16  (.D(net56),
    .GATE(net81),
    .Q(\ConfigBits[398] ),
    .Q_N(\ConfigBits_N[398] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit17  (.D(net57),
    .GATE(net81),
    .Q(\ConfigBits[399] ),
    .Q_N(\ConfigBits_N[399] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit18  (.D(net58),
    .GATE(net81),
    .Q(\ConfigBits[400] ),
    .Q_N(\ConfigBits_N[400] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit19  (.D(net59),
    .GATE(net81),
    .Q(\ConfigBits[401] ),
    .Q_N(\ConfigBits_N[401] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit2  (.D(net71),
    .GATE(net81),
    .Q(\ConfigBits[384] ),
    .Q_N(\ConfigBits_N[384] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit20  (.D(net61),
    .GATE(net81),
    .Q(\ConfigBits[402] ),
    .Q_N(\ConfigBits_N[402] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit21  (.D(net62),
    .GATE(net81),
    .Q(\ConfigBits[403] ),
    .Q_N(\ConfigBits_N[403] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit22  (.D(net63),
    .GATE(net81),
    .Q(\ConfigBits[404] ),
    .Q_N(\ConfigBits_N[404] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit23  (.D(net64),
    .GATE(net81),
    .Q(\ConfigBits[405] ),
    .Q_N(\ConfigBits_N[405] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit24  (.D(net65),
    .GATE(net81),
    .Q(\ConfigBits[406] ),
    .Q_N(\ConfigBits_N[406] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit25  (.D(net66),
    .GATE(net81),
    .Q(\ConfigBits[407] ),
    .Q_N(\ConfigBits_N[407] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit26  (.D(net67),
    .GATE(net81),
    .Q(\ConfigBits[408] ),
    .Q_N(\ConfigBits_N[408] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit27  (.D(net68),
    .GATE(net81),
    .Q(\ConfigBits[409] ),
    .Q_N(\ConfigBits_N[409] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit28  (.D(net69),
    .GATE(net81),
    .Q(\ConfigBits[410] ),
    .Q_N(\ConfigBits_N[410] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit29  (.D(net70),
    .GATE(net81),
    .Q(\ConfigBits[411] ),
    .Q_N(\ConfigBits_N[411] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit3  (.D(net74),
    .GATE(net81),
    .Q(\ConfigBits[385] ),
    .Q_N(\ConfigBits_N[385] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit30  (.D(net72),
    .GATE(net81),
    .Q(\ConfigBits[412] ),
    .Q_N(\ConfigBits_N[412] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit31  (.D(net73),
    .GATE(net81),
    .Q(\ConfigBits[413] ),
    .Q_N(\ConfigBits_N[413] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit4  (.D(net75),
    .GATE(net81),
    .Q(\ConfigBits[386] ),
    .Q_N(\ConfigBits_N[386] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit5  (.D(net76),
    .GATE(net81),
    .Q(\ConfigBits[387] ),
    .Q_N(\ConfigBits_N[387] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit6  (.D(net77),
    .GATE(net81),
    .Q(\ConfigBits[388] ),
    .Q_N(\ConfigBits_N[388] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit7  (.D(net78),
    .GATE(net81),
    .Q(\ConfigBits[389] ),
    .Q_N(\ConfigBits_N[389] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit8  (.D(net79),
    .GATE(net81),
    .Q(\ConfigBits[390] ),
    .Q_N(\ConfigBits_N[390] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame0_bit9  (.D(net80),
    .GATE(net81),
    .Q(\ConfigBits[391] ),
    .Q_N(\ConfigBits_N[391] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit0  (.D(net49),
    .GATE(net82),
    .Q(\ConfigBits[62] ),
    .Q_N(\ConfigBits_N[62] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit1  (.D(net60),
    .GATE(net82),
    .Q(\ConfigBits[63] ),
    .Q_N(\ConfigBits_N[63] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit10  (.D(net50),
    .GATE(net82),
    .Q(\ConfigBits[72] ),
    .Q_N(\ConfigBits_N[72] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit11  (.D(net51),
    .GATE(net82),
    .Q(\ConfigBits[73] ),
    .Q_N(\ConfigBits_N[73] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit12  (.D(net52),
    .GATE(net82),
    .Q(\ConfigBits[74] ),
    .Q_N(\ConfigBits_N[74] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit13  (.D(net53),
    .GATE(net82),
    .Q(\ConfigBits[75] ),
    .Q_N(\ConfigBits_N[75] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit14  (.D(net54),
    .GATE(net82),
    .Q(\ConfigBits[76] ),
    .Q_N(\ConfigBits_N[76] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit15  (.D(net55),
    .GATE(net82),
    .Q(\ConfigBits[77] ),
    .Q_N(\ConfigBits_N[77] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit16  (.D(net56),
    .GATE(net82),
    .Q(\ConfigBits[78] ),
    .Q_N(\ConfigBits_N[78] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit17  (.D(net57),
    .GATE(net82),
    .Q(\ConfigBits[79] ),
    .Q_N(\ConfigBits_N[79] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit18  (.D(net58),
    .GATE(net82),
    .Q(\ConfigBits[80] ),
    .Q_N(\ConfigBits_N[80] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit19  (.D(net59),
    .GATE(net82),
    .Q(\ConfigBits[81] ),
    .Q_N(\ConfigBits_N[81] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit2  (.D(net71),
    .GATE(net82),
    .Q(\ConfigBits[64] ),
    .Q_N(\ConfigBits_N[64] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit20  (.D(net61),
    .GATE(net82),
    .Q(\ConfigBits[82] ),
    .Q_N(\ConfigBits_N[82] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit21  (.D(net62),
    .GATE(net82),
    .Q(\ConfigBits[83] ),
    .Q_N(\ConfigBits_N[83] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit22  (.D(net63),
    .GATE(net82),
    .Q(\ConfigBits[84] ),
    .Q_N(\ConfigBits_N[84] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit23  (.D(net64),
    .GATE(net82),
    .Q(\ConfigBits[85] ),
    .Q_N(\ConfigBits_N[85] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit24  (.D(net65),
    .GATE(net82),
    .Q(\ConfigBits[86] ),
    .Q_N(\ConfigBits_N[86] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit25  (.D(net66),
    .GATE(net82),
    .Q(\ConfigBits[87] ),
    .Q_N(\ConfigBits_N[87] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit26  (.D(net67),
    .GATE(net82),
    .Q(\ConfigBits[88] ),
    .Q_N(\ConfigBits_N[88] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit27  (.D(net68),
    .GATE(net82),
    .Q(\ConfigBits[89] ),
    .Q_N(\ConfigBits_N[89] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit28  (.D(net69),
    .GATE(net82),
    .Q(\ConfigBits[90] ),
    .Q_N(\ConfigBits_N[90] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit29  (.D(net70),
    .GATE(net82),
    .Q(\ConfigBits[91] ),
    .Q_N(\ConfigBits_N[91] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit3  (.D(net74),
    .GATE(net82),
    .Q(\ConfigBits[65] ),
    .Q_N(\ConfigBits_N[65] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit30  (.D(net72),
    .GATE(net82),
    .Q(\ConfigBits[92] ),
    .Q_N(\ConfigBits_N[92] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit31  (.D(net73),
    .GATE(net82),
    .Q(\ConfigBits[93] ),
    .Q_N(\ConfigBits_N[93] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit4  (.D(net75),
    .GATE(net82),
    .Q(\ConfigBits[66] ),
    .Q_N(\ConfigBits_N[66] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit5  (.D(net76),
    .GATE(net82),
    .Q(\ConfigBits[67] ),
    .Q_N(\ConfigBits_N[67] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit6  (.D(net77),
    .GATE(net82),
    .Q(\ConfigBits[68] ),
    .Q_N(\ConfigBits_N[68] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit7  (.D(net78),
    .GATE(net82),
    .Q(\ConfigBits[69] ),
    .Q_N(\ConfigBits_N[69] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit8  (.D(net79),
    .GATE(net82),
    .Q(\ConfigBits[70] ),
    .Q_N(\ConfigBits_N[70] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame10_bit9  (.D(net80),
    .GATE(net82),
    .Q(\ConfigBits[71] ),
    .Q_N(\ConfigBits_N[71] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit0  (.D(net49),
    .GATE(net83),
    .Q(\ConfigBits[30] ),
    .Q_N(\ConfigBits_N[30] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit1  (.D(net60),
    .GATE(net83),
    .Q(\ConfigBits[31] ),
    .Q_N(\ConfigBits_N[31] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit10  (.D(net50),
    .GATE(net83),
    .Q(\ConfigBits[40] ),
    .Q_N(\ConfigBits_N[40] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit11  (.D(net51),
    .GATE(net83),
    .Q(\ConfigBits[41] ),
    .Q_N(\ConfigBits_N[41] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit12  (.D(net52),
    .GATE(net83),
    .Q(\ConfigBits[42] ),
    .Q_N(\ConfigBits_N[42] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit13  (.D(net53),
    .GATE(net83),
    .Q(\ConfigBits[43] ),
    .Q_N(\ConfigBits_N[43] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit14  (.D(net54),
    .GATE(net83),
    .Q(\ConfigBits[44] ),
    .Q_N(\ConfigBits_N[44] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit15  (.D(net55),
    .GATE(net83),
    .Q(\ConfigBits[45] ),
    .Q_N(\ConfigBits_N[45] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit16  (.D(net56),
    .GATE(net83),
    .Q(\ConfigBits[46] ),
    .Q_N(\ConfigBits_N[46] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit17  (.D(net57),
    .GATE(net83),
    .Q(\ConfigBits[47] ),
    .Q_N(\ConfigBits_N[47] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit18  (.D(net58),
    .GATE(net83),
    .Q(\ConfigBits[48] ),
    .Q_N(\ConfigBits_N[48] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit19  (.D(net59),
    .GATE(net83),
    .Q(\ConfigBits[49] ),
    .Q_N(\ConfigBits_N[49] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit2  (.D(net71),
    .GATE(net83),
    .Q(\ConfigBits[32] ),
    .Q_N(\ConfigBits_N[32] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit20  (.D(net61),
    .GATE(net83),
    .Q(\ConfigBits[50] ),
    .Q_N(\ConfigBits_N[50] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit21  (.D(net62),
    .GATE(net83),
    .Q(\ConfigBits[51] ),
    .Q_N(\ConfigBits_N[51] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit22  (.D(net63),
    .GATE(net83),
    .Q(\ConfigBits[52] ),
    .Q_N(\ConfigBits_N[52] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit23  (.D(net64),
    .GATE(net83),
    .Q(\ConfigBits[53] ),
    .Q_N(\ConfigBits_N[53] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit24  (.D(net65),
    .GATE(net83),
    .Q(\ConfigBits[54] ),
    .Q_N(\ConfigBits_N[54] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit25  (.D(net66),
    .GATE(net83),
    .Q(\ConfigBits[55] ),
    .Q_N(\ConfigBits_N[55] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit26  (.D(net67),
    .GATE(net83),
    .Q(\ConfigBits[56] ),
    .Q_N(\ConfigBits_N[56] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit27  (.D(net68),
    .GATE(net83),
    .Q(\ConfigBits[57] ),
    .Q_N(\ConfigBits_N[57] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit28  (.D(net69),
    .GATE(net83),
    .Q(\ConfigBits[58] ),
    .Q_N(\ConfigBits_N[58] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit29  (.D(net70),
    .GATE(net83),
    .Q(\ConfigBits[59] ),
    .Q_N(\ConfigBits_N[59] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit3  (.D(net74),
    .GATE(net83),
    .Q(\ConfigBits[33] ),
    .Q_N(\ConfigBits_N[33] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit30  (.D(net72),
    .GATE(net83),
    .Q(\ConfigBits[60] ),
    .Q_N(\ConfigBits_N[60] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit31  (.D(net73),
    .GATE(net83),
    .Q(\ConfigBits[61] ),
    .Q_N(\ConfigBits_N[61] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit4  (.D(net75),
    .GATE(net83),
    .Q(\ConfigBits[34] ),
    .Q_N(\ConfigBits_N[34] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit5  (.D(net76),
    .GATE(net83),
    .Q(\ConfigBits[35] ),
    .Q_N(\ConfigBits_N[35] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit6  (.D(net77),
    .GATE(net83),
    .Q(\ConfigBits[36] ),
    .Q_N(\ConfigBits_N[36] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit7  (.D(net78),
    .GATE(net83),
    .Q(\ConfigBits[37] ),
    .Q_N(\ConfigBits_N[37] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit8  (.D(net79),
    .GATE(net83),
    .Q(\ConfigBits[38] ),
    .Q_N(\ConfigBits_N[38] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame11_bit9  (.D(net80),
    .GATE(net83),
    .Q(\ConfigBits[39] ),
    .Q_N(\ConfigBits_N[39] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit10  (.D(net50),
    .GATE(net84),
    .Q(\ConfigBits[8] ),
    .Q_N(\ConfigBits_N[8] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit11  (.D(net51),
    .GATE(net84),
    .Q(\ConfigBits[9] ),
    .Q_N(\ConfigBits_N[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit12  (.D(net52),
    .GATE(net84),
    .Q(\ConfigBits[10] ),
    .Q_N(\ConfigBits_N[10] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit13  (.D(net53),
    .GATE(net84),
    .Q(\ConfigBits[11] ),
    .Q_N(\ConfigBits_N[11] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit14  (.D(net54),
    .GATE(net84),
    .Q(\ConfigBits[12] ),
    .Q_N(\ConfigBits_N[12] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit15  (.D(net55),
    .GATE(net84),
    .Q(\ConfigBits[13] ),
    .Q_N(\ConfigBits_N[13] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit16  (.D(net56),
    .GATE(net84),
    .Q(\ConfigBits[14] ),
    .Q_N(\ConfigBits_N[14] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit17  (.D(net57),
    .GATE(net84),
    .Q(\ConfigBits[15] ),
    .Q_N(\ConfigBits_N[15] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit18  (.D(net58),
    .GATE(net84),
    .Q(\ConfigBits[16] ),
    .Q_N(\ConfigBits_N[16] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit19  (.D(net59),
    .GATE(net84),
    .Q(\ConfigBits[17] ),
    .Q_N(\ConfigBits_N[17] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit2  (.D(net71),
    .GATE(net84),
    .Q(\ConfigBits[0] ),
    .Q_N(\ConfigBits_N[0] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit20  (.D(net61),
    .GATE(net84),
    .Q(\ConfigBits[18] ),
    .Q_N(\ConfigBits_N[18] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit21  (.D(net62),
    .GATE(net84),
    .Q(\ConfigBits[19] ),
    .Q_N(\ConfigBits_N[19] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit22  (.D(net63),
    .GATE(net84),
    .Q(\ConfigBits[20] ),
    .Q_N(\ConfigBits_N[20] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit23  (.D(net64),
    .GATE(net84),
    .Q(\ConfigBits[21] ),
    .Q_N(\ConfigBits_N[21] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit24  (.D(net65),
    .GATE(net84),
    .Q(\ConfigBits[22] ),
    .Q_N(\ConfigBits_N[22] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit25  (.D(net66),
    .GATE(net84),
    .Q(\ConfigBits[23] ),
    .Q_N(\ConfigBits_N[23] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit26  (.D(net67),
    .GATE(net84),
    .Q(\ConfigBits[24] ),
    .Q_N(\ConfigBits_N[24] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit27  (.D(net68),
    .GATE(net84),
    .Q(\ConfigBits[25] ),
    .Q_N(\ConfigBits_N[25] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit28  (.D(net69),
    .GATE(net84),
    .Q(\ConfigBits[26] ),
    .Q_N(\ConfigBits_N[26] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit29  (.D(net70),
    .GATE(net84),
    .Q(\ConfigBits[27] ),
    .Q_N(\ConfigBits_N[27] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit3  (.D(net74),
    .GATE(net84),
    .Q(\ConfigBits[1] ),
    .Q_N(\ConfigBits_N[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit30  (.D(net72),
    .GATE(net84),
    .Q(\ConfigBits[28] ),
    .Q_N(\ConfigBits_N[28] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit31  (.D(net73),
    .GATE(net84),
    .Q(\ConfigBits[29] ),
    .Q_N(\ConfigBits_N[29] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit4  (.D(net75),
    .GATE(net84),
    .Q(\ConfigBits[2] ),
    .Q_N(\ConfigBits_N[2] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit5  (.D(net76),
    .GATE(net84),
    .Q(\ConfigBits[3] ),
    .Q_N(\ConfigBits_N[3] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit6  (.D(net77),
    .GATE(net84),
    .Q(\ConfigBits[4] ),
    .Q_N(\ConfigBits_N[4] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit7  (.D(net78),
    .GATE(net84),
    .Q(\ConfigBits[5] ),
    .Q_N(\ConfigBits_N[5] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit8  (.D(net79),
    .GATE(net84),
    .Q(\ConfigBits[6] ),
    .Q_N(\ConfigBits_N[6] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame12_bit9  (.D(net80),
    .GATE(net84),
    .Q(\ConfigBits[7] ),
    .Q_N(\ConfigBits_N[7] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit0  (.D(net49),
    .GATE(net92),
    .Q(\ConfigBits[350] ),
    .Q_N(\ConfigBits_N[350] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit1  (.D(net60),
    .GATE(net92),
    .Q(\ConfigBits[351] ),
    .Q_N(\ConfigBits_N[351] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit10  (.D(net50),
    .GATE(net92),
    .Q(\ConfigBits[360] ),
    .Q_N(\ConfigBits_N[360] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit11  (.D(net51),
    .GATE(net92),
    .Q(\ConfigBits[361] ),
    .Q_N(\ConfigBits_N[361] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit12  (.D(net52),
    .GATE(net92),
    .Q(\ConfigBits[362] ),
    .Q_N(\ConfigBits_N[362] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit13  (.D(net53),
    .GATE(net92),
    .Q(\ConfigBits[363] ),
    .Q_N(\ConfigBits_N[363] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit14  (.D(net54),
    .GATE(net92),
    .Q(\ConfigBits[364] ),
    .Q_N(\ConfigBits_N[364] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit15  (.D(net55),
    .GATE(net92),
    .Q(\ConfigBits[365] ),
    .Q_N(\ConfigBits_N[365] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit16  (.D(net56),
    .GATE(net92),
    .Q(\ConfigBits[366] ),
    .Q_N(\ConfigBits_N[366] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit17  (.D(net57),
    .GATE(net92),
    .Q(\ConfigBits[367] ),
    .Q_N(\ConfigBits_N[367] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit18  (.D(net58),
    .GATE(net92),
    .Q(\ConfigBits[368] ),
    .Q_N(\ConfigBits_N[368] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit19  (.D(net59),
    .GATE(net92),
    .Q(\ConfigBits[369] ),
    .Q_N(\ConfigBits_N[369] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit2  (.D(net71),
    .GATE(net92),
    .Q(\ConfigBits[352] ),
    .Q_N(\ConfigBits_N[352] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit20  (.D(net61),
    .GATE(net92),
    .Q(\ConfigBits[370] ),
    .Q_N(\ConfigBits_N[370] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit21  (.D(net62),
    .GATE(net92),
    .Q(\ConfigBits[371] ),
    .Q_N(\ConfigBits_N[371] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit22  (.D(net63),
    .GATE(net92),
    .Q(\ConfigBits[372] ),
    .Q_N(\ConfigBits_N[372] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit23  (.D(net64),
    .GATE(net92),
    .Q(\ConfigBits[373] ),
    .Q_N(\ConfigBits_N[373] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit24  (.D(net65),
    .GATE(net92),
    .Q(\ConfigBits[374] ),
    .Q_N(\ConfigBits_N[374] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit25  (.D(net66),
    .GATE(net92),
    .Q(\ConfigBits[375] ),
    .Q_N(\ConfigBits_N[375] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit26  (.D(net67),
    .GATE(net92),
    .Q(\ConfigBits[376] ),
    .Q_N(\ConfigBits_N[376] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit27  (.D(net68),
    .GATE(net92),
    .Q(\ConfigBits[377] ),
    .Q_N(\ConfigBits_N[377] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit28  (.D(net69),
    .GATE(net92),
    .Q(\ConfigBits[378] ),
    .Q_N(\ConfigBits_N[378] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit29  (.D(net70),
    .GATE(net92),
    .Q(\ConfigBits[379] ),
    .Q_N(\ConfigBits_N[379] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit3  (.D(net74),
    .GATE(net92),
    .Q(\ConfigBits[353] ),
    .Q_N(\ConfigBits_N[353] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit30  (.D(net72),
    .GATE(net92),
    .Q(\ConfigBits[380] ),
    .Q_N(\ConfigBits_N[380] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit31  (.D(net73),
    .GATE(net92),
    .Q(\ConfigBits[381] ),
    .Q_N(\ConfigBits_N[381] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit4  (.D(net75),
    .GATE(net92),
    .Q(\ConfigBits[354] ),
    .Q_N(\ConfigBits_N[354] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit5  (.D(net76),
    .GATE(net92),
    .Q(\ConfigBits[355] ),
    .Q_N(\ConfigBits_N[355] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit6  (.D(net77),
    .GATE(net92),
    .Q(\ConfigBits[356] ),
    .Q_N(\ConfigBits_N[356] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit7  (.D(net78),
    .GATE(net92),
    .Q(\ConfigBits[357] ),
    .Q_N(\ConfigBits_N[357] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit8  (.D(net79),
    .GATE(net92),
    .Q(\ConfigBits[358] ),
    .Q_N(\ConfigBits_N[358] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame1_bit9  (.D(net80),
    .GATE(net92),
    .Q(\ConfigBits[359] ),
    .Q_N(\ConfigBits_N[359] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit0  (.D(net49),
    .GATE(net93),
    .Q(\ConfigBits[318] ),
    .Q_N(\ConfigBits_N[318] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit1  (.D(net60),
    .GATE(net93),
    .Q(\ConfigBits[319] ),
    .Q_N(\ConfigBits_N[319] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit10  (.D(net50),
    .GATE(net93),
    .Q(\ConfigBits[328] ),
    .Q_N(\ConfigBits_N[328] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit11  (.D(net51),
    .GATE(net93),
    .Q(\ConfigBits[329] ),
    .Q_N(\ConfigBits_N[329] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit12  (.D(net52),
    .GATE(net93),
    .Q(\ConfigBits[330] ),
    .Q_N(\ConfigBits_N[330] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit13  (.D(net53),
    .GATE(net93),
    .Q(\ConfigBits[331] ),
    .Q_N(\ConfigBits_N[331] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit14  (.D(net54),
    .GATE(net93),
    .Q(\ConfigBits[332] ),
    .Q_N(\ConfigBits_N[332] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit15  (.D(net55),
    .GATE(net93),
    .Q(\ConfigBits[333] ),
    .Q_N(\ConfigBits_N[333] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit16  (.D(net56),
    .GATE(net93),
    .Q(\ConfigBits[334] ),
    .Q_N(\ConfigBits_N[334] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit17  (.D(net57),
    .GATE(net93),
    .Q(\ConfigBits[335] ),
    .Q_N(\ConfigBits_N[335] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit18  (.D(net58),
    .GATE(net93),
    .Q(\ConfigBits[336] ),
    .Q_N(\ConfigBits_N[336] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit19  (.D(net59),
    .GATE(net93),
    .Q(\ConfigBits[337] ),
    .Q_N(\ConfigBits_N[337] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit2  (.D(net71),
    .GATE(net93),
    .Q(\ConfigBits[320] ),
    .Q_N(\ConfigBits_N[320] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit20  (.D(net61),
    .GATE(net93),
    .Q(\ConfigBits[338] ),
    .Q_N(\ConfigBits_N[338] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit21  (.D(net62),
    .GATE(net93),
    .Q(\ConfigBits[339] ),
    .Q_N(\ConfigBits_N[339] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit22  (.D(net63),
    .GATE(net93),
    .Q(\ConfigBits[340] ),
    .Q_N(\ConfigBits_N[340] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit23  (.D(net64),
    .GATE(net93),
    .Q(\ConfigBits[341] ),
    .Q_N(\ConfigBits_N[341] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit24  (.D(net65),
    .GATE(net93),
    .Q(\ConfigBits[342] ),
    .Q_N(\ConfigBits_N[342] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit25  (.D(net66),
    .GATE(net93),
    .Q(\ConfigBits[343] ),
    .Q_N(\ConfigBits_N[343] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit26  (.D(net67),
    .GATE(net93),
    .Q(\ConfigBits[344] ),
    .Q_N(\ConfigBits_N[344] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit27  (.D(net68),
    .GATE(net93),
    .Q(\ConfigBits[345] ),
    .Q_N(\ConfigBits_N[345] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit28  (.D(net69),
    .GATE(net93),
    .Q(\ConfigBits[346] ),
    .Q_N(\ConfigBits_N[346] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit29  (.D(net70),
    .GATE(net93),
    .Q(\ConfigBits[347] ),
    .Q_N(\ConfigBits_N[347] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit3  (.D(net74),
    .GATE(net93),
    .Q(\ConfigBits[321] ),
    .Q_N(\ConfigBits_N[321] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit30  (.D(net72),
    .GATE(net93),
    .Q(\ConfigBits[348] ),
    .Q_N(\ConfigBits_N[348] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit31  (.D(net73),
    .GATE(net93),
    .Q(\ConfigBits[349] ),
    .Q_N(\ConfigBits_N[349] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit4  (.D(net75),
    .GATE(net93),
    .Q(\ConfigBits[322] ),
    .Q_N(\ConfigBits_N[322] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit5  (.D(net76),
    .GATE(net93),
    .Q(\ConfigBits[323] ),
    .Q_N(\ConfigBits_N[323] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit6  (.D(net77),
    .GATE(net93),
    .Q(\ConfigBits[324] ),
    .Q_N(\ConfigBits_N[324] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit7  (.D(net78),
    .GATE(net93),
    .Q(\ConfigBits[325] ),
    .Q_N(\ConfigBits_N[325] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit8  (.D(net79),
    .GATE(net93),
    .Q(\ConfigBits[326] ),
    .Q_N(\ConfigBits_N[326] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame2_bit9  (.D(net80),
    .GATE(net93),
    .Q(\ConfigBits[327] ),
    .Q_N(\ConfigBits_N[327] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit0  (.D(net49),
    .GATE(net94),
    .Q(\ConfigBits[286] ),
    .Q_N(\ConfigBits_N[286] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit1  (.D(net60),
    .GATE(net94),
    .Q(\ConfigBits[287] ),
    .Q_N(\ConfigBits_N[287] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit10  (.D(net50),
    .GATE(net94),
    .Q(\ConfigBits[296] ),
    .Q_N(\ConfigBits_N[296] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit11  (.D(net51),
    .GATE(net94),
    .Q(\ConfigBits[297] ),
    .Q_N(\ConfigBits_N[297] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit12  (.D(net52),
    .GATE(net94),
    .Q(\ConfigBits[298] ),
    .Q_N(\ConfigBits_N[298] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit13  (.D(net53),
    .GATE(net94),
    .Q(\ConfigBits[299] ),
    .Q_N(\ConfigBits_N[299] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit14  (.D(net54),
    .GATE(net94),
    .Q(\ConfigBits[300] ),
    .Q_N(\ConfigBits_N[300] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit15  (.D(net55),
    .GATE(net94),
    .Q(\ConfigBits[301] ),
    .Q_N(\ConfigBits_N[301] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit16  (.D(net56),
    .GATE(net94),
    .Q(\ConfigBits[302] ),
    .Q_N(\ConfigBits_N[302] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit17  (.D(net57),
    .GATE(net94),
    .Q(\ConfigBits[303] ),
    .Q_N(\ConfigBits_N[303] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit18  (.D(net58),
    .GATE(net94),
    .Q(\ConfigBits[304] ),
    .Q_N(\ConfigBits_N[304] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit19  (.D(net59),
    .GATE(net94),
    .Q(\ConfigBits[305] ),
    .Q_N(\ConfigBits_N[305] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit2  (.D(net71),
    .GATE(net94),
    .Q(\ConfigBits[288] ),
    .Q_N(\ConfigBits_N[288] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit20  (.D(net61),
    .GATE(net94),
    .Q(\ConfigBits[306] ),
    .Q_N(\ConfigBits_N[306] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit21  (.D(net62),
    .GATE(net94),
    .Q(\ConfigBits[307] ),
    .Q_N(\ConfigBits_N[307] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit22  (.D(net63),
    .GATE(net94),
    .Q(\ConfigBits[308] ),
    .Q_N(\ConfigBits_N[308] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit23  (.D(net64),
    .GATE(net94),
    .Q(\ConfigBits[309] ),
    .Q_N(\ConfigBits_N[309] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit24  (.D(net65),
    .GATE(net94),
    .Q(\ConfigBits[310] ),
    .Q_N(\ConfigBits_N[310] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit25  (.D(net66),
    .GATE(net94),
    .Q(\ConfigBits[311] ),
    .Q_N(\ConfigBits_N[311] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit26  (.D(net67),
    .GATE(net94),
    .Q(\ConfigBits[312] ),
    .Q_N(\ConfigBits_N[312] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit27  (.D(net68),
    .GATE(net94),
    .Q(\ConfigBits[313] ),
    .Q_N(\ConfigBits_N[313] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit28  (.D(net69),
    .GATE(net94),
    .Q(\ConfigBits[314] ),
    .Q_N(\ConfigBits_N[314] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit29  (.D(net70),
    .GATE(net94),
    .Q(\ConfigBits[315] ),
    .Q_N(\ConfigBits_N[315] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit3  (.D(net74),
    .GATE(net94),
    .Q(\ConfigBits[289] ),
    .Q_N(\ConfigBits_N[289] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit30  (.D(net72),
    .GATE(net94),
    .Q(\ConfigBits[316] ),
    .Q_N(\ConfigBits_N[316] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit31  (.D(net73),
    .GATE(net94),
    .Q(\ConfigBits[317] ),
    .Q_N(\ConfigBits_N[317] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit4  (.D(net75),
    .GATE(net94),
    .Q(\ConfigBits[290] ),
    .Q_N(\ConfigBits_N[290] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit5  (.D(net76),
    .GATE(net94),
    .Q(\ConfigBits[291] ),
    .Q_N(\ConfigBits_N[291] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit6  (.D(net77),
    .GATE(net94),
    .Q(\ConfigBits[292] ),
    .Q_N(\ConfigBits_N[292] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit7  (.D(net78),
    .GATE(net94),
    .Q(\ConfigBits[293] ),
    .Q_N(\ConfigBits_N[293] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit8  (.D(net79),
    .GATE(net94),
    .Q(\ConfigBits[294] ),
    .Q_N(\ConfigBits_N[294] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame3_bit9  (.D(net80),
    .GATE(net94),
    .Q(\ConfigBits[295] ),
    .Q_N(\ConfigBits_N[295] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit0  (.D(net49),
    .GATE(net95),
    .Q(\ConfigBits[254] ),
    .Q_N(\ConfigBits_N[254] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit1  (.D(net60),
    .GATE(net95),
    .Q(\ConfigBits[255] ),
    .Q_N(\ConfigBits_N[255] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit10  (.D(net50),
    .GATE(net95),
    .Q(\ConfigBits[264] ),
    .Q_N(\ConfigBits_N[264] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit11  (.D(net51),
    .GATE(net95),
    .Q(\ConfigBits[265] ),
    .Q_N(\ConfigBits_N[265] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit12  (.D(net52),
    .GATE(net95),
    .Q(\ConfigBits[266] ),
    .Q_N(\ConfigBits_N[266] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit13  (.D(net53),
    .GATE(net95),
    .Q(\ConfigBits[267] ),
    .Q_N(\ConfigBits_N[267] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit14  (.D(net54),
    .GATE(net95),
    .Q(\ConfigBits[268] ),
    .Q_N(\ConfigBits_N[268] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit15  (.D(net55),
    .GATE(net95),
    .Q(\ConfigBits[269] ),
    .Q_N(\ConfigBits_N[269] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit16  (.D(net56),
    .GATE(net95),
    .Q(\ConfigBits[270] ),
    .Q_N(\ConfigBits_N[270] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit17  (.D(net57),
    .GATE(net95),
    .Q(\ConfigBits[271] ),
    .Q_N(\ConfigBits_N[271] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit18  (.D(net58),
    .GATE(net95),
    .Q(\ConfigBits[272] ),
    .Q_N(\ConfigBits_N[272] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit19  (.D(net59),
    .GATE(net95),
    .Q(\ConfigBits[273] ),
    .Q_N(\ConfigBits_N[273] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit2  (.D(net71),
    .GATE(net95),
    .Q(\ConfigBits[256] ),
    .Q_N(\ConfigBits_N[256] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit20  (.D(net61),
    .GATE(net95),
    .Q(\ConfigBits[274] ),
    .Q_N(\ConfigBits_N[274] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit21  (.D(net62),
    .GATE(net95),
    .Q(\ConfigBits[275] ),
    .Q_N(\ConfigBits_N[275] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit22  (.D(net63),
    .GATE(net95),
    .Q(\ConfigBits[276] ),
    .Q_N(\ConfigBits_N[276] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit23  (.D(net64),
    .GATE(net95),
    .Q(\ConfigBits[277] ),
    .Q_N(\ConfigBits_N[277] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit24  (.D(net65),
    .GATE(net95),
    .Q(\ConfigBits[278] ),
    .Q_N(\ConfigBits_N[278] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit25  (.D(net66),
    .GATE(net95),
    .Q(\ConfigBits[279] ),
    .Q_N(\ConfigBits_N[279] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit26  (.D(net67),
    .GATE(net95),
    .Q(\ConfigBits[280] ),
    .Q_N(\ConfigBits_N[280] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit27  (.D(net68),
    .GATE(net95),
    .Q(\ConfigBits[281] ),
    .Q_N(\ConfigBits_N[281] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit28  (.D(net69),
    .GATE(net95),
    .Q(\ConfigBits[282] ),
    .Q_N(\ConfigBits_N[282] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit29  (.D(net70),
    .GATE(net95),
    .Q(\ConfigBits[283] ),
    .Q_N(\ConfigBits_N[283] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit3  (.D(net74),
    .GATE(net95),
    .Q(\ConfigBits[257] ),
    .Q_N(\ConfigBits_N[257] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit30  (.D(net72),
    .GATE(net95),
    .Q(\ConfigBits[284] ),
    .Q_N(\ConfigBits_N[284] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit31  (.D(net73),
    .GATE(net95),
    .Q(\ConfigBits[285] ),
    .Q_N(\ConfigBits_N[285] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit4  (.D(net75),
    .GATE(net95),
    .Q(\ConfigBits[258] ),
    .Q_N(\ConfigBits_N[258] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit5  (.D(net76),
    .GATE(net95),
    .Q(\ConfigBits[259] ),
    .Q_N(\ConfigBits_N[259] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit6  (.D(net77),
    .GATE(net95),
    .Q(\ConfigBits[260] ),
    .Q_N(\ConfigBits_N[260] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit7  (.D(net78),
    .GATE(net95),
    .Q(\ConfigBits[261] ),
    .Q_N(\ConfigBits_N[261] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit8  (.D(net79),
    .GATE(net95),
    .Q(\ConfigBits[262] ),
    .Q_N(\ConfigBits_N[262] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame4_bit9  (.D(net80),
    .GATE(net95),
    .Q(\ConfigBits[263] ),
    .Q_N(\ConfigBits_N[263] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit0  (.D(net49),
    .GATE(net96),
    .Q(\ConfigBits[222] ),
    .Q_N(\ConfigBits_N[222] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit1  (.D(net60),
    .GATE(net96),
    .Q(\ConfigBits[223] ),
    .Q_N(\ConfigBits_N[223] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit10  (.D(net50),
    .GATE(net96),
    .Q(\ConfigBits[232] ),
    .Q_N(\ConfigBits_N[232] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit11  (.D(net51),
    .GATE(net96),
    .Q(\ConfigBits[233] ),
    .Q_N(\ConfigBits_N[233] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit12  (.D(net52),
    .GATE(net96),
    .Q(\ConfigBits[234] ),
    .Q_N(\ConfigBits_N[234] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit13  (.D(net53),
    .GATE(net96),
    .Q(\ConfigBits[235] ),
    .Q_N(\ConfigBits_N[235] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit14  (.D(net54),
    .GATE(net96),
    .Q(\ConfigBits[236] ),
    .Q_N(\ConfigBits_N[236] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit15  (.D(net55),
    .GATE(net96),
    .Q(\ConfigBits[237] ),
    .Q_N(\ConfigBits_N[237] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit16  (.D(net56),
    .GATE(net96),
    .Q(\ConfigBits[238] ),
    .Q_N(\ConfigBits_N[238] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit17  (.D(net57),
    .GATE(net96),
    .Q(\ConfigBits[239] ),
    .Q_N(\ConfigBits_N[239] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit18  (.D(net58),
    .GATE(net96),
    .Q(\ConfigBits[240] ),
    .Q_N(\ConfigBits_N[240] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit19  (.D(net59),
    .GATE(net96),
    .Q(\ConfigBits[241] ),
    .Q_N(\ConfigBits_N[241] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit2  (.D(net71),
    .GATE(net96),
    .Q(\ConfigBits[224] ),
    .Q_N(\ConfigBits_N[224] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit20  (.D(net61),
    .GATE(net96),
    .Q(\ConfigBits[242] ),
    .Q_N(\ConfigBits_N[242] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit21  (.D(net62),
    .GATE(net96),
    .Q(\ConfigBits[243] ),
    .Q_N(\ConfigBits_N[243] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit22  (.D(net63),
    .GATE(net96),
    .Q(\ConfigBits[244] ),
    .Q_N(\ConfigBits_N[244] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit23  (.D(net64),
    .GATE(net96),
    .Q(\ConfigBits[245] ),
    .Q_N(\ConfigBits_N[245] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit24  (.D(net65),
    .GATE(net96),
    .Q(\ConfigBits[246] ),
    .Q_N(\ConfigBits_N[246] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit25  (.D(net66),
    .GATE(net96),
    .Q(\ConfigBits[247] ),
    .Q_N(\ConfigBits_N[247] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit26  (.D(net67),
    .GATE(net96),
    .Q(\ConfigBits[248] ),
    .Q_N(\ConfigBits_N[248] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit27  (.D(net68),
    .GATE(net96),
    .Q(\ConfigBits[249] ),
    .Q_N(\ConfigBits_N[249] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit28  (.D(net69),
    .GATE(net96),
    .Q(\ConfigBits[250] ),
    .Q_N(\ConfigBits_N[250] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit29  (.D(net70),
    .GATE(net96),
    .Q(\ConfigBits[251] ),
    .Q_N(\ConfigBits_N[251] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit3  (.D(net74),
    .GATE(net96),
    .Q(\ConfigBits[225] ),
    .Q_N(\ConfigBits_N[225] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit30  (.D(net72),
    .GATE(net96),
    .Q(\ConfigBits[252] ),
    .Q_N(\ConfigBits_N[252] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit31  (.D(net73),
    .GATE(net96),
    .Q(\ConfigBits[253] ),
    .Q_N(\ConfigBits_N[253] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit4  (.D(net75),
    .GATE(net96),
    .Q(\ConfigBits[226] ),
    .Q_N(\ConfigBits_N[226] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit5  (.D(net76),
    .GATE(net96),
    .Q(\ConfigBits[227] ),
    .Q_N(\ConfigBits_N[227] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit6  (.D(net77),
    .GATE(net96),
    .Q(\ConfigBits[228] ),
    .Q_N(\ConfigBits_N[228] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit7  (.D(net78),
    .GATE(net96),
    .Q(\ConfigBits[229] ),
    .Q_N(\ConfigBits_N[229] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit8  (.D(net79),
    .GATE(net96),
    .Q(\ConfigBits[230] ),
    .Q_N(\ConfigBits_N[230] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame5_bit9  (.D(net80),
    .GATE(net96),
    .Q(\ConfigBits[231] ),
    .Q_N(\ConfigBits_N[231] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit0  (.D(net49),
    .GATE(net97),
    .Q(\ConfigBits[190] ),
    .Q_N(\ConfigBits_N[190] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit1  (.D(net60),
    .GATE(net97),
    .Q(\ConfigBits[191] ),
    .Q_N(\ConfigBits_N[191] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit10  (.D(net50),
    .GATE(net97),
    .Q(\ConfigBits[200] ),
    .Q_N(\ConfigBits_N[200] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit11  (.D(net51),
    .GATE(net97),
    .Q(\ConfigBits[201] ),
    .Q_N(\ConfigBits_N[201] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit12  (.D(net52),
    .GATE(net97),
    .Q(\ConfigBits[202] ),
    .Q_N(\ConfigBits_N[202] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit13  (.D(net53),
    .GATE(net97),
    .Q(\ConfigBits[203] ),
    .Q_N(\ConfigBits_N[203] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit14  (.D(net54),
    .GATE(net97),
    .Q(\ConfigBits[204] ),
    .Q_N(\ConfigBits_N[204] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit15  (.D(net55),
    .GATE(net97),
    .Q(\ConfigBits[205] ),
    .Q_N(\ConfigBits_N[205] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit16  (.D(net56),
    .GATE(net97),
    .Q(\ConfigBits[206] ),
    .Q_N(\ConfigBits_N[206] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit17  (.D(net57),
    .GATE(net97),
    .Q(\ConfigBits[207] ),
    .Q_N(\ConfigBits_N[207] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit18  (.D(net58),
    .GATE(net97),
    .Q(\ConfigBits[208] ),
    .Q_N(\ConfigBits_N[208] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit19  (.D(net59),
    .GATE(net97),
    .Q(\ConfigBits[209] ),
    .Q_N(\ConfigBits_N[209] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit2  (.D(net71),
    .GATE(net97),
    .Q(\ConfigBits[192] ),
    .Q_N(\ConfigBits_N[192] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit20  (.D(net61),
    .GATE(net97),
    .Q(\ConfigBits[210] ),
    .Q_N(\ConfigBits_N[210] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit21  (.D(net62),
    .GATE(net97),
    .Q(\ConfigBits[211] ),
    .Q_N(\ConfigBits_N[211] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit22  (.D(net63),
    .GATE(net97),
    .Q(\ConfigBits[212] ),
    .Q_N(\ConfigBits_N[212] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit23  (.D(net64),
    .GATE(net97),
    .Q(\ConfigBits[213] ),
    .Q_N(\ConfigBits_N[213] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit24  (.D(net65),
    .GATE(net97),
    .Q(\ConfigBits[214] ),
    .Q_N(\ConfigBits_N[214] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit25  (.D(net66),
    .GATE(net97),
    .Q(\ConfigBits[215] ),
    .Q_N(\ConfigBits_N[215] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit26  (.D(net67),
    .GATE(net97),
    .Q(\ConfigBits[216] ),
    .Q_N(\ConfigBits_N[216] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit27  (.D(net68),
    .GATE(net97),
    .Q(\ConfigBits[217] ),
    .Q_N(\ConfigBits_N[217] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit28  (.D(net69),
    .GATE(net97),
    .Q(\ConfigBits[218] ),
    .Q_N(\ConfigBits_N[218] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit29  (.D(net70),
    .GATE(net97),
    .Q(\ConfigBits[219] ),
    .Q_N(\ConfigBits_N[219] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit3  (.D(net74),
    .GATE(net97),
    .Q(\ConfigBits[193] ),
    .Q_N(\ConfigBits_N[193] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit30  (.D(net72),
    .GATE(net97),
    .Q(\ConfigBits[220] ),
    .Q_N(\ConfigBits_N[220] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit31  (.D(net73),
    .GATE(net97),
    .Q(\ConfigBits[221] ),
    .Q_N(\ConfigBits_N[221] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit4  (.D(net75),
    .GATE(net97),
    .Q(\ConfigBits[194] ),
    .Q_N(\ConfigBits_N[194] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit5  (.D(net76),
    .GATE(net97),
    .Q(\ConfigBits[195] ),
    .Q_N(\ConfigBits_N[195] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit6  (.D(net77),
    .GATE(net97),
    .Q(\ConfigBits[196] ),
    .Q_N(\ConfigBits_N[196] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit7  (.D(net78),
    .GATE(net97),
    .Q(\ConfigBits[197] ),
    .Q_N(\ConfigBits_N[197] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit8  (.D(net79),
    .GATE(net97),
    .Q(\ConfigBits[198] ),
    .Q_N(\ConfigBits_N[198] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame6_bit9  (.D(net80),
    .GATE(net97),
    .Q(\ConfigBits[199] ),
    .Q_N(\ConfigBits_N[199] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit0  (.D(net49),
    .GATE(net98),
    .Q(\ConfigBits[158] ),
    .Q_N(\ConfigBits_N[158] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit1  (.D(net60),
    .GATE(net98),
    .Q(\ConfigBits[159] ),
    .Q_N(\ConfigBits_N[159] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit10  (.D(net50),
    .GATE(net98),
    .Q(\ConfigBits[168] ),
    .Q_N(\ConfigBits_N[168] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit11  (.D(net51),
    .GATE(net98),
    .Q(\ConfigBits[169] ),
    .Q_N(\ConfigBits_N[169] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit12  (.D(net52),
    .GATE(net98),
    .Q(\ConfigBits[170] ),
    .Q_N(\ConfigBits_N[170] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit13  (.D(net53),
    .GATE(net98),
    .Q(\ConfigBits[171] ),
    .Q_N(\ConfigBits_N[171] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit14  (.D(net54),
    .GATE(net98),
    .Q(\ConfigBits[172] ),
    .Q_N(\ConfigBits_N[172] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit15  (.D(net55),
    .GATE(net98),
    .Q(\ConfigBits[173] ),
    .Q_N(\ConfigBits_N[173] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit16  (.D(net56),
    .GATE(net98),
    .Q(\ConfigBits[174] ),
    .Q_N(\ConfigBits_N[174] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit17  (.D(net57),
    .GATE(net98),
    .Q(\ConfigBits[175] ),
    .Q_N(\ConfigBits_N[175] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit18  (.D(net58),
    .GATE(net98),
    .Q(\ConfigBits[176] ),
    .Q_N(\ConfigBits_N[176] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit19  (.D(net59),
    .GATE(net98),
    .Q(\ConfigBits[177] ),
    .Q_N(\ConfigBits_N[177] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit2  (.D(net71),
    .GATE(net98),
    .Q(\ConfigBits[160] ),
    .Q_N(\ConfigBits_N[160] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit20  (.D(net61),
    .GATE(net98),
    .Q(\ConfigBits[178] ),
    .Q_N(\ConfigBits_N[178] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit21  (.D(net62),
    .GATE(net98),
    .Q(\ConfigBits[179] ),
    .Q_N(\ConfigBits_N[179] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit22  (.D(net63),
    .GATE(net98),
    .Q(\ConfigBits[180] ),
    .Q_N(\ConfigBits_N[180] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit23  (.D(net64),
    .GATE(net98),
    .Q(\ConfigBits[181] ),
    .Q_N(\ConfigBits_N[181] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit24  (.D(net65),
    .GATE(net98),
    .Q(\ConfigBits[182] ),
    .Q_N(\ConfigBits_N[182] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit25  (.D(net66),
    .GATE(net98),
    .Q(\ConfigBits[183] ),
    .Q_N(\ConfigBits_N[183] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit26  (.D(net67),
    .GATE(net98),
    .Q(\ConfigBits[184] ),
    .Q_N(\ConfigBits_N[184] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit27  (.D(net68),
    .GATE(net98),
    .Q(\ConfigBits[185] ),
    .Q_N(\ConfigBits_N[185] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit28  (.D(net69),
    .GATE(net98),
    .Q(\ConfigBits[186] ),
    .Q_N(\ConfigBits_N[186] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit29  (.D(net70),
    .GATE(net98),
    .Q(\ConfigBits[187] ),
    .Q_N(\ConfigBits_N[187] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit3  (.D(net74),
    .GATE(net98),
    .Q(\ConfigBits[161] ),
    .Q_N(\ConfigBits_N[161] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit30  (.D(net72),
    .GATE(net98),
    .Q(\ConfigBits[188] ),
    .Q_N(\ConfigBits_N[188] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit31  (.D(net73),
    .GATE(net98),
    .Q(\ConfigBits[189] ),
    .Q_N(\ConfigBits_N[189] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit4  (.D(net75),
    .GATE(net98),
    .Q(\ConfigBits[162] ),
    .Q_N(\ConfigBits_N[162] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit5  (.D(net76),
    .GATE(net98),
    .Q(\ConfigBits[163] ),
    .Q_N(\ConfigBits_N[163] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit6  (.D(net77),
    .GATE(net98),
    .Q(\ConfigBits[164] ),
    .Q_N(\ConfigBits_N[164] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit7  (.D(net78),
    .GATE(net98),
    .Q(\ConfigBits[165] ),
    .Q_N(\ConfigBits_N[165] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit8  (.D(net79),
    .GATE(net98),
    .Q(\ConfigBits[166] ),
    .Q_N(\ConfigBits_N[166] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame7_bit9  (.D(net80),
    .GATE(net98),
    .Q(\ConfigBits[167] ),
    .Q_N(\ConfigBits_N[167] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit0  (.D(net49),
    .GATE(net99),
    .Q(\ConfigBits[126] ),
    .Q_N(\ConfigBits_N[126] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit1  (.D(net60),
    .GATE(net99),
    .Q(\ConfigBits[127] ),
    .Q_N(\ConfigBits_N[127] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit10  (.D(net50),
    .GATE(net99),
    .Q(\ConfigBits[136] ),
    .Q_N(\ConfigBits_N[136] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit11  (.D(net51),
    .GATE(net99),
    .Q(\ConfigBits[137] ),
    .Q_N(\ConfigBits_N[137] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit12  (.D(net52),
    .GATE(net99),
    .Q(\ConfigBits[138] ),
    .Q_N(\ConfigBits_N[138] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit13  (.D(net53),
    .GATE(net99),
    .Q(\ConfigBits[139] ),
    .Q_N(\ConfigBits_N[139] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit14  (.D(net54),
    .GATE(net99),
    .Q(\ConfigBits[140] ),
    .Q_N(\ConfigBits_N[140] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit15  (.D(net55),
    .GATE(net99),
    .Q(\ConfigBits[141] ),
    .Q_N(\ConfigBits_N[141] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit16  (.D(net56),
    .GATE(net99),
    .Q(\ConfigBits[142] ),
    .Q_N(\ConfigBits_N[142] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit17  (.D(net57),
    .GATE(net99),
    .Q(\ConfigBits[143] ),
    .Q_N(\ConfigBits_N[143] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit18  (.D(net58),
    .GATE(net99),
    .Q(\ConfigBits[144] ),
    .Q_N(\ConfigBits_N[144] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit19  (.D(net59),
    .GATE(net99),
    .Q(\ConfigBits[145] ),
    .Q_N(\ConfigBits_N[145] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit2  (.D(net71),
    .GATE(net99),
    .Q(\ConfigBits[128] ),
    .Q_N(\ConfigBits_N[128] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit20  (.D(net61),
    .GATE(net99),
    .Q(\ConfigBits[146] ),
    .Q_N(\ConfigBits_N[146] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit21  (.D(net62),
    .GATE(net99),
    .Q(\ConfigBits[147] ),
    .Q_N(\ConfigBits_N[147] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit22  (.D(net63),
    .GATE(net99),
    .Q(\ConfigBits[148] ),
    .Q_N(\ConfigBits_N[148] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit23  (.D(net64),
    .GATE(net99),
    .Q(\ConfigBits[149] ),
    .Q_N(\ConfigBits_N[149] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit24  (.D(net65),
    .GATE(net99),
    .Q(\ConfigBits[150] ),
    .Q_N(\ConfigBits_N[150] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit25  (.D(net66),
    .GATE(net99),
    .Q(\ConfigBits[151] ),
    .Q_N(\ConfigBits_N[151] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit26  (.D(net67),
    .GATE(net99),
    .Q(\ConfigBits[152] ),
    .Q_N(\ConfigBits_N[152] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit27  (.D(net68),
    .GATE(net99),
    .Q(\ConfigBits[153] ),
    .Q_N(\ConfigBits_N[153] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit28  (.D(net69),
    .GATE(net99),
    .Q(\ConfigBits[154] ),
    .Q_N(\ConfigBits_N[154] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit29  (.D(net70),
    .GATE(net99),
    .Q(\ConfigBits[155] ),
    .Q_N(\ConfigBits_N[155] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit3  (.D(net74),
    .GATE(net99),
    .Q(\ConfigBits[129] ),
    .Q_N(\ConfigBits_N[129] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit30  (.D(net72),
    .GATE(net99),
    .Q(\ConfigBits[156] ),
    .Q_N(\ConfigBits_N[156] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit31  (.D(net73),
    .GATE(net99),
    .Q(\ConfigBits[157] ),
    .Q_N(\ConfigBits_N[157] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit4  (.D(net75),
    .GATE(net99),
    .Q(\ConfigBits[130] ),
    .Q_N(\ConfigBits_N[130] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit5  (.D(net76),
    .GATE(net99),
    .Q(\ConfigBits[131] ),
    .Q_N(\ConfigBits_N[131] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit6  (.D(net77),
    .GATE(net99),
    .Q(\ConfigBits[132] ),
    .Q_N(\ConfigBits_N[132] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit7  (.D(net78),
    .GATE(net99),
    .Q(\ConfigBits[133] ),
    .Q_N(\ConfigBits_N[133] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit8  (.D(net79),
    .GATE(net99),
    .Q(\ConfigBits[134] ),
    .Q_N(\ConfigBits_N[134] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame8_bit9  (.D(net80),
    .GATE(net99),
    .Q(\ConfigBits[135] ),
    .Q_N(\ConfigBits_N[135] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit0  (.D(net49),
    .GATE(net100),
    .Q(\ConfigBits[94] ),
    .Q_N(\ConfigBits_N[94] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit1  (.D(net60),
    .GATE(net100),
    .Q(\ConfigBits[95] ),
    .Q_N(\ConfigBits_N[95] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit10  (.D(net50),
    .GATE(net100),
    .Q(\ConfigBits[104] ),
    .Q_N(\ConfigBits_N[104] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit11  (.D(net51),
    .GATE(net100),
    .Q(\ConfigBits[105] ),
    .Q_N(\ConfigBits_N[105] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit12  (.D(net52),
    .GATE(net100),
    .Q(\ConfigBits[106] ),
    .Q_N(\ConfigBits_N[106] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit13  (.D(net53),
    .GATE(net100),
    .Q(\ConfigBits[107] ),
    .Q_N(\ConfigBits_N[107] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit14  (.D(net54),
    .GATE(net100),
    .Q(\ConfigBits[108] ),
    .Q_N(\ConfigBits_N[108] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit15  (.D(net55),
    .GATE(net100),
    .Q(\ConfigBits[109] ),
    .Q_N(\ConfigBits_N[109] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit16  (.D(net56),
    .GATE(net100),
    .Q(\ConfigBits[110] ),
    .Q_N(\ConfigBits_N[110] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit17  (.D(net57),
    .GATE(net100),
    .Q(\ConfigBits[111] ),
    .Q_N(\ConfigBits_N[111] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit18  (.D(net58),
    .GATE(net100),
    .Q(\ConfigBits[112] ),
    .Q_N(\ConfigBits_N[112] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit19  (.D(net59),
    .GATE(net100),
    .Q(\ConfigBits[113] ),
    .Q_N(\ConfigBits_N[113] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit2  (.D(net71),
    .GATE(net100),
    .Q(\ConfigBits[96] ),
    .Q_N(\ConfigBits_N[96] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit20  (.D(net61),
    .GATE(net100),
    .Q(\ConfigBits[114] ),
    .Q_N(\ConfigBits_N[114] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit21  (.D(net62),
    .GATE(net100),
    .Q(\ConfigBits[115] ),
    .Q_N(\ConfigBits_N[115] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit22  (.D(net63),
    .GATE(net100),
    .Q(\ConfigBits[116] ),
    .Q_N(\ConfigBits_N[116] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit23  (.D(net64),
    .GATE(net100),
    .Q(\ConfigBits[117] ),
    .Q_N(\ConfigBits_N[117] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit24  (.D(net65),
    .GATE(net100),
    .Q(\ConfigBits[118] ),
    .Q_N(\ConfigBits_N[118] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit25  (.D(net66),
    .GATE(net100),
    .Q(\ConfigBits[119] ),
    .Q_N(\ConfigBits_N[119] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit26  (.D(net67),
    .GATE(net100),
    .Q(\ConfigBits[120] ),
    .Q_N(\ConfigBits_N[120] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit27  (.D(net68),
    .GATE(net100),
    .Q(\ConfigBits[121] ),
    .Q_N(\ConfigBits_N[121] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit28  (.D(net69),
    .GATE(net100),
    .Q(\ConfigBits[122] ),
    .Q_N(\ConfigBits_N[122] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit29  (.D(net70),
    .GATE(net100),
    .Q(\ConfigBits[123] ),
    .Q_N(\ConfigBits_N[123] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit3  (.D(net74),
    .GATE(net100),
    .Q(\ConfigBits[97] ),
    .Q_N(\ConfigBits_N[97] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit30  (.D(net72),
    .GATE(net100),
    .Q(\ConfigBits[124] ),
    .Q_N(\ConfigBits_N[124] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit31  (.D(net73),
    .GATE(net100),
    .Q(\ConfigBits[125] ),
    .Q_N(\ConfigBits_N[125] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit4  (.D(net75),
    .GATE(net100),
    .Q(\ConfigBits[98] ),
    .Q_N(\ConfigBits_N[98] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit5  (.D(net76),
    .GATE(net100),
    .Q(\ConfigBits[99] ),
    .Q_N(\ConfigBits_N[99] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit6  (.D(net77),
    .GATE(net100),
    .Q(\ConfigBits[100] ),
    .Q_N(\ConfigBits_N[100] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit7  (.D(net78),
    .GATE(net100),
    .Q(\ConfigBits[101] ),
    .Q_N(\ConfigBits_N[101] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit8  (.D(net79),
    .GATE(net100),
    .Q(\ConfigBits[102] ),
    .Q_N(\ConfigBits_N[102] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RegFile_ConfigMem/Inst_frame9_bit9  (.D(net80),
    .GATE(net100),
    .Q(\ConfigBits[103] ),
    .Q_N(\ConfigBits_N[103] ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_switch_matrix/_00_  (.A(\JE2BEG[0] ),
    .X(net258));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/_01_  (.A(\JE2BEG[1] ),
    .X(net259));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/_02_  (.A(\JE2BEG[2] ),
    .X(net260));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/_03_  (.A(\JE2BEG[3] ),
    .X(net261));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/_04_  (.A(\JE2BEG[4] ),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_switch_matrix/_05_  (.A(\JE2BEG[5] ),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_switch_matrix/_06_  (.A(\JE2BEG[6] ),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_switch_matrix/_07_  (.A(\JE2BEG[7] ),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_switch_matrix/_08_  (.A(net13),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_switch_matrix/_09_  (.A(net14),
    .X(net267));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/_10_  (.A(net15),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_switch_matrix/_11_  (.A(net16),
    .X(net269));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/_12_  (.A(net17),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_switch_matrix/_13_  (.A(net18),
    .X(net271));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/_14_  (.A(net19),
    .X(net272));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/_15_  (.A(net20),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_16_  (.A(\JN2BEG[0] ),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_17_  (.A(\JN2BEG[1] ),
    .X(net359));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/_18_  (.A(\JN2BEG[2] ),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_19_  (.A(\JN2BEG[3] ),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_20_  (.A(\JN2BEG[4] ),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_21_  (.A(\JN2BEG[5] ),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_22_  (.A(\JN2BEG[6] ),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_23_  (.A(\JN2BEG[7] ),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_24_  (.A(net113),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_switch_matrix/_25_  (.A(net114),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_26_  (.A(net115),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RegFile_switch_matrix/_27_  (.A(net116),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_28_  (.A(net117),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_29_  (.A(net118),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_30_  (.A(net119),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_31_  (.A(net120),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_32_  (.A(\JS2BEG[0] ),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_33_  (.A(\JS2BEG[1] ),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_34_  (.A(\JS2BEG[2] ),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_35_  (.A(\JS2BEG[3] ),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_36_  (.A(\JS2BEG[4] ),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_37_  (.A(\JS2BEG[5] ),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_38_  (.A(\JS2BEG[6] ),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_39_  (.A(\JS2BEG[7] ),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_40_  (.A(net165),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_41_  (.A(net166),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_42_  (.A(net167),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_43_  (.A(net168),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_44_  (.A(net169),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_45_  (.A(net170),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_46_  (.A(net171),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_47_  (.A(net172),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_48_  (.A(\JW2BEG[0] ),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_49_  (.A(\JW2BEG[1] ),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_50_  (.A(\JW2BEG[2] ),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_51_  (.A(\JW2BEG[3] ),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_52_  (.A(\JW2BEG[4] ),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_53_  (.A(\JW2BEG[5] ),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_54_  (.A(\JW2BEG[6] ),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_55_  (.A(\JW2BEG[7] ),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_56_  (.A(net218),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_57_  (.A(net219),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_58_  (.A(net220),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_59_  (.A(net221),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_60_  (.A(net222),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_61_  (.A(net223),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/_62_  (.A(net224),
    .X(net477));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/_63_  (.A(net225),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst0  (.A0(net137),
    .A1(net4),
    .A2(net189),
    .A3(net209),
    .S0(\ConfigBits[50] ),
    .S1(\ConfigBits[51] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst1  (.A0(AD0),
    .A1(AD1),
    .A2(AD2),
    .A3(AD3),
    .S0(\ConfigBits[50] ),
    .S1(\ConfigBits[51] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst2  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[50] ),
    .S1(\ConfigBits[51] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst3  (.A0(\J2MID_ABb_BEG[1] ),
    .A1(\J2MID_CDb_BEG[1] ),
    .A2(\J2MID_EFb_BEG[1] ),
    .A3(\J2MID_GHb_BEG[1] ),
    .S0(\ConfigBits[50] ),
    .S1(\ConfigBits[51] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[52] ),
    .S1(\ConfigBits[53] ),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst0  (.A0(net146),
    .A1(net3),
    .A2(net198),
    .A3(net208),
    .S0(\ConfigBits[54] ),
    .S1(\ConfigBits[55] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst1  (.A0(AD0),
    .A1(AD1),
    .A2(AD2),
    .A3(AD3),
    .S0(\ConfigBits[54] ),
    .S1(\ConfigBits[55] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst2  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[54] ),
    .S1(\ConfigBits[55] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst3  (.A0(\J2MID_ABa_BEG[2] ),
    .A1(\J2MID_CDa_BEG[2] ),
    .A2(\J2MID_EFa_BEG[2] ),
    .A3(\J2MID_GHa_BEG[2] ),
    .S0(\ConfigBits[54] ),
    .S1(\ConfigBits[55] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[56] ),
    .S1(\ConfigBits[57] ),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net106),
    .A2(net128),
    .A3(net137),
    .S0(\ConfigBits[286] ),
    .S1(\ConfigBits[287] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst1  (.A0(net6),
    .A1(net24),
    .A2(net158),
    .A3(net211),
    .S0(\ConfigBits[286] ),
    .S1(\ConfigBits[287] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst2  (.A0(net229),
    .A1(AD1),
    .A2(AD2),
    .A3(AD3),
    .S0(\ConfigBits[286] ),
    .S1(\ConfigBits[287] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[286] ),
    .S1(\ConfigBits[287] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[288] ),
    .S1(\ConfigBits[289] ),
    .X(\JE2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst0  (.A0(net101),
    .A1(net107),
    .A2(net129),
    .A3(net144),
    .S0(\ConfigBits[290] ),
    .S1(\ConfigBits[291] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst1  (.A0(net7),
    .A1(net21),
    .A2(net159),
    .A3(net212),
    .S0(\ConfigBits[290] ),
    .S1(\ConfigBits[291] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst2  (.A0(net226),
    .A1(AD0),
    .A2(AD2),
    .A3(AD3),
    .S0(\ConfigBits[290] ),
    .S1(\ConfigBits[291] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[290] ),
    .S1(\ConfigBits[291] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[292] ),
    .S1(\ConfigBits[293] ),
    .X(\JE2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net108),
    .A2(net130),
    .A3(net8),
    .S0(\ConfigBits[294] ),
    .S1(\ConfigBits[295] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst1  (.A0(net24),
    .A1(net160),
    .A2(net197),
    .A3(net213),
    .S0(\ConfigBits[294] ),
    .S1(\ConfigBits[295] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst2  (.A0(net229),
    .A1(AD0),
    .A2(AD1),
    .A3(AD3),
    .S0(\ConfigBits[294] ),
    .S1(\ConfigBits[295] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[294] ),
    .S1(\ConfigBits[295] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[296] ),
    .S1(\ConfigBits[297] ),
    .X(\JE2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net109),
    .A2(net121),
    .A3(net9),
    .S0(\ConfigBits[298] ),
    .S1(\ConfigBits[299] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst1  (.A0(net21),
    .A1(net161),
    .A2(net198),
    .A3(net214),
    .S0(\ConfigBits[298] ),
    .S1(\ConfigBits[299] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst2  (.A0(net226),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[298] ),
    .S1(\ConfigBits[299] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[298] ),
    .S1(\ConfigBits[299] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[300] ),
    .S1(\ConfigBits[301] ),
    .X(\JE2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net110),
    .A2(net2),
    .A3(net10),
    .S0(\ConfigBits[302] ),
    .S1(\ConfigBits[303] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst1  (.A0(net42),
    .A1(net154),
    .A2(net156),
    .A3(net162),
    .S0(\ConfigBits[302] ),
    .S1(\ConfigBits[303] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst2  (.A0(net207),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[302] ),
    .S1(\ConfigBits[303] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[302] ),
    .S1(\ConfigBits[303] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[304] ),
    .S1(\ConfigBits[305] ),
    .X(\JE2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net111),
    .A2(net3),
    .A3(net11),
    .S0(\ConfigBits[306] ),
    .S1(\ConfigBits[307] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst1  (.A0(net41),
    .A1(net153),
    .A2(net155),
    .A3(net163),
    .S0(\ConfigBits[306] ),
    .S1(\ConfigBits[307] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst2  (.A0(net208),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[306] ),
    .S1(\ConfigBits[307] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD0),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[306] ),
    .S1(\ConfigBits[307] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[308] ),
    .S1(\ConfigBits[309] ),
    .X(\JE2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net112),
    .A2(net4),
    .A3(net12),
    .S0(\ConfigBits[310] ),
    .S1(\ConfigBits[311] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst1  (.A0(net40),
    .A1(net154),
    .A2(net156),
    .A3(net164),
    .S0(\ConfigBits[310] ),
    .S1(\ConfigBits[311] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst2  (.A0(net209),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[310] ),
    .S1(\ConfigBits[311] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD0),
    .A2(BD1),
    .A3(BD3),
    .S0(\ConfigBits[310] ),
    .S1(\ConfigBits[311] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[312] ),
    .S1(\ConfigBits[313] ),
    .X(\JE2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst0  (.A0(net101),
    .A1(net105),
    .A2(net1),
    .A3(net5),
    .S0(\ConfigBits[314] ),
    .S1(\ConfigBits[315] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst1  (.A0(net33),
    .A1(net153),
    .A2(net155),
    .A3(net157),
    .S0(\ConfigBits[314] ),
    .S1(\ConfigBits[315] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst2  (.A0(net206),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[314] ),
    .S1(\ConfigBits[315] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD0),
    .A2(BD1),
    .A3(BD2),
    .S0(\ConfigBits[314] ),
    .S1(\ConfigBits[315] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[316] ),
    .S1(\ConfigBits[317] ),
    .X(\JE2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst0  (.A0(net106),
    .A1(net128),
    .A2(net4),
    .A3(net6),
    .S0(\ConfigBits[254] ),
    .S1(\ConfigBits[255] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst1  (.A0(net33),
    .A1(net24),
    .A2(net158),
    .A3(net211),
    .S0(\ConfigBits[254] ),
    .S1(\ConfigBits[255] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst2  (.A0(net229),
    .A1(AD1),
    .A2(AD2),
    .A3(AD3),
    .S0(\ConfigBits[254] ),
    .S1(\ConfigBits[255] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[254] ),
    .S1(\ConfigBits[255] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[256] ),
    .S1(\ConfigBits[257] ),
    .X(\JN2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst0  (.A0(net107),
    .A1(net129),
    .A2(net1),
    .A3(net7),
    .S0(\ConfigBits[258] ),
    .S1(\ConfigBits[259] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst1  (.A0(net40),
    .A1(net21),
    .A2(net159),
    .A3(net212),
    .S0(\ConfigBits[258] ),
    .S1(\ConfigBits[259] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst2  (.A0(net226),
    .A1(AD0),
    .A2(AD2),
    .A3(AD3),
    .S0(\ConfigBits[258] ),
    .S1(\ConfigBits[259] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[258] ),
    .S1(\ConfigBits[259] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[260] ),
    .S1(\ConfigBits[261] ),
    .X(\JN2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst0  (.A0(net108),
    .A1(net130),
    .A2(net2),
    .A3(net8),
    .S0(\ConfigBits[262] ),
    .S1(\ConfigBits[263] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst1  (.A0(net24),
    .A1(net160),
    .A2(net213),
    .A3(net246),
    .S0(\ConfigBits[262] ),
    .S1(\ConfigBits[263] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst2  (.A0(net229),
    .A1(AD0),
    .A2(AD1),
    .A3(AD3),
    .S0(\ConfigBits[262] ),
    .S1(\ConfigBits[263] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[262] ),
    .S1(\ConfigBits[263] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[264] ),
    .S1(\ConfigBits[265] ),
    .X(\JN2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst0  (.A0(net109),
    .A1(net121),
    .A2(net3),
    .A3(net9),
    .S0(\ConfigBits[266] ),
    .S1(\ConfigBits[267] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst1  (.A0(net21),
    .A1(net161),
    .A2(net214),
    .A3(net247),
    .S0(\ConfigBits[266] ),
    .S1(\ConfigBits[267] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst2  (.A0(net226),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[266] ),
    .S1(\ConfigBits[267] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[266] ),
    .S1(\ConfigBits[267] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[268] ),
    .S1(\ConfigBits[269] ),
    .X(\JN2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net110),
    .A2(net146),
    .A3(net2),
    .S0(\ConfigBits[270] ),
    .S1(\ConfigBits[271] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst1  (.A0(net10),
    .A1(net154),
    .A2(net162),
    .A3(net207),
    .S0(\ConfigBits[270] ),
    .S1(\ConfigBits[271] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst2  (.A0(net209),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[270] ),
    .S1(\ConfigBits[271] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[270] ),
    .S1(\ConfigBits[271] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[272] ),
    .S1(\ConfigBits[273] ),
    .X(\JN2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net111),
    .A2(net145),
    .A3(net3),
    .S0(\ConfigBits[274] ),
    .S1(\ConfigBits[275] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst1  (.A0(net11),
    .A1(net155),
    .A2(net163),
    .A3(net206),
    .S0(\ConfigBits[274] ),
    .S1(\ConfigBits[275] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst2  (.A0(net208),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[274] ),
    .S1(\ConfigBits[275] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD0),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[274] ),
    .S1(\ConfigBits[275] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[276] ),
    .S1(\ConfigBits[277] ),
    .X(\JN2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net112),
    .A2(net144),
    .A3(net4),
    .S0(\ConfigBits[278] ),
    .S1(\ConfigBits[279] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst1  (.A0(net12),
    .A1(net156),
    .A2(net164),
    .A3(net207),
    .S0(\ConfigBits[278] ),
    .S1(\ConfigBits[279] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst2  (.A0(net209),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[278] ),
    .S1(\ConfigBits[279] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD0),
    .A2(BD1),
    .A3(BD3),
    .S0(\ConfigBits[278] ),
    .S1(\ConfigBits[279] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[280] ),
    .S1(\ConfigBits[281] ),
    .X(\JN2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst0  (.A0(net101),
    .A1(net105),
    .A2(net137),
    .A3(net1),
    .S0(\ConfigBits[282] ),
    .S1(\ConfigBits[283] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst1  (.A0(net5),
    .A1(net153),
    .A2(net157),
    .A3(net206),
    .S0(\ConfigBits[282] ),
    .S1(\ConfigBits[283] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst2  (.A0(net208),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[282] ),
    .S1(\ConfigBits[283] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD0),
    .A2(BD1),
    .A3(BD2),
    .S0(\ConfigBits[282] ),
    .S1(\ConfigBits[283] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[284] ),
    .S1(\ConfigBits[285] ),
    .X(\JN2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst0  (.A0(net106),
    .A1(net4),
    .A2(net6),
    .A3(net24),
    .S0(\ConfigBits[318] ),
    .S1(\ConfigBits[319] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst1  (.A0(net158),
    .A1(net180),
    .A2(net211),
    .A3(net238),
    .S0(\ConfigBits[318] ),
    .S1(\ConfigBits[319] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst2  (.A0(net229),
    .A1(AD1),
    .A2(AD2),
    .A3(AD3),
    .S0(\ConfigBits[318] ),
    .S1(\ConfigBits[319] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[318] ),
    .S1(\ConfigBits[319] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[320] ),
    .S1(\ConfigBits[321] ),
    .X(\JS2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst0  (.A0(net107),
    .A1(net1),
    .A2(net7),
    .A3(net21),
    .S0(\ConfigBits[322] ),
    .S1(\ConfigBits[323] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst1  (.A0(net159),
    .A1(net181),
    .A2(net212),
    .A3(net245),
    .S0(\ConfigBits[322] ),
    .S1(\ConfigBits[323] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst2  (.A0(net226),
    .A1(AD0),
    .A2(AD2),
    .A3(AD3),
    .S0(\ConfigBits[322] ),
    .S1(\ConfigBits[323] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[322] ),
    .S1(\ConfigBits[323] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[324] ),
    .S1(\ConfigBits[325] ),
    .X(\JS2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst0  (.A0(net108),
    .A1(net2),
    .A2(net8),
    .A3(net41),
    .S0(\ConfigBits[326] ),
    .S1(\ConfigBits[327] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst1  (.A0(net24),
    .A1(net160),
    .A2(net182),
    .A3(net213),
    .S0(\ConfigBits[326] ),
    .S1(\ConfigBits[327] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst2  (.A0(net229),
    .A1(AD0),
    .A2(AD1),
    .A3(AD3),
    .S0(\ConfigBits[326] ),
    .S1(\ConfigBits[327] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[326] ),
    .S1(\ConfigBits[327] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[328] ),
    .S1(\ConfigBits[329] ),
    .X(\JS2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst0  (.A0(net109),
    .A1(net3),
    .A2(net9),
    .A3(net42),
    .S0(\ConfigBits[330] ),
    .S1(\ConfigBits[331] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst1  (.A0(net21),
    .A1(net161),
    .A2(net173),
    .A3(net214),
    .S0(\ConfigBits[330] ),
    .S1(\ConfigBits[331] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst2  (.A0(net226),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[330] ),
    .S1(\ConfigBits[331] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[330] ),
    .S1(\ConfigBits[331] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[332] ),
    .S1(\ConfigBits[333] ),
    .X(\JS2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net110),
    .A2(net2),
    .A3(net10),
    .S0(\ConfigBits[334] ),
    .S1(\ConfigBits[335] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst1  (.A0(net154),
    .A1(net162),
    .A2(net198),
    .A3(net207),
    .S0(\ConfigBits[334] ),
    .S1(\ConfigBits[335] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst2  (.A0(net209),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[334] ),
    .S1(\ConfigBits[335] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[334] ),
    .S1(\ConfigBits[335] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[336] ),
    .S1(\ConfigBits[337] ),
    .X(\JS2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net111),
    .A2(net3),
    .A3(net11),
    .S0(\ConfigBits[338] ),
    .S1(\ConfigBits[339] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst1  (.A0(net155),
    .A1(net163),
    .A2(net197),
    .A3(net206),
    .S0(\ConfigBits[338] ),
    .S1(\ConfigBits[339] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst2  (.A0(net208),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[338] ),
    .S1(\ConfigBits[339] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD0),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[338] ),
    .S1(\ConfigBits[339] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[340] ),
    .S1(\ConfigBits[341] ),
    .X(\JS2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net112),
    .A2(net4),
    .A3(net12),
    .S0(\ConfigBits[342] ),
    .S1(\ConfigBits[343] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst1  (.A0(net156),
    .A1(net164),
    .A2(net196),
    .A3(net207),
    .S0(\ConfigBits[342] ),
    .S1(\ConfigBits[343] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst2  (.A0(net209),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[342] ),
    .S1(\ConfigBits[343] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD0),
    .A2(BD1),
    .A3(BD3),
    .S0(\ConfigBits[342] ),
    .S1(\ConfigBits[343] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[344] ),
    .S1(\ConfigBits[345] ),
    .X(\JS2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst0  (.A0(net101),
    .A1(net105),
    .A2(net1),
    .A3(net5),
    .S0(\ConfigBits[346] ),
    .S1(\ConfigBits[347] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst1  (.A0(net153),
    .A1(net157),
    .A2(net189),
    .A3(net206),
    .S0(\ConfigBits[346] ),
    .S1(\ConfigBits[347] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst2  (.A0(net208),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[346] ),
    .S1(\ConfigBits[347] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD0),
    .A2(BD1),
    .A3(BD2),
    .S0(\ConfigBits[346] ),
    .S1(\ConfigBits[347] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[348] ),
    .S1(\ConfigBits[349] ),
    .X(\JS2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net106),
    .A2(net6),
    .A3(net24),
    .S0(\ConfigBits[350] ),
    .S1(\ConfigBits[351] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst1  (.A0(net158),
    .A1(net180),
    .A2(net189),
    .A3(net211),
    .S0(\ConfigBits[350] ),
    .S1(\ConfigBits[351] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst2  (.A0(net229),
    .A1(AD1),
    .A2(AD2),
    .A3(AD3),
    .S0(\ConfigBits[350] ),
    .S1(\ConfigBits[351] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[350] ),
    .S1(\ConfigBits[351] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[352] ),
    .S1(\ConfigBits[353] ),
    .X(\JW2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst0  (.A0(net101),
    .A1(net107),
    .A2(net7),
    .A3(net21),
    .S0(\ConfigBits[354] ),
    .S1(\ConfigBits[355] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst1  (.A0(net159),
    .A1(net181),
    .A2(net196),
    .A3(net212),
    .S0(\ConfigBits[354] ),
    .S1(\ConfigBits[355] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst2  (.A0(net226),
    .A1(AD0),
    .A2(AD2),
    .A3(AD3),
    .S0(\ConfigBits[354] ),
    .S1(\ConfigBits[355] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[354] ),
    .S1(\ConfigBits[355] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[356] ),
    .S1(\ConfigBits[357] ),
    .X(\JW2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net108),
    .A2(net145),
    .A3(net8),
    .S0(\ConfigBits[358] ),
    .S1(\ConfigBits[359] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst1  (.A0(net24),
    .A1(net160),
    .A2(net182),
    .A3(net213),
    .S0(\ConfigBits[358] ),
    .S1(\ConfigBits[359] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst2  (.A0(net229),
    .A1(AD0),
    .A2(AD1),
    .A3(AD3),
    .S0(\ConfigBits[358] ),
    .S1(\ConfigBits[359] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[358] ),
    .S1(\ConfigBits[359] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[360] ),
    .S1(\ConfigBits[361] ),
    .X(\JW2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net109),
    .A2(net146),
    .A3(net9),
    .S0(\ConfigBits[362] ),
    .S1(\ConfigBits[363] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst1  (.A0(net21),
    .A1(net161),
    .A2(net173),
    .A3(net214),
    .S0(\ConfigBits[362] ),
    .S1(\ConfigBits[363] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst2  (.A0(net226),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[362] ),
    .S1(\ConfigBits[363] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst3  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[362] ),
    .S1(\ConfigBits[363] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[364] ),
    .S1(\ConfigBits[365] ),
    .X(\JW2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net110),
    .A2(net2),
    .A3(net10),
    .S0(\ConfigBits[366] ),
    .S1(\ConfigBits[367] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst1  (.A0(net154),
    .A1(net156),
    .A2(net162),
    .A3(net207),
    .S0(\ConfigBits[366] ),
    .S1(\ConfigBits[367] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst2  (.A0(net247),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[366] ),
    .S1(\ConfigBits[367] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[366] ),
    .S1(\ConfigBits[367] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[368] ),
    .S1(\ConfigBits[369] ),
    .X(\JW2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net111),
    .A2(net3),
    .A3(net11),
    .S0(\ConfigBits[370] ),
    .S1(\ConfigBits[371] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst1  (.A0(net153),
    .A1(net155),
    .A2(net163),
    .A3(net208),
    .S0(\ConfigBits[370] ),
    .S1(\ConfigBits[371] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst2  (.A0(net246),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[370] ),
    .S1(\ConfigBits[371] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD0),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[370] ),
    .S1(\ConfigBits[371] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[372] ),
    .S1(\ConfigBits[373] ),
    .X(\JW2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net112),
    .A2(net4),
    .A3(net12),
    .S0(\ConfigBits[374] ),
    .S1(\ConfigBits[375] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst1  (.A0(net154),
    .A1(net156),
    .A2(net164),
    .A3(net209),
    .S0(\ConfigBits[374] ),
    .S1(\ConfigBits[375] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst2  (.A0(net245),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[374] ),
    .S1(\ConfigBits[375] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD0),
    .A2(BD1),
    .A3(BD3),
    .S0(\ConfigBits[374] ),
    .S1(\ConfigBits[375] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[376] ),
    .S1(\ConfigBits[377] ),
    .X(\JW2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst0  (.A0(net101),
    .A1(net105),
    .A2(net1),
    .A3(net5),
    .S0(\ConfigBits[378] ),
    .S1(\ConfigBits[379] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst1  (.A0(net153),
    .A1(net155),
    .A2(net157),
    .A3(net206),
    .S0(\ConfigBits[378] ),
    .S1(\ConfigBits[379] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst2  (.A0(net238),
    .A1(AD0),
    .A2(AD1),
    .A3(AD2),
    .S0(\ConfigBits[378] ),
    .S1(\ConfigBits[379] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst3  (.A0(AD3),
    .A1(BD0),
    .A2(BD1),
    .A3(BD2),
    .S0(\ConfigBits[378] ),
    .S1(\ConfigBits[379] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[380] ),
    .S1(\ConfigBits[381] ),
    .X(\JW2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst0  (.A0(net144),
    .A1(net4),
    .A2(net196),
    .A3(net209),
    .S0(\ConfigBits[106] ),
    .S1(\ConfigBits[107] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst1  (.A0(AD0),
    .A1(AD1),
    .A2(AD2),
    .A3(AD3),
    .S0(\ConfigBits[106] ),
    .S1(\ConfigBits[107] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst2  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[106] ),
    .S1(\ConfigBits[107] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst3  (.A0(\J2MID_ABb_BEG[1] ),
    .A1(\J2MID_CDb_BEG[1] ),
    .A2(\J2MID_EFb_BEG[1] ),
    .A3(\J2MID_GHb_BEG[1] ),
    .S0(\ConfigBits[106] ),
    .S1(\ConfigBits[107] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[108] ),
    .S1(\ConfigBits[109] ),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst0  (.A0(net145),
    .A1(net3),
    .A2(net197),
    .A3(net208),
    .S0(\ConfigBits[110] ),
    .S1(\ConfigBits[111] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst1  (.A0(AD0),
    .A1(AD1),
    .A2(AD2),
    .A3(AD3),
    .S0(\ConfigBits[110] ),
    .S1(\ConfigBits[111] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst2  (.A0(BD0),
    .A1(BD1),
    .A2(BD2),
    .A3(BD3),
    .S0(\ConfigBits[110] ),
    .S1(\ConfigBits[111] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst3  (.A0(\J2MID_ABa_BEG[2] ),
    .A1(\J2MID_CDa_BEG[2] ),
    .A2(\J2MID_EFa_BEG[2] ),
    .A3(\J2MID_GHa_BEG[2] ),
    .S0(\ConfigBits[110] ),
    .S1(\ConfigBits[111] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst4  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ),
    .A2(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ),
    .A3(\Inst_RegFile_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[112] ),
    .S1(\ConfigBits[113] ),
    .X(net481));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_A_ADR0  (.A0(\J2MID_EFa_BEG[0] ),
    .A1(\J2MID_EFb_BEG[0] ),
    .A2(\J2END_EF_BEG[0] ),
    .A3(\J_l_EF_BEG[0] ),
    .S0(\ConfigBits[114] ),
    .S1(\ConfigBits[115] ),
    .X(A_ADR0));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_A_ADR1  (.A0(\J2MID_EFa_BEG[1] ),
    .A1(\J2MID_EFb_BEG[1] ),
    .A2(\J2END_EF_BEG[1] ),
    .A3(\J_l_EF_BEG[1] ),
    .S0(\ConfigBits[116] ),
    .S1(\ConfigBits[117] ),
    .X(A_ADR1));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_A_ADR2  (.A0(\J2MID_EFa_BEG[2] ),
    .A1(\J2MID_EFb_BEG[2] ),
    .A2(\J2END_EF_BEG[2] ),
    .A3(\J_l_EF_BEG[2] ),
    .S0(\ConfigBits[118] ),
    .S1(\ConfigBits[119] ),
    .X(A_ADR2));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_A_ADR3  (.A0(\J2MID_EFa_BEG[3] ),
    .A1(\J2MID_EFb_BEG[3] ),
    .A2(\J2END_EF_BEG[3] ),
    .A3(\J_l_EF_BEG[3] ),
    .S0(\ConfigBits[120] ),
    .S1(\ConfigBits[121] ),
    .X(A_ADR3));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_B_ADR0  (.A0(\J2MID_GHa_BEG[0] ),
    .A1(\J2MID_GHb_BEG[0] ),
    .A2(\J2END_GH_BEG[0] ),
    .A3(\J_l_GH_BEG[0] ),
    .S0(\ConfigBits[125] ),
    .S1(\ConfigBits[126] ),
    .X(B_ADR0));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_B_ADR1  (.A0(\J2MID_GHa_BEG[1] ),
    .A1(\J2MID_GHb_BEG[1] ),
    .A2(\J2END_GH_BEG[1] ),
    .A3(\J_l_GH_BEG[1] ),
    .S0(\ConfigBits[127] ),
    .S1(\ConfigBits[128] ),
    .X(B_ADR1));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_B_ADR2  (.A0(\J2MID_GHa_BEG[2] ),
    .A1(\J2MID_GHb_BEG[2] ),
    .A2(\J2END_GH_BEG[2] ),
    .A3(\J_l_GH_BEG[2] ),
    .S0(\ConfigBits[129] ),
    .S1(\ConfigBits[130] ),
    .X(B_ADR2));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_B_ADR3  (.A0(\J2MID_GHa_BEG[3] ),
    .A1(\J2MID_GHb_BEG[3] ),
    .A2(\J2END_GH_BEG[3] ),
    .A3(\J_l_GH_BEG[3] ),
    .S0(\ConfigBits[131] ),
    .S1(\ConfigBits[132] ),
    .X(B_ADR3));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_D0  (.A0(\J2MID_ABa_BEG[0] ),
    .A1(\J2MID_ABb_BEG[0] ),
    .A2(\J2END_AB_BEG[0] ),
    .A3(\J_l_AB_BEG[0] ),
    .S0(\ConfigBits[136] ),
    .S1(\ConfigBits[137] ),
    .X(D0));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_D1  (.A0(\J2MID_ABa_BEG[1] ),
    .A1(\J2MID_ABb_BEG[1] ),
    .A2(\J2END_AB_BEG[1] ),
    .A3(\J_l_AB_BEG[1] ),
    .S0(\ConfigBits[138] ),
    .S1(\ConfigBits[139] ),
    .X(D1));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_D2  (.A0(\J2MID_ABa_BEG[2] ),
    .A1(\J2MID_ABb_BEG[2] ),
    .A2(\J2END_AB_BEG[2] ),
    .A3(\J_l_AB_BEG[2] ),
    .S0(\ConfigBits[140] ),
    .S1(\ConfigBits[141] ),
    .X(D2));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_D3  (.A0(\J2MID_ABa_BEG[3] ),
    .A1(\J2MID_ABb_BEG[3] ),
    .A2(\J2END_AB_BEG[3] ),
    .A3(\J_l_AB_BEG[3] ),
    .S0(\ConfigBits[142] ),
    .S1(\ConfigBits[143] ),
    .X(D3));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_E1BEG0  (.A0(AD3),
    .A1(\J2MID_CDb_BEG[3] ),
    .A2(\JN2BEG[3] ),
    .A3(\J_l_CD_BEG[1] ),
    .S0(\ConfigBits[30] ),
    .S1(\ConfigBits[31] ),
    .X(net254));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_E1BEG1  (.A0(BD0),
    .A1(\J2MID_EFb_BEG[0] ),
    .A2(\JN2BEG[0] ),
    .A3(\J_l_EF_BEG[2] ),
    .S0(\ConfigBits[32] ),
    .S1(\ConfigBits[33] ),
    .X(net255));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_E1BEG2  (.A0(BD1),
    .A1(\J2MID_GHb_BEG[1] ),
    .A2(\JN2BEG[1] ),
    .A3(\J_l_GH_BEG[3] ),
    .S0(\ConfigBits[34] ),
    .S1(\ConfigBits[35] ),
    .X(net256));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_E1BEG3  (.A0(BD2),
    .A1(\J2MID_ABb_BEG[2] ),
    .A2(\JN2BEG[2] ),
    .A3(\J_l_AB_BEG[0] ),
    .S0(\ConfigBits[36] ),
    .S1(\ConfigBits[37] ),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG0  (.A0(net111),
    .A1(net11),
    .A2(net198),
    .A3(net216),
    .S0(\ConfigBits[222] ),
    .S1(\ConfigBits[223] ),
    .X(\J2END_AB_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG1  (.A0(net137),
    .A1(net7),
    .A2(net159),
    .A3(net212),
    .S0(\ConfigBits[224] ),
    .S1(\ConfigBits[225] ),
    .X(\J2END_AB_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG2  (.A0(net109),
    .A1(net33),
    .A2(net161),
    .A3(net214),
    .S0(\ConfigBits[226] ),
    .S1(\ConfigBits[227] ),
    .X(\J2END_AB_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG3  (.A0(net105),
    .A1(net5),
    .A2(net157),
    .A3(net247),
    .S0(\ConfigBits[228] ),
    .S1(\ConfigBits[229] ),
    .X(\J2END_AB_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG0  (.A0(net146),
    .A1(net11),
    .A2(net163),
    .A3(net216),
    .S0(\ConfigBits[230] ),
    .S1(\ConfigBits[231] ),
    .X(\J2END_CD_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG1  (.A0(net107),
    .A1(net7),
    .A2(net159),
    .A3(net246),
    .S0(\ConfigBits[232] ),
    .S1(\ConfigBits[233] ),
    .X(\J2END_CD_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG2  (.A0(net109),
    .A1(net9),
    .A2(net197),
    .A3(net214),
    .S0(\ConfigBits[234] ),
    .S1(\ConfigBits[235] ),
    .X(\J2END_CD_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG3  (.A0(net105),
    .A1(net40),
    .A2(net157),
    .A3(net210),
    .S0(\ConfigBits[236] ),
    .S1(\ConfigBits[237] ),
    .X(\J2END_CD_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG0  (.A0(net112),
    .A1(net41),
    .A2(net164),
    .A3(net217),
    .S0(\ConfigBits[238] ),
    .S1(\ConfigBits[239] ),
    .X(\J2END_EF_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG1  (.A0(net108),
    .A1(net8),
    .A2(net160),
    .A3(net245),
    .S0(\ConfigBits[240] ),
    .S1(\ConfigBits[241] ),
    .X(\J2END_EF_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG2  (.A0(net110),
    .A1(net10),
    .A2(net196),
    .A3(net215),
    .S0(\ConfigBits[242] ),
    .S1(\ConfigBits[243] ),
    .X(\J2END_EF_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG3  (.A0(net145),
    .A1(net6),
    .A2(net158),
    .A3(net211),
    .S0(\ConfigBits[244] ),
    .S1(\ConfigBits[245] ),
    .X(\J2END_EF_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG0  (.A0(net112),
    .A1(net12),
    .A2(net164),
    .A3(net238),
    .S0(\ConfigBits[246] ),
    .S1(\ConfigBits[247] ),
    .X(\J2END_GH_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG1  (.A0(net108),
    .A1(net8),
    .A2(net189),
    .A3(net213),
    .S0(\ConfigBits[248] ),
    .S1(\ConfigBits[249] ),
    .X(\J2END_GH_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG2  (.A0(net144),
    .A1(net10),
    .A2(net162),
    .A3(net215),
    .S0(\ConfigBits[250] ),
    .S1(\ConfigBits[251] ),
    .X(\J2END_GH_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG3  (.A0(net106),
    .A1(net42),
    .A2(net158),
    .A3(net211),
    .S0(\ConfigBits[252] ),
    .S1(\ConfigBits[253] ),
    .X(\J2END_GH_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG0  (.A0(net119),
    .A1(net171),
    .A2(net224),
    .A3(\JN2BEG[3] ),
    .S0(\ConfigBits[158] ),
    .S1(\ConfigBits[159] ),
    .X(\J2MID_ABa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG1  (.A0(net15),
    .A1(net167),
    .A2(net220),
    .A3(\JE2BEG[3] ),
    .S0(\ConfigBits[160] ),
    .S1(\ConfigBits[161] ),
    .X(\J2MID_ABa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG2  (.A0(net117),
    .A1(net17),
    .A2(net222),
    .A3(\JS2BEG[3] ),
    .S0(\ConfigBits[162] ),
    .S1(\ConfigBits[163] ),
    .X(\J2MID_ABa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG3  (.A0(net113),
    .A1(net13),
    .A2(net165),
    .A3(\JW2BEG[3] ),
    .S0(\ConfigBits[164] ),
    .S1(\ConfigBits[165] ),
    .X(\J2MID_ABa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG0  (.A0(net120),
    .A1(net20),
    .A2(net172),
    .A3(net225),
    .S0(\ConfigBits[190] ),
    .S1(\ConfigBits[191] ),
    .X(\J2MID_ABb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG1  (.A0(net116),
    .A1(net16),
    .A2(net168),
    .A3(net221),
    .S0(\ConfigBits[192] ),
    .S1(\ConfigBits[193] ),
    .X(\J2MID_ABb_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG2  (.A0(net118),
    .A1(net18),
    .A2(net170),
    .A3(net223),
    .S0(\ConfigBits[194] ),
    .S1(\ConfigBits[195] ),
    .X(\J2MID_ABb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG3  (.A0(net114),
    .A1(net14),
    .A2(net166),
    .A3(net219),
    .S0(\ConfigBits[196] ),
    .S1(\ConfigBits[197] ),
    .X(\J2MID_ABb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG0  (.A0(net19),
    .A1(net171),
    .A2(net224),
    .A3(\JN2BEG[4] ),
    .S0(\ConfigBits[166] ),
    .S1(\ConfigBits[167] ),
    .X(\J2MID_CDa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG1  (.A0(net115),
    .A1(net15),
    .A2(net220),
    .A3(\JE2BEG[4] ),
    .S0(\ConfigBits[168] ),
    .S1(\ConfigBits[169] ),
    .X(\J2MID_CDa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG2  (.A0(net117),
    .A1(net17),
    .A2(net169),
    .A3(\JS2BEG[4] ),
    .S0(\ConfigBits[170] ),
    .S1(\ConfigBits[171] ),
    .X(\J2MID_CDa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG3  (.A0(net113),
    .A1(net165),
    .A2(net218),
    .A3(\JW2BEG[4] ),
    .S0(\ConfigBits[172] ),
    .S1(\ConfigBits[173] ),
    .X(\J2MID_CDa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG0  (.A0(net120),
    .A1(net20),
    .A2(net172),
    .A3(net225),
    .S0(\ConfigBits[198] ),
    .S1(\ConfigBits[199] ),
    .X(\J2MID_CDb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG1  (.A0(net116),
    .A1(net16),
    .A2(net168),
    .A3(net221),
    .S0(\ConfigBits[200] ),
    .S1(\ConfigBits[201] ),
    .X(\J2MID_CDb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG2  (.A0(net118),
    .A1(net18),
    .A2(net170),
    .A3(net223),
    .S0(\ConfigBits[202] ),
    .S1(\ConfigBits[203] ),
    .X(\J2MID_CDb_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG3  (.A0(net114),
    .A1(net14),
    .A2(net166),
    .A3(net219),
    .S0(\ConfigBits[204] ),
    .S1(\ConfigBits[205] ),
    .X(\J2MID_CDb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG0  (.A0(net119),
    .A1(net19),
    .A2(net224),
    .A3(\JN2BEG[5] ),
    .S0(\ConfigBits[174] ),
    .S1(\ConfigBits[175] ),
    .X(\J2MID_EFa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG1  (.A0(net115),
    .A1(net15),
    .A2(net167),
    .A3(\JE2BEG[5] ),
    .S0(\ConfigBits[176] ),
    .S1(\ConfigBits[177] ),
    .X(\J2MID_EFa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG2  (.A0(net117),
    .A1(net169),
    .A2(net222),
    .A3(\JS2BEG[5] ),
    .S0(\ConfigBits[178] ),
    .S1(\ConfigBits[179] ),
    .X(\J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG3  (.A0(net13),
    .A1(net165),
    .A2(net218),
    .A3(\JW2BEG[5] ),
    .S0(\ConfigBits[180] ),
    .S1(\ConfigBits[181] ),
    .X(\J2MID_EFa_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG0  (.A0(net120),
    .A1(net20),
    .A2(net172),
    .A3(net225),
    .S0(\ConfigBits[206] ),
    .S1(\ConfigBits[207] ),
    .X(\J2MID_EFb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG1  (.A0(net116),
    .A1(net16),
    .A2(net168),
    .A3(net221),
    .S0(\ConfigBits[208] ),
    .S1(\ConfigBits[209] ),
    .X(\J2MID_EFb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG2  (.A0(net118),
    .A1(net18),
    .A2(net170),
    .A3(net223),
    .S0(\ConfigBits[210] ),
    .S1(\ConfigBits[211] ),
    .X(\J2MID_EFb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG3  (.A0(net114),
    .A1(net14),
    .A2(net166),
    .A3(net219),
    .S0(\ConfigBits[212] ),
    .S1(\ConfigBits[213] ),
    .X(\J2MID_EFb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG0  (.A0(net119),
    .A1(net19),
    .A2(net171),
    .A3(\JN2BEG[6] ),
    .S0(\ConfigBits[182] ),
    .S1(\ConfigBits[183] ),
    .X(\J2MID_GHa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG1  (.A0(net115),
    .A1(net167),
    .A2(net220),
    .A3(\JE2BEG[6] ),
    .S0(\ConfigBits[184] ),
    .S1(\ConfigBits[185] ),
    .X(\J2MID_GHa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG2  (.A0(net17),
    .A1(net169),
    .A2(net222),
    .A3(\JS2BEG[6] ),
    .S0(\ConfigBits[186] ),
    .S1(\ConfigBits[187] ),
    .X(\J2MID_GHa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG3  (.A0(net113),
    .A1(net13),
    .A2(net218),
    .A3(\JW2BEG[6] ),
    .S0(\ConfigBits[188] ),
    .S1(\ConfigBits[189] ),
    .X(\J2MID_GHa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG0  (.A0(net120),
    .A1(net20),
    .A2(net172),
    .A3(net225),
    .S0(\ConfigBits[214] ),
    .S1(\ConfigBits[215] ),
    .X(\J2MID_GHb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG1  (.A0(net116),
    .A1(net16),
    .A2(net168),
    .A3(net221),
    .S0(\ConfigBits[216] ),
    .S1(\ConfigBits[217] ),
    .X(\J2MID_GHb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG2  (.A0(net118),
    .A1(net18),
    .A2(net170),
    .A3(net223),
    .S0(\ConfigBits[218] ),
    .S1(\ConfigBits[219] ),
    .X(\J2MID_GHb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG3  (.A0(net114),
    .A1(net14),
    .A2(net166),
    .A3(net219),
    .S0(\ConfigBits[220] ),
    .S1(\ConfigBits[221] ),
    .X(\J2MID_GHb_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG0  (.A0(net146),
    .A1(net182),
    .A2(net238),
    .A3(\JN2BEG[1] ),
    .S0(\ConfigBits[382] ),
    .S1(\ConfigBits[383] ),
    .X(\J_l_AB_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG1  (.A0(net41),
    .A1(net181),
    .A2(net217),
    .A3(\JE2BEG[1] ),
    .S0(\ConfigBits[384] ),
    .S1(\ConfigBits[385] ),
    .X(\J_l_AB_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG2  (.A0(net128),
    .A1(net24),
    .A2(net229),
    .A3(\JS2BEG[1] ),
    .S0(\ConfigBits[386] ),
    .S1(\ConfigBits[387] ),
    .X(\J_l_AB_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG3  (.A0(net121),
    .A1(net21),
    .A2(net173),
    .A3(\JW2BEG[1] ),
    .S0(\ConfigBits[388] ),
    .S1(\ConfigBits[389] ),
    .X(\J_l_AB_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG0  (.A0(net8),
    .A1(net198),
    .A2(net246),
    .A3(\JN2BEG[2] ),
    .S0(\ConfigBits[390] ),
    .S1(\ConfigBits[391] ),
    .X(\J_l_CD_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG1  (.A0(net129),
    .A1(net7),
    .A2(net217),
    .A3(\JE2BEG[2] ),
    .S0(\ConfigBits[392] ),
    .S1(\ConfigBits[393] ),
    .X(\J_l_CD_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG2  (.A0(net144),
    .A1(net40),
    .A2(net180),
    .A3(\JS2BEG[2] ),
    .S0(\ConfigBits[394] ),
    .S1(\ConfigBits[395] ),
    .X(\J_l_CD_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG3  (.A0(net121),
    .A1(net189),
    .A2(net226),
    .A3(\JW2BEG[2] ),
    .S0(\ConfigBits[396] ),
    .S1(\ConfigBits[397] ),
    .X(\J_l_CD_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG0  (.A0(net130),
    .A1(net8),
    .A2(net213),
    .A3(\JN2BEG[3] ),
    .S0(\ConfigBits[398] ),
    .S1(\ConfigBits[399] ),
    .X(\J_l_EF_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG1  (.A0(net145),
    .A1(net7),
    .A2(net181),
    .A3(\JE2BEG[3] ),
    .S0(\ConfigBits[400] ),
    .S1(\ConfigBits[401] ),
    .X(\J_l_EF_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG2  (.A0(net128),
    .A1(net196),
    .A2(net214),
    .A3(\JS2BEG[3] ),
    .S0(\ConfigBits[402] ),
    .S1(\ConfigBits[403] ),
    .X(\J_l_EF_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG3  (.A0(net42),
    .A1(net173),
    .A2(net245),
    .A3(\JW2BEG[3] ),
    .S0(\ConfigBits[404] ),
    .S1(\ConfigBits[405] ),
    .X(\J_l_EF_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG0  (.A0(net130),
    .A1(net33),
    .A2(net182),
    .A3(\JN2BEG[4] ),
    .S0(\ConfigBits[406] ),
    .S1(\ConfigBits[407] ),
    .X(\J_l_GH_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG1  (.A0(net129),
    .A1(net197),
    .A2(net212),
    .A3(\JE2BEG[4] ),
    .S0(\ConfigBits[408] ),
    .S1(\ConfigBits[409] ),
    .X(\J_l_GH_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG2  (.A0(net24),
    .A1(net180),
    .A2(net247),
    .A3(\JS2BEG[4] ),
    .S0(\ConfigBits[410] ),
    .S1(\ConfigBits[411] ),
    .X(\J_l_GH_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG3  (.A0(net137),
    .A1(net21),
    .A2(net210),
    .A3(\JW2BEG[4] ),
    .S0(\ConfigBits[412] ),
    .S1(\ConfigBits[413] ),
    .X(\J_l_GH_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_N1BEG0  (.A0(AD2),
    .A1(\J2MID_CDb_BEG[3] ),
    .A2(\JW2BEG[3] ),
    .A3(\J_l_CD_BEG[1] ),
    .S0(\ConfigBits[2] ),
    .S1(\ConfigBits[3] ),
    .X(net354));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_N1BEG1  (.A0(AD3),
    .A1(\J2MID_EFb_BEG[0] ),
    .A2(\JW2BEG[0] ),
    .A3(\J_l_EF_BEG[2] ),
    .S0(\ConfigBits[4] ),
    .S1(\ConfigBits[5] ),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_N1BEG2  (.A0(BD0),
    .A1(\J2MID_GHb_BEG[1] ),
    .A2(\JW2BEG[1] ),
    .A3(\J_l_GH_BEG[3] ),
    .S0(\ConfigBits[6] ),
    .S1(\ConfigBits[7] ),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_N1BEG3  (.A0(BD1),
    .A1(\J2MID_ABb_BEG[2] ),
    .A2(\JW2BEG[2] ),
    .A3(\J_l_AB_BEG[0] ),
    .S0(\ConfigBits[8] ),
    .S1(\ConfigBits[9] ),
    .X(net357));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_N4BEG0  (.A0(net107),
    .A1(net128),
    .A2(net24),
    .A3(BD0),
    .S0(\ConfigBits[10] ),
    .S1(\ConfigBits[11] ),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_N4BEG1  (.A0(net108),
    .A1(net129),
    .A2(net21),
    .A3(BD1),
    .S0(\ConfigBits[12] ),
    .S1(\ConfigBits[13] ),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_N4BEG2  (.A0(net105),
    .A1(net130),
    .A2(net229),
    .A3(BD2),
    .S0(\ConfigBits[14] ),
    .S1(\ConfigBits[15] ),
    .X(net379));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_N4BEG3  (.A0(net106),
    .A1(net121),
    .A2(net226),
    .A3(BD3),
    .S0(\ConfigBits[16] ),
    .S1(\ConfigBits[17] ),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_S1BEG0  (.A0(BD0),
    .A1(\J2MID_CDb_BEG[3] ),
    .A2(\JE2BEG[3] ),
    .A3(\J_l_CD_BEG[1] ),
    .S0(\ConfigBits[58] ),
    .S1(\ConfigBits[59] ),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_S1BEG1  (.A0(BD1),
    .A1(\J2MID_EFb_BEG[0] ),
    .A2(\JE2BEG[0] ),
    .A3(\J_l_EF_BEG[2] ),
    .S0(\ConfigBits[60] ),
    .S1(\ConfigBits[61] ),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_S1BEG2  (.A0(BD2),
    .A1(\J2MID_GHb_BEG[1] ),
    .A2(\JE2BEG[1] ),
    .A3(\J_l_GH_BEG[3] ),
    .S0(\ConfigBits[62] ),
    .S1(\ConfigBits[63] ),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_S1BEG3  (.A0(BD3),
    .A1(\J2MID_ABb_BEG[2] ),
    .A2(\JE2BEG[2] ),
    .A3(\J_l_AB_BEG[0] ),
    .S0(\ConfigBits[64] ),
    .S1(\ConfigBits[65] ),
    .X(net409));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_S4BEG0  (.A0(net24),
    .A1(net159),
    .A2(net180),
    .A3(AD0),
    .S0(\ConfigBits[66] ),
    .S1(\ConfigBits[67] ),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_S4BEG1  (.A0(net21),
    .A1(net160),
    .A2(net181),
    .A3(AD1),
    .S0(\ConfigBits[68] ),
    .S1(\ConfigBits[69] ),
    .X(net430));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_S4BEG2  (.A0(net157),
    .A1(net182),
    .A2(net229),
    .A3(AD2),
    .S0(\ConfigBits[70] ),
    .S1(\ConfigBits[71] ),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_S4BEG3  (.A0(net158),
    .A1(net173),
    .A2(net226),
    .A3(AD3),
    .S0(\ConfigBits[72] ),
    .S1(\ConfigBits[73] ),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_W1BEG0  (.A0(BD1),
    .A1(\J2MID_CDb_BEG[3] ),
    .A2(\JS2BEG[3] ),
    .A3(\J_l_CD_BEG[1] ),
    .S0(\ConfigBits[86] ),
    .S1(\ConfigBits[87] ),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_W1BEG1  (.A0(BD2),
    .A1(\J2MID_EFb_BEG[0] ),
    .A2(\JS2BEG[0] ),
    .A3(\J_l_EF_BEG[2] ),
    .S0(\ConfigBits[88] ),
    .S1(\ConfigBits[89] ),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_W1BEG2  (.A0(BD3),
    .A1(\J2MID_GHb_BEG[1] ),
    .A2(\JS2BEG[1] ),
    .A3(\J_l_GH_BEG[3] ),
    .S0(\ConfigBits[90] ),
    .S1(\ConfigBits[91] ),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_W1BEG3  (.A0(AD0),
    .A1(\J2MID_ABb_BEG[2] ),
    .A2(\JS2BEG[2] ),
    .A3(\J_l_AB_BEG[0] ),
    .S0(\ConfigBits[92] ),
    .S1(\ConfigBits[93] ),
    .X(net462));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_W_ADR0  (.A0(\J2MID_CDa_BEG[0] ),
    .A1(\J2MID_CDb_BEG[0] ),
    .A2(\J2END_CD_BEG[0] ),
    .A3(\J_l_CD_BEG[0] ),
    .S0(\ConfigBits[144] ),
    .S1(\ConfigBits[145] ),
    .X(W_ADR0));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_W_ADR1  (.A0(\J2MID_CDa_BEG[1] ),
    .A1(\J2MID_CDb_BEG[1] ),
    .A2(\J2END_CD_BEG[1] ),
    .A3(\J_l_CD_BEG[1] ),
    .S0(\ConfigBits[146] ),
    .S1(\ConfigBits[147] ),
    .X(W_ADR1));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_W_ADR2  (.A0(\J2MID_CDa_BEG[2] ),
    .A1(\J2MID_CDb_BEG[2] ),
    .A2(\J2END_CD_BEG[2] ),
    .A3(\J_l_CD_BEG[2] ),
    .S0(\ConfigBits[148] ),
    .S1(\ConfigBits[149] ),
    .X(W_ADR2));
 sky130_fd_sc_hd__mux4_2 \Inst_RegFile_switch_matrix/inst_cus_mux41_buf_W_ADR3  (.A0(\J2MID_CDa_BEG[3] ),
    .A1(\J2MID_CDb_BEG[3] ),
    .A2(\J2END_CD_BEG[3] ),
    .A3(\J_l_CD_BEG[3] ),
    .S0(\ConfigBits[150] ),
    .S1(\ConfigBits[151] ),
    .X(W_ADR3));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/cus_mux41_buf_inst0  (.A0(net106),
    .A1(net158),
    .A2(\J2MID_GHa_BEG[1] ),
    .A3(\J2MID_GHb_BEG[2] ),
    .S0(\ConfigBits[122] ),
    .S1(\ConfigBits[123] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/cus_mux41_buf_inst1  (.A0(\J2END_CD_BEG[3] ),
    .A1(\JN2BEG[5] ),
    .A2(\JS2BEG[5] ),
    .A3(\JW2BEG[5] ),
    .S0(\ConfigBits[122] ),
    .S1(\ConfigBits[123] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/cus_mux41_buf_out1 ),
    .S(\ConfigBits[124] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_A_ADR4/my_mux2_inst/_0_ ),
    .X(A_ADR4));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/cus_mux41_buf_inst0  (.A0(net107),
    .A1(net159),
    .A2(\J2MID_ABa_BEG[1] ),
    .A3(\J2MID_ABb_BEG[2] ),
    .S0(\ConfigBits[133] ),
    .S1(\ConfigBits[134] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/cus_mux41_buf_inst1  (.A0(\J2END_EF_BEG[3] ),
    .A1(\JN2BEG[6] ),
    .A2(\JS2BEG[6] ),
    .A3(\JW2BEG[6] ),
    .S0(\ConfigBits[133] ),
    .S1(\ConfigBits[134] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/cus_mux41_buf_out1 ),
    .S(\ConfigBits[135] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_B_ADR4/my_mux2_inst/_0_ ),
    .X(B_ADR4));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net3),
    .A2(net155),
    .A3(AD1),
    .S0(\ConfigBits[38] ),
    .S1(\ConfigBits[39] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst1  (.A0(BD1),
    .A1(\J2MID_ABb_BEG[1] ),
    .A2(\J2MID_CDb_BEG[1] ),
    .A3(\J2END_GH_BEG[0] ),
    .S0(\ConfigBits[38] ),
    .S1(\ConfigBits[39] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ),
    .S(\ConfigBits[40] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net4),
    .A2(net156),
    .A3(AD2),
    .S0(\ConfigBits[41] ),
    .S1(\ConfigBits[42] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst1  (.A0(BD2),
    .A1(\J2MID_ABa_BEG[2] ),
    .A2(\J2MID_CDa_BEG[2] ),
    .A3(\J2END_EF_BEG[0] ),
    .S0(\ConfigBits[41] ),
    .S1(\ConfigBits[42] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ),
    .S(\ConfigBits[43] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst0  (.A0(net101),
    .A1(net1),
    .A2(net153),
    .A3(AD3),
    .S0(\ConfigBits[44] ),
    .S1(\ConfigBits[45] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst1  (.A0(BD3),
    .A1(\J2MID_EFb_BEG[1] ),
    .A2(\J2MID_GHb_BEG[1] ),
    .A3(\J2END_CD_BEG[0] ),
    .S0(\ConfigBits[44] ),
    .S1(\ConfigBits[45] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ),
    .S(\ConfigBits[46] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net2),
    .A2(net154),
    .A3(AD0),
    .S0(\ConfigBits[47] ),
    .S1(\ConfigBits[48] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst1  (.A0(BD0),
    .A1(\J2MID_EFa_BEG[2] ),
    .A2(\J2MID_GHa_BEG[2] ),
    .A3(\J2END_AB_BEG[0] ),
    .S0(\ConfigBits[47] ),
    .S1(\ConfigBits[48] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ),
    .S(\ConfigBits[49] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net3),
    .A2(net208),
    .A3(AD1),
    .S0(\ConfigBits[18] ),
    .S1(\ConfigBits[19] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst1  (.A0(BD1),
    .A1(\J2MID_ABb_BEG[1] ),
    .A2(\J2MID_CDb_BEG[1] ),
    .A3(\J2END_GH_BEG[1] ),
    .S0(\ConfigBits[18] ),
    .S1(\ConfigBits[19] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ),
    .S(\ConfigBits[20] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net4),
    .A2(net209),
    .A3(AD2),
    .S0(\ConfigBits[21] ),
    .S1(\ConfigBits[22] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst1  (.A0(BD2),
    .A1(\J2MID_ABa_BEG[2] ),
    .A2(\J2MID_CDa_BEG[2] ),
    .A3(\J2END_EF_BEG[1] ),
    .S0(\ConfigBits[21] ),
    .S1(\ConfigBits[22] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ),
    .S(\ConfigBits[23] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst0  (.A0(net101),
    .A1(net1),
    .A2(net206),
    .A3(AD3),
    .S0(\ConfigBits[24] ),
    .S1(\ConfigBits[25] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst1  (.A0(BD3),
    .A1(\J2MID_EFb_BEG[1] ),
    .A2(\J2MID_GHb_BEG[1] ),
    .A3(\J2END_CD_BEG[1] ),
    .S0(\ConfigBits[24] ),
    .S1(\ConfigBits[25] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ),
    .S(\ConfigBits[26] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net2),
    .A2(net207),
    .A3(AD0),
    .S0(\ConfigBits[27] ),
    .S1(\ConfigBits[28] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst1  (.A0(BD0),
    .A1(\J2MID_EFa_BEG[2] ),
    .A2(\J2MID_GHa_BEG[2] ),
    .A3(\J2END_AB_BEG[1] ),
    .S0(\ConfigBits[27] ),
    .S1(\ConfigBits[28] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ),
    .S(\ConfigBits[29] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net3),
    .A2(net208),
    .A3(AD1),
    .S0(\ConfigBits[74] ),
    .S1(\ConfigBits[75] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst1  (.A0(BD1),
    .A1(\J2MID_ABb_BEG[1] ),
    .A2(\J2MID_CDb_BEG[1] ),
    .A3(\J2END_GH_BEG[3] ),
    .S0(\ConfigBits[74] ),
    .S1(\ConfigBits[75] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ),
    .S(\ConfigBits[76] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ),
    .X(net445));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net4),
    .A2(net209),
    .A3(AD2),
    .S0(\ConfigBits[77] ),
    .S1(\ConfigBits[78] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst1  (.A0(BD2),
    .A1(\J2MID_ABa_BEG[2] ),
    .A2(\J2MID_CDa_BEG[2] ),
    .A3(\J2END_EF_BEG[3] ),
    .S0(\ConfigBits[77] ),
    .S1(\ConfigBits[78] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ),
    .S(\ConfigBits[79] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst0  (.A0(net101),
    .A1(net1),
    .A2(net206),
    .A3(AD3),
    .S0(\ConfigBits[80] ),
    .S1(\ConfigBits[81] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst1  (.A0(BD3),
    .A1(\J2MID_EFb_BEG[1] ),
    .A2(\J2MID_GHb_BEG[1] ),
    .A3(\J2END_CD_BEG[3] ),
    .S0(\ConfigBits[80] ),
    .S1(\ConfigBits[81] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ),
    .S(\ConfigBits[82] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ),
    .X(net447));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net2),
    .A2(net207),
    .A3(AD0),
    .S0(\ConfigBits[83] ),
    .S1(\ConfigBits[84] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst1  (.A0(BD0),
    .A1(\J2MID_EFa_BEG[2] ),
    .A2(\J2MID_GHa_BEG[2] ),
    .A3(\J2END_AB_BEG[3] ),
    .S0(\ConfigBits[83] ),
    .S1(\ConfigBits[84] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ),
    .S(\ConfigBits[85] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ),
    .X(net448));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net155),
    .A2(net208),
    .A3(AD1),
    .S0(\ConfigBits[94] ),
    .S1(\ConfigBits[95] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst1  (.A0(BD1),
    .A1(\J2MID_ABb_BEG[1] ),
    .A2(\J2MID_CDb_BEG[1] ),
    .A3(\J2END_GH_BEG[2] ),
    .S0(\ConfigBits[94] ),
    .S1(\ConfigBits[95] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ),
    .S(\ConfigBits[96] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net156),
    .A2(net209),
    .A3(AD2),
    .S0(\ConfigBits[97] ),
    .S1(\ConfigBits[98] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst1  (.A0(BD2),
    .A1(\J2MID_ABa_BEG[2] ),
    .A2(\J2MID_CDa_BEG[2] ),
    .A3(\J2END_EF_BEG[2] ),
    .S0(\ConfigBits[97] ),
    .S1(\ConfigBits[98] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ),
    .S(\ConfigBits[99] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst0  (.A0(net101),
    .A1(net153),
    .A2(net206),
    .A3(AD3),
    .S0(\ConfigBits[100] ),
    .S1(\ConfigBits[101] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst1  (.A0(BD3),
    .A1(\J2MID_EFb_BEG[1] ),
    .A2(\J2MID_GHb_BEG[1] ),
    .A3(\J2END_CD_BEG[2] ),
    .S0(\ConfigBits[100] ),
    .S1(\ConfigBits[101] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ),
    .S(\ConfigBits[102] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net154),
    .A2(net207),
    .A3(AD0),
    .S0(\ConfigBits[103] ),
    .S1(\ConfigBits[104] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst1  (.A0(BD0),
    .A1(\J2MID_EFa_BEG[2] ),
    .A2(\J2MID_GHa_BEG[2] ),
    .A3(\J2END_AB_BEG[2] ),
    .S0(\ConfigBits[103] ),
    .S1(\ConfigBits[104] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ),
    .S(\ConfigBits[105] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/cus_mux41_buf_inst0  (.A0(net105),
    .A1(net157),
    .A2(\J2MID_EFa_BEG[1] ),
    .A3(\J2MID_EFb_BEG[2] ),
    .S0(\ConfigBits[152] ),
    .S1(\ConfigBits[153] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/cus_mux41_buf_inst1  (.A0(\J2END_AB_BEG[3] ),
    .A1(\JN2BEG[7] ),
    .A2(\JS2BEG[7] ),
    .A3(\JW2BEG[7] ),
    .S0(\ConfigBits[152] ),
    .S1(\ConfigBits[153] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/cus_mux41_buf_out1 ),
    .S(\ConfigBits[154] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__buf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_ADR4/my_mux2_inst/_0_ ),
    .X(W_ADR4));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/cus_mux41_buf_inst0  (.A0(net108),
    .A1(net160),
    .A2(\J2MID_CDa_BEG[1] ),
    .A3(\J2MID_CDb_BEG[2] ),
    .S0(\ConfigBits[155] ),
    .S1(\ConfigBits[156] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/cus_mux41_buf_inst1  (.A0(\J2END_GH_BEG[3] ),
    .A1(\JN2BEG[0] ),
    .A2(\JS2BEG[0] ),
    .A3(\JW2BEG[0] ),
    .S0(\ConfigBits[155] ),
    .S1(\ConfigBits[156] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/my_mux2_inst/_1_  (.A0(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/cus_mux41_buf_out0 ),
    .A1(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/cus_mux41_buf_out1 ),
    .S(\ConfigBits[157] ),
    .X(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/my_mux2_inst/_2_  (.A(\Inst_RegFile_switch_matrix/inst_cus_mux81_buf_W_en/my_mux2_inst/_0_ ),
    .X(W_en));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_0/_0_  (.A(\N4BEG_i[0] ),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_1/_0_  (.A(\N4BEG_i[1] ),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_10/_0_  (.A(\N4BEG_i[10] ),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_11/_0_  (.A(\N4BEG_i[11] ),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_2/_0_  (.A(\N4BEG_i[2] ),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_3/_0_  (.A(\N4BEG_i[3] ),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_4/_0_  (.A(\N4BEG_i[4] ),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_5/_0_  (.A(\N4BEG_i[5] ),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_6/_0_  (.A(\N4BEG_i[6] ),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_7/_0_  (.A(\N4BEG_i[7] ),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_8/_0_  (.A(\N4BEG_i[8] ),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_9/_0_  (.A(\N4BEG_i[9] ),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_0/_0_  (.A(net131),
    .X(\N4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_1/_0_  (.A(net132),
    .X(\N4BEG_i[1] ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_10/_0_  (.A(net126),
    .X(\N4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_11/_0_  (.A(net127),
    .X(\N4BEG_i[11] ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_2/_0_  (.A(net133),
    .X(\N4BEG_i[2] ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_3/_0_  (.A(net134),
    .X(\N4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_4 \N4END_inbuf_4/_0_  (.A(net135),
    .X(\N4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_5/_0_  (.A(net136),
    .X(\N4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_6/_0_  (.A(net122),
    .X(\N4BEG_i[6] ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_7/_0_  (.A(net123),
    .X(\N4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_8/_0_  (.A(net124),
    .X(\N4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_9/_0_  (.A(net125),
    .X(\N4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_0/_0_  (.A(\NN4BEG_i[0] ),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_1/_0_  (.A(\NN4BEG_i[1] ),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_10/_0_  (.A(\NN4BEG_i[10] ),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_11/_0_  (.A(\NN4BEG_i[11] ),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_2/_0_  (.A(\NN4BEG_i[2] ),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_3/_0_  (.A(\NN4BEG_i[3] ),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_4/_0_  (.A(\NN4BEG_i[4] ),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_5/_0_  (.A(\NN4BEG_i[5] ),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_6/_0_  (.A(\NN4BEG_i[6] ),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_7/_0_  (.A(\NN4BEG_i[7] ),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_8/_0_  (.A(\NN4BEG_i[8] ),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_9/_0_  (.A(\NN4BEG_i[9] ),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_0/_0_  (.A(net147),
    .X(\NN4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_1/_0_  (.A(net148),
    .X(\NN4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_10/_0_  (.A(net142),
    .X(\NN4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_4 \NN4END_inbuf_11/_0_  (.A(net143),
    .X(\NN4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_2/_0_  (.A(net149),
    .X(\NN4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_3/_0_  (.A(net150),
    .X(\NN4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_4/_0_  (.A(net151),
    .X(\NN4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_5/_0_  (.A(net152),
    .X(\NN4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_6/_0_  (.A(net138),
    .X(\NN4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_7/_0_  (.A(net139),
    .X(\NN4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_8/_0_  (.A(net140),
    .X(\NN4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_9/_0_  (.A(net141),
    .X(\NN4BEG_i[9] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_0/_0_  (.A(\S4BEG_i[0] ),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_1/_0_  (.A(\S4BEG_i[1] ),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_10/_0_  (.A(\S4BEG_i[10] ),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_11/_0_  (.A(\S4BEG_i[11] ),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_2/_0_  (.A(\S4BEG_i[2] ),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_3/_0_  (.A(\S4BEG_i[3] ),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_4/_0_  (.A(\S4BEG_i[4] ),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_5/_0_  (.A(\S4BEG_i[5] ),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_6/_0_  (.A(\S4BEG_i[6] ),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_7/_0_  (.A(\S4BEG_i[7] ),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_8/_0_  (.A(\S4BEG_i[8] ),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_9/_0_  (.A(\S4BEG_i[9] ),
    .X(net441));
 sky130_fd_sc_hd__buf_2 \S4END_inbuf_0/_0_  (.A(net183),
    .X(\S4BEG_i[0] ));
 sky130_fd_sc_hd__buf_2 \S4END_inbuf_1/_0_  (.A(net184),
    .X(\S4BEG_i[1] ));
 sky130_fd_sc_hd__buf_2 \S4END_inbuf_10/_0_  (.A(net178),
    .X(\S4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_11/_0_  (.A(net179),
    .X(\S4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_2/_0_  (.A(net185),
    .X(\S4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_3/_0_  (.A(net186),
    .X(\S4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_4/_0_  (.A(net187),
    .X(\S4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_5/_0_  (.A(net188),
    .X(\S4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_6/_0_  (.A(net174),
    .X(\S4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_7/_0_  (.A(net175),
    .X(\S4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_8/_0_  (.A(net176),
    .X(\S4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_9/_0_  (.A(net177),
    .X(\S4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_0/_0_  (.A(\SS4BEG_i[0] ),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_1/_0_  (.A(\SS4BEG_i[1] ),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_10/_0_  (.A(\SS4BEG_i[10] ),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_11/_0_  (.A(\SS4BEG_i[11] ),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_2/_0_  (.A(\SS4BEG_i[2] ),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_3/_0_  (.A(\SS4BEG_i[3] ),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_4/_0_  (.A(\SS4BEG_i[4] ),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_5/_0_  (.A(\SS4BEG_i[5] ),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_6/_0_  (.A(\SS4BEG_i[6] ),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_7/_0_  (.A(\SS4BEG_i[7] ),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_8/_0_  (.A(\SS4BEG_i[8] ),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_9/_0_  (.A(\SS4BEG_i[9] ),
    .X(net457));
 sky130_fd_sc_hd__buf_2 \SS4END_inbuf_0/_0_  (.A(net199),
    .X(\SS4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_1/_0_  (.A(net200),
    .X(\SS4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_10/_0_  (.A(net194),
    .X(\SS4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_11/_0_  (.A(net195),
    .X(\SS4BEG_i[11] ));
 sky130_fd_sc_hd__buf_2 \SS4END_inbuf_2/_0_  (.A(net201),
    .X(\SS4BEG_i[2] ));
 sky130_fd_sc_hd__buf_2 \SS4END_inbuf_3/_0_  (.A(net202),
    .X(\SS4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_4/_0_  (.A(net203),
    .X(\SS4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_5/_0_  (.A(net204),
    .X(\SS4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_6/_0_  (.A(net190),
    .X(\SS4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_7/_0_  (.A(net191),
    .X(\SS4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_8/_0_  (.A(net192),
    .X(\SS4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_9/_0_  (.A(net193),
    .X(\SS4BEG_i[9] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_0/_0_  (.A(\W6BEG_i[0] ),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_1/_0_  (.A(\W6BEG_i[1] ),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_2/_0_  (.A(\W6BEG_i[2] ),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_3/_0_  (.A(\W6BEG_i[3] ),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_4/_0_  (.A(\W6BEG_i[4] ),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_5/_0_  (.A(\W6BEG_i[5] ),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_6/_0_  (.A(\W6BEG_i[6] ),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_7/_0_  (.A(\W6BEG_i[7] ),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_8/_0_  (.A(\W6BEG_i[8] ),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_9/_0_  (.A(\W6BEG_i[9] ),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_0/_0_  (.A(net230),
    .X(\W6BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_1/_0_  (.A(net231),
    .X(\W6BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_2/_0_  (.A(net232),
    .X(\W6BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_3/_0_  (.A(net233),
    .X(\W6BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_4/_0_  (.A(net234),
    .X(\W6BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_5/_0_  (.A(net235),
    .X(\W6BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_6/_0_  (.A(net236),
    .X(\W6BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_7/_0_  (.A(net237),
    .X(\W6BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_8/_0_  (.A(net227),
    .X(\W6BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_9/_0_  (.A(net228),
    .X(\W6BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_0/_0_  (.A(\WW4BEG_i[0] ),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_1/_0_  (.A(\WW4BEG_i[1] ),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_10/_0_  (.A(\WW4BEG_i[10] ),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_11/_0_  (.A(\WW4BEG_i[11] ),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_2/_0_  (.A(\WW4BEG_i[2] ),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_3/_0_  (.A(\WW4BEG_i[3] ),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_4/_0_  (.A(\WW4BEG_i[4] ),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_5/_0_  (.A(\WW4BEG_i[5] ),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_6/_0_  (.A(\WW4BEG_i[6] ),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_7/_0_  (.A(\WW4BEG_i[7] ),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_8/_0_  (.A(\WW4BEG_i[8] ),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_9/_0_  (.A(\WW4BEG_i[9] ),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_0/_0_  (.A(net248),
    .X(\WW4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_1/_0_  (.A(net249),
    .X(\WW4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_10/_0_  (.A(net243),
    .X(\WW4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_11/_0_  (.A(net244),
    .X(\WW4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_2/_0_  (.A(net250),
    .X(\WW4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_3/_0_  (.A(net251),
    .X(\WW4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_4/_0_  (.A(net252),
    .X(\WW4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_5/_0_  (.A(net253),
    .X(\WW4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_6/_0_  (.A(net239),
    .X(\WW4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_7/_0_  (.A(net240),
    .X(\WW4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_8/_0_  (.A(net241),
    .X(\WW4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_9/_0_  (.A(net242),
    .X(\WW4BEG_i[9] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_0/_0_  (.A(net49),
    .X(\FrameData_O_i[0] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_1/_0_  (.A(net60),
    .X(\FrameData_O_i[1] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_10/_0_  (.A(net50),
    .X(\FrameData_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_11/_0_  (.A(net51),
    .X(\FrameData_O_i[11] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_12/_0_  (.A(net52),
    .X(\FrameData_O_i[12] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_13/_0_  (.A(net53),
    .X(\FrameData_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_14/_0_  (.A(net54),
    .X(\FrameData_O_i[14] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_15/_0_  (.A(net55),
    .X(\FrameData_O_i[15] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_16/_0_  (.A(net56),
    .X(\FrameData_O_i[16] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_17/_0_  (.A(net57),
    .X(\FrameData_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_18/_0_  (.A(net58),
    .X(\FrameData_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_19/_0_  (.A(net59),
    .X(\FrameData_O_i[19] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_2/_0_  (.A(net71),
    .X(\FrameData_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_20/_0_  (.A(net61),
    .X(\FrameData_O_i[20] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_21/_0_  (.A(net62),
    .X(\FrameData_O_i[21] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_22/_0_  (.A(net63),
    .X(\FrameData_O_i[22] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_23/_0_  (.A(net64),
    .X(\FrameData_O_i[23] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_24/_0_  (.A(net65),
    .X(\FrameData_O_i[24] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_25/_0_  (.A(net66),
    .X(\FrameData_O_i[25] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_26/_0_  (.A(net67),
    .X(\FrameData_O_i[26] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_27/_0_  (.A(net68),
    .X(\FrameData_O_i[27] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_28/_0_  (.A(net69),
    .X(\FrameData_O_i[28] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_29/_0_  (.A(net70),
    .X(\FrameData_O_i[29] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_3/_0_  (.A(net74),
    .X(\FrameData_O_i[3] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_30/_0_  (.A(net72),
    .X(\FrameData_O_i[30] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_31/_0_  (.A(net73),
    .X(\FrameData_O_i[31] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_4/_0_  (.A(net75),
    .X(\FrameData_O_i[4] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_5/_0_  (.A(net76),
    .X(\FrameData_O_i[5] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_6/_0_  (.A(net77),
    .X(\FrameData_O_i[6] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_7/_0_  (.A(net78),
    .X(\FrameData_O_i[7] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_8/_0_  (.A(net79),
    .X(\FrameData_O_i[8] ));
 sky130_fd_sc_hd__buf_1 \data_inbuf_9/_0_  (.A(net80),
    .X(\FrameData_O_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_0/_0_  (.A(\FrameData_O_i[0] ),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_1/_0_  (.A(\FrameData_O_i[1] ),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_10/_0_  (.A(\FrameData_O_i[10] ),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_11/_0_  (.A(\FrameData_O_i[11] ),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_12/_0_  (.A(\FrameData_O_i[12] ),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_13/_0_  (.A(\FrameData_O_i[13] ),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_14/_0_  (.A(\FrameData_O_i[14] ),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_15/_0_  (.A(\FrameData_O_i[15] ),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_16/_0_  (.A(\FrameData_O_i[16] ),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_17/_0_  (.A(\FrameData_O_i[17] ),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_18/_0_  (.A(\FrameData_O_i[18] ),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_19/_0_  (.A(\FrameData_O_i[19] ),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_2/_0_  (.A(\FrameData_O_i[2] ),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_20/_0_  (.A(\FrameData_O_i[20] ),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_21/_0_  (.A(\FrameData_O_i[21] ),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_22/_0_  (.A(\FrameData_O_i[22] ),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_23/_0_  (.A(\FrameData_O_i[23] ),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_24/_0_  (.A(\FrameData_O_i[24] ),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_25/_0_  (.A(\FrameData_O_i[25] ),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_26/_0_  (.A(\FrameData_O_i[26] ),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_27/_0_  (.A(\FrameData_O_i[27] ),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_28/_0_  (.A(\FrameData_O_i[28] ),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_29/_0_  (.A(\FrameData_O_i[29] ),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_3/_0_  (.A(\FrameData_O_i[3] ),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_30/_0_  (.A(\FrameData_O_i[30] ),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_31/_0_  (.A(\FrameData_O_i[31] ),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_4/_0_  (.A(\FrameData_O_i[4] ),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_5/_0_  (.A(\FrameData_O_i[5] ),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_6/_0_  (.A(\FrameData_O_i[6] ),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_7/_0_  (.A(\FrameData_O_i[7] ),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_8/_0_  (.A(\FrameData_O_i[8] ),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_9/_0_  (.A(\FrameData_O_i[9] ),
    .X(net333));
 sky130_fd_sc_hd__buf_4 input1 (.A(E1END[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(E2END[5]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_16 input100 (.A(FrameStrobe[9]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_8 input101 (.A(N1END[0]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_8 input102 (.A(N1END[1]),
    .X(net102));
 sky130_fd_sc_hd__buf_4 input103 (.A(N1END[2]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_8 input104 (.A(N1END[3]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 input105 (.A(N2END[0]),
    .X(net105));
 sky130_fd_sc_hd__buf_2 input106 (.A(N2END[1]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 input107 (.A(N2END[2]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 input108 (.A(N2END[3]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(N2END[4]),
    .X(net109));
 sky130_fd_sc_hd__buf_2 input11 (.A(E2END[6]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input110 (.A(N2END[5]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 input111 (.A(N2END[6]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 input112 (.A(N2END[7]),
    .X(net112));
 sky130_fd_sc_hd__buf_2 input113 (.A(N2MID[0]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(N2MID[1]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 input115 (.A(N2MID[2]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(N2MID[3]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_4 input117 (.A(N2MID[4]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 input118 (.A(N2MID[5]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 input119 (.A(N2MID[6]),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input12 (.A(E2END[7]),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input120 (.A(N2MID[7]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(N4END[0]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(N4END[10]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(N4END[11]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(N4END[12]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(N4END[13]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(N4END[14]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(N4END[15]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(N4END[1]),
    .X(net128));
 sky130_fd_sc_hd__buf_2 input129 (.A(N4END[2]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(E2MID[0]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input130 (.A(N4END[3]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(N4END[4]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(N4END[5]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(N4END[6]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(N4END[7]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(N4END[8]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(N4END[9]),
    .X(net136));
 sky130_fd_sc_hd__buf_2 input137 (.A(NN4END[0]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(NN4END[10]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(NN4END[11]),
    .X(net139));
 sky130_fd_sc_hd__buf_2 input14 (.A(E2MID[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(NN4END[12]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(NN4END[13]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 input142 (.A(NN4END[14]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(NN4END[15]),
    .X(net143));
 sky130_fd_sc_hd__buf_2 input144 (.A(NN4END[1]),
    .X(net144));
 sky130_fd_sc_hd__buf_2 input145 (.A(NN4END[2]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_4 input146 (.A(NN4END[3]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(NN4END[4]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(NN4END[5]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(NN4END[6]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(E2MID[2]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(NN4END[7]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(NN4END[8]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(NN4END[9]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 input153 (.A(S1END[0]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 input154 (.A(S1END[1]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 input155 (.A(S1END[2]),
    .X(net155));
 sky130_fd_sc_hd__buf_4 input156 (.A(S1END[3]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 input157 (.A(S2END[0]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 input158 (.A(S2END[1]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 input159 (.A(S2END[2]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(E2MID[3]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input160 (.A(S2END[3]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 input161 (.A(S2END[4]),
    .X(net161));
 sky130_fd_sc_hd__buf_2 input162 (.A(S2END[5]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 input163 (.A(S2END[6]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_4 input164 (.A(S2END[7]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 input165 (.A(S2MID[0]),
    .X(net165));
 sky130_fd_sc_hd__buf_2 input166 (.A(S2MID[1]),
    .X(net166));
 sky130_fd_sc_hd__buf_2 input167 (.A(S2MID[2]),
    .X(net167));
 sky130_fd_sc_hd__buf_4 input168 (.A(S2MID[3]),
    .X(net168));
 sky130_fd_sc_hd__buf_2 input169 (.A(S2MID[4]),
    .X(net169));
 sky130_fd_sc_hd__buf_2 input17 (.A(E2MID[4]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input170 (.A(S2MID[5]),
    .X(net170));
 sky130_fd_sc_hd__buf_2 input171 (.A(S2MID[6]),
    .X(net171));
 sky130_fd_sc_hd__buf_2 input172 (.A(S2MID[7]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 input173 (.A(S4END[0]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(S4END[10]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(S4END[11]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(S4END[12]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(S4END[13]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(S4END[14]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(S4END[15]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(E2MID[5]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input180 (.A(S4END[1]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 input181 (.A(S4END[2]),
    .X(net181));
 sky130_fd_sc_hd__buf_2 input182 (.A(S4END[3]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(S4END[4]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(S4END[5]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(S4END[6]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(S4END[7]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(S4END[8]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(S4END[9]),
    .X(net188));
 sky130_fd_sc_hd__buf_2 input189 (.A(SS4END[0]),
    .X(net189));
 sky130_fd_sc_hd__buf_2 input19 (.A(E2MID[6]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(SS4END[10]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(SS4END[11]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(SS4END[12]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(SS4END[13]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(SS4END[14]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(SS4END[15]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_4 input196 (.A(SS4END[1]),
    .X(net196));
 sky130_fd_sc_hd__buf_2 input197 (.A(SS4END[2]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_4 input198 (.A(SS4END[3]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 input199 (.A(SS4END[4]),
    .X(net199));
 sky130_fd_sc_hd__buf_4 input2 (.A(E1END[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(E2MID[7]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input200 (.A(SS4END[5]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 input201 (.A(SS4END[6]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 input202 (.A(SS4END[7]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(SS4END[8]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 input204 (.A(SS4END[9]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_16 input205 (.A(UserCLK),
    .X(net205));
 sky130_fd_sc_hd__buf_4 input206 (.A(W1END[0]),
    .X(net206));
 sky130_fd_sc_hd__buf_4 input207 (.A(W1END[1]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_8 input208 (.A(W1END[2]),
    .X(net208));
 sky130_fd_sc_hd__buf_4 input209 (.A(W1END[3]),
    .X(net209));
 sky130_fd_sc_hd__buf_4 input21 (.A(E6END[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input210 (.A(W2END[0]),
    .X(net210));
 sky130_fd_sc_hd__buf_2 input211 (.A(W2END[1]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_4 input212 (.A(W2END[2]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 input213 (.A(W2END[3]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 input214 (.A(W2END[4]),
    .X(net214));
 sky130_fd_sc_hd__buf_2 input215 (.A(W2END[5]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 input216 (.A(W2END[6]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 input217 (.A(W2END[7]),
    .X(net217));
 sky130_fd_sc_hd__buf_2 input218 (.A(W2MID[0]),
    .X(net218));
 sky130_fd_sc_hd__buf_2 input219 (.A(W2MID[1]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(E6END[10]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input220 (.A(W2MID[2]),
    .X(net220));
 sky130_fd_sc_hd__buf_2 input221 (.A(W2MID[3]),
    .X(net221));
 sky130_fd_sc_hd__buf_2 input222 (.A(W2MID[4]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_4 input223 (.A(W2MID[5]),
    .X(net223));
 sky130_fd_sc_hd__buf_4 input224 (.A(W2MID[6]),
    .X(net224));
 sky130_fd_sc_hd__buf_2 input225 (.A(W2MID[7]),
    .X(net225));
 sky130_fd_sc_hd__buf_4 input226 (.A(W6END[0]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 input227 (.A(W6END[10]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 input228 (.A(W6END[11]),
    .X(net228));
 sky130_fd_sc_hd__buf_4 input229 (.A(W6END[1]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(E6END[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input230 (.A(W6END[2]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 input231 (.A(W6END[3]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 input232 (.A(W6END[4]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 input233 (.A(W6END[5]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 input234 (.A(W6END[6]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 input235 (.A(W6END[7]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 input236 (.A(W6END[8]),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 input237 (.A(W6END[9]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_4 input238 (.A(WW4END[0]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 input239 (.A(WW4END[10]),
    .X(net239));
 sky130_fd_sc_hd__buf_4 input24 (.A(E6END[1]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input240 (.A(WW4END[11]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 input241 (.A(WW4END[12]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 input242 (.A(WW4END[13]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 input243 (.A(WW4END[14]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 input244 (.A(WW4END[15]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_4 input245 (.A(WW4END[1]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 input246 (.A(WW4END[2]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_4 input247 (.A(WW4END[3]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 input248 (.A(WW4END[4]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 input249 (.A(WW4END[5]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(E6END[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input250 (.A(WW4END[6]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 input251 (.A(WW4END[7]),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 input252 (.A(WW4END[8]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 input253 (.A(WW4END[9]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(E6END[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(E6END[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(E6END[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(E6END[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input3 (.A(E1END[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(E6END[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(E6END[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(E6END[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(EE4END[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(EE4END[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(EE4END[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(EE4END[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(EE4END[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(EE4END[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(EE4END[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input4 (.A(E1END[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(EE4END[1]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(EE4END[2]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(EE4END[3]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(EE4END[4]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(EE4END[5]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(EE4END[6]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(EE4END[7]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(EE4END[8]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(EE4END[9]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_8 input49 (.A(FrameData[0]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(E2END[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_8 input50 (.A(FrameData[10]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_8 input51 (.A(FrameData[11]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_8 input52 (.A(FrameData[12]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_8 input53 (.A(FrameData[13]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_8 input54 (.A(FrameData[14]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_8 input55 (.A(FrameData[15]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_8 input56 (.A(FrameData[16]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_8 input57 (.A(FrameData[17]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_8 input58 (.A(FrameData[18]),
    .X(net58));
 sky130_fd_sc_hd__buf_6 input59 (.A(FrameData[19]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(E2END[1]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input60 (.A(FrameData[1]),
    .X(net60));
 sky130_fd_sc_hd__buf_6 input61 (.A(FrameData[20]),
    .X(net61));
 sky130_fd_sc_hd__buf_6 input62 (.A(FrameData[21]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_8 input63 (.A(FrameData[22]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_8 input64 (.A(FrameData[23]),
    .X(net64));
 sky130_fd_sc_hd__buf_6 input65 (.A(FrameData[24]),
    .X(net65));
 sky130_fd_sc_hd__buf_6 input66 (.A(FrameData[25]),
    .X(net66));
 sky130_fd_sc_hd__buf_6 input67 (.A(FrameData[26]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_8 input68 (.A(FrameData[27]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_8 input69 (.A(FrameData[28]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(E2END[2]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_8 input70 (.A(FrameData[29]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_8 input71 (.A(FrameData[2]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_8 input72 (.A(FrameData[30]),
    .X(net72));
 sky130_fd_sc_hd__buf_6 input73 (.A(FrameData[31]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_8 input74 (.A(FrameData[3]),
    .X(net74));
 sky130_fd_sc_hd__buf_6 input75 (.A(FrameData[4]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_8 input76 (.A(FrameData[5]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_8 input77 (.A(FrameData[6]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_8 input78 (.A(FrameData[7]),
    .X(net78));
 sky130_fd_sc_hd__buf_4 input79 (.A(FrameData[8]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(E2END[3]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input80 (.A(FrameData[9]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_16 input81 (.A(FrameStrobe[0]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_16 input82 (.A(FrameStrobe[10]),
    .X(net82));
 sky130_fd_sc_hd__buf_8 input83 (.A(FrameStrobe[11]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_16 input84 (.A(FrameStrobe[12]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(FrameStrobe[13]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(FrameStrobe[14]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(FrameStrobe[15]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(FrameStrobe[16]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(FrameStrobe[17]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(E2END[4]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(FrameStrobe[18]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(FrameStrobe[19]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_16 input92 (.A(FrameStrobe[1]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_16 input93 (.A(FrameStrobe[2]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_16 input94 (.A(FrameStrobe[3]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_16 input95 (.A(FrameStrobe[4]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_16 input96 (.A(FrameStrobe[5]),
    .X(net96));
 sky130_fd_sc_hd__buf_12 input97 (.A(FrameStrobe[6]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_16 input98 (.A(FrameStrobe[7]),
    .X(net98));
 sky130_fd_sc_hd__buf_12 input99 (.A(FrameStrobe[8]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 inst_clk_buf (.A(net205),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_4 output254 (.A(net254),
    .X(E1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output255 (.A(net255),
    .X(E1BEG[1]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(E1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output257 (.A(net257),
    .X(E1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output258 (.A(net258),
    .X(E2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output259 (.A(net259),
    .X(E2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output260 (.A(net260),
    .X(E2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output261 (.A(net261),
    .X(E2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output262 (.A(net262),
    .X(E2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output263 (.A(net263),
    .X(E2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output264 (.A(net264),
    .X(E2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output265 (.A(net265),
    .X(E2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output266 (.A(net266),
    .X(E2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output267 (.A(net267),
    .X(E2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output268 (.A(net268),
    .X(E2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output269 (.A(net269),
    .X(E2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output270 (.A(net270),
    .X(E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(E2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output272 (.A(net272),
    .X(E2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output273 (.A(net273),
    .X(E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(E6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output275 (.A(net275),
    .X(E6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output276 (.A(net276),
    .X(E6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output277 (.A(net277),
    .X(E6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output278 (.A(net278),
    .X(E6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output279 (.A(net279),
    .X(E6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output280 (.A(net280),
    .X(E6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output281 (.A(net281),
    .X(E6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output282 (.A(net282),
    .X(E6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output283 (.A(net283),
    .X(E6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output284 (.A(net284),
    .X(E6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output285 (.A(net285),
    .X(E6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output286 (.A(net286),
    .X(EE4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output287 (.A(net287),
    .X(EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(EE4BEG[11]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(EE4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output290 (.A(net290),
    .X(EE4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output291 (.A(net291),
    .X(EE4BEG[14]));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(EE4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output293 (.A(net293),
    .X(EE4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output294 (.A(net294),
    .X(EE4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output295 (.A(net295),
    .X(EE4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output296 (.A(net296),
    .X(EE4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output297 (.A(net297),
    .X(EE4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output298 (.A(net298),
    .X(EE4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output299 (.A(net299),
    .X(EE4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output300 (.A(net300),
    .X(EE4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output301 (.A(net301),
    .X(EE4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output302 (.A(net302),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output303 (.A(net303),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output304 (.A(net304),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output305 (.A(net305),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output306 (.A(net306),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output307 (.A(net307),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output308 (.A(net308),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output309 (.A(net309),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output310 (.A(net310),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output311 (.A(net311),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output313 (.A(net313),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__clkbuf_4 output314 (.A(net314),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__clkbuf_4 output315 (.A(net315),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__clkbuf_4 output316 (.A(net316),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output318 (.A(net318),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__clkbuf_4 output319 (.A(net319),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__clkbuf_4 output320 (.A(net320),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__clkbuf_4 output321 (.A(net321),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__clkbuf_4 output323 (.A(net323),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__clkbuf_4 output324 (.A(net324),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output325 (.A(net325),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__clkbuf_4 output326 (.A(net326),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output329 (.A(net329),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output330 (.A(net330),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output331 (.A(net331),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output332 (.A(net332),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output333 (.A(net333),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output334 (.A(net334),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output335 (.A(net335),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output336 (.A(net336),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output337 (.A(net337),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output338 (.A(net338),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output339 (.A(net339),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output340 (.A(net340),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output341 (.A(net341),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output342 (.A(net342),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output343 (.A(net343),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output344 (.A(net344),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output345 (.A(net345),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output346 (.A(net346),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output347 (.A(net347),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__clkbuf_4 output348 (.A(net348),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output349 (.A(net349),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output350 (.A(net350),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output351 (.A(net351),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__clkbuf_4 output352 (.A(net352),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output353 (.A(net353),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output354 (.A(net354),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output355 (.A(net355),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output356 (.A(net356),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__buf_2 output357 (.A(net357),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output358 (.A(net358),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output359 (.A(net359),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net360),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__buf_2 output361 (.A(net361),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output362 (.A(net362),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output363 (.A(net363),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__buf_2 output364 (.A(net364),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net365),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output366 (.A(net366),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output367 (.A(net367),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output368 (.A(net368),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output369 (.A(net369),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output370 (.A(net370),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output371 (.A(net371),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output372 (.A(net372),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output373 (.A(net373),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output374 (.A(net374),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output375 (.A(net375),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output376 (.A(net376),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output377 (.A(net377),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__buf_2 output378 (.A(net378),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output379 (.A(net379),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output380 (.A(net380),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output381 (.A(net381),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output382 (.A(net382),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output383 (.A(net383),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output384 (.A(net384),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output385 (.A(net385),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output386 (.A(net386),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output387 (.A(net387),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output388 (.A(net388),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output389 (.A(net389),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output390 (.A(net390),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output391 (.A(net391),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output392 (.A(net392),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__buf_2 output393 (.A(net393),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output394 (.A(net394),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output395 (.A(net395),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__buf_2 output396 (.A(net396),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__buf_2 output397 (.A(net397),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output398 (.A(net398),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output399 (.A(net399),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output400 (.A(net400),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__buf_2 output401 (.A(net401),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output402 (.A(net402),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output403 (.A(net403),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output404 (.A(net404),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__buf_2 output405 (.A(net405),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__buf_2 output406 (.A(net406),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__buf_2 output407 (.A(net407),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output408 (.A(net408),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__buf_2 output409 (.A(net409),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output410 (.A(net410),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__buf_2 output411 (.A(net411),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__buf_2 output412 (.A(net412),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output413 (.A(net413),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output414 (.A(net414),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__buf_2 output415 (.A(net415),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__buf_2 output416 (.A(net416),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output417 (.A(net417),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output418 (.A(net418),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output419 (.A(net419),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output420 (.A(net420),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output421 (.A(net421),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output422 (.A(net422),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output423 (.A(net423),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output424 (.A(net424),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output425 (.A(net425),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output426 (.A(net426),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output427 (.A(net427),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output428 (.A(net428),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__buf_2 output429 (.A(net429),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output430 (.A(net430),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output431 (.A(net431),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__buf_2 output432 (.A(net432),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output433 (.A(net433),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output434 (.A(net434),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output435 (.A(net435),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output436 (.A(net436),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output437 (.A(net437),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output438 (.A(net438),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output439 (.A(net439),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__buf_2 output440 (.A(net440),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output441 (.A(net441),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output442 (.A(net442),
    .X(SS4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output443 (.A(net443),
    .X(SS4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output444 (.A(net444),
    .X(SS4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output445 (.A(net445),
    .X(SS4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output446 (.A(net446),
    .X(SS4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output447 (.A(net447),
    .X(SS4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output448 (.A(net448),
    .X(SS4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output449 (.A(net449),
    .X(SS4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output450 (.A(net450),
    .X(SS4BEG[2]));
 sky130_fd_sc_hd__buf_2 output451 (.A(net451),
    .X(SS4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output452 (.A(net452),
    .X(SS4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output453 (.A(net453),
    .X(SS4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output454 (.A(net454),
    .X(SS4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output455 (.A(net455),
    .X(SS4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output456 (.A(net456),
    .X(SS4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output457 (.A(net457),
    .X(SS4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output458 (.A(net458),
    .X(UserCLKo));
 sky130_fd_sc_hd__clkbuf_4 output459 (.A(net459),
    .X(W1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output460 (.A(net460),
    .X(W1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output461 (.A(net461),
    .X(W1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output462 (.A(net462),
    .X(W1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output463 (.A(net463),
    .X(W2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output464 (.A(net464),
    .X(W2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output465 (.A(net465),
    .X(W2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output466 (.A(net466),
    .X(W2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output467 (.A(net467),
    .X(W2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output468 (.A(net468),
    .X(W2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output469 (.A(net469),
    .X(W2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output470 (.A(net470),
    .X(W2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output471 (.A(net471),
    .X(W2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output472 (.A(net472),
    .X(W2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output473 (.A(net473),
    .X(W2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output474 (.A(net474),
    .X(W2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output475 (.A(net475),
    .X(W2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output476 (.A(net476),
    .X(W2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output477 (.A(net477),
    .X(W2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output478 (.A(net478),
    .X(W2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output479 (.A(net479),
    .X(W6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output480 (.A(net480),
    .X(W6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output481 (.A(net481),
    .X(W6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output482 (.A(net482),
    .X(W6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output483 (.A(net483),
    .X(W6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output484 (.A(net484),
    .X(W6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output485 (.A(net485),
    .X(W6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output486 (.A(net486),
    .X(W6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output487 (.A(net487),
    .X(W6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output488 (.A(net488),
    .X(W6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output489 (.A(net489),
    .X(W6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output490 (.A(net490),
    .X(W6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output491 (.A(net491),
    .X(WW4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output492 (.A(net492),
    .X(WW4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output493 (.A(net493),
    .X(WW4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output494 (.A(net494),
    .X(WW4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output495 (.A(net495),
    .X(WW4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output496 (.A(net496),
    .X(WW4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output497 (.A(net497),
    .X(WW4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output498 (.A(net498),
    .X(WW4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output499 (.A(net499),
    .X(WW4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output500 (.A(net500),
    .X(WW4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output501 (.A(net501),
    .X(WW4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output502 (.A(net502),
    .X(WW4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output503 (.A(net503),
    .X(WW4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output504 (.A(net504),
    .X(WW4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output505 (.A(net505),
    .X(WW4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output506 (.A(net506),
    .X(WW4BEG[9]));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_0/_0_  (.A(net81),
    .X(\FrameStrobe_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_1/_0_  (.A(net92),
    .X(\FrameStrobe_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_10/_0_  (.A(net82),
    .X(\FrameStrobe_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_11/_0_  (.A(net83),
    .X(\FrameStrobe_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_12/_0_  (.A(net84),
    .X(\FrameStrobe_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_13/_0_  (.A(net85),
    .X(\FrameStrobe_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_14/_0_  (.A(net86),
    .X(\FrameStrobe_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_15/_0_  (.A(net87),
    .X(\FrameStrobe_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_16/_0_  (.A(net88),
    .X(\FrameStrobe_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_17/_0_  (.A(net89),
    .X(\FrameStrobe_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_18/_0_  (.A(net90),
    .X(\FrameStrobe_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_19/_0_  (.A(net91),
    .X(\FrameStrobe_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_2/_0_  (.A(net93),
    .X(\FrameStrobe_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_3/_0_  (.A(net94),
    .X(\FrameStrobe_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_4/_0_  (.A(net95),
    .X(\FrameStrobe_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_5/_0_  (.A(net96),
    .X(\FrameStrobe_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_6/_0_  (.A(net97),
    .X(\FrameStrobe_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_7/_0_  (.A(net98),
    .X(\FrameStrobe_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_8/_0_  (.A(net99),
    .X(\FrameStrobe_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_9/_0_  (.A(net100),
    .X(\FrameStrobe_O_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_0/_0_  (.A(\FrameStrobe_O_i[0] ),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_1/_0_  (.A(\FrameStrobe_O_i[1] ),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_10/_0_  (.A(\FrameStrobe_O_i[10] ),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_11/_0_  (.A(\FrameStrobe_O_i[11] ),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_12/_0_  (.A(\FrameStrobe_O_i[12] ),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_13/_0_  (.A(\FrameStrobe_O_i[13] ),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_14/_0_  (.A(\FrameStrobe_O_i[14] ),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_15/_0_  (.A(\FrameStrobe_O_i[15] ),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_16/_0_  (.A(\FrameStrobe_O_i[16] ),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_17/_0_  (.A(\FrameStrobe_O_i[17] ),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_18/_0_  (.A(\FrameStrobe_O_i[18] ),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_19/_0_  (.A(\FrameStrobe_O_i[19] ),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_2/_0_  (.A(\FrameStrobe_O_i[2] ),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_3/_0_  (.A(\FrameStrobe_O_i[3] ),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_4/_0_  (.A(\FrameStrobe_O_i[4] ),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_5/_0_  (.A(\FrameStrobe_O_i[5] ),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_6/_0_  (.A(\FrameStrobe_O_i[6] ),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_7/_0_  (.A(\FrameStrobe_O_i[7] ),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_8/_0_  (.A(\FrameStrobe_O_i[8] ),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_9/_0_  (.A(\FrameStrobe_O_i[9] ),
    .X(net353));
endmodule

