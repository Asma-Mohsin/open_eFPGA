magic
tech sky130A
magscale 1 2
timestamp 1733394398
<< viali >>
rect 3893 8585 3927 8619
rect 6009 8585 6043 8619
rect 8033 8585 8067 8619
rect 10425 8585 10459 8619
rect 12633 8585 12667 8619
rect 14841 8585 14875 8619
rect 17049 8585 17083 8619
rect 19349 8585 19383 8619
rect 21465 8585 21499 8619
rect 23673 8585 23707 8619
rect 25881 8585 25915 8619
rect 28089 8585 28123 8619
rect 30113 8585 30147 8619
rect 32505 8585 32539 8619
rect 34989 8585 35023 8619
rect 36921 8585 36955 8619
rect 39129 8585 39163 8619
rect 41153 8585 41187 8619
rect 43545 8585 43579 8619
rect 45385 8585 45419 8619
rect 1409 8517 1443 8551
rect 1777 8517 1811 8551
rect 4077 8449 4111 8483
rect 6193 8449 6227 8483
rect 8309 8449 8343 8483
rect 10609 8449 10643 8483
rect 12725 8449 12759 8483
rect 15025 8449 15059 8483
rect 17233 8449 17267 8483
rect 19625 8449 19659 8483
rect 21649 8449 21683 8483
rect 23765 8449 23799 8483
rect 26065 8449 26099 8483
rect 28273 8449 28307 8483
rect 30389 8449 30423 8483
rect 32689 8449 32723 8483
rect 35081 8449 35115 8483
rect 37105 8449 37139 8483
rect 39313 8449 39347 8483
rect 41429 8449 41463 8483
rect 43729 8449 43763 8483
rect 45109 8449 45143 8483
rect 17417 2601 17451 2635
rect 22753 2601 22787 2635
rect 23029 2601 23063 2635
rect 23305 2601 23339 2635
rect 23581 2601 23615 2635
rect 23949 2601 23983 2635
rect 28273 2601 28307 2635
rect 32689 2601 32723 2635
rect 35081 2601 35115 2635
rect 37105 2601 37139 2635
rect 39497 2601 39531 2635
rect 41613 2601 41647 2635
rect 44005 2601 44039 2635
rect 44833 2601 44867 2635
rect 18705 2533 18739 2567
rect 19625 2533 19659 2567
rect 21373 2533 21407 2567
rect 24409 2533 24443 2567
rect 26065 2533 26099 2567
rect 26525 2533 26559 2567
rect 30297 2533 30331 2567
rect 17601 2397 17635 2431
rect 18521 2397 18555 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 19717 2397 19751 2431
rect 20269 2397 20303 2431
rect 20453 2397 20487 2431
rect 20913 2397 20947 2431
rect 21189 2397 21223 2431
rect 21833 2397 21867 2431
rect 21925 2397 21959 2431
rect 22385 2397 22419 2431
rect 22477 2397 22511 2431
rect 22937 2397 22971 2431
rect 23213 2397 23247 2431
rect 23489 2397 23523 2431
rect 23765 2397 23799 2431
rect 24593 2397 24627 2431
rect 26249 2397 26283 2431
rect 26341 2397 26375 2431
rect 26617 2397 26651 2431
rect 26893 2397 26927 2431
rect 27353 2397 27387 2431
rect 27445 2397 27479 2431
rect 27905 2397 27939 2431
rect 28457 2397 28491 2431
rect 30113 2397 30147 2431
rect 30665 2397 30699 2431
rect 30757 2397 30791 2431
rect 31125 2397 31159 2431
rect 31401 2397 31435 2431
rect 32137 2397 32171 2431
rect 32873 2397 32907 2431
rect 33425 2397 33459 2431
rect 34897 2397 34931 2431
rect 37289 2397 37323 2431
rect 39681 2397 39715 2431
rect 41797 2397 41831 2431
rect 44189 2397 44223 2431
rect 44649 2397 44683 2431
rect 45201 2397 45235 2431
rect 45477 2397 45511 2431
rect 24041 2329 24075 2363
rect 19073 2261 19107 2295
rect 19901 2261 19935 2295
rect 20085 2261 20119 2295
rect 20637 2261 20671 2295
rect 21097 2261 21131 2295
rect 21649 2261 21683 2295
rect 22109 2261 22143 2295
rect 22201 2261 22235 2295
rect 22661 2261 22695 2295
rect 26801 2261 26835 2295
rect 27077 2261 27111 2295
rect 27169 2261 27203 2295
rect 27629 2261 27663 2295
rect 28089 2261 28123 2295
rect 30481 2261 30515 2295
rect 30941 2261 30975 2295
rect 31309 2261 31343 2295
rect 31585 2261 31619 2295
rect 32321 2261 32355 2295
rect 33241 2261 33275 2295
rect 45017 2261 45051 2295
rect 45293 2261 45327 2295
rect 1869 2057 1903 2091
rect 2789 2057 2823 2091
rect 3157 2057 3191 2091
rect 9413 2057 9447 2091
rect 9781 2057 9815 2091
rect 15945 2057 15979 2091
rect 16221 2057 16255 2091
rect 16497 2057 16531 2091
rect 17049 2057 17083 2091
rect 18981 2057 19015 2091
rect 19257 2057 19291 2091
rect 19809 2057 19843 2091
rect 22109 2057 22143 2091
rect 23029 2057 23063 2091
rect 23673 2057 23707 2091
rect 24777 2057 24811 2091
rect 25053 2057 25087 2091
rect 29929 2057 29963 2091
rect 30389 2057 30423 2091
rect 35173 2057 35207 2091
rect 37657 2057 37691 2091
rect 39405 2057 39439 2091
rect 39773 2057 39807 2091
rect 40969 2057 41003 2091
rect 42441 2057 42475 2091
rect 44649 2057 44683 2091
rect 44925 2057 44959 2091
rect 31033 1989 31067 2023
rect 32965 1989 32999 2023
rect 33609 1989 33643 2023
rect 34161 1989 34195 2023
rect 36185 1989 36219 2023
rect 39313 1989 39347 2023
rect 1409 1921 1443 1955
rect 1685 1921 1719 1955
rect 2605 1921 2639 1955
rect 2973 1921 3007 1955
rect 9229 1921 9263 1955
rect 9597 1921 9631 1955
rect 15209 1921 15243 1955
rect 15485 1921 15519 1955
rect 15761 1921 15795 1955
rect 16037 1921 16071 1955
rect 16313 1921 16347 1955
rect 16865 1921 16899 1955
rect 17141 1921 17175 1955
rect 17417 1921 17451 1955
rect 17693 1921 17727 1955
rect 17969 1921 18003 1955
rect 18245 1921 18279 1955
rect 18521 1921 18555 1955
rect 18797 1921 18831 1955
rect 19073 1921 19107 1955
rect 19349 1921 19383 1955
rect 19625 1921 19659 1955
rect 19901 1921 19935 1955
rect 20177 1921 20211 1955
rect 20453 1921 20487 1955
rect 20729 1921 20763 1955
rect 21005 1921 21039 1955
rect 21465 1921 21499 1955
rect 21925 1921 21959 1955
rect 22201 1921 22235 1955
rect 22465 1921 22499 1955
rect 22845 1921 22879 1955
rect 23121 1921 23155 1955
rect 23397 1921 23431 1955
rect 23857 1921 23891 1955
rect 23949 1921 23983 1955
rect 24501 1921 24535 1955
rect 24961 1921 24995 1955
rect 25237 1921 25271 1955
rect 25329 1921 25363 1955
rect 25789 1921 25823 1955
rect 26157 1921 26191 1955
rect 26433 1921 26467 1955
rect 26985 1921 27019 1955
rect 27721 1921 27755 1955
rect 27905 1921 27939 1955
rect 28457 1921 28491 1955
rect 28825 1921 28859 1955
rect 29101 1921 29135 1955
rect 29377 1921 29411 1955
rect 29653 1921 29687 1955
rect 30113 1921 30147 1955
rect 30205 1921 30239 1955
rect 30481 1921 30515 1955
rect 31585 1921 31619 1955
rect 32137 1921 32171 1955
rect 32597 1921 32631 1955
rect 35357 1921 35391 1955
rect 35541 1921 35575 1955
rect 36737 1921 36771 1955
rect 37841 1921 37875 1955
rect 38117 1921 38151 1955
rect 38761 1921 38795 1955
rect 39957 1921 39991 1955
rect 40601 1921 40635 1955
rect 40877 1921 40911 1955
rect 41153 1921 41187 1955
rect 41613 1921 41647 1955
rect 42625 1921 42659 1955
rect 44833 1921 44867 1955
rect 45109 1921 45143 1955
rect 45477 1921 45511 1955
rect 27537 1853 27571 1887
rect 31309 1853 31343 1887
rect 31861 1853 31895 1887
rect 41337 1853 41371 1887
rect 15393 1785 15427 1819
rect 17325 1785 17359 1819
rect 17877 1785 17911 1819
rect 18429 1785 18463 1819
rect 19533 1785 19567 1819
rect 21649 1785 21683 1819
rect 24685 1785 24719 1819
rect 26617 1785 26651 1819
rect 29009 1785 29043 1819
rect 29837 1785 29871 1819
rect 30665 1785 30699 1819
rect 32321 1785 32355 1819
rect 32413 1785 32447 1819
rect 33149 1785 33183 1819
rect 40693 1785 40727 1819
rect 45293 1785 45327 1819
rect 1593 1717 1627 1751
rect 15669 1717 15703 1751
rect 17601 1717 17635 1751
rect 18153 1717 18187 1751
rect 18705 1717 18739 1751
rect 20085 1717 20119 1751
rect 20361 1717 20395 1751
rect 20637 1717 20671 1751
rect 20913 1717 20947 1751
rect 21189 1717 21223 1751
rect 22385 1717 22419 1751
rect 22661 1717 22695 1751
rect 23305 1717 23339 1751
rect 23581 1717 23615 1751
rect 24133 1717 24167 1751
rect 25513 1717 25547 1751
rect 25973 1717 26007 1751
rect 26341 1717 26375 1751
rect 27169 1717 27203 1751
rect 28089 1717 28123 1751
rect 28641 1717 28675 1751
rect 29285 1717 29319 1751
rect 29561 1717 29595 1751
rect 33701 1717 33735 1751
rect 34253 1717 34287 1751
rect 35633 1717 35667 1751
rect 36277 1717 36311 1751
rect 36829 1717 36863 1751
rect 38209 1717 38243 1751
rect 38853 1717 38887 1751
rect 40417 1717 40451 1751
rect 6837 1513 6871 1547
rect 14289 1513 14323 1547
rect 15117 1513 15151 1547
rect 15393 1513 15427 1547
rect 15669 1513 15703 1547
rect 15945 1513 15979 1547
rect 16221 1513 16255 1547
rect 16497 1513 16531 1547
rect 16957 1513 16991 1547
rect 17509 1513 17543 1547
rect 17969 1513 18003 1547
rect 18337 1513 18371 1547
rect 18613 1513 18647 1547
rect 19257 1513 19291 1547
rect 22293 1513 22327 1547
rect 26341 1513 26375 1547
rect 27169 1513 27203 1547
rect 27905 1513 27939 1547
rect 28457 1513 28491 1547
rect 29745 1513 29779 1547
rect 30297 1513 30331 1547
rect 30849 1513 30883 1547
rect 32873 1513 32907 1547
rect 33425 1513 33459 1547
rect 35449 1513 35483 1547
rect 36553 1513 36587 1547
rect 38025 1513 38059 1547
rect 39129 1513 39163 1547
rect 40049 1513 40083 1547
rect 43453 1513 43487 1547
rect 45293 1513 45327 1547
rect 20913 1445 20947 1479
rect 32413 1445 32447 1479
rect 38669 1445 38703 1479
rect 39497 1445 39531 1479
rect 45017 1445 45051 1479
rect 28917 1377 28951 1411
rect 35081 1377 35115 1411
rect 37657 1377 37691 1411
rect 1501 1309 1535 1343
rect 1869 1309 1903 1343
rect 2237 1309 2271 1343
rect 2513 1309 2547 1343
rect 3341 1309 3375 1343
rect 3801 1309 3835 1343
rect 4077 1309 4111 1343
rect 4445 1309 4479 1343
rect 4813 1309 4847 1343
rect 5181 1309 5215 1343
rect 5549 1309 5583 1343
rect 5917 1309 5951 1343
rect 6377 1309 6411 1343
rect 6653 1309 6687 1343
rect 7021 1309 7055 1343
rect 7389 1309 7423 1343
rect 7757 1309 7791 1343
rect 8125 1309 8159 1343
rect 8585 1309 8619 1343
rect 8953 1309 8987 1343
rect 9229 1309 9263 1343
rect 9965 1309 9999 1343
rect 10333 1309 10367 1343
rect 10701 1309 10735 1343
rect 11069 1309 11103 1343
rect 11529 1309 11563 1343
rect 11805 1309 11839 1343
rect 12173 1309 12207 1343
rect 12541 1309 12575 1343
rect 12909 1309 12943 1343
rect 13277 1309 13311 1343
rect 13645 1309 13679 1343
rect 14105 1309 14139 1343
rect 14381 1309 14415 1343
rect 14657 1309 14691 1343
rect 14933 1309 14967 1343
rect 15209 1309 15243 1343
rect 15485 1309 15519 1343
rect 15761 1309 15795 1343
rect 16037 1309 16071 1343
rect 16313 1309 16347 1343
rect 16773 1309 16807 1343
rect 17049 1309 17083 1343
rect 17693 1309 17727 1343
rect 17785 1309 17819 1343
rect 18061 1309 18095 1343
rect 18521 1309 18555 1343
rect 18797 1309 18831 1343
rect 18889 1309 18923 1343
rect 19441 1309 19475 1343
rect 19533 1309 19567 1343
rect 19901 1309 19935 1343
rect 20269 1309 20303 1343
rect 21373 1309 21407 1343
rect 21833 1309 21867 1343
rect 22845 1309 22879 1343
rect 23213 1309 23247 1343
rect 24777 1309 24811 1343
rect 25789 1309 25823 1343
rect 26249 1309 26283 1343
rect 27077 1309 27111 1343
rect 27813 1309 27847 1343
rect 28365 1309 28399 1343
rect 29193 1309 29227 1343
rect 30205 1309 30239 1343
rect 31309 1309 31343 1343
rect 32229 1309 32263 1343
rect 33333 1309 33367 1343
rect 33885 1309 33919 1343
rect 37381 1309 37415 1343
rect 37933 1309 37967 1343
rect 38485 1309 38519 1343
rect 39037 1309 39071 1343
rect 39681 1309 39715 1343
rect 40601 1309 40635 1343
rect 40877 1309 40911 1343
rect 40969 1309 41003 1343
rect 41245 1309 41279 1343
rect 42073 1309 42107 1343
rect 42625 1309 42659 1343
rect 42901 1309 42935 1343
rect 43269 1309 43303 1343
rect 43637 1309 43671 1343
rect 44005 1309 44039 1343
rect 44373 1309 44407 1343
rect 44741 1309 44775 1343
rect 45201 1309 45235 1343
rect 45477 1309 45511 1343
rect 20729 1241 20763 1275
rect 22201 1241 22235 1275
rect 23673 1241 23707 1275
rect 25329 1241 25363 1275
rect 29653 1241 29687 1275
rect 30757 1241 30791 1275
rect 32781 1241 32815 1275
rect 34805 1241 34839 1275
rect 35357 1241 35391 1275
rect 35909 1241 35943 1275
rect 36461 1241 36495 1275
rect 39957 1241 39991 1275
rect 1685 1173 1719 1207
rect 2053 1173 2087 1207
rect 3525 1173 3559 1207
rect 3985 1173 4019 1207
rect 4261 1173 4295 1207
rect 4629 1173 4663 1207
rect 4997 1173 5031 1207
rect 5365 1173 5399 1207
rect 5733 1173 5767 1207
rect 6101 1173 6135 1207
rect 6561 1173 6595 1207
rect 7205 1173 7239 1207
rect 7573 1173 7607 1207
rect 7941 1173 7975 1207
rect 8309 1173 8343 1207
rect 8769 1173 8803 1207
rect 10149 1173 10183 1207
rect 10517 1173 10551 1207
rect 10885 1173 10919 1207
rect 11253 1173 11287 1207
rect 11713 1173 11747 1207
rect 11989 1173 12023 1207
rect 12357 1173 12391 1207
rect 12725 1173 12759 1207
rect 13093 1173 13127 1207
rect 13461 1173 13495 1207
rect 13829 1173 13863 1207
rect 14565 1173 14599 1207
rect 14841 1173 14875 1207
rect 17233 1173 17267 1207
rect 18245 1173 18279 1207
rect 19073 1173 19107 1207
rect 19717 1173 19751 1207
rect 20085 1173 20119 1207
rect 20453 1173 20487 1207
rect 21557 1173 21591 1207
rect 22017 1173 22051 1207
rect 23029 1173 23063 1207
rect 23397 1173 23431 1207
rect 23765 1173 23799 1207
rect 24869 1173 24903 1207
rect 25421 1173 25455 1207
rect 25973 1173 26007 1207
rect 31401 1173 31435 1207
rect 33977 1173 34011 1207
rect 36001 1173 36035 1207
rect 40417 1173 40451 1207
rect 40693 1173 40727 1207
rect 41889 1173 41923 1207
rect 42441 1173 42475 1207
rect 42717 1173 42751 1207
rect 43085 1173 43119 1207
rect 43821 1173 43855 1207
rect 44189 1173 44223 1207
rect 44557 1173 44591 1207
<< metal1 >>
rect 14918 8984 14924 9036
rect 14976 9024 14982 9036
rect 23014 9024 23020 9036
rect 14976 8996 23020 9024
rect 14976 8984 14982 8996
rect 23014 8984 23020 8996
rect 23072 8984 23078 9036
rect 22738 8956 22744 8968
rect 6196 8928 22744 8956
rect 6196 8832 6224 8928
rect 22738 8916 22744 8928
rect 22796 8916 22802 8968
rect 23934 8888 23940 8900
rect 6886 8860 23940 8888
rect 6178 8780 6184 8832
rect 6236 8780 6242 8832
rect 6270 8780 6276 8832
rect 6328 8820 6334 8832
rect 6886 8820 6914 8860
rect 23934 8848 23940 8860
rect 23992 8848 23998 8900
rect 6328 8792 6914 8820
rect 6328 8780 6334 8792
rect 10134 8780 10140 8832
rect 10192 8820 10198 8832
rect 27522 8820 27528 8832
rect 10192 8792 27528 8820
rect 10192 8780 10198 8792
rect 27522 8780 27528 8792
rect 27580 8780 27586 8832
rect 1104 8730 45976 8752
rect 1104 8678 12128 8730
rect 12180 8678 12192 8730
rect 12244 8678 12256 8730
rect 12308 8678 12320 8730
rect 12372 8678 12384 8730
rect 12436 8678 23306 8730
rect 23358 8678 23370 8730
rect 23422 8678 23434 8730
rect 23486 8678 23498 8730
rect 23550 8678 23562 8730
rect 23614 8678 34484 8730
rect 34536 8678 34548 8730
rect 34600 8678 34612 8730
rect 34664 8678 34676 8730
rect 34728 8678 34740 8730
rect 34792 8678 45662 8730
rect 45714 8678 45726 8730
rect 45778 8678 45790 8730
rect 45842 8678 45854 8730
rect 45906 8678 45918 8730
rect 45970 8678 45976 8730
rect 1104 8656 45976 8678
rect 3602 8576 3608 8628
rect 3660 8616 3666 8628
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 3660 8588 3893 8616
rect 3660 8576 3666 8588
rect 3881 8585 3893 8588
rect 3927 8585 3939 8619
rect 3881 8579 3939 8585
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 5997 8619 6055 8625
rect 5997 8616 6009 8619
rect 5868 8588 6009 8616
rect 5868 8576 5874 8588
rect 5997 8585 6009 8588
rect 6043 8585 6055 8619
rect 5997 8579 6055 8585
rect 8018 8576 8024 8628
rect 8076 8576 8082 8628
rect 10134 8576 10140 8628
rect 10192 8576 10198 8628
rect 10226 8576 10232 8628
rect 10284 8616 10290 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 10284 8588 10425 8616
rect 10284 8576 10290 8588
rect 10413 8585 10425 8588
rect 10459 8585 10471 8619
rect 10413 8579 10471 8585
rect 12618 8576 12624 8628
rect 12676 8576 12682 8628
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 14829 8619 14887 8625
rect 14829 8616 14841 8619
rect 14700 8588 14841 8616
rect 14700 8576 14706 8588
rect 14829 8585 14841 8588
rect 14875 8585 14887 8619
rect 14829 8579 14887 8585
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 17037 8619 17095 8625
rect 17037 8616 17049 8619
rect 16908 8588 17049 8616
rect 16908 8576 16914 8588
rect 17037 8585 17049 8588
rect 17083 8585 17095 8619
rect 17037 8579 17095 8585
rect 19058 8576 19064 8628
rect 19116 8616 19122 8628
rect 19337 8619 19395 8625
rect 19337 8616 19349 8619
rect 19116 8588 19349 8616
rect 19116 8576 19122 8588
rect 19337 8585 19349 8588
rect 19383 8585 19395 8619
rect 19337 8579 19395 8585
rect 21266 8576 21272 8628
rect 21324 8616 21330 8628
rect 21453 8619 21511 8625
rect 21453 8616 21465 8619
rect 21324 8588 21465 8616
rect 21324 8576 21330 8588
rect 21453 8585 21465 8588
rect 21499 8585 21511 8619
rect 21453 8579 21511 8585
rect 23658 8576 23664 8628
rect 23716 8576 23722 8628
rect 25682 8576 25688 8628
rect 25740 8616 25746 8628
rect 25869 8619 25927 8625
rect 25869 8616 25881 8619
rect 25740 8588 25881 8616
rect 25740 8576 25746 8588
rect 25869 8585 25881 8588
rect 25915 8585 25927 8619
rect 25869 8579 25927 8585
rect 27890 8576 27896 8628
rect 27948 8616 27954 8628
rect 28077 8619 28135 8625
rect 28077 8616 28089 8619
rect 27948 8588 28089 8616
rect 27948 8576 27954 8588
rect 28077 8585 28089 8588
rect 28123 8585 28135 8619
rect 28077 8579 28135 8585
rect 30098 8576 30104 8628
rect 30156 8576 30162 8628
rect 32306 8576 32312 8628
rect 32364 8616 32370 8628
rect 32493 8619 32551 8625
rect 32493 8616 32505 8619
rect 32364 8588 32505 8616
rect 32364 8576 32370 8588
rect 32493 8585 32505 8588
rect 32539 8585 32551 8619
rect 32493 8579 32551 8585
rect 34974 8576 34980 8628
rect 35032 8576 35038 8628
rect 36722 8576 36728 8628
rect 36780 8616 36786 8628
rect 36909 8619 36967 8625
rect 36909 8616 36921 8619
rect 36780 8588 36921 8616
rect 36780 8576 36786 8588
rect 36909 8585 36921 8588
rect 36955 8585 36967 8619
rect 36909 8579 36967 8585
rect 38930 8576 38936 8628
rect 38988 8616 38994 8628
rect 39117 8619 39175 8625
rect 39117 8616 39129 8619
rect 38988 8588 39129 8616
rect 38988 8576 38994 8588
rect 39117 8585 39129 8588
rect 39163 8585 39175 8619
rect 39117 8579 39175 8585
rect 41138 8576 41144 8628
rect 41196 8576 41202 8628
rect 43346 8576 43352 8628
rect 43404 8616 43410 8628
rect 43533 8619 43591 8625
rect 43533 8616 43545 8619
rect 43404 8588 43545 8616
rect 43404 8576 43410 8588
rect 43533 8585 43545 8588
rect 43579 8585 43591 8619
rect 43533 8579 43591 8585
rect 45373 8619 45431 8625
rect 45373 8585 45385 8619
rect 45419 8616 45431 8619
rect 45554 8616 45560 8628
rect 45419 8588 45560 8616
rect 45419 8585 45431 8588
rect 45373 8579 45431 8585
rect 45554 8576 45560 8588
rect 45612 8576 45618 8628
rect 1394 8508 1400 8560
rect 1452 8508 1458 8560
rect 1765 8551 1823 8557
rect 1765 8517 1777 8551
rect 1811 8548 1823 8551
rect 10152 8548 10180 8576
rect 23106 8548 23112 8560
rect 1811 8520 10180 8548
rect 10520 8520 23112 8548
rect 1811 8517 1823 8520
rect 1765 8511 1823 8517
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4080 8412 4108 8443
rect 6178 8440 6184 8492
rect 6236 8440 6242 8492
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 10520 8480 10548 8520
rect 23106 8508 23112 8520
rect 23164 8508 23170 8560
rect 8343 8452 10548 8480
rect 10597 8483 10655 8489
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 12713 8483 12771 8489
rect 12713 8449 12725 8483
rect 12759 8480 12771 8483
rect 14918 8480 14924 8492
rect 12759 8452 14924 8480
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 6270 8412 6276 8424
rect 4080 8384 6276 8412
rect 6270 8372 6276 8384
rect 6328 8372 6334 8424
rect 10612 8344 10640 8443
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 15028 8412 15056 8443
rect 17218 8440 17224 8492
rect 17276 8440 17282 8492
rect 19610 8440 19616 8492
rect 19668 8440 19674 8492
rect 21634 8440 21640 8492
rect 21692 8440 21698 8492
rect 23750 8440 23756 8492
rect 23808 8440 23814 8492
rect 26050 8440 26056 8492
rect 26108 8440 26114 8492
rect 28258 8440 28264 8492
rect 28316 8440 28322 8492
rect 30374 8440 30380 8492
rect 30432 8440 30438 8492
rect 32674 8440 32680 8492
rect 32732 8440 32738 8492
rect 35066 8440 35072 8492
rect 35124 8440 35130 8492
rect 37090 8440 37096 8492
rect 37148 8440 37154 8492
rect 39298 8440 39304 8492
rect 39356 8440 39362 8492
rect 41414 8440 41420 8492
rect 41472 8440 41478 8492
rect 43714 8440 43720 8492
rect 43772 8440 43778 8492
rect 45094 8440 45100 8492
rect 45152 8440 45158 8492
rect 19978 8412 19984 8424
rect 15028 8384 19984 8412
rect 19978 8372 19984 8384
rect 20036 8372 20042 8424
rect 23658 8344 23664 8356
rect 10612 8316 23664 8344
rect 23658 8304 23664 8316
rect 23716 8304 23722 8356
rect 1104 8186 45816 8208
rect 1104 8134 6539 8186
rect 6591 8134 6603 8186
rect 6655 8134 6667 8186
rect 6719 8134 6731 8186
rect 6783 8134 6795 8186
rect 6847 8134 17717 8186
rect 17769 8134 17781 8186
rect 17833 8134 17845 8186
rect 17897 8134 17909 8186
rect 17961 8134 17973 8186
rect 18025 8134 28895 8186
rect 28947 8134 28959 8186
rect 29011 8134 29023 8186
rect 29075 8134 29087 8186
rect 29139 8134 29151 8186
rect 29203 8134 40073 8186
rect 40125 8134 40137 8186
rect 40189 8134 40201 8186
rect 40253 8134 40265 8186
rect 40317 8134 40329 8186
rect 40381 8134 45816 8186
rect 1104 8112 45816 8134
rect 1104 7642 45976 7664
rect 1104 7590 12128 7642
rect 12180 7590 12192 7642
rect 12244 7590 12256 7642
rect 12308 7590 12320 7642
rect 12372 7590 12384 7642
rect 12436 7590 23306 7642
rect 23358 7590 23370 7642
rect 23422 7590 23434 7642
rect 23486 7590 23498 7642
rect 23550 7590 23562 7642
rect 23614 7590 34484 7642
rect 34536 7590 34548 7642
rect 34600 7590 34612 7642
rect 34664 7590 34676 7642
rect 34728 7590 34740 7642
rect 34792 7590 45662 7642
rect 45714 7590 45726 7642
rect 45778 7590 45790 7642
rect 45842 7590 45854 7642
rect 45906 7590 45918 7642
rect 45970 7590 45976 7642
rect 1104 7568 45976 7590
rect 1104 7098 45816 7120
rect 1104 7046 6539 7098
rect 6591 7046 6603 7098
rect 6655 7046 6667 7098
rect 6719 7046 6731 7098
rect 6783 7046 6795 7098
rect 6847 7046 17717 7098
rect 17769 7046 17781 7098
rect 17833 7046 17845 7098
rect 17897 7046 17909 7098
rect 17961 7046 17973 7098
rect 18025 7046 28895 7098
rect 28947 7046 28959 7098
rect 29011 7046 29023 7098
rect 29075 7046 29087 7098
rect 29139 7046 29151 7098
rect 29203 7046 40073 7098
rect 40125 7046 40137 7098
rect 40189 7046 40201 7098
rect 40253 7046 40265 7098
rect 40317 7046 40329 7098
rect 40381 7046 45816 7098
rect 1104 7024 45816 7046
rect 1104 6554 45976 6576
rect 1104 6502 12128 6554
rect 12180 6502 12192 6554
rect 12244 6502 12256 6554
rect 12308 6502 12320 6554
rect 12372 6502 12384 6554
rect 12436 6502 23306 6554
rect 23358 6502 23370 6554
rect 23422 6502 23434 6554
rect 23486 6502 23498 6554
rect 23550 6502 23562 6554
rect 23614 6502 34484 6554
rect 34536 6502 34548 6554
rect 34600 6502 34612 6554
rect 34664 6502 34676 6554
rect 34728 6502 34740 6554
rect 34792 6502 45662 6554
rect 45714 6502 45726 6554
rect 45778 6502 45790 6554
rect 45842 6502 45854 6554
rect 45906 6502 45918 6554
rect 45970 6502 45976 6554
rect 1104 6480 45976 6502
rect 1104 6010 45816 6032
rect 1104 5958 6539 6010
rect 6591 5958 6603 6010
rect 6655 5958 6667 6010
rect 6719 5958 6731 6010
rect 6783 5958 6795 6010
rect 6847 5958 17717 6010
rect 17769 5958 17781 6010
rect 17833 5958 17845 6010
rect 17897 5958 17909 6010
rect 17961 5958 17973 6010
rect 18025 5958 28895 6010
rect 28947 5958 28959 6010
rect 29011 5958 29023 6010
rect 29075 5958 29087 6010
rect 29139 5958 29151 6010
rect 29203 5958 40073 6010
rect 40125 5958 40137 6010
rect 40189 5958 40201 6010
rect 40253 5958 40265 6010
rect 40317 5958 40329 6010
rect 40381 5958 45816 6010
rect 1104 5936 45816 5958
rect 1104 5466 45976 5488
rect 1104 5414 12128 5466
rect 12180 5414 12192 5466
rect 12244 5414 12256 5466
rect 12308 5414 12320 5466
rect 12372 5414 12384 5466
rect 12436 5414 23306 5466
rect 23358 5414 23370 5466
rect 23422 5414 23434 5466
rect 23486 5414 23498 5466
rect 23550 5414 23562 5466
rect 23614 5414 34484 5466
rect 34536 5414 34548 5466
rect 34600 5414 34612 5466
rect 34664 5414 34676 5466
rect 34728 5414 34740 5466
rect 34792 5414 45662 5466
rect 45714 5414 45726 5466
rect 45778 5414 45790 5466
rect 45842 5414 45854 5466
rect 45906 5414 45918 5466
rect 45970 5414 45976 5466
rect 1104 5392 45976 5414
rect 1104 4922 45816 4944
rect 1104 4870 6539 4922
rect 6591 4870 6603 4922
rect 6655 4870 6667 4922
rect 6719 4870 6731 4922
rect 6783 4870 6795 4922
rect 6847 4870 17717 4922
rect 17769 4870 17781 4922
rect 17833 4870 17845 4922
rect 17897 4870 17909 4922
rect 17961 4870 17973 4922
rect 18025 4870 28895 4922
rect 28947 4870 28959 4922
rect 29011 4870 29023 4922
rect 29075 4870 29087 4922
rect 29139 4870 29151 4922
rect 29203 4870 40073 4922
rect 40125 4870 40137 4922
rect 40189 4870 40201 4922
rect 40253 4870 40265 4922
rect 40317 4870 40329 4922
rect 40381 4870 45816 4922
rect 1104 4848 45816 4870
rect 4982 4496 4988 4548
rect 5040 4536 5046 4548
rect 26142 4536 26148 4548
rect 5040 4508 26148 4536
rect 5040 4496 5046 4508
rect 26142 4496 26148 4508
rect 26200 4496 26206 4548
rect 9398 4428 9404 4480
rect 9456 4468 9462 4480
rect 32122 4468 32128 4480
rect 9456 4440 32128 4468
rect 9456 4428 9462 4440
rect 32122 4428 32128 4440
rect 32180 4428 32186 4480
rect 1104 4378 45976 4400
rect 1104 4326 12128 4378
rect 12180 4326 12192 4378
rect 12244 4326 12256 4378
rect 12308 4326 12320 4378
rect 12372 4326 12384 4378
rect 12436 4326 23306 4378
rect 23358 4326 23370 4378
rect 23422 4326 23434 4378
rect 23486 4326 23498 4378
rect 23550 4326 23562 4378
rect 23614 4326 34484 4378
rect 34536 4326 34548 4378
rect 34600 4326 34612 4378
rect 34664 4326 34676 4378
rect 34728 4326 34740 4378
rect 34792 4326 45662 4378
rect 45714 4326 45726 4378
rect 45778 4326 45790 4378
rect 45842 4326 45854 4378
rect 45906 4326 45918 4378
rect 45970 4326 45976 4378
rect 1104 4304 45976 4326
rect 18782 4224 18788 4276
rect 18840 4264 18846 4276
rect 41598 4264 41604 4276
rect 18840 4236 41604 4264
rect 18840 4224 18846 4236
rect 41598 4224 41604 4236
rect 41656 4224 41662 4276
rect 2774 4156 2780 4208
rect 2832 4196 2838 4208
rect 26418 4196 26424 4208
rect 2832 4168 26424 4196
rect 2832 4156 2838 4168
rect 26418 4156 26424 4168
rect 26476 4156 26482 4208
rect 1104 3834 45816 3856
rect 1104 3782 6539 3834
rect 6591 3782 6603 3834
rect 6655 3782 6667 3834
rect 6719 3782 6731 3834
rect 6783 3782 6795 3834
rect 6847 3782 17717 3834
rect 17769 3782 17781 3834
rect 17833 3782 17845 3834
rect 17897 3782 17909 3834
rect 17961 3782 17973 3834
rect 18025 3782 28895 3834
rect 28947 3782 28959 3834
rect 29011 3782 29023 3834
rect 29075 3782 29087 3834
rect 29139 3782 29151 3834
rect 29203 3782 40073 3834
rect 40125 3782 40137 3834
rect 40189 3782 40201 3834
rect 40253 3782 40265 3834
rect 40317 3782 40329 3834
rect 40381 3782 45816 3834
rect 1104 3760 45816 3782
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 22462 3584 22468 3596
rect 6972 3556 22468 3584
rect 6972 3544 6978 3556
rect 22462 3544 22468 3556
rect 22520 3544 22526 3596
rect 17126 3476 17132 3528
rect 17184 3516 17190 3528
rect 36630 3516 36636 3528
rect 17184 3488 36636 3516
rect 17184 3476 17190 3488
rect 36630 3476 36636 3488
rect 36688 3476 36694 3528
rect 21818 3408 21824 3460
rect 21876 3448 21882 3460
rect 31754 3448 31760 3460
rect 21876 3420 31760 3448
rect 21876 3408 21882 3420
rect 31754 3408 31760 3420
rect 31812 3408 31818 3460
rect 19150 3340 19156 3392
rect 19208 3380 19214 3392
rect 38654 3380 38660 3392
rect 19208 3352 38660 3380
rect 19208 3340 19214 3352
rect 38654 3340 38660 3352
rect 38712 3340 38718 3392
rect 1104 3290 45976 3312
rect 1104 3238 12128 3290
rect 12180 3238 12192 3290
rect 12244 3238 12256 3290
rect 12308 3238 12320 3290
rect 12372 3238 12384 3290
rect 12436 3238 23306 3290
rect 23358 3238 23370 3290
rect 23422 3238 23434 3290
rect 23486 3238 23498 3290
rect 23550 3238 23562 3290
rect 23614 3238 34484 3290
rect 34536 3238 34548 3290
rect 34600 3238 34612 3290
rect 34664 3238 34676 3290
rect 34728 3238 34740 3290
rect 34792 3238 45662 3290
rect 45714 3238 45726 3290
rect 45778 3238 45790 3290
rect 45842 3238 45854 3290
rect 45906 3238 45918 3290
rect 45970 3238 45976 3290
rect 1104 3216 45976 3238
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 24486 3176 24492 3188
rect 11204 3148 24492 3176
rect 11204 3136 11210 3148
rect 24486 3136 24492 3148
rect 24544 3136 24550 3188
rect 11422 3068 11428 3120
rect 11480 3108 11486 3120
rect 26326 3108 26332 3120
rect 11480 3080 26332 3108
rect 11480 3068 11486 3080
rect 26326 3068 26332 3080
rect 26384 3068 26390 3120
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 23198 3040 23204 3052
rect 8536 3012 23204 3040
rect 8536 3000 8542 3012
rect 23198 3000 23204 3012
rect 23256 3000 23262 3052
rect 23842 3000 23848 3052
rect 23900 3040 23906 3052
rect 35526 3040 35532 3052
rect 23900 3012 35532 3040
rect 23900 3000 23906 3012
rect 35526 3000 35532 3012
rect 35584 3000 35590 3052
rect 16482 2932 16488 2984
rect 16540 2972 16546 2984
rect 35710 2972 35716 2984
rect 16540 2944 35716 2972
rect 16540 2932 16546 2944
rect 35710 2932 35716 2944
rect 35768 2932 35774 2984
rect 5626 2864 5632 2916
rect 5684 2904 5690 2916
rect 20530 2904 20536 2916
rect 5684 2876 20536 2904
rect 5684 2864 5690 2876
rect 20530 2864 20536 2876
rect 20588 2864 20594 2916
rect 34330 2904 34336 2916
rect 30024 2876 34336 2904
rect 30024 2848 30052 2876
rect 34330 2864 34336 2876
rect 34388 2864 34394 2916
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 19242 2836 19248 2848
rect 14608 2808 19248 2836
rect 14608 2796 14614 2808
rect 19242 2796 19248 2808
rect 19300 2796 19306 2848
rect 26694 2796 26700 2848
rect 26752 2836 26758 2848
rect 27706 2836 27712 2848
rect 26752 2808 27712 2836
rect 26752 2796 26758 2808
rect 27706 2796 27712 2808
rect 27764 2796 27770 2848
rect 30006 2796 30012 2848
rect 30064 2796 30070 2848
rect 30098 2796 30104 2848
rect 30156 2836 30162 2848
rect 31846 2836 31852 2848
rect 30156 2808 31852 2836
rect 30156 2796 30162 2808
rect 31846 2796 31852 2808
rect 31904 2796 31910 2848
rect 32582 2796 32588 2848
rect 32640 2836 32646 2848
rect 37458 2836 37464 2848
rect 32640 2808 37464 2836
rect 32640 2796 32646 2808
rect 37458 2796 37464 2808
rect 37516 2796 37522 2848
rect 1104 2746 45816 2768
rect 1104 2694 6539 2746
rect 6591 2694 6603 2746
rect 6655 2694 6667 2746
rect 6719 2694 6731 2746
rect 6783 2694 6795 2746
rect 6847 2694 17717 2746
rect 17769 2694 17781 2746
rect 17833 2694 17845 2746
rect 17897 2694 17909 2746
rect 17961 2694 17973 2746
rect 18025 2694 28895 2746
rect 28947 2694 28959 2746
rect 29011 2694 29023 2746
rect 29075 2694 29087 2746
rect 29139 2694 29151 2746
rect 29203 2694 40073 2746
rect 40125 2694 40137 2746
rect 40189 2694 40201 2746
rect 40253 2694 40265 2746
rect 40317 2694 40329 2746
rect 40381 2694 45816 2746
rect 1104 2672 45816 2694
rect 17218 2592 17224 2644
rect 17276 2632 17282 2644
rect 17405 2635 17463 2641
rect 17405 2632 17417 2635
rect 17276 2604 17417 2632
rect 17276 2592 17282 2604
rect 17405 2601 17417 2604
rect 17451 2601 17463 2635
rect 17405 2595 17463 2601
rect 19168 2604 22692 2632
rect 18693 2567 18751 2573
rect 18693 2533 18705 2567
rect 18739 2564 18751 2567
rect 19168 2564 19196 2604
rect 18739 2536 19196 2564
rect 18739 2533 18751 2536
rect 18693 2527 18751 2533
rect 19610 2524 19616 2576
rect 19668 2524 19674 2576
rect 20438 2524 20444 2576
rect 20496 2524 20502 2576
rect 21361 2567 21419 2573
rect 21361 2533 21373 2567
rect 21407 2564 21419 2567
rect 22186 2564 22192 2576
rect 21407 2536 22192 2564
rect 21407 2533 21419 2536
rect 21361 2527 21419 2533
rect 22186 2524 22192 2536
rect 22244 2524 22250 2576
rect 22664 2564 22692 2604
rect 22738 2592 22744 2644
rect 22796 2592 22802 2644
rect 23014 2592 23020 2644
rect 23072 2592 23078 2644
rect 23106 2592 23112 2644
rect 23164 2632 23170 2644
rect 23293 2635 23351 2641
rect 23293 2632 23305 2635
rect 23164 2604 23305 2632
rect 23164 2592 23170 2604
rect 23293 2601 23305 2604
rect 23339 2601 23351 2635
rect 23293 2595 23351 2601
rect 23569 2635 23627 2641
rect 23569 2601 23581 2635
rect 23615 2632 23627 2635
rect 23658 2632 23664 2644
rect 23615 2604 23664 2632
rect 23615 2601 23627 2604
rect 23569 2595 23627 2601
rect 23658 2592 23664 2604
rect 23716 2592 23722 2644
rect 23750 2592 23756 2644
rect 23808 2592 23814 2644
rect 23934 2592 23940 2644
rect 23992 2592 23998 2644
rect 24026 2592 24032 2644
rect 24084 2632 24090 2644
rect 26878 2632 26884 2644
rect 24084 2604 26884 2632
rect 24084 2592 24090 2604
rect 26878 2592 26884 2604
rect 26936 2592 26942 2644
rect 27540 2604 27752 2632
rect 23768 2564 23796 2592
rect 24397 2567 24455 2573
rect 24397 2564 24409 2567
rect 22664 2536 23336 2564
rect 23768 2536 24409 2564
rect 15010 2456 15016 2508
rect 15068 2496 15074 2508
rect 20456 2496 20484 2524
rect 15068 2468 20208 2496
rect 20456 2468 21956 2496
rect 15068 2456 15074 2468
rect 14734 2388 14740 2440
rect 14792 2428 14798 2440
rect 17494 2428 17500 2440
rect 14792 2400 17500 2428
rect 14792 2388 14798 2400
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 17586 2388 17592 2440
rect 17644 2388 17650 2440
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18509 2431 18567 2437
rect 18509 2428 18521 2431
rect 18104 2400 18521 2428
rect 18104 2388 18110 2400
rect 18509 2397 18521 2400
rect 18555 2397 18567 2431
rect 18509 2391 18567 2397
rect 18690 2388 18696 2440
rect 18748 2428 18754 2440
rect 18877 2431 18935 2437
rect 18877 2428 18889 2431
rect 18748 2400 18889 2428
rect 18748 2388 18754 2400
rect 18877 2397 18889 2400
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 18966 2388 18972 2440
rect 19024 2428 19030 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19024 2400 19441 2428
rect 19024 2388 19030 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 19702 2388 19708 2440
rect 19760 2388 19766 2440
rect 20070 2428 20076 2440
rect 19812 2400 20076 2428
rect 14274 2320 14280 2372
rect 14332 2360 14338 2372
rect 19628 2360 19656 2388
rect 14332 2332 19656 2360
rect 14332 2320 14338 2332
rect 12618 2252 12624 2304
rect 12676 2292 12682 2304
rect 17678 2292 17684 2304
rect 12676 2264 17684 2292
rect 12676 2252 12682 2264
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 19058 2252 19064 2304
rect 19116 2252 19122 2304
rect 19242 2252 19248 2304
rect 19300 2292 19306 2304
rect 19812 2292 19840 2400
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 19978 2320 19984 2372
rect 20036 2360 20042 2372
rect 20036 2332 20116 2360
rect 20036 2320 20042 2332
rect 19300 2264 19840 2292
rect 19300 2252 19306 2264
rect 19886 2252 19892 2304
rect 19944 2252 19950 2304
rect 20088 2301 20116 2332
rect 20180 2304 20208 2468
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 20272 2304 20300 2391
rect 20346 2388 20352 2440
rect 20404 2428 20410 2440
rect 20441 2431 20499 2437
rect 20441 2428 20453 2431
rect 20404 2400 20453 2428
rect 20404 2388 20410 2400
rect 20441 2397 20453 2400
rect 20487 2397 20499 2431
rect 20441 2391 20499 2397
rect 20898 2388 20904 2440
rect 20956 2388 20962 2440
rect 21174 2388 21180 2440
rect 21232 2388 21238 2440
rect 21634 2388 21640 2440
rect 21692 2388 21698 2440
rect 21928 2437 21956 2468
rect 22646 2456 22652 2508
rect 22704 2496 22710 2508
rect 23308 2496 23336 2536
rect 24397 2533 24409 2536
rect 24443 2533 24455 2567
rect 24397 2527 24455 2533
rect 26050 2524 26056 2576
rect 26108 2524 26114 2576
rect 26513 2567 26571 2573
rect 26513 2533 26525 2567
rect 26559 2564 26571 2567
rect 27540 2564 27568 2604
rect 26559 2536 27568 2564
rect 27724 2564 27752 2604
rect 28258 2592 28264 2644
rect 28316 2592 28322 2644
rect 31478 2632 31484 2644
rect 30208 2604 31484 2632
rect 30208 2564 30236 2604
rect 31478 2592 31484 2604
rect 31536 2592 31542 2644
rect 31662 2592 31668 2644
rect 31720 2632 31726 2644
rect 31720 2604 32628 2632
rect 31720 2592 31726 2604
rect 27724 2536 30236 2564
rect 30285 2567 30343 2573
rect 26559 2533 26571 2536
rect 26513 2527 26571 2533
rect 30285 2533 30297 2567
rect 30331 2564 30343 2567
rect 31938 2564 31944 2576
rect 30331 2536 31944 2564
rect 30331 2533 30343 2536
rect 30285 2527 30343 2533
rect 31938 2524 31944 2536
rect 31996 2524 32002 2576
rect 32600 2564 32628 2604
rect 32674 2592 32680 2644
rect 32732 2592 32738 2644
rect 35066 2592 35072 2644
rect 35124 2592 35130 2644
rect 36906 2592 36912 2644
rect 36964 2632 36970 2644
rect 37093 2635 37151 2641
rect 37093 2632 37105 2635
rect 36964 2604 37105 2632
rect 36964 2592 36970 2604
rect 37093 2601 37105 2604
rect 37139 2601 37151 2635
rect 37093 2595 37151 2601
rect 37182 2592 37188 2644
rect 37240 2632 37246 2644
rect 37550 2632 37556 2644
rect 37240 2604 37556 2632
rect 37240 2592 37246 2604
rect 37550 2592 37556 2604
rect 37608 2592 37614 2644
rect 39482 2592 39488 2644
rect 39540 2592 39546 2644
rect 39684 2604 41368 2632
rect 33134 2564 33140 2576
rect 32600 2536 33140 2564
rect 33134 2524 33140 2536
rect 33192 2524 33198 2576
rect 34330 2524 34336 2576
rect 34388 2564 34394 2576
rect 39574 2564 39580 2576
rect 34388 2536 39580 2564
rect 34388 2524 34394 2536
rect 39574 2524 39580 2536
rect 39632 2524 39638 2576
rect 24118 2496 24124 2508
rect 22704 2468 23244 2496
rect 23308 2468 24124 2496
rect 22704 2456 22710 2468
rect 21821 2431 21879 2437
rect 21821 2397 21833 2431
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 21913 2431 21971 2437
rect 21913 2397 21925 2431
rect 21959 2397 21971 2431
rect 21913 2391 21971 2397
rect 20073 2295 20131 2301
rect 20073 2261 20085 2295
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 20162 2252 20168 2304
rect 20220 2252 20226 2304
rect 20254 2252 20260 2304
rect 20312 2252 20318 2304
rect 20622 2252 20628 2304
rect 20680 2252 20686 2304
rect 21082 2252 21088 2304
rect 21140 2252 21146 2304
rect 21652 2301 21680 2388
rect 21836 2360 21864 2391
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 22373 2431 22431 2437
rect 22373 2428 22385 2431
rect 22336 2400 22385 2428
rect 22336 2388 22342 2400
rect 22373 2397 22385 2400
rect 22419 2397 22431 2431
rect 22373 2391 22431 2397
rect 22462 2388 22468 2440
rect 22520 2388 22526 2440
rect 22922 2388 22928 2440
rect 22980 2388 22986 2440
rect 23014 2388 23020 2440
rect 23072 2428 23078 2440
rect 23216 2437 23244 2468
rect 24118 2456 24124 2468
rect 24176 2456 24182 2508
rect 26528 2468 27200 2496
rect 23201 2431 23259 2437
rect 23072 2400 23152 2428
rect 23072 2388 23078 2400
rect 23124 2360 23152 2400
rect 23201 2397 23213 2431
rect 23247 2397 23259 2431
rect 23201 2391 23259 2397
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 23492 2360 23520 2391
rect 23750 2388 23756 2440
rect 23808 2388 23814 2440
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 26237 2431 26295 2437
rect 26237 2397 26249 2431
rect 26283 2397 26295 2431
rect 26237 2391 26295 2397
rect 21836 2332 22232 2360
rect 23124 2332 23520 2360
rect 24029 2363 24087 2369
rect 21637 2295 21695 2301
rect 21637 2261 21649 2295
rect 21683 2261 21695 2295
rect 21637 2255 21695 2261
rect 22094 2252 22100 2304
rect 22152 2252 22158 2304
rect 22204 2301 22232 2332
rect 24029 2329 24041 2363
rect 24075 2360 24087 2363
rect 25038 2360 25044 2372
rect 24075 2332 25044 2360
rect 24075 2329 24087 2332
rect 24029 2323 24087 2329
rect 25038 2320 25044 2332
rect 25096 2320 25102 2372
rect 26252 2360 26280 2391
rect 26326 2388 26332 2440
rect 26384 2388 26390 2440
rect 26528 2360 26556 2468
rect 26602 2388 26608 2440
rect 26660 2388 26666 2440
rect 26878 2388 26884 2440
rect 26936 2388 26942 2440
rect 26252 2332 26556 2360
rect 22189 2295 22247 2301
rect 22189 2261 22201 2295
rect 22235 2261 22247 2295
rect 22189 2255 22247 2261
rect 22649 2295 22707 2301
rect 22649 2261 22661 2295
rect 22695 2292 22707 2295
rect 22738 2292 22744 2304
rect 22695 2264 22744 2292
rect 22695 2261 22707 2264
rect 22649 2255 22707 2261
rect 22738 2252 22744 2264
rect 22796 2252 22802 2304
rect 26786 2252 26792 2304
rect 26844 2252 26850 2304
rect 27062 2252 27068 2304
rect 27120 2252 27126 2304
rect 27172 2301 27200 2468
rect 27706 2456 27712 2508
rect 27764 2496 27770 2508
rect 30926 2496 30932 2508
rect 27764 2468 30932 2496
rect 27764 2456 27770 2468
rect 30926 2456 30932 2468
rect 30984 2456 30990 2508
rect 31478 2456 31484 2508
rect 31536 2456 31542 2508
rect 31754 2456 31760 2508
rect 31812 2496 31818 2508
rect 39684 2496 39712 2604
rect 41340 2564 41368 2604
rect 41414 2592 41420 2644
rect 41472 2632 41478 2644
rect 41601 2635 41659 2641
rect 41601 2632 41613 2635
rect 41472 2604 41613 2632
rect 41472 2592 41478 2604
rect 41601 2601 41613 2604
rect 41647 2601 41659 2635
rect 41601 2595 41659 2601
rect 43714 2592 43720 2644
rect 43772 2632 43778 2644
rect 43993 2635 44051 2641
rect 43993 2632 44005 2635
rect 43772 2604 44005 2632
rect 43772 2592 43778 2604
rect 43993 2601 44005 2604
rect 44039 2601 44051 2635
rect 43993 2595 44051 2601
rect 44821 2635 44879 2641
rect 44821 2601 44833 2635
rect 44867 2632 44879 2635
rect 45094 2632 45100 2644
rect 44867 2604 45100 2632
rect 44867 2601 44879 2604
rect 44821 2595 44879 2601
rect 45094 2592 45100 2604
rect 45152 2592 45158 2644
rect 41340 2536 41414 2564
rect 31812 2468 32444 2496
rect 31812 2456 31818 2468
rect 27341 2431 27399 2437
rect 27341 2397 27353 2431
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 27356 2360 27384 2391
rect 27430 2388 27436 2440
rect 27488 2388 27494 2440
rect 27614 2388 27620 2440
rect 27672 2428 27678 2440
rect 27893 2431 27951 2437
rect 27893 2428 27905 2431
rect 27672 2400 27905 2428
rect 27672 2388 27678 2400
rect 27893 2397 27905 2400
rect 27939 2397 27951 2431
rect 27893 2391 27951 2397
rect 28442 2388 28448 2440
rect 28500 2388 28506 2440
rect 29822 2388 29828 2440
rect 29880 2428 29886 2440
rect 30101 2431 30159 2437
rect 30101 2428 30113 2431
rect 29880 2400 30113 2428
rect 29880 2388 29886 2400
rect 30101 2397 30113 2400
rect 30147 2397 30159 2431
rect 30101 2391 30159 2397
rect 30653 2431 30711 2437
rect 30653 2397 30665 2431
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 28810 2360 28816 2372
rect 27356 2332 28816 2360
rect 28810 2320 28816 2332
rect 28868 2320 28874 2372
rect 28902 2320 28908 2372
rect 28960 2360 28966 2372
rect 30282 2360 30288 2372
rect 28960 2332 30288 2360
rect 28960 2320 28966 2332
rect 30282 2320 30288 2332
rect 30340 2320 30346 2372
rect 30668 2360 30696 2391
rect 30742 2388 30748 2440
rect 30800 2388 30806 2440
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 31113 2431 31171 2437
rect 31113 2428 31125 2431
rect 30892 2400 31125 2428
rect 30892 2388 30898 2400
rect 31113 2397 31125 2400
rect 31159 2397 31171 2431
rect 31113 2391 31171 2397
rect 31386 2388 31392 2440
rect 31444 2388 31450 2440
rect 31496 2428 31524 2456
rect 32030 2428 32036 2440
rect 31496 2400 32036 2428
rect 32030 2388 32036 2400
rect 32088 2388 32094 2440
rect 32125 2431 32183 2437
rect 32125 2397 32137 2431
rect 32171 2428 32183 2431
rect 32214 2428 32220 2440
rect 32171 2400 32220 2428
rect 32171 2397 32183 2400
rect 32125 2391 32183 2397
rect 32214 2388 32220 2400
rect 32272 2388 32278 2440
rect 32306 2388 32312 2440
rect 32364 2388 32370 2440
rect 32324 2360 32352 2388
rect 30668 2332 32352 2360
rect 32416 2360 32444 2468
rect 35360 2468 39712 2496
rect 41386 2496 41414 2536
rect 44450 2496 44456 2508
rect 41386 2468 44456 2496
rect 35360 2440 35388 2468
rect 44450 2456 44456 2468
rect 44508 2456 44514 2508
rect 32861 2431 32919 2437
rect 32861 2397 32873 2431
rect 32907 2428 32919 2431
rect 33226 2428 33232 2440
rect 32907 2400 33232 2428
rect 32907 2397 32919 2400
rect 32861 2391 32919 2397
rect 33226 2388 33232 2400
rect 33284 2388 33290 2440
rect 33413 2431 33471 2437
rect 33413 2397 33425 2431
rect 33459 2397 33471 2431
rect 33413 2391 33471 2397
rect 33428 2360 33456 2391
rect 34882 2388 34888 2440
rect 34940 2388 34946 2440
rect 35342 2388 35348 2440
rect 35400 2388 35406 2440
rect 37182 2388 37188 2440
rect 37240 2388 37246 2440
rect 37277 2431 37335 2437
rect 37277 2397 37289 2431
rect 37323 2424 37335 2431
rect 37323 2397 37412 2424
rect 37277 2396 37412 2397
rect 37277 2391 37335 2396
rect 37200 2360 37228 2388
rect 32416 2332 33364 2360
rect 33428 2332 37228 2360
rect 27157 2295 27215 2301
rect 27157 2261 27169 2295
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 27617 2295 27675 2301
rect 27617 2261 27629 2295
rect 27663 2292 27675 2295
rect 27982 2292 27988 2304
rect 27663 2264 27988 2292
rect 27663 2261 27675 2264
rect 27617 2255 27675 2261
rect 27982 2252 27988 2264
rect 28040 2252 28046 2304
rect 28074 2252 28080 2304
rect 28132 2252 28138 2304
rect 30466 2252 30472 2304
rect 30524 2252 30530 2304
rect 30926 2252 30932 2304
rect 30984 2252 30990 2304
rect 31294 2252 31300 2304
rect 31352 2252 31358 2304
rect 31573 2295 31631 2301
rect 31573 2261 31585 2295
rect 31619 2292 31631 2295
rect 31754 2292 31760 2304
rect 31619 2264 31760 2292
rect 31619 2261 31631 2264
rect 31573 2255 31631 2261
rect 31754 2252 31760 2264
rect 31812 2252 31818 2304
rect 32309 2295 32367 2301
rect 32309 2261 32321 2295
rect 32355 2292 32367 2295
rect 32950 2292 32956 2304
rect 32355 2264 32956 2292
rect 32355 2261 32367 2264
rect 32309 2255 32367 2261
rect 32950 2252 32956 2264
rect 33008 2252 33014 2304
rect 33226 2252 33232 2304
rect 33284 2252 33290 2304
rect 33336 2292 33364 2332
rect 37384 2304 37412 2396
rect 37458 2388 37464 2440
rect 37516 2428 37522 2440
rect 38838 2428 38844 2440
rect 37516 2400 38844 2428
rect 37516 2388 37522 2400
rect 38838 2388 38844 2400
rect 38896 2388 38902 2440
rect 39666 2388 39672 2440
rect 39724 2388 39730 2440
rect 39758 2388 39764 2440
rect 39816 2428 39822 2440
rect 41506 2428 41512 2440
rect 39816 2400 41512 2428
rect 39816 2388 39822 2400
rect 41506 2388 41512 2400
rect 41564 2388 41570 2440
rect 41782 2388 41788 2440
rect 41840 2388 41846 2440
rect 44174 2388 44180 2440
rect 44232 2388 44238 2440
rect 44637 2431 44695 2437
rect 44637 2397 44649 2431
rect 44683 2428 44695 2431
rect 44910 2428 44916 2440
rect 44683 2400 44916 2428
rect 44683 2397 44695 2400
rect 44637 2391 44695 2397
rect 44910 2388 44916 2400
rect 44968 2388 44974 2440
rect 45186 2388 45192 2440
rect 45244 2388 45250 2440
rect 45465 2431 45523 2437
rect 45465 2397 45477 2431
rect 45511 2428 45523 2431
rect 45922 2428 45928 2440
rect 45511 2400 45928 2428
rect 45511 2397 45523 2400
rect 45465 2391 45523 2397
rect 45922 2388 45928 2400
rect 45980 2388 45986 2440
rect 37550 2320 37556 2372
rect 37608 2360 37614 2372
rect 41414 2360 41420 2372
rect 37608 2332 41420 2360
rect 37608 2320 37614 2332
rect 41414 2320 41420 2332
rect 41472 2320 41478 2372
rect 37182 2292 37188 2304
rect 33336 2264 37188 2292
rect 37182 2252 37188 2264
rect 37240 2252 37246 2304
rect 37366 2252 37372 2304
rect 37424 2252 37430 2304
rect 37826 2252 37832 2304
rect 37884 2292 37890 2304
rect 44266 2292 44272 2304
rect 37884 2264 44272 2292
rect 37884 2252 37890 2264
rect 44266 2252 44272 2264
rect 44324 2252 44330 2304
rect 45002 2252 45008 2304
rect 45060 2252 45066 2304
rect 45278 2252 45284 2304
rect 45336 2252 45342 2304
rect 1104 2202 45976 2224
rect 1104 2150 12128 2202
rect 12180 2150 12192 2202
rect 12244 2150 12256 2202
rect 12308 2150 12320 2202
rect 12372 2150 12384 2202
rect 12436 2150 23306 2202
rect 23358 2150 23370 2202
rect 23422 2150 23434 2202
rect 23486 2150 23498 2202
rect 23550 2150 23562 2202
rect 23614 2150 34484 2202
rect 34536 2150 34548 2202
rect 34600 2150 34612 2202
rect 34664 2150 34676 2202
rect 34728 2150 34740 2202
rect 34792 2150 45662 2202
rect 45714 2150 45726 2202
rect 45778 2150 45790 2202
rect 45842 2150 45854 2202
rect 45906 2150 45918 2202
rect 45970 2150 45976 2202
rect 1104 2128 45976 2150
rect 1857 2091 1915 2097
rect 1857 2057 1869 2091
rect 1903 2057 1915 2091
rect 1857 2051 1915 2057
rect 1872 2020 1900 2051
rect 2774 2048 2780 2100
rect 2832 2048 2838 2100
rect 3145 2091 3203 2097
rect 3145 2057 3157 2091
rect 3191 2088 3203 2091
rect 4982 2088 4988 2100
rect 3191 2060 4988 2088
rect 3191 2057 3203 2060
rect 3145 2051 3203 2057
rect 4982 2048 4988 2060
rect 5040 2048 5046 2100
rect 9398 2048 9404 2100
rect 9456 2048 9462 2100
rect 9582 2048 9588 2100
rect 9640 2048 9646 2100
rect 9769 2091 9827 2097
rect 9769 2057 9781 2091
rect 9815 2088 9827 2091
rect 13722 2088 13728 2100
rect 9815 2060 13728 2088
rect 9815 2057 9827 2060
rect 9769 2051 9827 2057
rect 13722 2048 13728 2060
rect 13780 2048 13786 2100
rect 15933 2091 15991 2097
rect 15933 2057 15945 2091
rect 15979 2057 15991 2091
rect 15933 2051 15991 2057
rect 9600 2020 9628 2048
rect 1872 1992 9628 2020
rect 15948 2020 15976 2051
rect 16206 2048 16212 2100
rect 16264 2048 16270 2100
rect 16482 2048 16488 2100
rect 16540 2048 16546 2100
rect 17037 2091 17095 2097
rect 17037 2057 17049 2091
rect 17083 2088 17095 2091
rect 17586 2088 17592 2100
rect 17083 2060 17592 2088
rect 17083 2057 17095 2060
rect 17037 2051 17095 2057
rect 17586 2048 17592 2060
rect 17644 2048 17650 2100
rect 18966 2048 18972 2100
rect 19024 2048 19030 2100
rect 19242 2048 19248 2100
rect 19300 2048 19306 2100
rect 19610 2048 19616 2100
rect 19668 2048 19674 2100
rect 19797 2091 19855 2097
rect 19797 2057 19809 2091
rect 19843 2088 19855 2091
rect 20070 2088 20076 2100
rect 19843 2060 20076 2088
rect 19843 2057 19855 2060
rect 19797 2051 19855 2057
rect 20070 2048 20076 2060
rect 20128 2048 20134 2100
rect 20622 2048 20628 2100
rect 20680 2048 20686 2100
rect 21082 2048 21088 2100
rect 21140 2048 21146 2100
rect 22097 2091 22155 2097
rect 22097 2057 22109 2091
rect 22143 2088 22155 2091
rect 22922 2088 22928 2100
rect 22143 2060 22928 2088
rect 22143 2057 22155 2060
rect 22097 2051 22155 2057
rect 22922 2048 22928 2060
rect 22980 2048 22986 2100
rect 23014 2048 23020 2100
rect 23072 2048 23078 2100
rect 23661 2091 23719 2097
rect 23661 2057 23673 2091
rect 23707 2088 23719 2091
rect 23750 2088 23756 2100
rect 23707 2060 23756 2088
rect 23707 2057 23719 2060
rect 23661 2051 23719 2057
rect 23750 2048 23756 2060
rect 23808 2048 23814 2100
rect 24578 2048 24584 2100
rect 24636 2088 24642 2100
rect 24765 2091 24823 2097
rect 24765 2088 24777 2091
rect 24636 2060 24777 2088
rect 24636 2048 24642 2060
rect 24765 2057 24777 2060
rect 24811 2057 24823 2091
rect 24765 2051 24823 2057
rect 25038 2048 25044 2100
rect 25096 2048 25102 2100
rect 25130 2048 25136 2100
rect 25188 2048 25194 2100
rect 25406 2048 25412 2100
rect 25464 2088 25470 2100
rect 25464 2060 28028 2088
rect 25464 2048 25470 2060
rect 17310 2020 17316 2032
rect 15948 1992 17316 2020
rect 17310 1980 17316 1992
rect 17368 1980 17374 2032
rect 17494 1980 17500 2032
rect 17552 2020 17558 2032
rect 19628 2020 19656 2048
rect 17552 1992 19656 2020
rect 17552 1980 17558 1992
rect 19702 1980 19708 2032
rect 19760 2020 19766 2032
rect 20640 2020 20668 2048
rect 21100 2020 21128 2048
rect 25148 2020 25176 2048
rect 26694 2020 26700 2032
rect 19760 1992 20024 2020
rect 19760 1980 19766 1992
rect 658 1912 664 1964
rect 716 1952 722 1964
rect 1397 1955 1455 1961
rect 1397 1952 1409 1955
rect 716 1924 1409 1952
rect 716 1912 722 1924
rect 1397 1921 1409 1924
rect 1443 1921 1455 1955
rect 1397 1915 1455 1921
rect 1673 1955 1731 1961
rect 1673 1921 1685 1955
rect 1719 1921 1731 1955
rect 1673 1915 1731 1921
rect 1026 1844 1032 1896
rect 1084 1884 1090 1896
rect 1688 1884 1716 1915
rect 2590 1912 2596 1964
rect 2648 1912 2654 1964
rect 2958 1912 2964 1964
rect 3016 1912 3022 1964
rect 9214 1912 9220 1964
rect 9272 1912 9278 1964
rect 9582 1912 9588 1964
rect 9640 1912 9646 1964
rect 15102 1912 15108 1964
rect 15160 1952 15166 1964
rect 15197 1955 15255 1961
rect 15197 1952 15209 1955
rect 15160 1924 15209 1952
rect 15160 1912 15166 1924
rect 15197 1921 15209 1924
rect 15243 1921 15255 1955
rect 15197 1915 15255 1921
rect 15470 1912 15476 1964
rect 15528 1912 15534 1964
rect 15746 1912 15752 1964
rect 15804 1912 15810 1964
rect 16022 1912 16028 1964
rect 16080 1912 16086 1964
rect 16298 1912 16304 1964
rect 16356 1912 16362 1964
rect 16850 1912 16856 1964
rect 16908 1912 16914 1964
rect 17126 1912 17132 1964
rect 17184 1912 17190 1964
rect 17402 1912 17408 1964
rect 17460 1912 17466 1964
rect 17678 1912 17684 1964
rect 17736 1912 17742 1964
rect 17957 1955 18015 1961
rect 17957 1921 17969 1955
rect 18003 1952 18015 1955
rect 18138 1952 18144 1964
rect 18003 1924 18144 1952
rect 18003 1921 18015 1924
rect 17957 1915 18015 1921
rect 18138 1912 18144 1924
rect 18196 1912 18202 1964
rect 18233 1955 18291 1961
rect 18233 1921 18245 1955
rect 18279 1921 18291 1955
rect 18233 1915 18291 1921
rect 1084 1856 1716 1884
rect 1084 1844 1090 1856
rect 16758 1844 16764 1896
rect 16816 1844 16822 1896
rect 16942 1844 16948 1896
rect 17000 1884 17006 1896
rect 18248 1884 18276 1915
rect 18506 1912 18512 1964
rect 18564 1912 18570 1964
rect 18782 1912 18788 1964
rect 18840 1912 18846 1964
rect 19058 1912 19064 1964
rect 19116 1912 19122 1964
rect 19334 1912 19340 1964
rect 19392 1912 19398 1964
rect 19610 1912 19616 1964
rect 19668 1912 19674 1964
rect 19889 1956 19947 1961
rect 19812 1955 19947 1956
rect 19812 1928 19901 1955
rect 17000 1856 18276 1884
rect 17000 1844 17006 1856
rect 18322 1844 18328 1896
rect 18380 1884 18386 1896
rect 19812 1884 19840 1928
rect 19889 1921 19901 1928
rect 19935 1921 19947 1955
rect 19889 1915 19947 1921
rect 18380 1856 19840 1884
rect 19996 1884 20024 1992
rect 20272 1992 20576 2020
rect 20640 1992 21036 2020
rect 21100 1992 22508 2020
rect 20272 1964 20300 1992
rect 20070 1912 20076 1964
rect 20128 1952 20134 1964
rect 20165 1955 20223 1961
rect 20165 1952 20177 1955
rect 20128 1924 20177 1952
rect 20128 1912 20134 1924
rect 20165 1921 20177 1924
rect 20211 1921 20223 1955
rect 20165 1915 20223 1921
rect 20254 1912 20260 1964
rect 20312 1912 20318 1964
rect 20441 1955 20499 1961
rect 20441 1921 20453 1955
rect 20487 1921 20499 1955
rect 20548 1952 20576 1992
rect 21008 1961 21036 1992
rect 20717 1955 20775 1961
rect 20717 1952 20729 1955
rect 20548 1924 20729 1952
rect 20441 1915 20499 1921
rect 20717 1921 20729 1924
rect 20763 1921 20775 1955
rect 20717 1915 20775 1921
rect 20993 1955 21051 1961
rect 20993 1921 21005 1955
rect 21039 1921 21051 1955
rect 20993 1915 21051 1921
rect 21453 1955 21511 1961
rect 21453 1921 21465 1955
rect 21499 1921 21511 1955
rect 21453 1915 21511 1921
rect 20456 1884 20484 1915
rect 19996 1856 20484 1884
rect 18380 1844 18386 1856
rect 20530 1844 20536 1896
rect 20588 1884 20594 1896
rect 21468 1884 21496 1915
rect 21726 1912 21732 1964
rect 21784 1952 21790 1964
rect 21913 1955 21971 1961
rect 21913 1952 21925 1955
rect 21784 1924 21925 1952
rect 21784 1912 21790 1924
rect 21913 1921 21925 1924
rect 21959 1921 21971 1955
rect 21913 1915 21971 1921
rect 22002 1912 22008 1964
rect 22060 1952 22066 1964
rect 22480 1961 22508 1992
rect 24136 1992 25176 2020
rect 25240 1992 26700 2020
rect 22189 1955 22247 1961
rect 22189 1952 22201 1955
rect 22060 1924 22201 1952
rect 22060 1912 22066 1924
rect 22189 1921 22201 1924
rect 22235 1921 22247 1955
rect 22189 1915 22247 1921
rect 22453 1955 22511 1961
rect 22453 1921 22465 1955
rect 22499 1921 22511 1955
rect 22453 1915 22511 1921
rect 22830 1912 22836 1964
rect 22888 1912 22894 1964
rect 22922 1912 22928 1964
rect 22980 1952 22986 1964
rect 23109 1955 23167 1961
rect 23109 1952 23121 1955
rect 22980 1924 23121 1952
rect 22980 1912 22986 1924
rect 23109 1921 23121 1924
rect 23155 1921 23167 1955
rect 23109 1915 23167 1921
rect 23382 1912 23388 1964
rect 23440 1912 23446 1964
rect 23842 1912 23848 1964
rect 23900 1912 23906 1964
rect 23937 1955 23995 1961
rect 23937 1921 23949 1955
rect 23983 1921 23995 1955
rect 23937 1915 23995 1921
rect 23952 1884 23980 1915
rect 20588 1856 21496 1884
rect 22020 1856 23980 1884
rect 20588 1844 20594 1856
rect 15381 1819 15439 1825
rect 15381 1785 15393 1819
rect 15427 1816 15439 1819
rect 16776 1816 16804 1844
rect 15427 1788 16804 1816
rect 17313 1819 17371 1825
rect 15427 1785 15439 1788
rect 15381 1779 15439 1785
rect 17313 1785 17325 1819
rect 17359 1816 17371 1819
rect 17865 1819 17923 1825
rect 17359 1788 17816 1816
rect 17359 1785 17371 1788
rect 17313 1779 17371 1785
rect 1578 1708 1584 1760
rect 1636 1708 1642 1760
rect 15654 1708 15660 1760
rect 15712 1708 15718 1760
rect 17494 1708 17500 1760
rect 17552 1748 17558 1760
rect 17589 1751 17647 1757
rect 17589 1748 17601 1751
rect 17552 1720 17601 1748
rect 17552 1708 17558 1720
rect 17589 1717 17601 1720
rect 17635 1717 17647 1751
rect 17788 1748 17816 1788
rect 17865 1785 17877 1819
rect 17911 1816 17923 1819
rect 18230 1816 18236 1828
rect 17911 1788 18236 1816
rect 17911 1785 17923 1788
rect 17865 1779 17923 1785
rect 18230 1776 18236 1788
rect 18288 1776 18294 1828
rect 18417 1819 18475 1825
rect 18417 1785 18429 1819
rect 18463 1816 18475 1819
rect 19334 1816 19340 1828
rect 18463 1788 19340 1816
rect 18463 1785 18475 1788
rect 18417 1779 18475 1785
rect 19334 1776 19340 1788
rect 19392 1776 19398 1828
rect 19521 1819 19579 1825
rect 19521 1785 19533 1819
rect 19567 1816 19579 1819
rect 20714 1816 20720 1828
rect 19567 1788 20720 1816
rect 19567 1785 19579 1788
rect 19521 1779 19579 1785
rect 20714 1776 20720 1788
rect 20772 1776 20778 1828
rect 21637 1819 21695 1825
rect 21637 1785 21649 1819
rect 21683 1816 21695 1819
rect 22020 1816 22048 1856
rect 21683 1788 22048 1816
rect 21683 1785 21695 1788
rect 21637 1779 21695 1785
rect 23474 1776 23480 1828
rect 23532 1816 23538 1828
rect 24136 1816 24164 1992
rect 24486 1912 24492 1964
rect 24544 1912 24550 1964
rect 24949 1955 25007 1961
rect 24949 1921 24961 1955
rect 24995 1952 25007 1955
rect 25130 1952 25136 1964
rect 24995 1924 25136 1952
rect 24995 1921 25007 1924
rect 24949 1915 25007 1921
rect 25130 1912 25136 1924
rect 25188 1912 25194 1964
rect 25240 1961 25268 1992
rect 26694 1980 26700 1992
rect 26752 1980 26758 2032
rect 26786 1980 26792 2032
rect 26844 2020 26850 2032
rect 28000 2020 28028 2060
rect 28442 2048 28448 2100
rect 28500 2088 28506 2100
rect 29917 2091 29975 2097
rect 29917 2088 29929 2091
rect 28500 2060 29929 2088
rect 28500 2048 28506 2060
rect 29917 2057 29929 2060
rect 29963 2057 29975 2091
rect 29917 2051 29975 2057
rect 30374 2048 30380 2100
rect 30432 2048 30438 2100
rect 30926 2048 30932 2100
rect 30984 2048 30990 2100
rect 31294 2048 31300 2100
rect 31352 2088 31358 2100
rect 31352 2060 31984 2088
rect 31352 2048 31358 2060
rect 30944 2020 30972 2048
rect 31021 2023 31079 2029
rect 31021 2020 31033 2023
rect 26844 1992 27936 2020
rect 28000 1992 28856 2020
rect 26844 1980 26850 1992
rect 25225 1955 25283 1961
rect 25225 1921 25237 1955
rect 25271 1921 25283 1955
rect 25225 1915 25283 1921
rect 25314 1912 25320 1964
rect 25372 1912 25378 1964
rect 25777 1955 25835 1961
rect 25777 1921 25789 1955
rect 25823 1921 25835 1955
rect 25777 1915 25835 1921
rect 25792 1884 25820 1915
rect 26142 1912 26148 1964
rect 26200 1912 26206 1964
rect 26418 1912 26424 1964
rect 26476 1912 26482 1964
rect 27908 1961 27936 1992
rect 26973 1955 27031 1961
rect 26973 1952 26985 1955
rect 26620 1924 26985 1952
rect 24688 1856 25820 1884
rect 24688 1825 24716 1856
rect 23532 1788 24164 1816
rect 24673 1819 24731 1825
rect 23532 1776 23538 1788
rect 24673 1785 24685 1819
rect 24719 1785 24731 1819
rect 24673 1779 24731 1785
rect 25314 1776 25320 1828
rect 25372 1816 25378 1828
rect 26620 1825 26648 1924
rect 26973 1921 26985 1924
rect 27019 1921 27031 1955
rect 26973 1915 27031 1921
rect 27709 1955 27767 1961
rect 27709 1921 27721 1955
rect 27755 1921 27767 1955
rect 27709 1915 27767 1921
rect 27893 1955 27951 1961
rect 27893 1921 27905 1955
rect 27939 1921 27951 1955
rect 27893 1915 27951 1921
rect 27522 1844 27528 1896
rect 27580 1844 27586 1896
rect 27724 1884 27752 1915
rect 28074 1912 28080 1964
rect 28132 1952 28138 1964
rect 28445 1955 28503 1961
rect 28445 1952 28457 1955
rect 28132 1924 28457 1952
rect 28132 1912 28138 1924
rect 28445 1921 28457 1924
rect 28491 1921 28503 1955
rect 28445 1915 28503 1921
rect 28534 1912 28540 1964
rect 28592 1952 28598 1964
rect 28828 1961 28856 1992
rect 28920 1992 29408 2020
rect 30944 1992 31033 2020
rect 28813 1955 28871 1961
rect 28592 1924 28764 1952
rect 28592 1912 28598 1924
rect 28350 1884 28356 1896
rect 27724 1856 28356 1884
rect 28350 1844 28356 1856
rect 28408 1844 28414 1896
rect 28736 1884 28764 1924
rect 28813 1921 28825 1955
rect 28859 1921 28871 1955
rect 28813 1915 28871 1921
rect 28920 1884 28948 1992
rect 29380 1961 29408 1992
rect 31021 1989 31033 1992
rect 31067 1989 31079 2023
rect 31956 2020 31984 2060
rect 32030 2048 32036 2100
rect 32088 2088 32094 2100
rect 32088 2060 34192 2088
rect 32088 2048 32094 2060
rect 32953 2023 33011 2029
rect 32953 2020 32965 2023
rect 31956 1992 32965 2020
rect 31021 1983 31079 1989
rect 32953 1989 32965 1992
rect 32999 1989 33011 2023
rect 32953 1983 33011 1989
rect 33134 1980 33140 2032
rect 33192 2020 33198 2032
rect 34164 2029 34192 2060
rect 34882 2048 34888 2100
rect 34940 2088 34946 2100
rect 35161 2091 35219 2097
rect 35161 2088 35173 2091
rect 34940 2060 35173 2088
rect 34940 2048 34946 2060
rect 35161 2057 35173 2060
rect 35207 2057 35219 2091
rect 35161 2051 35219 2057
rect 35268 2060 35388 2088
rect 33597 2023 33655 2029
rect 33597 2020 33609 2023
rect 33192 1992 33609 2020
rect 33192 1980 33198 1992
rect 33597 1989 33609 1992
rect 33643 1989 33655 2023
rect 33597 1983 33655 1989
rect 34149 2023 34207 2029
rect 34149 1989 34161 2023
rect 34195 1989 34207 2023
rect 34149 1983 34207 1989
rect 34238 1980 34244 2032
rect 34296 2020 34302 2032
rect 35268 2020 35296 2060
rect 34296 1992 35296 2020
rect 35360 2020 35388 2060
rect 35526 2048 35532 2100
rect 35584 2088 35590 2100
rect 35584 2060 37228 2088
rect 35584 2048 35590 2060
rect 35360 1992 35664 2020
rect 34296 1980 34302 1992
rect 29089 1955 29147 1961
rect 29089 1921 29101 1955
rect 29135 1921 29147 1955
rect 29089 1915 29147 1921
rect 29365 1955 29423 1961
rect 29365 1921 29377 1955
rect 29411 1921 29423 1955
rect 29365 1915 29423 1921
rect 28736 1856 28948 1884
rect 29104 1884 29132 1915
rect 29638 1912 29644 1964
rect 29696 1912 29702 1964
rect 30006 1912 30012 1964
rect 30064 1952 30070 1964
rect 30101 1955 30159 1961
rect 30101 1952 30113 1955
rect 30064 1924 30113 1952
rect 30064 1912 30070 1924
rect 30101 1921 30113 1924
rect 30147 1921 30159 1955
rect 30101 1915 30159 1921
rect 30190 1912 30196 1964
rect 30248 1912 30254 1964
rect 30466 1912 30472 1964
rect 30524 1912 30530 1964
rect 31573 1955 31631 1961
rect 31573 1921 31585 1955
rect 31619 1921 31631 1955
rect 31573 1915 31631 1921
rect 29104 1856 29684 1884
rect 29656 1828 29684 1856
rect 31294 1844 31300 1896
rect 31352 1844 31358 1896
rect 26605 1819 26663 1825
rect 25372 1788 26004 1816
rect 25372 1776 25378 1788
rect 17954 1748 17960 1760
rect 17788 1720 17960 1748
rect 17589 1711 17647 1717
rect 17954 1708 17960 1720
rect 18012 1708 18018 1760
rect 18141 1751 18199 1757
rect 18141 1717 18153 1751
rect 18187 1748 18199 1751
rect 18598 1748 18604 1760
rect 18187 1720 18604 1748
rect 18187 1717 18199 1720
rect 18141 1711 18199 1717
rect 18598 1708 18604 1720
rect 18656 1708 18662 1760
rect 18693 1751 18751 1757
rect 18693 1717 18705 1751
rect 18739 1748 18751 1751
rect 19978 1748 19984 1760
rect 18739 1720 19984 1748
rect 18739 1717 18751 1720
rect 18693 1711 18751 1717
rect 19978 1708 19984 1720
rect 20036 1708 20042 1760
rect 20073 1751 20131 1757
rect 20073 1717 20085 1751
rect 20119 1748 20131 1751
rect 20254 1748 20260 1760
rect 20119 1720 20260 1748
rect 20119 1717 20131 1720
rect 20073 1711 20131 1717
rect 20254 1708 20260 1720
rect 20312 1708 20318 1760
rect 20346 1708 20352 1760
rect 20404 1708 20410 1760
rect 20622 1708 20628 1760
rect 20680 1708 20686 1760
rect 20901 1751 20959 1757
rect 20901 1717 20913 1751
rect 20947 1748 20959 1751
rect 21082 1748 21088 1760
rect 20947 1720 21088 1748
rect 20947 1717 20959 1720
rect 20901 1711 20959 1717
rect 21082 1708 21088 1720
rect 21140 1708 21146 1760
rect 21174 1708 21180 1760
rect 21232 1708 21238 1760
rect 22370 1708 22376 1760
rect 22428 1708 22434 1760
rect 22554 1708 22560 1760
rect 22612 1748 22618 1760
rect 22649 1751 22707 1757
rect 22649 1748 22661 1751
rect 22612 1720 22661 1748
rect 22612 1708 22618 1720
rect 22649 1717 22661 1720
rect 22695 1717 22707 1751
rect 22649 1711 22707 1717
rect 23290 1708 23296 1760
rect 23348 1708 23354 1760
rect 23566 1708 23572 1760
rect 23624 1708 23630 1760
rect 23842 1708 23848 1760
rect 23900 1748 23906 1760
rect 24121 1751 24179 1757
rect 24121 1748 24133 1751
rect 23900 1720 24133 1748
rect 23900 1708 23906 1720
rect 24121 1717 24133 1720
rect 24167 1717 24179 1751
rect 24121 1711 24179 1717
rect 25501 1751 25559 1757
rect 25501 1717 25513 1751
rect 25547 1748 25559 1751
rect 25866 1748 25872 1760
rect 25547 1720 25872 1748
rect 25547 1717 25559 1720
rect 25501 1711 25559 1717
rect 25866 1708 25872 1720
rect 25924 1708 25930 1760
rect 25976 1757 26004 1788
rect 26605 1785 26617 1819
rect 26651 1785 26663 1819
rect 26605 1779 26663 1785
rect 26878 1776 26884 1828
rect 26936 1816 26942 1828
rect 27614 1816 27620 1828
rect 26936 1788 27620 1816
rect 26936 1776 26942 1788
rect 27614 1776 27620 1788
rect 27672 1776 27678 1828
rect 27890 1776 27896 1828
rect 27948 1816 27954 1828
rect 28997 1819 29055 1825
rect 27948 1788 28672 1816
rect 27948 1776 27954 1788
rect 25961 1751 26019 1757
rect 25961 1717 25973 1751
rect 26007 1717 26019 1751
rect 25961 1711 26019 1717
rect 26326 1708 26332 1760
rect 26384 1708 26390 1760
rect 26418 1708 26424 1760
rect 26476 1748 26482 1760
rect 27157 1751 27215 1757
rect 27157 1748 27169 1751
rect 26476 1720 27169 1748
rect 26476 1708 26482 1720
rect 27157 1717 27169 1720
rect 27203 1717 27215 1751
rect 27157 1711 27215 1717
rect 27246 1708 27252 1760
rect 27304 1748 27310 1760
rect 28644 1757 28672 1788
rect 28997 1785 29009 1819
rect 29043 1816 29055 1819
rect 29362 1816 29368 1828
rect 29043 1788 29368 1816
rect 29043 1785 29055 1788
rect 28997 1779 29055 1785
rect 29362 1776 29368 1788
rect 29420 1776 29426 1828
rect 29638 1776 29644 1828
rect 29696 1776 29702 1828
rect 29825 1819 29883 1825
rect 29825 1785 29837 1819
rect 29871 1816 29883 1819
rect 30466 1816 30472 1828
rect 29871 1788 30472 1816
rect 29871 1785 29883 1788
rect 29825 1779 29883 1785
rect 30466 1776 30472 1788
rect 30524 1776 30530 1828
rect 30653 1819 30711 1825
rect 30653 1785 30665 1819
rect 30699 1816 30711 1819
rect 31588 1816 31616 1915
rect 32122 1912 32128 1964
rect 32180 1912 32186 1964
rect 32582 1912 32588 1964
rect 32640 1912 32646 1964
rect 35342 1912 35348 1964
rect 35400 1912 35406 1964
rect 35529 1955 35587 1961
rect 35529 1921 35541 1955
rect 35575 1921 35587 1955
rect 35636 1952 35664 1992
rect 35710 1980 35716 2032
rect 35768 2020 35774 2032
rect 36173 2023 36231 2029
rect 36173 2020 36185 2023
rect 35768 1992 36185 2020
rect 35768 1980 35774 1992
rect 36173 1989 36185 1992
rect 36219 1989 36231 2023
rect 36173 1983 36231 1989
rect 36725 1955 36783 1961
rect 36725 1952 36737 1955
rect 35636 1924 36737 1952
rect 35529 1915 35587 1921
rect 36725 1921 36737 1924
rect 36771 1921 36783 1955
rect 36725 1915 36783 1921
rect 31846 1844 31852 1896
rect 31904 1844 31910 1896
rect 35544 1884 35572 1915
rect 37090 1884 37096 1896
rect 32508 1856 35572 1884
rect 35636 1856 37096 1884
rect 30699 1788 31616 1816
rect 30699 1785 30711 1788
rect 30653 1779 30711 1785
rect 32306 1776 32312 1828
rect 32364 1776 32370 1828
rect 32398 1776 32404 1828
rect 32456 1776 32462 1828
rect 28077 1751 28135 1757
rect 28077 1748 28089 1751
rect 27304 1720 28089 1748
rect 27304 1708 27310 1720
rect 28077 1717 28089 1720
rect 28123 1717 28135 1751
rect 28077 1711 28135 1717
rect 28629 1751 28687 1757
rect 28629 1717 28641 1751
rect 28675 1717 28687 1751
rect 28629 1711 28687 1717
rect 29270 1708 29276 1760
rect 29328 1708 29334 1760
rect 29546 1708 29552 1760
rect 29604 1708 29610 1760
rect 30282 1708 30288 1760
rect 30340 1748 30346 1760
rect 32508 1748 32536 1856
rect 32582 1776 32588 1828
rect 32640 1816 32646 1828
rect 33137 1819 33195 1825
rect 33137 1816 33149 1819
rect 32640 1788 33149 1816
rect 32640 1776 32646 1788
rect 33137 1785 33149 1788
rect 33183 1785 33195 1819
rect 33137 1779 33195 1785
rect 33244 1788 34284 1816
rect 30340 1720 32536 1748
rect 30340 1708 30346 1720
rect 33042 1708 33048 1760
rect 33100 1748 33106 1760
rect 33244 1748 33272 1788
rect 33100 1720 33272 1748
rect 33100 1708 33106 1720
rect 33410 1708 33416 1760
rect 33468 1748 33474 1760
rect 34256 1757 34284 1788
rect 34330 1776 34336 1828
rect 34388 1816 34394 1828
rect 35636 1816 35664 1856
rect 37090 1844 37096 1856
rect 37148 1844 37154 1896
rect 34388 1788 35664 1816
rect 34388 1776 34394 1788
rect 35710 1776 35716 1828
rect 35768 1816 35774 1828
rect 37200 1816 37228 2060
rect 37274 2048 37280 2100
rect 37332 2048 37338 2100
rect 37366 2048 37372 2100
rect 37424 2088 37430 2100
rect 37645 2091 37703 2097
rect 37645 2088 37657 2091
rect 37424 2060 37657 2088
rect 37424 2048 37430 2060
rect 37645 2057 37657 2060
rect 37691 2057 37703 2091
rect 37645 2051 37703 2057
rect 38562 2048 38568 2100
rect 38620 2088 38626 2100
rect 39393 2091 39451 2097
rect 39393 2088 39405 2091
rect 38620 2060 39405 2088
rect 38620 2048 38626 2060
rect 39393 2057 39405 2060
rect 39439 2057 39451 2091
rect 39393 2051 39451 2057
rect 39666 2048 39672 2100
rect 39724 2088 39730 2100
rect 39761 2091 39819 2097
rect 39761 2088 39773 2091
rect 39724 2060 39773 2088
rect 39724 2048 39730 2060
rect 39761 2057 39773 2060
rect 39807 2057 39819 2091
rect 40957 2091 41015 2097
rect 40957 2088 40969 2091
rect 39761 2051 39819 2057
rect 39868 2060 40969 2088
rect 37292 1884 37320 2048
rect 38654 1980 38660 2032
rect 38712 2020 38718 2032
rect 39301 2023 39359 2029
rect 39301 2020 39313 2023
rect 38712 1992 39313 2020
rect 38712 1980 38718 1992
rect 39301 1989 39313 1992
rect 39347 1989 39359 2023
rect 39301 1983 39359 1989
rect 37826 1912 37832 1964
rect 37884 1912 37890 1964
rect 38102 1912 38108 1964
rect 38160 1912 38166 1964
rect 38746 1912 38752 1964
rect 38804 1912 38810 1964
rect 39868 1884 39896 2060
rect 40957 2057 40969 2060
rect 41003 2057 41015 2091
rect 40957 2051 41015 2057
rect 41782 2048 41788 2100
rect 41840 2088 41846 2100
rect 42429 2091 42487 2097
rect 42429 2088 42441 2091
rect 41840 2060 42441 2088
rect 41840 2048 41846 2060
rect 42429 2057 42441 2060
rect 42475 2057 42487 2091
rect 42429 2051 42487 2057
rect 44174 2048 44180 2100
rect 44232 2088 44238 2100
rect 44637 2091 44695 2097
rect 44637 2088 44649 2091
rect 44232 2060 44649 2088
rect 44232 2048 44238 2060
rect 44637 2057 44649 2060
rect 44683 2057 44695 2091
rect 44637 2051 44695 2057
rect 44910 2048 44916 2100
rect 44968 2048 44974 2100
rect 45002 2048 45008 2100
rect 45060 2048 45066 2100
rect 45278 2048 45284 2100
rect 45336 2048 45342 2100
rect 45020 2020 45048 2048
rect 39960 1992 42564 2020
rect 39960 1961 39988 1992
rect 39945 1955 40003 1961
rect 39945 1921 39957 1955
rect 39991 1921 40003 1955
rect 39945 1915 40003 1921
rect 40586 1912 40592 1964
rect 40644 1912 40650 1964
rect 40678 1912 40684 1964
rect 40736 1952 40742 1964
rect 40865 1955 40923 1961
rect 40865 1952 40877 1955
rect 40736 1924 40877 1952
rect 40736 1912 40742 1924
rect 40865 1921 40877 1924
rect 40911 1921 40923 1955
rect 40865 1915 40923 1921
rect 41141 1955 41199 1961
rect 41141 1921 41153 1955
rect 41187 1921 41199 1955
rect 41141 1915 41199 1921
rect 37292 1856 39896 1884
rect 40770 1844 40776 1896
rect 40828 1884 40834 1896
rect 41156 1884 41184 1915
rect 41598 1912 41604 1964
rect 41656 1912 41662 1964
rect 40828 1856 41184 1884
rect 41325 1887 41383 1893
rect 40828 1844 40834 1856
rect 41325 1853 41337 1887
rect 41371 1853 41383 1887
rect 42536 1884 42564 1992
rect 42628 1992 45048 2020
rect 42628 1961 42656 1992
rect 42613 1955 42671 1961
rect 42613 1921 42625 1955
rect 42659 1921 42671 1955
rect 42613 1915 42671 1921
rect 44821 1955 44879 1961
rect 44821 1921 44833 1955
rect 44867 1921 44879 1955
rect 44821 1915 44879 1921
rect 45097 1955 45155 1961
rect 45097 1921 45109 1955
rect 45143 1952 45155 1955
rect 45296 1952 45324 2048
rect 45143 1924 45324 1952
rect 45143 1921 45155 1924
rect 45097 1915 45155 1921
rect 44174 1884 44180 1896
rect 42536 1856 44180 1884
rect 41325 1847 41383 1853
rect 40681 1819 40739 1825
rect 40681 1816 40693 1819
rect 35768 1788 36860 1816
rect 37200 1788 40693 1816
rect 35768 1776 35774 1788
rect 33689 1751 33747 1757
rect 33689 1748 33701 1751
rect 33468 1720 33701 1748
rect 33468 1708 33474 1720
rect 33689 1717 33701 1720
rect 33735 1717 33747 1751
rect 33689 1711 33747 1717
rect 34241 1751 34299 1757
rect 34241 1717 34253 1751
rect 34287 1717 34299 1751
rect 34241 1711 34299 1717
rect 34882 1708 34888 1760
rect 34940 1748 34946 1760
rect 35621 1751 35679 1757
rect 35621 1748 35633 1751
rect 34940 1720 35633 1748
rect 34940 1708 34946 1720
rect 35621 1717 35633 1720
rect 35667 1717 35679 1751
rect 35621 1711 35679 1717
rect 36262 1708 36268 1760
rect 36320 1708 36326 1760
rect 36832 1757 36860 1788
rect 40681 1785 40693 1788
rect 40727 1785 40739 1819
rect 41340 1816 41368 1847
rect 44174 1844 44180 1856
rect 44232 1844 44238 1896
rect 44836 1884 44864 1915
rect 45462 1912 45468 1964
rect 45520 1912 45526 1964
rect 44836 1856 45324 1884
rect 41874 1816 41880 1828
rect 41340 1788 41880 1816
rect 40681 1779 40739 1785
rect 41874 1776 41880 1788
rect 41932 1776 41938 1828
rect 45296 1825 45324 1856
rect 45281 1819 45339 1825
rect 45281 1785 45293 1819
rect 45327 1785 45339 1819
rect 45281 1779 45339 1785
rect 36817 1751 36875 1757
rect 36817 1717 36829 1751
rect 36863 1717 36875 1751
rect 36817 1711 36875 1717
rect 37274 1708 37280 1760
rect 37332 1748 37338 1760
rect 38197 1751 38255 1757
rect 38197 1748 38209 1751
rect 37332 1720 38209 1748
rect 37332 1708 37338 1720
rect 38197 1717 38209 1720
rect 38243 1717 38255 1751
rect 38197 1711 38255 1717
rect 38470 1708 38476 1760
rect 38528 1748 38534 1760
rect 38841 1751 38899 1757
rect 38841 1748 38853 1751
rect 38528 1720 38853 1748
rect 38528 1708 38534 1720
rect 38841 1717 38853 1720
rect 38887 1717 38899 1751
rect 38841 1711 38899 1717
rect 38930 1708 38936 1760
rect 38988 1748 38994 1760
rect 40405 1751 40463 1757
rect 40405 1748 40417 1751
rect 38988 1720 40417 1748
rect 38988 1708 38994 1720
rect 40405 1717 40417 1720
rect 40451 1717 40463 1751
rect 40405 1711 40463 1717
rect 1104 1658 45816 1680
rect 1104 1606 6539 1658
rect 6591 1606 6603 1658
rect 6655 1606 6667 1658
rect 6719 1606 6731 1658
rect 6783 1606 6795 1658
rect 6847 1606 17717 1658
rect 17769 1606 17781 1658
rect 17833 1606 17845 1658
rect 17897 1606 17909 1658
rect 17961 1606 17973 1658
rect 18025 1606 28895 1658
rect 28947 1606 28959 1658
rect 29011 1606 29023 1658
rect 29075 1606 29087 1658
rect 29139 1606 29151 1658
rect 29203 1606 40073 1658
rect 40125 1606 40137 1658
rect 40189 1606 40201 1658
rect 40253 1606 40265 1658
rect 40317 1606 40329 1658
rect 40381 1606 45816 1658
rect 1104 1584 45816 1606
rect 1578 1504 1584 1556
rect 1636 1544 1642 1556
rect 6825 1547 6883 1553
rect 1636 1516 2774 1544
rect 1636 1504 1642 1516
rect 2746 1476 2774 1516
rect 6825 1513 6837 1547
rect 6871 1544 6883 1547
rect 9674 1544 9680 1556
rect 6871 1516 9680 1544
rect 6871 1513 6883 1516
rect 6825 1507 6883 1513
rect 9674 1504 9680 1516
rect 9732 1504 9738 1556
rect 14274 1504 14280 1556
rect 14332 1504 14338 1556
rect 15102 1504 15108 1556
rect 15160 1504 15166 1556
rect 15381 1547 15439 1553
rect 15381 1513 15393 1547
rect 15427 1544 15439 1547
rect 15470 1544 15476 1556
rect 15427 1516 15476 1544
rect 15427 1513 15439 1516
rect 15381 1507 15439 1513
rect 15470 1504 15476 1516
rect 15528 1504 15534 1556
rect 15657 1547 15715 1553
rect 15657 1513 15669 1547
rect 15703 1544 15715 1547
rect 15746 1544 15752 1556
rect 15703 1516 15752 1544
rect 15703 1513 15715 1516
rect 15657 1507 15715 1513
rect 15746 1504 15752 1516
rect 15804 1504 15810 1556
rect 15933 1547 15991 1553
rect 15933 1513 15945 1547
rect 15979 1544 15991 1547
rect 16022 1544 16028 1556
rect 15979 1516 16028 1544
rect 15979 1513 15991 1516
rect 15933 1507 15991 1513
rect 16022 1504 16028 1516
rect 16080 1504 16086 1556
rect 16209 1547 16267 1553
rect 16209 1513 16221 1547
rect 16255 1544 16267 1547
rect 16298 1544 16304 1556
rect 16255 1516 16304 1544
rect 16255 1513 16267 1516
rect 16209 1507 16267 1513
rect 16298 1504 16304 1516
rect 16356 1504 16362 1556
rect 16482 1504 16488 1556
rect 16540 1504 16546 1556
rect 16945 1547 17003 1553
rect 16945 1513 16957 1547
rect 16991 1544 17003 1547
rect 17126 1544 17132 1556
rect 16991 1516 17132 1544
rect 16991 1513 17003 1516
rect 16945 1507 17003 1513
rect 17126 1504 17132 1516
rect 17184 1504 17190 1556
rect 17402 1504 17408 1556
rect 17460 1544 17466 1556
rect 17497 1547 17555 1553
rect 17497 1544 17509 1547
rect 17460 1516 17509 1544
rect 17460 1504 17466 1516
rect 17497 1513 17509 1516
rect 17543 1513 17555 1547
rect 17497 1507 17555 1513
rect 17957 1547 18015 1553
rect 17957 1513 17969 1547
rect 18003 1544 18015 1547
rect 18046 1544 18052 1556
rect 18003 1516 18052 1544
rect 18003 1513 18015 1516
rect 17957 1507 18015 1513
rect 18046 1504 18052 1516
rect 18104 1504 18110 1556
rect 18138 1504 18144 1556
rect 18196 1544 18202 1556
rect 18325 1547 18383 1553
rect 18325 1544 18337 1547
rect 18196 1516 18337 1544
rect 18196 1504 18202 1516
rect 18325 1513 18337 1516
rect 18371 1513 18383 1547
rect 18325 1507 18383 1513
rect 18506 1504 18512 1556
rect 18564 1544 18570 1556
rect 18601 1547 18659 1553
rect 18601 1544 18613 1547
rect 18564 1516 18613 1544
rect 18564 1504 18570 1516
rect 18601 1513 18613 1516
rect 18647 1513 18659 1547
rect 18601 1507 18659 1513
rect 19058 1504 19064 1556
rect 19116 1544 19122 1556
rect 19245 1547 19303 1553
rect 19245 1544 19257 1547
rect 19116 1516 19257 1544
rect 19116 1504 19122 1516
rect 19245 1513 19257 1516
rect 19291 1513 19303 1547
rect 19245 1507 19303 1513
rect 19610 1504 19616 1556
rect 19668 1544 19674 1556
rect 19668 1516 21036 1544
rect 19668 1504 19674 1516
rect 17586 1476 17592 1488
rect 2746 1448 17592 1476
rect 17586 1436 17592 1448
rect 17644 1436 17650 1488
rect 18230 1436 18236 1488
rect 18288 1476 18294 1488
rect 18288 1448 19288 1476
rect 18288 1436 18294 1448
rect 18322 1408 18328 1420
rect 5460 1380 7144 1408
rect 1486 1300 1492 1352
rect 1544 1300 1550 1352
rect 1854 1300 1860 1352
rect 1912 1300 1918 1352
rect 2222 1300 2228 1352
rect 2280 1300 2286 1352
rect 2501 1343 2559 1349
rect 2501 1309 2513 1343
rect 2547 1340 2559 1343
rect 3234 1340 3240 1352
rect 2547 1312 3240 1340
rect 2547 1309 2559 1312
rect 2501 1303 2559 1309
rect 3234 1300 3240 1312
rect 3292 1300 3298 1352
rect 3326 1300 3332 1352
rect 3384 1300 3390 1352
rect 3786 1300 3792 1352
rect 3844 1300 3850 1352
rect 4062 1300 4068 1352
rect 4120 1300 4126 1352
rect 4430 1300 4436 1352
rect 4488 1300 4494 1352
rect 4798 1300 4804 1352
rect 4856 1300 4862 1352
rect 5166 1300 5172 1352
rect 5224 1300 5230 1352
rect 5460 1272 5488 1380
rect 5534 1300 5540 1352
rect 5592 1300 5598 1352
rect 5626 1300 5632 1352
rect 5684 1300 5690 1352
rect 5902 1300 5908 1352
rect 5960 1300 5966 1352
rect 6362 1300 6368 1352
rect 6420 1300 6426 1352
rect 6638 1300 6644 1352
rect 6696 1300 6702 1352
rect 6914 1300 6920 1352
rect 6972 1300 6978 1352
rect 7006 1300 7012 1352
rect 7064 1300 7070 1352
rect 4264 1244 5488 1272
rect 1673 1207 1731 1213
rect 1673 1173 1685 1207
rect 1719 1204 1731 1207
rect 1946 1204 1952 1216
rect 1719 1176 1952 1204
rect 1719 1173 1731 1176
rect 1673 1167 1731 1173
rect 1946 1164 1952 1176
rect 2004 1164 2010 1216
rect 2038 1164 2044 1216
rect 2096 1164 2102 1216
rect 3510 1164 3516 1216
rect 3568 1164 3574 1216
rect 3973 1207 4031 1213
rect 3973 1173 3985 1207
rect 4019 1204 4031 1207
rect 4154 1204 4160 1216
rect 4019 1176 4160 1204
rect 4019 1173 4031 1176
rect 3973 1167 4031 1173
rect 4154 1164 4160 1176
rect 4212 1164 4218 1216
rect 4264 1213 4292 1244
rect 4249 1207 4307 1213
rect 4249 1173 4261 1207
rect 4295 1173 4307 1207
rect 4249 1167 4307 1173
rect 4614 1164 4620 1216
rect 4672 1164 4678 1216
rect 4982 1164 4988 1216
rect 5040 1164 5046 1216
rect 5353 1207 5411 1213
rect 5353 1173 5365 1207
rect 5399 1204 5411 1207
rect 5644 1204 5672 1300
rect 6932 1272 6960 1300
rect 5736 1244 6960 1272
rect 7116 1272 7144 1380
rect 12452 1380 12664 1408
rect 7374 1300 7380 1352
rect 7432 1300 7438 1352
rect 7742 1300 7748 1352
rect 7800 1300 7806 1352
rect 8110 1300 8116 1352
rect 8168 1300 8174 1352
rect 8478 1340 8484 1352
rect 8220 1312 8484 1340
rect 8220 1272 8248 1312
rect 8478 1300 8484 1312
rect 8536 1300 8542 1352
rect 8570 1300 8576 1352
rect 8628 1300 8634 1352
rect 8941 1343 8999 1349
rect 8941 1309 8953 1343
rect 8987 1309 8999 1343
rect 8941 1303 8999 1309
rect 9217 1343 9275 1349
rect 9217 1309 9229 1343
rect 9263 1340 9275 1343
rect 9490 1340 9496 1352
rect 9263 1312 9496 1340
rect 9263 1309 9275 1312
rect 9217 1303 9275 1309
rect 7116 1244 8248 1272
rect 5736 1213 5764 1244
rect 8386 1232 8392 1284
rect 8444 1272 8450 1284
rect 8956 1272 8984 1303
rect 9490 1300 9496 1312
rect 9548 1300 9554 1352
rect 9950 1300 9956 1352
rect 10008 1300 10014 1352
rect 10318 1300 10324 1352
rect 10376 1300 10382 1352
rect 10686 1300 10692 1352
rect 10744 1300 10750 1352
rect 11054 1300 11060 1352
rect 11112 1300 11118 1352
rect 11514 1300 11520 1352
rect 11572 1300 11578 1352
rect 11790 1300 11796 1352
rect 11848 1300 11854 1352
rect 12158 1300 12164 1352
rect 12216 1300 12222 1352
rect 12452 1340 12480 1380
rect 12268 1312 12480 1340
rect 11422 1272 11428 1284
rect 8444 1244 8984 1272
rect 10520 1244 11428 1272
rect 8444 1232 8450 1244
rect 5399 1176 5672 1204
rect 5721 1207 5779 1213
rect 5399 1173 5411 1176
rect 5353 1167 5411 1173
rect 5721 1173 5733 1207
rect 5767 1173 5779 1207
rect 5721 1167 5779 1173
rect 6086 1164 6092 1216
rect 6144 1164 6150 1216
rect 6546 1164 6552 1216
rect 6604 1164 6610 1216
rect 7190 1164 7196 1216
rect 7248 1164 7254 1216
rect 7558 1164 7564 1216
rect 7616 1164 7622 1216
rect 7926 1164 7932 1216
rect 7984 1164 7990 1216
rect 8294 1164 8300 1216
rect 8352 1164 8358 1216
rect 8754 1164 8760 1216
rect 8812 1164 8818 1216
rect 10134 1164 10140 1216
rect 10192 1164 10198 1216
rect 10520 1213 10548 1244
rect 11422 1232 11428 1244
rect 11480 1232 11486 1284
rect 10505 1207 10563 1213
rect 10505 1173 10517 1207
rect 10551 1173 10563 1207
rect 10505 1167 10563 1173
rect 10870 1164 10876 1216
rect 10928 1164 10934 1216
rect 11238 1164 11244 1216
rect 11296 1164 11302 1216
rect 11701 1207 11759 1213
rect 11701 1173 11713 1207
rect 11747 1204 11759 1207
rect 11882 1204 11888 1216
rect 11747 1176 11888 1204
rect 11747 1173 11759 1176
rect 11701 1167 11759 1173
rect 11882 1164 11888 1176
rect 11940 1164 11946 1216
rect 11977 1207 12035 1213
rect 11977 1173 11989 1207
rect 12023 1204 12035 1207
rect 12268 1204 12296 1312
rect 12526 1300 12532 1352
rect 12584 1300 12590 1352
rect 12636 1340 12664 1380
rect 14568 1380 18328 1408
rect 12802 1340 12808 1352
rect 12636 1312 12808 1340
rect 12802 1300 12808 1312
rect 12860 1300 12866 1352
rect 12894 1300 12900 1352
rect 12952 1300 12958 1352
rect 13262 1300 13268 1352
rect 13320 1300 13326 1352
rect 13630 1300 13636 1352
rect 13688 1300 13694 1352
rect 14090 1300 14096 1352
rect 14148 1300 14154 1352
rect 14366 1300 14372 1352
rect 14424 1300 14430 1352
rect 12360 1244 14504 1272
rect 12360 1213 12388 1244
rect 14476 1216 14504 1244
rect 12023 1176 12296 1204
rect 12345 1207 12403 1213
rect 12023 1173 12035 1176
rect 11977 1167 12035 1173
rect 12345 1173 12357 1207
rect 12391 1173 12403 1207
rect 12345 1167 12403 1173
rect 12710 1164 12716 1216
rect 12768 1164 12774 1216
rect 13081 1207 13139 1213
rect 13081 1173 13093 1207
rect 13127 1204 13139 1207
rect 13354 1204 13360 1216
rect 13127 1176 13360 1204
rect 13127 1173 13139 1176
rect 13081 1167 13139 1173
rect 13354 1164 13360 1176
rect 13412 1164 13418 1216
rect 13446 1164 13452 1216
rect 13504 1164 13510 1216
rect 13814 1164 13820 1216
rect 13872 1164 13878 1216
rect 14458 1164 14464 1216
rect 14516 1164 14522 1216
rect 14568 1213 14596 1380
rect 18322 1368 18328 1380
rect 18380 1368 18386 1420
rect 18708 1380 18920 1408
rect 14642 1300 14648 1352
rect 14700 1300 14706 1352
rect 14918 1300 14924 1352
rect 14976 1300 14982 1352
rect 15194 1300 15200 1352
rect 15252 1300 15258 1352
rect 15470 1300 15476 1352
rect 15528 1300 15534 1352
rect 15749 1343 15807 1349
rect 15749 1309 15761 1343
rect 15795 1309 15807 1343
rect 15749 1303 15807 1309
rect 16025 1343 16083 1349
rect 16025 1309 16037 1343
rect 16071 1340 16083 1343
rect 16206 1340 16212 1352
rect 16071 1312 16212 1340
rect 16071 1309 16083 1312
rect 16025 1303 16083 1309
rect 15764 1272 15792 1303
rect 16206 1300 16212 1312
rect 16264 1300 16270 1352
rect 16301 1343 16359 1349
rect 16301 1309 16313 1343
rect 16347 1340 16359 1343
rect 16574 1340 16580 1352
rect 16347 1312 16580 1340
rect 16347 1309 16359 1312
rect 16301 1303 16359 1309
rect 16574 1300 16580 1312
rect 16632 1300 16638 1352
rect 16758 1300 16764 1352
rect 16816 1300 16822 1352
rect 17037 1343 17095 1349
rect 17037 1309 17049 1343
rect 17083 1309 17095 1343
rect 17037 1303 17095 1309
rect 16114 1272 16120 1284
rect 15764 1244 16120 1272
rect 16114 1232 16120 1244
rect 16172 1232 16178 1284
rect 16482 1232 16488 1284
rect 16540 1272 16546 1284
rect 17052 1272 17080 1303
rect 17678 1300 17684 1352
rect 17736 1300 17742 1352
rect 17770 1300 17776 1352
rect 17828 1300 17834 1352
rect 18046 1300 18052 1352
rect 18104 1300 18110 1352
rect 18506 1300 18512 1352
rect 18564 1300 18570 1352
rect 18708 1340 18736 1380
rect 18616 1312 18736 1340
rect 18616 1272 18644 1312
rect 18782 1300 18788 1352
rect 18840 1300 18846 1352
rect 18892 1349 18920 1380
rect 18877 1343 18935 1349
rect 18877 1309 18889 1343
rect 18923 1309 18935 1343
rect 18877 1303 18935 1309
rect 19150 1300 19156 1352
rect 19208 1300 19214 1352
rect 16540 1244 17080 1272
rect 17144 1244 18644 1272
rect 16540 1232 16546 1244
rect 14553 1207 14611 1213
rect 14553 1173 14565 1207
rect 14599 1173 14611 1207
rect 14553 1167 14611 1173
rect 14829 1207 14887 1213
rect 14829 1173 14841 1207
rect 14875 1204 14887 1207
rect 17144 1204 17172 1244
rect 18690 1232 18696 1284
rect 18748 1232 18754 1284
rect 14875 1176 17172 1204
rect 14875 1173 14887 1176
rect 14829 1167 14887 1173
rect 17218 1164 17224 1216
rect 17276 1164 17282 1216
rect 18233 1207 18291 1213
rect 18233 1173 18245 1207
rect 18279 1204 18291 1207
rect 18708 1204 18736 1232
rect 18279 1176 18736 1204
rect 19061 1207 19119 1213
rect 18279 1173 18291 1176
rect 18233 1167 18291 1173
rect 19061 1173 19073 1207
rect 19107 1204 19119 1207
rect 19168 1204 19196 1300
rect 19260 1272 19288 1448
rect 19978 1436 19984 1488
rect 20036 1436 20042 1488
rect 20898 1436 20904 1488
rect 20956 1436 20962 1488
rect 21008 1476 21036 1516
rect 21910 1504 21916 1556
rect 21968 1544 21974 1556
rect 22281 1547 22339 1553
rect 22281 1544 22293 1547
rect 21968 1516 22293 1544
rect 21968 1504 21974 1516
rect 22281 1513 22293 1516
rect 22327 1513 22339 1547
rect 22281 1507 22339 1513
rect 22370 1504 22376 1556
rect 22428 1544 22434 1556
rect 23934 1544 23940 1556
rect 22428 1516 23940 1544
rect 22428 1504 22434 1516
rect 23934 1504 23940 1516
rect 23992 1504 23998 1556
rect 24412 1516 25544 1544
rect 24412 1476 24440 1516
rect 21008 1448 24440 1476
rect 25516 1476 25544 1516
rect 26234 1504 26240 1556
rect 26292 1544 26298 1556
rect 26329 1547 26387 1553
rect 26329 1544 26341 1547
rect 26292 1516 26341 1544
rect 26292 1504 26298 1516
rect 26329 1513 26341 1516
rect 26375 1513 26387 1547
rect 26329 1507 26387 1513
rect 26602 1504 26608 1556
rect 26660 1544 26666 1556
rect 27157 1547 27215 1553
rect 27157 1544 27169 1547
rect 26660 1516 27169 1544
rect 26660 1504 26666 1516
rect 27157 1513 27169 1516
rect 27203 1513 27215 1547
rect 27157 1507 27215 1513
rect 27614 1504 27620 1556
rect 27672 1544 27678 1556
rect 27893 1547 27951 1553
rect 27893 1544 27905 1547
rect 27672 1516 27905 1544
rect 27672 1504 27678 1516
rect 27893 1513 27905 1516
rect 27939 1513 27951 1547
rect 27893 1507 27951 1513
rect 28445 1547 28503 1553
rect 28445 1513 28457 1547
rect 28491 1513 28503 1547
rect 28445 1507 28503 1513
rect 25516 1448 27292 1476
rect 19996 1408 20024 1436
rect 23474 1408 23480 1420
rect 19352 1380 19932 1408
rect 19996 1380 23480 1408
rect 19352 1352 19380 1380
rect 19334 1300 19340 1352
rect 19392 1300 19398 1352
rect 19426 1300 19432 1352
rect 19484 1300 19490 1352
rect 19904 1349 19932 1380
rect 23474 1368 23480 1380
rect 23532 1368 23538 1420
rect 23566 1368 23572 1420
rect 23624 1408 23630 1420
rect 23624 1380 25636 1408
rect 23624 1368 23630 1380
rect 19521 1343 19579 1349
rect 19521 1309 19533 1343
rect 19567 1309 19579 1343
rect 19521 1303 19579 1309
rect 19889 1343 19947 1349
rect 19889 1309 19901 1343
rect 19935 1309 19947 1343
rect 19889 1303 19947 1309
rect 19536 1272 19564 1303
rect 19978 1300 19984 1352
rect 20036 1340 20042 1352
rect 20257 1343 20315 1349
rect 20257 1340 20269 1343
rect 20036 1312 20269 1340
rect 20036 1300 20042 1312
rect 20257 1309 20269 1312
rect 20303 1309 20315 1343
rect 20257 1303 20315 1309
rect 20346 1300 20352 1352
rect 20404 1340 20410 1352
rect 21361 1343 21419 1349
rect 21361 1340 21373 1343
rect 20404 1312 21373 1340
rect 20404 1300 20410 1312
rect 21361 1309 21373 1312
rect 21407 1309 21419 1343
rect 21361 1303 21419 1309
rect 21818 1300 21824 1352
rect 21876 1300 21882 1352
rect 22094 1300 22100 1352
rect 22152 1340 22158 1352
rect 22833 1343 22891 1349
rect 22833 1340 22845 1343
rect 22152 1312 22845 1340
rect 22152 1300 22158 1312
rect 22833 1309 22845 1312
rect 22879 1309 22891 1343
rect 22833 1303 22891 1309
rect 23198 1300 23204 1352
rect 23256 1300 23262 1352
rect 23290 1300 23296 1352
rect 23348 1340 23354 1352
rect 24765 1343 24823 1349
rect 24765 1340 24777 1343
rect 23348 1312 24777 1340
rect 23348 1300 23354 1312
rect 24765 1309 24777 1312
rect 24811 1309 24823 1343
rect 24765 1303 24823 1309
rect 24946 1300 24952 1352
rect 25004 1340 25010 1352
rect 25608 1340 25636 1380
rect 26142 1368 26148 1420
rect 26200 1408 26206 1420
rect 26602 1408 26608 1420
rect 26200 1380 26608 1408
rect 26200 1368 26206 1380
rect 26602 1368 26608 1380
rect 26660 1368 26666 1420
rect 27264 1408 27292 1448
rect 27706 1436 27712 1488
rect 27764 1476 27770 1488
rect 28460 1476 28488 1507
rect 28626 1504 28632 1556
rect 28684 1544 28690 1556
rect 29733 1547 29791 1553
rect 29733 1544 29745 1547
rect 28684 1516 29745 1544
rect 28684 1504 28690 1516
rect 29733 1513 29745 1516
rect 29779 1513 29791 1547
rect 29733 1507 29791 1513
rect 30285 1547 30343 1553
rect 30285 1513 30297 1547
rect 30331 1513 30343 1547
rect 30285 1507 30343 1513
rect 30837 1547 30895 1553
rect 30837 1513 30849 1547
rect 30883 1513 30895 1547
rect 30837 1507 30895 1513
rect 27764 1448 28488 1476
rect 27764 1436 27770 1448
rect 28994 1436 29000 1488
rect 29052 1476 29058 1488
rect 30300 1476 30328 1507
rect 29052 1448 30328 1476
rect 29052 1436 29058 1448
rect 28074 1408 28080 1420
rect 27264 1380 28080 1408
rect 28074 1368 28080 1380
rect 28132 1368 28138 1420
rect 28258 1368 28264 1420
rect 28316 1408 28322 1420
rect 28905 1411 28963 1417
rect 28905 1408 28917 1411
rect 28316 1380 28917 1408
rect 28316 1368 28322 1380
rect 28905 1377 28917 1380
rect 28951 1377 28963 1411
rect 28905 1371 28963 1377
rect 29454 1368 29460 1420
rect 29512 1408 29518 1420
rect 30852 1408 30880 1507
rect 31662 1504 31668 1556
rect 31720 1544 31726 1556
rect 32861 1547 32919 1553
rect 32861 1544 32873 1547
rect 31720 1516 32873 1544
rect 31720 1504 31726 1516
rect 32861 1513 32873 1516
rect 32907 1513 32919 1547
rect 32861 1507 32919 1513
rect 33413 1547 33471 1553
rect 33413 1513 33425 1547
rect 33459 1513 33471 1547
rect 33413 1507 33471 1513
rect 31018 1436 31024 1488
rect 31076 1476 31082 1488
rect 32401 1479 32459 1485
rect 32401 1476 32413 1479
rect 31076 1448 32413 1476
rect 31076 1436 31082 1448
rect 32401 1445 32413 1448
rect 32447 1445 32459 1479
rect 32401 1439 32459 1445
rect 29512 1380 30880 1408
rect 29512 1368 29518 1380
rect 31662 1368 31668 1420
rect 31720 1408 31726 1420
rect 33428 1408 33456 1507
rect 34330 1504 34336 1556
rect 34388 1544 34394 1556
rect 35437 1547 35495 1553
rect 35437 1544 35449 1547
rect 34388 1516 35449 1544
rect 34388 1504 34394 1516
rect 35437 1513 35449 1516
rect 35483 1513 35495 1547
rect 35437 1507 35495 1513
rect 36541 1547 36599 1553
rect 36541 1513 36553 1547
rect 36587 1513 36599 1547
rect 36541 1507 36599 1513
rect 34974 1436 34980 1488
rect 35032 1476 35038 1488
rect 36556 1476 36584 1507
rect 36906 1504 36912 1556
rect 36964 1544 36970 1556
rect 38013 1547 38071 1553
rect 38013 1544 38025 1547
rect 36964 1516 38025 1544
rect 36964 1504 36970 1516
rect 38013 1513 38025 1516
rect 38059 1513 38071 1547
rect 38013 1507 38071 1513
rect 38102 1504 38108 1556
rect 38160 1544 38166 1556
rect 39117 1547 39175 1553
rect 39117 1544 39129 1547
rect 38160 1516 39129 1544
rect 38160 1504 38166 1516
rect 39117 1513 39129 1516
rect 39163 1513 39175 1547
rect 39117 1507 39175 1513
rect 40037 1547 40095 1553
rect 40037 1513 40049 1547
rect 40083 1513 40095 1547
rect 40037 1507 40095 1513
rect 35032 1448 36584 1476
rect 35032 1436 35038 1448
rect 37090 1436 37096 1488
rect 37148 1476 37154 1488
rect 38657 1479 38715 1485
rect 38657 1476 38669 1479
rect 37148 1448 38669 1476
rect 37148 1436 37154 1448
rect 38657 1445 38669 1448
rect 38703 1445 38715 1479
rect 38657 1439 38715 1445
rect 39482 1436 39488 1488
rect 39540 1436 39546 1488
rect 35069 1411 35127 1417
rect 35069 1408 35081 1411
rect 31720 1380 33456 1408
rect 33520 1380 35081 1408
rect 31720 1368 31726 1380
rect 25777 1343 25835 1349
rect 25777 1340 25789 1343
rect 25004 1312 25544 1340
rect 25608 1312 25789 1340
rect 25004 1300 25010 1312
rect 19260 1244 19564 1272
rect 20714 1232 20720 1284
rect 20772 1232 20778 1284
rect 22186 1232 22192 1284
rect 22244 1232 22250 1284
rect 22462 1232 22468 1284
rect 22520 1232 22526 1284
rect 22738 1232 22744 1284
rect 22796 1272 22802 1284
rect 23661 1275 23719 1281
rect 23661 1272 23673 1275
rect 22796 1244 23673 1272
rect 22796 1232 22802 1244
rect 23661 1241 23673 1244
rect 23707 1241 23719 1275
rect 23661 1235 23719 1241
rect 23934 1232 23940 1284
rect 23992 1272 23998 1284
rect 25317 1275 25375 1281
rect 25317 1272 25329 1275
rect 23992 1244 25329 1272
rect 23992 1232 23998 1244
rect 25317 1241 25329 1244
rect 25363 1241 25375 1275
rect 25516 1272 25544 1312
rect 25777 1309 25789 1312
rect 25823 1309 25835 1343
rect 25777 1303 25835 1309
rect 25866 1300 25872 1352
rect 25924 1340 25930 1352
rect 26237 1343 26295 1349
rect 26237 1340 26249 1343
rect 25924 1312 26249 1340
rect 25924 1300 25930 1312
rect 26237 1309 26249 1312
rect 26283 1309 26295 1343
rect 26237 1303 26295 1309
rect 26326 1300 26332 1352
rect 26384 1340 26390 1352
rect 27065 1343 27123 1349
rect 27065 1340 27077 1343
rect 26384 1312 27077 1340
rect 26384 1300 26390 1312
rect 27065 1309 27077 1312
rect 27111 1309 27123 1343
rect 27065 1303 27123 1309
rect 27154 1300 27160 1352
rect 27212 1340 27218 1352
rect 27801 1343 27859 1349
rect 27801 1340 27813 1343
rect 27212 1312 27813 1340
rect 27212 1300 27218 1312
rect 27801 1309 27813 1312
rect 27847 1309 27859 1343
rect 27801 1303 27859 1309
rect 27982 1300 27988 1352
rect 28040 1340 28046 1352
rect 28353 1343 28411 1349
rect 28353 1340 28365 1343
rect 28040 1312 28365 1340
rect 28040 1300 28046 1312
rect 28353 1309 28365 1312
rect 28399 1309 28411 1343
rect 28353 1303 28411 1309
rect 29181 1343 29239 1349
rect 29181 1309 29193 1343
rect 29227 1340 29239 1343
rect 29362 1340 29368 1352
rect 29227 1312 29368 1340
rect 29227 1309 29239 1312
rect 29181 1303 29239 1309
rect 29362 1300 29368 1312
rect 29420 1300 29426 1352
rect 29546 1300 29552 1352
rect 29604 1340 29610 1352
rect 30193 1343 30251 1349
rect 30193 1340 30205 1343
rect 29604 1312 30205 1340
rect 29604 1300 29610 1312
rect 30193 1309 30205 1312
rect 30239 1309 30251 1343
rect 30193 1303 30251 1309
rect 30374 1300 30380 1352
rect 30432 1340 30438 1352
rect 31297 1343 31355 1349
rect 31297 1340 31309 1343
rect 30432 1312 31309 1340
rect 30432 1300 30438 1312
rect 31297 1309 31309 1312
rect 31343 1309 31355 1343
rect 31297 1303 31355 1309
rect 31754 1300 31760 1352
rect 31812 1300 31818 1352
rect 31938 1300 31944 1352
rect 31996 1340 32002 1352
rect 32217 1343 32275 1349
rect 32217 1340 32229 1343
rect 31996 1312 32229 1340
rect 31996 1300 32002 1312
rect 32217 1309 32229 1312
rect 32263 1309 32275 1343
rect 32217 1303 32275 1309
rect 32306 1300 32312 1352
rect 32364 1340 32370 1352
rect 33321 1343 33379 1349
rect 33321 1340 33333 1343
rect 32364 1312 33333 1340
rect 32364 1300 32370 1312
rect 33321 1309 33333 1312
rect 33367 1309 33379 1343
rect 33321 1303 33379 1309
rect 25516 1244 26004 1272
rect 25317 1235 25375 1241
rect 19107 1176 19196 1204
rect 19107 1173 19119 1176
rect 19061 1167 19119 1173
rect 19702 1164 19708 1216
rect 19760 1164 19766 1216
rect 20070 1164 20076 1216
rect 20128 1164 20134 1216
rect 20438 1164 20444 1216
rect 20496 1164 20502 1216
rect 21542 1164 21548 1216
rect 21600 1164 21606 1216
rect 22005 1207 22063 1213
rect 22005 1173 22017 1207
rect 22051 1204 22063 1207
rect 22480 1204 22508 1232
rect 22051 1176 22508 1204
rect 22051 1173 22063 1176
rect 22005 1167 22063 1173
rect 23014 1164 23020 1216
rect 23072 1164 23078 1216
rect 23106 1164 23112 1216
rect 23164 1204 23170 1216
rect 23385 1207 23443 1213
rect 23385 1204 23397 1207
rect 23164 1176 23397 1204
rect 23164 1164 23170 1176
rect 23385 1173 23397 1176
rect 23431 1173 23443 1207
rect 23385 1167 23443 1173
rect 23750 1164 23756 1216
rect 23808 1164 23814 1216
rect 24762 1164 24768 1216
rect 24820 1204 24826 1216
rect 24857 1207 24915 1213
rect 24857 1204 24869 1207
rect 24820 1176 24869 1204
rect 24820 1164 24826 1176
rect 24857 1173 24869 1176
rect 24903 1173 24915 1207
rect 24857 1167 24915 1173
rect 25038 1164 25044 1216
rect 25096 1204 25102 1216
rect 25976 1213 26004 1244
rect 29270 1232 29276 1284
rect 29328 1272 29334 1284
rect 29641 1275 29699 1281
rect 29641 1272 29653 1275
rect 29328 1244 29653 1272
rect 29328 1232 29334 1244
rect 29641 1241 29653 1244
rect 29687 1241 29699 1275
rect 29641 1235 29699 1241
rect 30466 1232 30472 1284
rect 30524 1272 30530 1284
rect 30745 1275 30803 1281
rect 30745 1272 30757 1275
rect 30524 1244 30757 1272
rect 30524 1232 30530 1244
rect 30745 1241 30757 1244
rect 30791 1241 30803 1275
rect 31772 1272 31800 1300
rect 32769 1275 32827 1281
rect 32769 1272 32781 1275
rect 31772 1244 32781 1272
rect 30745 1235 30803 1241
rect 32769 1241 32781 1244
rect 32815 1241 32827 1275
rect 32769 1235 32827 1241
rect 33042 1232 33048 1284
rect 33100 1272 33106 1284
rect 33520 1272 33548 1380
rect 35069 1377 35081 1380
rect 35115 1377 35127 1411
rect 35069 1371 35127 1377
rect 35710 1368 35716 1420
rect 35768 1408 35774 1420
rect 37645 1411 37703 1417
rect 37645 1408 37657 1411
rect 35768 1380 37657 1408
rect 35768 1368 35774 1380
rect 37645 1377 37657 1380
rect 37691 1377 37703 1411
rect 37645 1371 37703 1377
rect 38378 1368 38384 1420
rect 38436 1408 38442 1420
rect 40052 1408 40080 1507
rect 41414 1504 41420 1556
rect 41472 1504 41478 1556
rect 41506 1504 41512 1556
rect 41564 1544 41570 1556
rect 43441 1547 43499 1553
rect 43441 1544 43453 1547
rect 41564 1516 43453 1544
rect 41564 1504 41570 1516
rect 43441 1513 43453 1516
rect 43487 1513 43499 1547
rect 43441 1507 43499 1513
rect 44174 1504 44180 1556
rect 44232 1544 44238 1556
rect 45281 1547 45339 1553
rect 45281 1544 45293 1547
rect 44232 1516 45293 1544
rect 44232 1504 44238 1516
rect 45281 1513 45293 1516
rect 45327 1513 45339 1547
rect 45281 1507 45339 1513
rect 38436 1380 40080 1408
rect 41432 1408 41460 1504
rect 44266 1436 44272 1488
rect 44324 1476 44330 1488
rect 45005 1479 45063 1485
rect 45005 1476 45017 1479
rect 44324 1448 45017 1476
rect 44324 1436 44330 1448
rect 45005 1445 45017 1448
rect 45051 1445 45063 1479
rect 45005 1439 45063 1445
rect 41432 1380 43760 1408
rect 38436 1368 38442 1380
rect 33594 1300 33600 1352
rect 33652 1340 33658 1352
rect 33873 1343 33931 1349
rect 33873 1340 33885 1343
rect 33652 1312 33885 1340
rect 33652 1300 33658 1312
rect 33873 1309 33885 1312
rect 33919 1309 33931 1343
rect 33873 1303 33931 1309
rect 36630 1300 36636 1352
rect 36688 1340 36694 1352
rect 37369 1343 37427 1349
rect 37369 1340 37381 1343
rect 36688 1312 37381 1340
rect 36688 1300 36694 1312
rect 37369 1309 37381 1312
rect 37415 1309 37427 1343
rect 37369 1303 37427 1309
rect 37734 1300 37740 1352
rect 37792 1340 37798 1352
rect 37921 1343 37979 1349
rect 37921 1340 37933 1343
rect 37792 1312 37933 1340
rect 37792 1300 37798 1312
rect 37921 1309 37933 1312
rect 37967 1309 37979 1343
rect 37921 1303 37979 1309
rect 38194 1300 38200 1352
rect 38252 1340 38258 1352
rect 38473 1343 38531 1349
rect 38473 1340 38485 1343
rect 38252 1312 38485 1340
rect 38252 1300 38258 1312
rect 38473 1309 38485 1312
rect 38519 1309 38531 1343
rect 38473 1303 38531 1309
rect 39022 1300 39028 1352
rect 39080 1300 39086 1352
rect 39298 1300 39304 1352
rect 39356 1340 39362 1352
rect 39669 1343 39727 1349
rect 39669 1340 39681 1343
rect 39356 1312 39681 1340
rect 39356 1300 39362 1312
rect 39669 1309 39681 1312
rect 39715 1309 39727 1343
rect 39669 1303 39727 1309
rect 40034 1300 40040 1352
rect 40092 1340 40098 1352
rect 40589 1343 40647 1349
rect 40589 1340 40601 1343
rect 40092 1312 40601 1340
rect 40092 1300 40098 1312
rect 40589 1309 40601 1312
rect 40635 1309 40647 1343
rect 40589 1303 40647 1309
rect 40865 1343 40923 1349
rect 40865 1309 40877 1343
rect 40911 1309 40923 1343
rect 40865 1303 40923 1309
rect 40957 1343 41015 1349
rect 40957 1309 40969 1343
rect 41003 1309 41015 1343
rect 40957 1303 41015 1309
rect 33100 1244 33548 1272
rect 33100 1232 33106 1244
rect 34146 1232 34152 1284
rect 34204 1272 34210 1284
rect 34793 1275 34851 1281
rect 34793 1272 34805 1275
rect 34204 1244 34805 1272
rect 34204 1232 34210 1244
rect 34793 1241 34805 1244
rect 34839 1241 34851 1275
rect 34793 1235 34851 1241
rect 35342 1232 35348 1284
rect 35400 1232 35406 1284
rect 35894 1232 35900 1284
rect 35952 1232 35958 1284
rect 36446 1232 36452 1284
rect 36504 1232 36510 1284
rect 36538 1232 36544 1284
rect 36596 1272 36602 1284
rect 39945 1275 40003 1281
rect 39945 1272 39957 1275
rect 36596 1244 39957 1272
rect 36596 1232 36602 1244
rect 39945 1241 39957 1244
rect 39991 1241 40003 1275
rect 39945 1235 40003 1241
rect 40218 1232 40224 1284
rect 40276 1272 40282 1284
rect 40880 1272 40908 1303
rect 40276 1244 40908 1272
rect 40972 1272 41000 1303
rect 41230 1300 41236 1352
rect 41288 1300 41294 1352
rect 41414 1300 41420 1352
rect 41472 1340 41478 1352
rect 42061 1343 42119 1349
rect 42061 1340 42073 1343
rect 41472 1312 42073 1340
rect 41472 1300 41478 1312
rect 42061 1309 42073 1312
rect 42107 1309 42119 1343
rect 42061 1303 42119 1309
rect 42242 1300 42248 1352
rect 42300 1340 42306 1352
rect 42613 1343 42671 1349
rect 42613 1340 42625 1343
rect 42300 1312 42625 1340
rect 42300 1300 42306 1312
rect 42613 1309 42625 1312
rect 42659 1309 42671 1343
rect 42613 1303 42671 1309
rect 42702 1300 42708 1352
rect 42760 1340 42766 1352
rect 42889 1343 42947 1349
rect 42889 1340 42901 1343
rect 42760 1312 42901 1340
rect 42760 1300 42766 1312
rect 42889 1309 42901 1312
rect 42935 1309 42947 1343
rect 42889 1303 42947 1309
rect 43254 1300 43260 1352
rect 43312 1300 43318 1352
rect 43622 1300 43628 1352
rect 43680 1300 43686 1352
rect 43732 1340 43760 1380
rect 43732 1312 43944 1340
rect 41322 1272 41328 1284
rect 40972 1244 41328 1272
rect 40276 1232 40282 1244
rect 41322 1232 41328 1244
rect 41380 1232 41386 1284
rect 41984 1244 43852 1272
rect 41984 1216 42012 1244
rect 25409 1207 25467 1213
rect 25409 1204 25421 1207
rect 25096 1176 25421 1204
rect 25096 1164 25102 1176
rect 25409 1173 25421 1176
rect 25455 1173 25467 1207
rect 25409 1167 25467 1173
rect 25961 1207 26019 1213
rect 25961 1173 25973 1207
rect 26007 1173 26019 1207
rect 25961 1167 26019 1173
rect 30006 1164 30012 1216
rect 30064 1204 30070 1216
rect 31389 1207 31447 1213
rect 31389 1204 31401 1207
rect 30064 1176 31401 1204
rect 30064 1164 30070 1176
rect 31389 1173 31401 1176
rect 31435 1173 31447 1207
rect 31389 1167 31447 1173
rect 32674 1164 32680 1216
rect 32732 1204 32738 1216
rect 33965 1207 34023 1213
rect 33965 1204 33977 1207
rect 32732 1176 33977 1204
rect 32732 1164 32738 1176
rect 33965 1173 33977 1176
rect 34011 1173 34023 1207
rect 33965 1167 34023 1173
rect 34238 1164 34244 1216
rect 34296 1204 34302 1216
rect 35989 1207 36047 1213
rect 35989 1204 36001 1207
rect 34296 1176 36001 1204
rect 34296 1164 34302 1176
rect 35989 1173 36001 1176
rect 36035 1173 36047 1207
rect 35989 1167 36047 1173
rect 37366 1164 37372 1216
rect 37424 1204 37430 1216
rect 40405 1207 40463 1213
rect 40405 1204 40417 1207
rect 37424 1176 40417 1204
rect 37424 1164 37430 1176
rect 40405 1173 40417 1176
rect 40451 1173 40463 1207
rect 40405 1167 40463 1173
rect 40494 1164 40500 1216
rect 40552 1204 40558 1216
rect 40681 1207 40739 1213
rect 40681 1204 40693 1207
rect 40552 1176 40693 1204
rect 40552 1164 40558 1176
rect 40681 1173 40693 1176
rect 40727 1173 40739 1207
rect 40681 1167 40739 1173
rect 40862 1164 40868 1216
rect 40920 1204 40926 1216
rect 41877 1207 41935 1213
rect 41877 1204 41889 1207
rect 40920 1176 41889 1204
rect 40920 1164 40926 1176
rect 41877 1173 41889 1176
rect 41923 1173 41935 1207
rect 41877 1167 41935 1173
rect 41966 1164 41972 1216
rect 42024 1164 42030 1216
rect 42426 1164 42432 1216
rect 42484 1164 42490 1216
rect 42702 1164 42708 1216
rect 42760 1164 42766 1216
rect 43070 1164 43076 1216
rect 43128 1164 43134 1216
rect 43824 1213 43852 1244
rect 43809 1207 43867 1213
rect 43809 1173 43821 1207
rect 43855 1173 43867 1207
rect 43916 1204 43944 1312
rect 43990 1300 43996 1352
rect 44048 1300 44054 1352
rect 44082 1300 44088 1352
rect 44140 1340 44146 1352
rect 44361 1343 44419 1349
rect 44361 1340 44373 1343
rect 44140 1312 44373 1340
rect 44140 1300 44146 1312
rect 44361 1309 44373 1312
rect 44407 1309 44419 1343
rect 44361 1303 44419 1309
rect 44726 1300 44732 1352
rect 44784 1300 44790 1352
rect 44818 1300 44824 1352
rect 44876 1340 44882 1352
rect 45189 1343 45247 1349
rect 45189 1340 45201 1343
rect 44876 1312 45201 1340
rect 44876 1300 44882 1312
rect 45189 1309 45201 1312
rect 45235 1309 45247 1343
rect 45189 1303 45247 1309
rect 45278 1300 45284 1352
rect 45336 1340 45342 1352
rect 45465 1343 45523 1349
rect 45465 1340 45477 1343
rect 45336 1312 45477 1340
rect 45336 1300 45342 1312
rect 45465 1309 45477 1312
rect 45511 1309 45523 1343
rect 45465 1303 45523 1309
rect 44450 1232 44456 1284
rect 44508 1232 44514 1284
rect 44177 1207 44235 1213
rect 44177 1204 44189 1207
rect 43916 1176 44189 1204
rect 43809 1167 43867 1173
rect 44177 1173 44189 1176
rect 44223 1173 44235 1207
rect 44468 1204 44496 1232
rect 44545 1207 44603 1213
rect 44545 1204 44557 1207
rect 44468 1176 44557 1204
rect 44177 1167 44235 1173
rect 44545 1173 44557 1176
rect 44591 1173 44603 1207
rect 44545 1167 44603 1173
rect 1104 1114 45976 1136
rect 1104 1062 12128 1114
rect 12180 1062 12192 1114
rect 12244 1062 12256 1114
rect 12308 1062 12320 1114
rect 12372 1062 12384 1114
rect 12436 1062 23306 1114
rect 23358 1062 23370 1114
rect 23422 1062 23434 1114
rect 23486 1062 23498 1114
rect 23550 1062 23562 1114
rect 23614 1062 34484 1114
rect 34536 1062 34548 1114
rect 34600 1062 34612 1114
rect 34664 1062 34676 1114
rect 34728 1062 34740 1114
rect 34792 1062 45662 1114
rect 45714 1062 45726 1114
rect 45778 1062 45790 1114
rect 45842 1062 45854 1114
rect 45906 1062 45918 1114
rect 45970 1062 45976 1114
rect 1104 1040 45976 1062
rect 6546 960 6552 1012
rect 6604 1000 6610 1012
rect 6604 972 12434 1000
rect 6604 960 6610 972
rect 4614 892 4620 944
rect 4672 892 4678 944
rect 6914 892 6920 944
rect 6972 932 6978 944
rect 7282 932 7288 944
rect 6972 904 7288 932
rect 6972 892 6978 904
rect 7282 892 7288 904
rect 7340 892 7346 944
rect 7926 892 7932 944
rect 7984 892 7990 944
rect 8294 892 8300 944
rect 8352 932 8358 944
rect 11330 932 11336 944
rect 8352 904 11336 932
rect 8352 892 8358 904
rect 11330 892 11336 904
rect 11388 892 11394 944
rect 12406 932 12434 972
rect 12802 960 12808 1012
rect 12860 1000 12866 1012
rect 12860 972 25728 1000
rect 12860 960 12866 972
rect 13722 932 13728 944
rect 12406 904 13728 932
rect 13722 892 13728 904
rect 13780 892 13786 944
rect 14458 892 14464 944
rect 14516 932 14522 944
rect 14516 904 25636 932
rect 14516 892 14522 904
rect 4632 796 4660 892
rect 7944 864 7972 892
rect 14550 864 14556 876
rect 7944 836 14556 864
rect 14550 824 14556 836
rect 14608 824 14614 876
rect 21082 824 21088 876
rect 21140 864 21146 876
rect 23198 864 23204 876
rect 21140 836 23204 864
rect 21140 824 21146 836
rect 23198 824 23204 836
rect 23256 824 23262 876
rect 4632 768 7328 796
rect 1946 688 1952 740
rect 2004 688 2010 740
rect 4982 688 4988 740
rect 5040 728 5046 740
rect 5040 700 7144 728
rect 5040 688 5046 700
rect 1964 592 1992 688
rect 6914 592 6920 604
rect 1964 564 6920 592
rect 6914 552 6920 564
rect 6972 552 6978 604
rect 6086 484 6092 536
rect 6144 484 6150 536
rect 6104 388 6132 484
rect 7116 456 7144 700
rect 7190 688 7196 740
rect 7248 688 7254 740
rect 7208 592 7236 688
rect 7300 660 7328 768
rect 8478 756 8484 808
rect 8536 796 8542 808
rect 12618 796 12624 808
rect 8536 768 12624 796
rect 8536 756 8542 768
rect 12618 756 12624 768
rect 12676 756 12682 808
rect 12710 756 12716 808
rect 12768 796 12774 808
rect 25406 796 25412 808
rect 12768 768 25412 796
rect 12768 756 12774 768
rect 25406 756 25412 768
rect 25464 756 25470 808
rect 10134 688 10140 740
rect 10192 728 10198 740
rect 10192 700 22094 728
rect 10192 688 10198 700
rect 22066 660 22094 700
rect 25498 660 25504 672
rect 7300 632 15424 660
rect 22066 632 25504 660
rect 14734 592 14740 604
rect 7208 564 14740 592
rect 14734 552 14740 564
rect 14792 552 14798 604
rect 7558 484 7564 536
rect 7616 524 7622 536
rect 15010 524 15016 536
rect 7616 496 15016 524
rect 7616 484 7622 496
rect 15010 484 15016 496
rect 15068 484 15074 536
rect 15396 524 15424 632
rect 25498 620 25504 632
rect 25556 620 25562 672
rect 25608 660 25636 904
rect 25700 864 25728 972
rect 27798 960 27804 1012
rect 27856 1000 27862 1012
rect 34146 1000 34152 1012
rect 27856 972 34152 1000
rect 27856 960 27862 972
rect 34146 960 34152 972
rect 34204 960 34210 1012
rect 35342 960 35348 1012
rect 35400 960 35406 1012
rect 35452 972 39344 1000
rect 28166 892 28172 944
rect 28224 932 28230 944
rect 35360 932 35388 960
rect 28224 904 35388 932
rect 28224 892 28230 904
rect 28534 864 28540 876
rect 25700 836 28540 864
rect 28534 824 28540 836
rect 28592 824 28598 876
rect 28810 824 28816 876
rect 28868 864 28874 876
rect 35452 864 35480 972
rect 28868 836 35480 864
rect 39316 864 39344 972
rect 39390 960 39396 1012
rect 39448 1000 39454 1012
rect 41230 1000 41236 1012
rect 39448 972 41236 1000
rect 39448 960 39454 972
rect 41230 960 41236 972
rect 41288 960 41294 1012
rect 43070 960 43076 1012
rect 43128 960 43134 1012
rect 43088 932 43116 960
rect 40972 904 43116 932
rect 40972 864 41000 904
rect 39316 836 41000 864
rect 28868 824 28874 836
rect 42426 824 42432 876
rect 42484 824 42490 876
rect 42702 824 42708 876
rect 42760 824 42766 876
rect 28074 756 28080 808
rect 28132 796 28138 808
rect 38746 796 38752 808
rect 28132 768 38752 796
rect 28132 756 28138 768
rect 38746 756 38752 768
rect 38804 756 38810 808
rect 38838 756 38844 808
rect 38896 796 38902 808
rect 38896 768 41414 796
rect 38896 756 38902 768
rect 28350 688 28356 740
rect 28408 728 28414 740
rect 39482 728 39488 740
rect 28408 700 39488 728
rect 28408 688 28414 700
rect 39482 688 39488 700
rect 39540 688 39546 740
rect 41386 728 41414 768
rect 41966 728 41972 740
rect 41386 700 41972 728
rect 41966 688 41972 700
rect 42024 688 42030 740
rect 29638 660 29644 672
rect 25608 632 29644 660
rect 29638 620 29644 632
rect 29696 620 29702 672
rect 29822 620 29828 672
rect 29880 660 29886 672
rect 42444 660 42472 824
rect 29880 632 42472 660
rect 29880 620 29886 632
rect 17494 552 17500 604
rect 17552 592 17558 604
rect 36446 592 36452 604
rect 17552 564 36452 592
rect 17552 552 17558 564
rect 36446 552 36452 564
rect 36504 552 36510 604
rect 38746 552 38752 604
rect 38804 592 38810 604
rect 40862 592 40868 604
rect 38804 564 40868 592
rect 38804 552 38810 564
rect 40862 552 40868 564
rect 40920 552 40926 604
rect 22922 524 22928 536
rect 15396 496 22928 524
rect 22922 484 22928 496
rect 22980 484 22986 536
rect 25130 484 25136 536
rect 25188 524 25194 536
rect 42720 524 42748 824
rect 25188 496 42748 524
rect 25188 484 25194 496
rect 7116 428 21128 456
rect 13078 388 13084 400
rect 6104 360 13084 388
rect 13078 348 13084 360
rect 13136 348 13142 400
rect 13446 348 13452 400
rect 13504 388 13510 400
rect 20622 388 20628 400
rect 13504 360 20628 388
rect 13504 348 13510 360
rect 20622 348 20628 360
rect 20680 348 20686 400
rect 21100 388 21128 428
rect 21726 416 21732 468
rect 21784 456 21790 468
rect 40494 456 40500 468
rect 21784 428 40500 456
rect 21784 416 21790 428
rect 40494 416 40500 428
rect 40552 416 40558 468
rect 22002 388 22008 400
rect 21100 360 22008 388
rect 22002 348 22008 360
rect 22060 348 22066 400
rect 30650 348 30656 400
rect 30708 348 30714 400
rect 31202 348 31208 400
rect 31260 388 31266 400
rect 35894 388 35900 400
rect 31260 360 35900 388
rect 31260 348 31266 360
rect 35894 348 35900 360
rect 35952 348 35958 400
rect 3510 280 3516 332
rect 3568 320 3574 332
rect 10410 320 10416 332
rect 3568 292 10416 320
rect 3568 280 3574 292
rect 10410 280 10416 292
rect 10468 280 10474 332
rect 11146 280 11152 332
rect 11204 280 11210 332
rect 13354 280 13360 332
rect 13412 280 13418 332
rect 22278 280 22284 332
rect 22336 320 22342 332
rect 22336 292 25452 320
rect 22336 280 22342 292
rect 4154 212 4160 264
rect 4212 252 4218 264
rect 11164 252 11192 280
rect 4212 224 11192 252
rect 4212 212 4218 224
rect 13372 116 13400 280
rect 13814 212 13820 264
rect 13872 252 13878 264
rect 24026 252 24032 264
rect 13872 224 24032 252
rect 13872 212 13878 224
rect 24026 212 24032 224
rect 24084 212 24090 264
rect 25424 252 25452 292
rect 25498 280 25504 332
rect 25556 320 25562 332
rect 30668 320 30696 348
rect 25556 292 30696 320
rect 25556 280 25562 292
rect 29822 252 29828 264
rect 25424 224 29828 252
rect 29822 212 29828 224
rect 29880 212 29886 264
rect 26878 184 26884 196
rect 19306 156 26884 184
rect 19306 116 19334 156
rect 26878 144 26884 156
rect 26936 144 26942 196
rect 27338 144 27344 196
rect 27396 144 27402 196
rect 13372 88 19334 116
rect 20622 76 20628 128
rect 20680 116 20686 128
rect 27356 116 27384 144
rect 20680 88 27384 116
rect 20680 76 20686 88
rect 11238 8 11244 60
rect 11296 48 11302 60
rect 30190 48 30196 60
rect 11296 20 30196 48
rect 11296 8 11302 20
rect 30190 8 30196 20
rect 30248 8 30254 60
<< via1 >>
rect 14924 8984 14976 9036
rect 23020 8984 23072 9036
rect 22744 8916 22796 8968
rect 6184 8780 6236 8832
rect 6276 8780 6328 8832
rect 23940 8848 23992 8900
rect 10140 8780 10192 8832
rect 27528 8780 27580 8832
rect 12128 8678 12180 8730
rect 12192 8678 12244 8730
rect 12256 8678 12308 8730
rect 12320 8678 12372 8730
rect 12384 8678 12436 8730
rect 23306 8678 23358 8730
rect 23370 8678 23422 8730
rect 23434 8678 23486 8730
rect 23498 8678 23550 8730
rect 23562 8678 23614 8730
rect 34484 8678 34536 8730
rect 34548 8678 34600 8730
rect 34612 8678 34664 8730
rect 34676 8678 34728 8730
rect 34740 8678 34792 8730
rect 45662 8678 45714 8730
rect 45726 8678 45778 8730
rect 45790 8678 45842 8730
rect 45854 8678 45906 8730
rect 45918 8678 45970 8730
rect 3608 8576 3660 8628
rect 5816 8576 5868 8628
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 10140 8576 10192 8628
rect 10232 8576 10284 8628
rect 12624 8619 12676 8628
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 14648 8576 14700 8628
rect 16856 8576 16908 8628
rect 19064 8576 19116 8628
rect 21272 8576 21324 8628
rect 23664 8619 23716 8628
rect 23664 8585 23673 8619
rect 23673 8585 23707 8619
rect 23707 8585 23716 8619
rect 23664 8576 23716 8585
rect 25688 8576 25740 8628
rect 27896 8576 27948 8628
rect 30104 8619 30156 8628
rect 30104 8585 30113 8619
rect 30113 8585 30147 8619
rect 30147 8585 30156 8619
rect 30104 8576 30156 8585
rect 32312 8576 32364 8628
rect 34980 8619 35032 8628
rect 34980 8585 34989 8619
rect 34989 8585 35023 8619
rect 35023 8585 35032 8619
rect 34980 8576 35032 8585
rect 36728 8576 36780 8628
rect 38936 8576 38988 8628
rect 41144 8619 41196 8628
rect 41144 8585 41153 8619
rect 41153 8585 41187 8619
rect 41187 8585 41196 8619
rect 41144 8576 41196 8585
rect 43352 8576 43404 8628
rect 45560 8576 45612 8628
rect 1400 8551 1452 8560
rect 1400 8517 1409 8551
rect 1409 8517 1443 8551
rect 1443 8517 1452 8551
rect 1400 8508 1452 8517
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 23112 8508 23164 8560
rect 6276 8372 6328 8424
rect 14924 8440 14976 8492
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 21640 8483 21692 8492
rect 21640 8449 21649 8483
rect 21649 8449 21683 8483
rect 21683 8449 21692 8483
rect 21640 8440 21692 8449
rect 23756 8483 23808 8492
rect 23756 8449 23765 8483
rect 23765 8449 23799 8483
rect 23799 8449 23808 8483
rect 23756 8440 23808 8449
rect 26056 8483 26108 8492
rect 26056 8449 26065 8483
rect 26065 8449 26099 8483
rect 26099 8449 26108 8483
rect 26056 8440 26108 8449
rect 28264 8483 28316 8492
rect 28264 8449 28273 8483
rect 28273 8449 28307 8483
rect 28307 8449 28316 8483
rect 28264 8440 28316 8449
rect 30380 8483 30432 8492
rect 30380 8449 30389 8483
rect 30389 8449 30423 8483
rect 30423 8449 30432 8483
rect 30380 8440 30432 8449
rect 32680 8483 32732 8492
rect 32680 8449 32689 8483
rect 32689 8449 32723 8483
rect 32723 8449 32732 8483
rect 32680 8440 32732 8449
rect 35072 8483 35124 8492
rect 35072 8449 35081 8483
rect 35081 8449 35115 8483
rect 35115 8449 35124 8483
rect 35072 8440 35124 8449
rect 37096 8483 37148 8492
rect 37096 8449 37105 8483
rect 37105 8449 37139 8483
rect 37139 8449 37148 8483
rect 37096 8440 37148 8449
rect 39304 8483 39356 8492
rect 39304 8449 39313 8483
rect 39313 8449 39347 8483
rect 39347 8449 39356 8483
rect 39304 8440 39356 8449
rect 41420 8483 41472 8492
rect 41420 8449 41429 8483
rect 41429 8449 41463 8483
rect 41463 8449 41472 8483
rect 41420 8440 41472 8449
rect 43720 8483 43772 8492
rect 43720 8449 43729 8483
rect 43729 8449 43763 8483
rect 43763 8449 43772 8483
rect 43720 8440 43772 8449
rect 45100 8483 45152 8492
rect 45100 8449 45109 8483
rect 45109 8449 45143 8483
rect 45143 8449 45152 8483
rect 45100 8440 45152 8449
rect 19984 8372 20036 8424
rect 23664 8304 23716 8356
rect 6539 8134 6591 8186
rect 6603 8134 6655 8186
rect 6667 8134 6719 8186
rect 6731 8134 6783 8186
rect 6795 8134 6847 8186
rect 17717 8134 17769 8186
rect 17781 8134 17833 8186
rect 17845 8134 17897 8186
rect 17909 8134 17961 8186
rect 17973 8134 18025 8186
rect 28895 8134 28947 8186
rect 28959 8134 29011 8186
rect 29023 8134 29075 8186
rect 29087 8134 29139 8186
rect 29151 8134 29203 8186
rect 40073 8134 40125 8186
rect 40137 8134 40189 8186
rect 40201 8134 40253 8186
rect 40265 8134 40317 8186
rect 40329 8134 40381 8186
rect 12128 7590 12180 7642
rect 12192 7590 12244 7642
rect 12256 7590 12308 7642
rect 12320 7590 12372 7642
rect 12384 7590 12436 7642
rect 23306 7590 23358 7642
rect 23370 7590 23422 7642
rect 23434 7590 23486 7642
rect 23498 7590 23550 7642
rect 23562 7590 23614 7642
rect 34484 7590 34536 7642
rect 34548 7590 34600 7642
rect 34612 7590 34664 7642
rect 34676 7590 34728 7642
rect 34740 7590 34792 7642
rect 45662 7590 45714 7642
rect 45726 7590 45778 7642
rect 45790 7590 45842 7642
rect 45854 7590 45906 7642
rect 45918 7590 45970 7642
rect 6539 7046 6591 7098
rect 6603 7046 6655 7098
rect 6667 7046 6719 7098
rect 6731 7046 6783 7098
rect 6795 7046 6847 7098
rect 17717 7046 17769 7098
rect 17781 7046 17833 7098
rect 17845 7046 17897 7098
rect 17909 7046 17961 7098
rect 17973 7046 18025 7098
rect 28895 7046 28947 7098
rect 28959 7046 29011 7098
rect 29023 7046 29075 7098
rect 29087 7046 29139 7098
rect 29151 7046 29203 7098
rect 40073 7046 40125 7098
rect 40137 7046 40189 7098
rect 40201 7046 40253 7098
rect 40265 7046 40317 7098
rect 40329 7046 40381 7098
rect 12128 6502 12180 6554
rect 12192 6502 12244 6554
rect 12256 6502 12308 6554
rect 12320 6502 12372 6554
rect 12384 6502 12436 6554
rect 23306 6502 23358 6554
rect 23370 6502 23422 6554
rect 23434 6502 23486 6554
rect 23498 6502 23550 6554
rect 23562 6502 23614 6554
rect 34484 6502 34536 6554
rect 34548 6502 34600 6554
rect 34612 6502 34664 6554
rect 34676 6502 34728 6554
rect 34740 6502 34792 6554
rect 45662 6502 45714 6554
rect 45726 6502 45778 6554
rect 45790 6502 45842 6554
rect 45854 6502 45906 6554
rect 45918 6502 45970 6554
rect 6539 5958 6591 6010
rect 6603 5958 6655 6010
rect 6667 5958 6719 6010
rect 6731 5958 6783 6010
rect 6795 5958 6847 6010
rect 17717 5958 17769 6010
rect 17781 5958 17833 6010
rect 17845 5958 17897 6010
rect 17909 5958 17961 6010
rect 17973 5958 18025 6010
rect 28895 5958 28947 6010
rect 28959 5958 29011 6010
rect 29023 5958 29075 6010
rect 29087 5958 29139 6010
rect 29151 5958 29203 6010
rect 40073 5958 40125 6010
rect 40137 5958 40189 6010
rect 40201 5958 40253 6010
rect 40265 5958 40317 6010
rect 40329 5958 40381 6010
rect 12128 5414 12180 5466
rect 12192 5414 12244 5466
rect 12256 5414 12308 5466
rect 12320 5414 12372 5466
rect 12384 5414 12436 5466
rect 23306 5414 23358 5466
rect 23370 5414 23422 5466
rect 23434 5414 23486 5466
rect 23498 5414 23550 5466
rect 23562 5414 23614 5466
rect 34484 5414 34536 5466
rect 34548 5414 34600 5466
rect 34612 5414 34664 5466
rect 34676 5414 34728 5466
rect 34740 5414 34792 5466
rect 45662 5414 45714 5466
rect 45726 5414 45778 5466
rect 45790 5414 45842 5466
rect 45854 5414 45906 5466
rect 45918 5414 45970 5466
rect 6539 4870 6591 4922
rect 6603 4870 6655 4922
rect 6667 4870 6719 4922
rect 6731 4870 6783 4922
rect 6795 4870 6847 4922
rect 17717 4870 17769 4922
rect 17781 4870 17833 4922
rect 17845 4870 17897 4922
rect 17909 4870 17961 4922
rect 17973 4870 18025 4922
rect 28895 4870 28947 4922
rect 28959 4870 29011 4922
rect 29023 4870 29075 4922
rect 29087 4870 29139 4922
rect 29151 4870 29203 4922
rect 40073 4870 40125 4922
rect 40137 4870 40189 4922
rect 40201 4870 40253 4922
rect 40265 4870 40317 4922
rect 40329 4870 40381 4922
rect 4988 4496 5040 4548
rect 26148 4496 26200 4548
rect 9404 4428 9456 4480
rect 32128 4428 32180 4480
rect 12128 4326 12180 4378
rect 12192 4326 12244 4378
rect 12256 4326 12308 4378
rect 12320 4326 12372 4378
rect 12384 4326 12436 4378
rect 23306 4326 23358 4378
rect 23370 4326 23422 4378
rect 23434 4326 23486 4378
rect 23498 4326 23550 4378
rect 23562 4326 23614 4378
rect 34484 4326 34536 4378
rect 34548 4326 34600 4378
rect 34612 4326 34664 4378
rect 34676 4326 34728 4378
rect 34740 4326 34792 4378
rect 45662 4326 45714 4378
rect 45726 4326 45778 4378
rect 45790 4326 45842 4378
rect 45854 4326 45906 4378
rect 45918 4326 45970 4378
rect 18788 4224 18840 4276
rect 41604 4224 41656 4276
rect 2780 4156 2832 4208
rect 26424 4156 26476 4208
rect 6539 3782 6591 3834
rect 6603 3782 6655 3834
rect 6667 3782 6719 3834
rect 6731 3782 6783 3834
rect 6795 3782 6847 3834
rect 17717 3782 17769 3834
rect 17781 3782 17833 3834
rect 17845 3782 17897 3834
rect 17909 3782 17961 3834
rect 17973 3782 18025 3834
rect 28895 3782 28947 3834
rect 28959 3782 29011 3834
rect 29023 3782 29075 3834
rect 29087 3782 29139 3834
rect 29151 3782 29203 3834
rect 40073 3782 40125 3834
rect 40137 3782 40189 3834
rect 40201 3782 40253 3834
rect 40265 3782 40317 3834
rect 40329 3782 40381 3834
rect 6920 3544 6972 3596
rect 22468 3544 22520 3596
rect 17132 3476 17184 3528
rect 36636 3476 36688 3528
rect 21824 3408 21876 3460
rect 31760 3408 31812 3460
rect 19156 3340 19208 3392
rect 38660 3340 38712 3392
rect 12128 3238 12180 3290
rect 12192 3238 12244 3290
rect 12256 3238 12308 3290
rect 12320 3238 12372 3290
rect 12384 3238 12436 3290
rect 23306 3238 23358 3290
rect 23370 3238 23422 3290
rect 23434 3238 23486 3290
rect 23498 3238 23550 3290
rect 23562 3238 23614 3290
rect 34484 3238 34536 3290
rect 34548 3238 34600 3290
rect 34612 3238 34664 3290
rect 34676 3238 34728 3290
rect 34740 3238 34792 3290
rect 45662 3238 45714 3290
rect 45726 3238 45778 3290
rect 45790 3238 45842 3290
rect 45854 3238 45906 3290
rect 45918 3238 45970 3290
rect 11152 3136 11204 3188
rect 24492 3136 24544 3188
rect 11428 3068 11480 3120
rect 26332 3068 26384 3120
rect 8484 3000 8536 3052
rect 23204 3000 23256 3052
rect 23848 3000 23900 3052
rect 35532 3000 35584 3052
rect 16488 2932 16540 2984
rect 35716 2932 35768 2984
rect 5632 2864 5684 2916
rect 20536 2864 20588 2916
rect 34336 2864 34388 2916
rect 14556 2796 14608 2848
rect 19248 2796 19300 2848
rect 26700 2796 26752 2848
rect 27712 2796 27764 2848
rect 30012 2796 30064 2848
rect 30104 2796 30156 2848
rect 31852 2796 31904 2848
rect 32588 2796 32640 2848
rect 37464 2796 37516 2848
rect 6539 2694 6591 2746
rect 6603 2694 6655 2746
rect 6667 2694 6719 2746
rect 6731 2694 6783 2746
rect 6795 2694 6847 2746
rect 17717 2694 17769 2746
rect 17781 2694 17833 2746
rect 17845 2694 17897 2746
rect 17909 2694 17961 2746
rect 17973 2694 18025 2746
rect 28895 2694 28947 2746
rect 28959 2694 29011 2746
rect 29023 2694 29075 2746
rect 29087 2694 29139 2746
rect 29151 2694 29203 2746
rect 40073 2694 40125 2746
rect 40137 2694 40189 2746
rect 40201 2694 40253 2746
rect 40265 2694 40317 2746
rect 40329 2694 40381 2746
rect 17224 2592 17276 2644
rect 19616 2567 19668 2576
rect 19616 2533 19625 2567
rect 19625 2533 19659 2567
rect 19659 2533 19668 2567
rect 19616 2524 19668 2533
rect 20444 2524 20496 2576
rect 22192 2524 22244 2576
rect 22744 2635 22796 2644
rect 22744 2601 22753 2635
rect 22753 2601 22787 2635
rect 22787 2601 22796 2635
rect 22744 2592 22796 2601
rect 23020 2635 23072 2644
rect 23020 2601 23029 2635
rect 23029 2601 23063 2635
rect 23063 2601 23072 2635
rect 23020 2592 23072 2601
rect 23112 2592 23164 2644
rect 23664 2592 23716 2644
rect 23756 2592 23808 2644
rect 23940 2635 23992 2644
rect 23940 2601 23949 2635
rect 23949 2601 23983 2635
rect 23983 2601 23992 2635
rect 23940 2592 23992 2601
rect 24032 2592 24084 2644
rect 26884 2592 26936 2644
rect 15016 2456 15068 2508
rect 14740 2388 14792 2440
rect 17500 2388 17552 2440
rect 17592 2431 17644 2440
rect 17592 2397 17601 2431
rect 17601 2397 17635 2431
rect 17635 2397 17644 2431
rect 17592 2388 17644 2397
rect 18052 2388 18104 2440
rect 18696 2388 18748 2440
rect 18972 2388 19024 2440
rect 19616 2388 19668 2440
rect 19708 2431 19760 2440
rect 19708 2397 19717 2431
rect 19717 2397 19751 2431
rect 19751 2397 19760 2431
rect 19708 2388 19760 2397
rect 14280 2320 14332 2372
rect 12624 2252 12676 2304
rect 17684 2252 17736 2304
rect 19064 2295 19116 2304
rect 19064 2261 19073 2295
rect 19073 2261 19107 2295
rect 19107 2261 19116 2295
rect 19064 2252 19116 2261
rect 19248 2252 19300 2304
rect 20076 2388 20128 2440
rect 19984 2320 20036 2372
rect 19892 2295 19944 2304
rect 19892 2261 19901 2295
rect 19901 2261 19935 2295
rect 19935 2261 19944 2295
rect 19892 2252 19944 2261
rect 20352 2388 20404 2440
rect 20904 2431 20956 2440
rect 20904 2397 20913 2431
rect 20913 2397 20947 2431
rect 20947 2397 20956 2431
rect 20904 2388 20956 2397
rect 21180 2431 21232 2440
rect 21180 2397 21189 2431
rect 21189 2397 21223 2431
rect 21223 2397 21232 2431
rect 21180 2388 21232 2397
rect 21640 2388 21692 2440
rect 22652 2456 22704 2508
rect 26056 2567 26108 2576
rect 26056 2533 26065 2567
rect 26065 2533 26099 2567
rect 26099 2533 26108 2567
rect 26056 2524 26108 2533
rect 28264 2635 28316 2644
rect 28264 2601 28273 2635
rect 28273 2601 28307 2635
rect 28307 2601 28316 2635
rect 28264 2592 28316 2601
rect 31484 2592 31536 2644
rect 31668 2592 31720 2644
rect 31944 2524 31996 2576
rect 32680 2635 32732 2644
rect 32680 2601 32689 2635
rect 32689 2601 32723 2635
rect 32723 2601 32732 2635
rect 32680 2592 32732 2601
rect 35072 2635 35124 2644
rect 35072 2601 35081 2635
rect 35081 2601 35115 2635
rect 35115 2601 35124 2635
rect 35072 2592 35124 2601
rect 36912 2592 36964 2644
rect 37188 2592 37240 2644
rect 37556 2592 37608 2644
rect 39488 2635 39540 2644
rect 39488 2601 39497 2635
rect 39497 2601 39531 2635
rect 39531 2601 39540 2635
rect 39488 2592 39540 2601
rect 33140 2524 33192 2576
rect 34336 2524 34388 2576
rect 39580 2524 39632 2576
rect 20168 2252 20220 2304
rect 20260 2252 20312 2304
rect 20628 2295 20680 2304
rect 20628 2261 20637 2295
rect 20637 2261 20671 2295
rect 20671 2261 20680 2295
rect 20628 2252 20680 2261
rect 21088 2295 21140 2304
rect 21088 2261 21097 2295
rect 21097 2261 21131 2295
rect 21131 2261 21140 2295
rect 21088 2252 21140 2261
rect 22284 2388 22336 2440
rect 22468 2431 22520 2440
rect 22468 2397 22477 2431
rect 22477 2397 22511 2431
rect 22511 2397 22520 2431
rect 22468 2388 22520 2397
rect 22928 2431 22980 2440
rect 22928 2397 22937 2431
rect 22937 2397 22971 2431
rect 22971 2397 22980 2431
rect 22928 2388 22980 2397
rect 23020 2388 23072 2440
rect 24124 2456 24176 2508
rect 23756 2431 23808 2440
rect 23756 2397 23765 2431
rect 23765 2397 23799 2431
rect 23799 2397 23808 2431
rect 23756 2388 23808 2397
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 22100 2295 22152 2304
rect 22100 2261 22109 2295
rect 22109 2261 22143 2295
rect 22143 2261 22152 2295
rect 22100 2252 22152 2261
rect 25044 2320 25096 2372
rect 26332 2431 26384 2440
rect 26332 2397 26341 2431
rect 26341 2397 26375 2431
rect 26375 2397 26384 2431
rect 26332 2388 26384 2397
rect 26608 2431 26660 2440
rect 26608 2397 26617 2431
rect 26617 2397 26651 2431
rect 26651 2397 26660 2431
rect 26608 2388 26660 2397
rect 26884 2431 26936 2440
rect 26884 2397 26893 2431
rect 26893 2397 26927 2431
rect 26927 2397 26936 2431
rect 26884 2388 26936 2397
rect 22744 2252 22796 2304
rect 26792 2295 26844 2304
rect 26792 2261 26801 2295
rect 26801 2261 26835 2295
rect 26835 2261 26844 2295
rect 26792 2252 26844 2261
rect 27068 2295 27120 2304
rect 27068 2261 27077 2295
rect 27077 2261 27111 2295
rect 27111 2261 27120 2295
rect 27068 2252 27120 2261
rect 27712 2456 27764 2508
rect 30932 2456 30984 2508
rect 31484 2456 31536 2508
rect 31760 2456 31812 2508
rect 41420 2592 41472 2644
rect 43720 2592 43772 2644
rect 45100 2592 45152 2644
rect 27436 2431 27488 2440
rect 27436 2397 27445 2431
rect 27445 2397 27479 2431
rect 27479 2397 27488 2431
rect 27436 2388 27488 2397
rect 27620 2388 27672 2440
rect 28448 2431 28500 2440
rect 28448 2397 28457 2431
rect 28457 2397 28491 2431
rect 28491 2397 28500 2431
rect 28448 2388 28500 2397
rect 29828 2388 29880 2440
rect 28816 2320 28868 2372
rect 28908 2320 28960 2372
rect 30288 2320 30340 2372
rect 30748 2431 30800 2440
rect 30748 2397 30757 2431
rect 30757 2397 30791 2431
rect 30791 2397 30800 2431
rect 30748 2388 30800 2397
rect 30840 2388 30892 2440
rect 31392 2431 31444 2440
rect 31392 2397 31401 2431
rect 31401 2397 31435 2431
rect 31435 2397 31444 2431
rect 31392 2388 31444 2397
rect 32036 2388 32088 2440
rect 32220 2388 32272 2440
rect 32312 2388 32364 2440
rect 44456 2456 44508 2508
rect 33232 2388 33284 2440
rect 34888 2431 34940 2440
rect 34888 2397 34897 2431
rect 34897 2397 34931 2431
rect 34931 2397 34940 2431
rect 34888 2388 34940 2397
rect 35348 2388 35400 2440
rect 37188 2388 37240 2440
rect 27988 2252 28040 2304
rect 28080 2295 28132 2304
rect 28080 2261 28089 2295
rect 28089 2261 28123 2295
rect 28123 2261 28132 2295
rect 28080 2252 28132 2261
rect 30472 2295 30524 2304
rect 30472 2261 30481 2295
rect 30481 2261 30515 2295
rect 30515 2261 30524 2295
rect 30472 2252 30524 2261
rect 30932 2295 30984 2304
rect 30932 2261 30941 2295
rect 30941 2261 30975 2295
rect 30975 2261 30984 2295
rect 30932 2252 30984 2261
rect 31300 2295 31352 2304
rect 31300 2261 31309 2295
rect 31309 2261 31343 2295
rect 31343 2261 31352 2295
rect 31300 2252 31352 2261
rect 31760 2252 31812 2304
rect 32956 2252 33008 2304
rect 33232 2295 33284 2304
rect 33232 2261 33241 2295
rect 33241 2261 33275 2295
rect 33275 2261 33284 2295
rect 33232 2252 33284 2261
rect 37464 2388 37516 2440
rect 38844 2388 38896 2440
rect 39672 2431 39724 2440
rect 39672 2397 39681 2431
rect 39681 2397 39715 2431
rect 39715 2397 39724 2431
rect 39672 2388 39724 2397
rect 39764 2388 39816 2440
rect 41512 2388 41564 2440
rect 41788 2431 41840 2440
rect 41788 2397 41797 2431
rect 41797 2397 41831 2431
rect 41831 2397 41840 2431
rect 41788 2388 41840 2397
rect 44180 2431 44232 2440
rect 44180 2397 44189 2431
rect 44189 2397 44223 2431
rect 44223 2397 44232 2431
rect 44180 2388 44232 2397
rect 44916 2388 44968 2440
rect 45192 2431 45244 2440
rect 45192 2397 45201 2431
rect 45201 2397 45235 2431
rect 45235 2397 45244 2431
rect 45192 2388 45244 2397
rect 45928 2388 45980 2440
rect 37556 2320 37608 2372
rect 41420 2320 41472 2372
rect 37188 2252 37240 2304
rect 37372 2252 37424 2304
rect 37832 2252 37884 2304
rect 44272 2252 44324 2304
rect 45008 2295 45060 2304
rect 45008 2261 45017 2295
rect 45017 2261 45051 2295
rect 45051 2261 45060 2295
rect 45008 2252 45060 2261
rect 45284 2295 45336 2304
rect 45284 2261 45293 2295
rect 45293 2261 45327 2295
rect 45327 2261 45336 2295
rect 45284 2252 45336 2261
rect 12128 2150 12180 2202
rect 12192 2150 12244 2202
rect 12256 2150 12308 2202
rect 12320 2150 12372 2202
rect 12384 2150 12436 2202
rect 23306 2150 23358 2202
rect 23370 2150 23422 2202
rect 23434 2150 23486 2202
rect 23498 2150 23550 2202
rect 23562 2150 23614 2202
rect 34484 2150 34536 2202
rect 34548 2150 34600 2202
rect 34612 2150 34664 2202
rect 34676 2150 34728 2202
rect 34740 2150 34792 2202
rect 45662 2150 45714 2202
rect 45726 2150 45778 2202
rect 45790 2150 45842 2202
rect 45854 2150 45906 2202
rect 45918 2150 45970 2202
rect 2780 2091 2832 2100
rect 2780 2057 2789 2091
rect 2789 2057 2823 2091
rect 2823 2057 2832 2091
rect 2780 2048 2832 2057
rect 4988 2048 5040 2100
rect 9404 2091 9456 2100
rect 9404 2057 9413 2091
rect 9413 2057 9447 2091
rect 9447 2057 9456 2091
rect 9404 2048 9456 2057
rect 9588 2048 9640 2100
rect 13728 2048 13780 2100
rect 16212 2091 16264 2100
rect 16212 2057 16221 2091
rect 16221 2057 16255 2091
rect 16255 2057 16264 2091
rect 16212 2048 16264 2057
rect 16488 2091 16540 2100
rect 16488 2057 16497 2091
rect 16497 2057 16531 2091
rect 16531 2057 16540 2091
rect 16488 2048 16540 2057
rect 17592 2048 17644 2100
rect 18972 2091 19024 2100
rect 18972 2057 18981 2091
rect 18981 2057 19015 2091
rect 19015 2057 19024 2091
rect 18972 2048 19024 2057
rect 19248 2091 19300 2100
rect 19248 2057 19257 2091
rect 19257 2057 19291 2091
rect 19291 2057 19300 2091
rect 19248 2048 19300 2057
rect 19616 2048 19668 2100
rect 20076 2048 20128 2100
rect 20628 2048 20680 2100
rect 21088 2048 21140 2100
rect 22928 2048 22980 2100
rect 23020 2091 23072 2100
rect 23020 2057 23029 2091
rect 23029 2057 23063 2091
rect 23063 2057 23072 2091
rect 23020 2048 23072 2057
rect 23756 2048 23808 2100
rect 24584 2048 24636 2100
rect 25044 2091 25096 2100
rect 25044 2057 25053 2091
rect 25053 2057 25087 2091
rect 25087 2057 25096 2091
rect 25044 2048 25096 2057
rect 25136 2048 25188 2100
rect 25412 2048 25464 2100
rect 17316 1980 17368 2032
rect 17500 1980 17552 2032
rect 19708 1980 19760 2032
rect 664 1912 716 1964
rect 1032 1844 1084 1896
rect 2596 1955 2648 1964
rect 2596 1921 2605 1955
rect 2605 1921 2639 1955
rect 2639 1921 2648 1955
rect 2596 1912 2648 1921
rect 2964 1955 3016 1964
rect 2964 1921 2973 1955
rect 2973 1921 3007 1955
rect 3007 1921 3016 1955
rect 2964 1912 3016 1921
rect 9220 1955 9272 1964
rect 9220 1921 9229 1955
rect 9229 1921 9263 1955
rect 9263 1921 9272 1955
rect 9220 1912 9272 1921
rect 9588 1955 9640 1964
rect 9588 1921 9597 1955
rect 9597 1921 9631 1955
rect 9631 1921 9640 1955
rect 9588 1912 9640 1921
rect 15108 1912 15160 1964
rect 15476 1955 15528 1964
rect 15476 1921 15485 1955
rect 15485 1921 15519 1955
rect 15519 1921 15528 1955
rect 15476 1912 15528 1921
rect 15752 1955 15804 1964
rect 15752 1921 15761 1955
rect 15761 1921 15795 1955
rect 15795 1921 15804 1955
rect 15752 1912 15804 1921
rect 16028 1955 16080 1964
rect 16028 1921 16037 1955
rect 16037 1921 16071 1955
rect 16071 1921 16080 1955
rect 16028 1912 16080 1921
rect 16304 1955 16356 1964
rect 16304 1921 16313 1955
rect 16313 1921 16347 1955
rect 16347 1921 16356 1955
rect 16304 1912 16356 1921
rect 16856 1955 16908 1964
rect 16856 1921 16865 1955
rect 16865 1921 16899 1955
rect 16899 1921 16908 1955
rect 16856 1912 16908 1921
rect 17132 1955 17184 1964
rect 17132 1921 17141 1955
rect 17141 1921 17175 1955
rect 17175 1921 17184 1955
rect 17132 1912 17184 1921
rect 17408 1955 17460 1964
rect 17408 1921 17417 1955
rect 17417 1921 17451 1955
rect 17451 1921 17460 1955
rect 17408 1912 17460 1921
rect 17684 1955 17736 1964
rect 17684 1921 17693 1955
rect 17693 1921 17727 1955
rect 17727 1921 17736 1955
rect 17684 1912 17736 1921
rect 18144 1912 18196 1964
rect 16764 1844 16816 1896
rect 16948 1844 17000 1896
rect 18512 1955 18564 1964
rect 18512 1921 18521 1955
rect 18521 1921 18555 1955
rect 18555 1921 18564 1955
rect 18512 1912 18564 1921
rect 18788 1955 18840 1964
rect 18788 1921 18797 1955
rect 18797 1921 18831 1955
rect 18831 1921 18840 1955
rect 18788 1912 18840 1921
rect 19064 1955 19116 1964
rect 19064 1921 19073 1955
rect 19073 1921 19107 1955
rect 19107 1921 19116 1955
rect 19064 1912 19116 1921
rect 19340 1955 19392 1964
rect 19340 1921 19349 1955
rect 19349 1921 19383 1955
rect 19383 1921 19392 1955
rect 19340 1912 19392 1921
rect 19616 1955 19668 1964
rect 19616 1921 19625 1955
rect 19625 1921 19659 1955
rect 19659 1921 19668 1955
rect 19616 1912 19668 1921
rect 18328 1844 18380 1896
rect 20076 1912 20128 1964
rect 20260 1912 20312 1964
rect 20536 1844 20588 1896
rect 21732 1912 21784 1964
rect 22008 1912 22060 1964
rect 22836 1955 22888 1964
rect 22836 1921 22845 1955
rect 22845 1921 22879 1955
rect 22879 1921 22888 1955
rect 22836 1912 22888 1921
rect 22928 1912 22980 1964
rect 23388 1955 23440 1964
rect 23388 1921 23397 1955
rect 23397 1921 23431 1955
rect 23431 1921 23440 1955
rect 23388 1912 23440 1921
rect 23848 1955 23900 1964
rect 23848 1921 23857 1955
rect 23857 1921 23891 1955
rect 23891 1921 23900 1955
rect 23848 1912 23900 1921
rect 1584 1751 1636 1760
rect 1584 1717 1593 1751
rect 1593 1717 1627 1751
rect 1627 1717 1636 1751
rect 1584 1708 1636 1717
rect 15660 1751 15712 1760
rect 15660 1717 15669 1751
rect 15669 1717 15703 1751
rect 15703 1717 15712 1751
rect 15660 1708 15712 1717
rect 17500 1708 17552 1760
rect 18236 1776 18288 1828
rect 19340 1776 19392 1828
rect 20720 1776 20772 1828
rect 23480 1776 23532 1828
rect 24492 1955 24544 1964
rect 24492 1921 24501 1955
rect 24501 1921 24535 1955
rect 24535 1921 24544 1955
rect 24492 1912 24544 1921
rect 25136 1912 25188 1964
rect 26700 1980 26752 2032
rect 26792 1980 26844 2032
rect 28448 2048 28500 2100
rect 30380 2091 30432 2100
rect 30380 2057 30389 2091
rect 30389 2057 30423 2091
rect 30423 2057 30432 2091
rect 30380 2048 30432 2057
rect 30932 2048 30984 2100
rect 31300 2048 31352 2100
rect 25320 1955 25372 1964
rect 25320 1921 25329 1955
rect 25329 1921 25363 1955
rect 25363 1921 25372 1955
rect 25320 1912 25372 1921
rect 26148 1955 26200 1964
rect 26148 1921 26157 1955
rect 26157 1921 26191 1955
rect 26191 1921 26200 1955
rect 26148 1912 26200 1921
rect 26424 1955 26476 1964
rect 26424 1921 26433 1955
rect 26433 1921 26467 1955
rect 26467 1921 26476 1955
rect 26424 1912 26476 1921
rect 25320 1776 25372 1828
rect 27528 1887 27580 1896
rect 27528 1853 27537 1887
rect 27537 1853 27571 1887
rect 27571 1853 27580 1887
rect 27528 1844 27580 1853
rect 28080 1912 28132 1964
rect 28540 1912 28592 1964
rect 28356 1844 28408 1896
rect 32036 2048 32088 2100
rect 33140 1980 33192 2032
rect 34888 2048 34940 2100
rect 34244 1980 34296 2032
rect 35532 2048 35584 2100
rect 29644 1955 29696 1964
rect 29644 1921 29653 1955
rect 29653 1921 29687 1955
rect 29687 1921 29696 1955
rect 29644 1912 29696 1921
rect 30012 1912 30064 1964
rect 30196 1955 30248 1964
rect 30196 1921 30205 1955
rect 30205 1921 30239 1955
rect 30239 1921 30248 1955
rect 30196 1912 30248 1921
rect 30472 1955 30524 1964
rect 30472 1921 30481 1955
rect 30481 1921 30515 1955
rect 30515 1921 30524 1955
rect 30472 1912 30524 1921
rect 31300 1887 31352 1896
rect 31300 1853 31309 1887
rect 31309 1853 31343 1887
rect 31343 1853 31352 1887
rect 31300 1844 31352 1853
rect 17960 1708 18012 1760
rect 18604 1708 18656 1760
rect 19984 1708 20036 1760
rect 20260 1708 20312 1760
rect 20352 1751 20404 1760
rect 20352 1717 20361 1751
rect 20361 1717 20395 1751
rect 20395 1717 20404 1751
rect 20352 1708 20404 1717
rect 20628 1751 20680 1760
rect 20628 1717 20637 1751
rect 20637 1717 20671 1751
rect 20671 1717 20680 1751
rect 20628 1708 20680 1717
rect 21088 1708 21140 1760
rect 21180 1751 21232 1760
rect 21180 1717 21189 1751
rect 21189 1717 21223 1751
rect 21223 1717 21232 1751
rect 21180 1708 21232 1717
rect 22376 1751 22428 1760
rect 22376 1717 22385 1751
rect 22385 1717 22419 1751
rect 22419 1717 22428 1751
rect 22376 1708 22428 1717
rect 22560 1708 22612 1760
rect 23296 1751 23348 1760
rect 23296 1717 23305 1751
rect 23305 1717 23339 1751
rect 23339 1717 23348 1751
rect 23296 1708 23348 1717
rect 23572 1751 23624 1760
rect 23572 1717 23581 1751
rect 23581 1717 23615 1751
rect 23615 1717 23624 1751
rect 23572 1708 23624 1717
rect 23848 1708 23900 1760
rect 25872 1708 25924 1760
rect 26884 1776 26936 1828
rect 27620 1776 27672 1828
rect 27896 1776 27948 1828
rect 26332 1751 26384 1760
rect 26332 1717 26341 1751
rect 26341 1717 26375 1751
rect 26375 1717 26384 1751
rect 26332 1708 26384 1717
rect 26424 1708 26476 1760
rect 27252 1708 27304 1760
rect 29368 1776 29420 1828
rect 29644 1776 29696 1828
rect 30472 1776 30524 1828
rect 32128 1955 32180 1964
rect 32128 1921 32137 1955
rect 32137 1921 32171 1955
rect 32171 1921 32180 1955
rect 32128 1912 32180 1921
rect 32588 1955 32640 1964
rect 32588 1921 32597 1955
rect 32597 1921 32631 1955
rect 32631 1921 32640 1955
rect 32588 1912 32640 1921
rect 35348 1955 35400 1964
rect 35348 1921 35357 1955
rect 35357 1921 35391 1955
rect 35391 1921 35400 1955
rect 35348 1912 35400 1921
rect 35716 1980 35768 2032
rect 31852 1887 31904 1896
rect 31852 1853 31861 1887
rect 31861 1853 31895 1887
rect 31895 1853 31904 1887
rect 31852 1844 31904 1853
rect 32312 1819 32364 1828
rect 32312 1785 32321 1819
rect 32321 1785 32355 1819
rect 32355 1785 32364 1819
rect 32312 1776 32364 1785
rect 32404 1819 32456 1828
rect 32404 1785 32413 1819
rect 32413 1785 32447 1819
rect 32447 1785 32456 1819
rect 32404 1776 32456 1785
rect 29276 1751 29328 1760
rect 29276 1717 29285 1751
rect 29285 1717 29319 1751
rect 29319 1717 29328 1751
rect 29276 1708 29328 1717
rect 29552 1751 29604 1760
rect 29552 1717 29561 1751
rect 29561 1717 29595 1751
rect 29595 1717 29604 1751
rect 29552 1708 29604 1717
rect 30288 1708 30340 1760
rect 32588 1776 32640 1828
rect 33048 1708 33100 1760
rect 33416 1708 33468 1760
rect 34336 1776 34388 1828
rect 37096 1844 37148 1896
rect 35716 1776 35768 1828
rect 37280 2048 37332 2100
rect 37372 2048 37424 2100
rect 38568 2048 38620 2100
rect 39672 2048 39724 2100
rect 38660 1980 38712 2032
rect 37832 1955 37884 1964
rect 37832 1921 37841 1955
rect 37841 1921 37875 1955
rect 37875 1921 37884 1955
rect 37832 1912 37884 1921
rect 38108 1955 38160 1964
rect 38108 1921 38117 1955
rect 38117 1921 38151 1955
rect 38151 1921 38160 1955
rect 38108 1912 38160 1921
rect 38752 1955 38804 1964
rect 38752 1921 38761 1955
rect 38761 1921 38795 1955
rect 38795 1921 38804 1955
rect 38752 1912 38804 1921
rect 41788 2048 41840 2100
rect 44180 2048 44232 2100
rect 44916 2091 44968 2100
rect 44916 2057 44925 2091
rect 44925 2057 44959 2091
rect 44959 2057 44968 2091
rect 44916 2048 44968 2057
rect 45008 2048 45060 2100
rect 45284 2048 45336 2100
rect 40592 1955 40644 1964
rect 40592 1921 40601 1955
rect 40601 1921 40635 1955
rect 40635 1921 40644 1955
rect 40592 1912 40644 1921
rect 40684 1912 40736 1964
rect 40776 1844 40828 1896
rect 41604 1955 41656 1964
rect 41604 1921 41613 1955
rect 41613 1921 41647 1955
rect 41647 1921 41656 1955
rect 41604 1912 41656 1921
rect 34888 1708 34940 1760
rect 36268 1751 36320 1760
rect 36268 1717 36277 1751
rect 36277 1717 36311 1751
rect 36311 1717 36320 1751
rect 36268 1708 36320 1717
rect 44180 1844 44232 1896
rect 45468 1955 45520 1964
rect 45468 1921 45477 1955
rect 45477 1921 45511 1955
rect 45511 1921 45520 1955
rect 45468 1912 45520 1921
rect 41880 1776 41932 1828
rect 37280 1708 37332 1760
rect 38476 1708 38528 1760
rect 38936 1708 38988 1760
rect 6539 1606 6591 1658
rect 6603 1606 6655 1658
rect 6667 1606 6719 1658
rect 6731 1606 6783 1658
rect 6795 1606 6847 1658
rect 17717 1606 17769 1658
rect 17781 1606 17833 1658
rect 17845 1606 17897 1658
rect 17909 1606 17961 1658
rect 17973 1606 18025 1658
rect 28895 1606 28947 1658
rect 28959 1606 29011 1658
rect 29023 1606 29075 1658
rect 29087 1606 29139 1658
rect 29151 1606 29203 1658
rect 40073 1606 40125 1658
rect 40137 1606 40189 1658
rect 40201 1606 40253 1658
rect 40265 1606 40317 1658
rect 40329 1606 40381 1658
rect 1584 1504 1636 1556
rect 9680 1504 9732 1556
rect 14280 1547 14332 1556
rect 14280 1513 14289 1547
rect 14289 1513 14323 1547
rect 14323 1513 14332 1547
rect 14280 1504 14332 1513
rect 15108 1547 15160 1556
rect 15108 1513 15117 1547
rect 15117 1513 15151 1547
rect 15151 1513 15160 1547
rect 15108 1504 15160 1513
rect 15476 1504 15528 1556
rect 15752 1504 15804 1556
rect 16028 1504 16080 1556
rect 16304 1504 16356 1556
rect 16488 1547 16540 1556
rect 16488 1513 16497 1547
rect 16497 1513 16531 1547
rect 16531 1513 16540 1547
rect 16488 1504 16540 1513
rect 17132 1504 17184 1556
rect 17408 1504 17460 1556
rect 18052 1504 18104 1556
rect 18144 1504 18196 1556
rect 18512 1504 18564 1556
rect 19064 1504 19116 1556
rect 19616 1504 19668 1556
rect 17592 1436 17644 1488
rect 18236 1436 18288 1488
rect 1492 1343 1544 1352
rect 1492 1309 1501 1343
rect 1501 1309 1535 1343
rect 1535 1309 1544 1343
rect 1492 1300 1544 1309
rect 1860 1343 1912 1352
rect 1860 1309 1869 1343
rect 1869 1309 1903 1343
rect 1903 1309 1912 1343
rect 1860 1300 1912 1309
rect 2228 1343 2280 1352
rect 2228 1309 2237 1343
rect 2237 1309 2271 1343
rect 2271 1309 2280 1343
rect 2228 1300 2280 1309
rect 3240 1300 3292 1352
rect 3332 1343 3384 1352
rect 3332 1309 3341 1343
rect 3341 1309 3375 1343
rect 3375 1309 3384 1343
rect 3332 1300 3384 1309
rect 3792 1343 3844 1352
rect 3792 1309 3801 1343
rect 3801 1309 3835 1343
rect 3835 1309 3844 1343
rect 3792 1300 3844 1309
rect 4068 1343 4120 1352
rect 4068 1309 4077 1343
rect 4077 1309 4111 1343
rect 4111 1309 4120 1343
rect 4068 1300 4120 1309
rect 4436 1343 4488 1352
rect 4436 1309 4445 1343
rect 4445 1309 4479 1343
rect 4479 1309 4488 1343
rect 4436 1300 4488 1309
rect 4804 1343 4856 1352
rect 4804 1309 4813 1343
rect 4813 1309 4847 1343
rect 4847 1309 4856 1343
rect 4804 1300 4856 1309
rect 5172 1343 5224 1352
rect 5172 1309 5181 1343
rect 5181 1309 5215 1343
rect 5215 1309 5224 1343
rect 5172 1300 5224 1309
rect 5540 1343 5592 1352
rect 5540 1309 5549 1343
rect 5549 1309 5583 1343
rect 5583 1309 5592 1343
rect 5540 1300 5592 1309
rect 5632 1300 5684 1352
rect 5908 1343 5960 1352
rect 5908 1309 5917 1343
rect 5917 1309 5951 1343
rect 5951 1309 5960 1343
rect 5908 1300 5960 1309
rect 6368 1343 6420 1352
rect 6368 1309 6377 1343
rect 6377 1309 6411 1343
rect 6411 1309 6420 1343
rect 6368 1300 6420 1309
rect 6644 1343 6696 1352
rect 6644 1309 6653 1343
rect 6653 1309 6687 1343
rect 6687 1309 6696 1343
rect 6644 1300 6696 1309
rect 6920 1300 6972 1352
rect 7012 1343 7064 1352
rect 7012 1309 7021 1343
rect 7021 1309 7055 1343
rect 7055 1309 7064 1343
rect 7012 1300 7064 1309
rect 1952 1164 2004 1216
rect 2044 1207 2096 1216
rect 2044 1173 2053 1207
rect 2053 1173 2087 1207
rect 2087 1173 2096 1207
rect 2044 1164 2096 1173
rect 3516 1207 3568 1216
rect 3516 1173 3525 1207
rect 3525 1173 3559 1207
rect 3559 1173 3568 1207
rect 3516 1164 3568 1173
rect 4160 1164 4212 1216
rect 4620 1207 4672 1216
rect 4620 1173 4629 1207
rect 4629 1173 4663 1207
rect 4663 1173 4672 1207
rect 4620 1164 4672 1173
rect 4988 1207 5040 1216
rect 4988 1173 4997 1207
rect 4997 1173 5031 1207
rect 5031 1173 5040 1207
rect 4988 1164 5040 1173
rect 7380 1343 7432 1352
rect 7380 1309 7389 1343
rect 7389 1309 7423 1343
rect 7423 1309 7432 1343
rect 7380 1300 7432 1309
rect 7748 1343 7800 1352
rect 7748 1309 7757 1343
rect 7757 1309 7791 1343
rect 7791 1309 7800 1343
rect 7748 1300 7800 1309
rect 8116 1343 8168 1352
rect 8116 1309 8125 1343
rect 8125 1309 8159 1343
rect 8159 1309 8168 1343
rect 8116 1300 8168 1309
rect 8484 1300 8536 1352
rect 8576 1343 8628 1352
rect 8576 1309 8585 1343
rect 8585 1309 8619 1343
rect 8619 1309 8628 1343
rect 8576 1300 8628 1309
rect 8392 1232 8444 1284
rect 9496 1300 9548 1352
rect 9956 1343 10008 1352
rect 9956 1309 9965 1343
rect 9965 1309 9999 1343
rect 9999 1309 10008 1343
rect 9956 1300 10008 1309
rect 10324 1343 10376 1352
rect 10324 1309 10333 1343
rect 10333 1309 10367 1343
rect 10367 1309 10376 1343
rect 10324 1300 10376 1309
rect 10692 1343 10744 1352
rect 10692 1309 10701 1343
rect 10701 1309 10735 1343
rect 10735 1309 10744 1343
rect 10692 1300 10744 1309
rect 11060 1343 11112 1352
rect 11060 1309 11069 1343
rect 11069 1309 11103 1343
rect 11103 1309 11112 1343
rect 11060 1300 11112 1309
rect 11520 1343 11572 1352
rect 11520 1309 11529 1343
rect 11529 1309 11563 1343
rect 11563 1309 11572 1343
rect 11520 1300 11572 1309
rect 11796 1343 11848 1352
rect 11796 1309 11805 1343
rect 11805 1309 11839 1343
rect 11839 1309 11848 1343
rect 11796 1300 11848 1309
rect 12164 1343 12216 1352
rect 12164 1309 12173 1343
rect 12173 1309 12207 1343
rect 12207 1309 12216 1343
rect 12164 1300 12216 1309
rect 6092 1207 6144 1216
rect 6092 1173 6101 1207
rect 6101 1173 6135 1207
rect 6135 1173 6144 1207
rect 6092 1164 6144 1173
rect 6552 1207 6604 1216
rect 6552 1173 6561 1207
rect 6561 1173 6595 1207
rect 6595 1173 6604 1207
rect 6552 1164 6604 1173
rect 7196 1207 7248 1216
rect 7196 1173 7205 1207
rect 7205 1173 7239 1207
rect 7239 1173 7248 1207
rect 7196 1164 7248 1173
rect 7564 1207 7616 1216
rect 7564 1173 7573 1207
rect 7573 1173 7607 1207
rect 7607 1173 7616 1207
rect 7564 1164 7616 1173
rect 7932 1207 7984 1216
rect 7932 1173 7941 1207
rect 7941 1173 7975 1207
rect 7975 1173 7984 1207
rect 7932 1164 7984 1173
rect 8300 1207 8352 1216
rect 8300 1173 8309 1207
rect 8309 1173 8343 1207
rect 8343 1173 8352 1207
rect 8300 1164 8352 1173
rect 8760 1207 8812 1216
rect 8760 1173 8769 1207
rect 8769 1173 8803 1207
rect 8803 1173 8812 1207
rect 8760 1164 8812 1173
rect 10140 1207 10192 1216
rect 10140 1173 10149 1207
rect 10149 1173 10183 1207
rect 10183 1173 10192 1207
rect 10140 1164 10192 1173
rect 11428 1232 11480 1284
rect 10876 1207 10928 1216
rect 10876 1173 10885 1207
rect 10885 1173 10919 1207
rect 10919 1173 10928 1207
rect 10876 1164 10928 1173
rect 11244 1207 11296 1216
rect 11244 1173 11253 1207
rect 11253 1173 11287 1207
rect 11287 1173 11296 1207
rect 11244 1164 11296 1173
rect 11888 1164 11940 1216
rect 12532 1343 12584 1352
rect 12532 1309 12541 1343
rect 12541 1309 12575 1343
rect 12575 1309 12584 1343
rect 12532 1300 12584 1309
rect 12808 1300 12860 1352
rect 12900 1343 12952 1352
rect 12900 1309 12909 1343
rect 12909 1309 12943 1343
rect 12943 1309 12952 1343
rect 12900 1300 12952 1309
rect 13268 1343 13320 1352
rect 13268 1309 13277 1343
rect 13277 1309 13311 1343
rect 13311 1309 13320 1343
rect 13268 1300 13320 1309
rect 13636 1343 13688 1352
rect 13636 1309 13645 1343
rect 13645 1309 13679 1343
rect 13679 1309 13688 1343
rect 13636 1300 13688 1309
rect 14096 1343 14148 1352
rect 14096 1309 14105 1343
rect 14105 1309 14139 1343
rect 14139 1309 14148 1343
rect 14096 1300 14148 1309
rect 14372 1343 14424 1352
rect 14372 1309 14381 1343
rect 14381 1309 14415 1343
rect 14415 1309 14424 1343
rect 14372 1300 14424 1309
rect 12716 1207 12768 1216
rect 12716 1173 12725 1207
rect 12725 1173 12759 1207
rect 12759 1173 12768 1207
rect 12716 1164 12768 1173
rect 13360 1164 13412 1216
rect 13452 1207 13504 1216
rect 13452 1173 13461 1207
rect 13461 1173 13495 1207
rect 13495 1173 13504 1207
rect 13452 1164 13504 1173
rect 13820 1207 13872 1216
rect 13820 1173 13829 1207
rect 13829 1173 13863 1207
rect 13863 1173 13872 1207
rect 13820 1164 13872 1173
rect 14464 1164 14516 1216
rect 18328 1368 18380 1420
rect 14648 1343 14700 1352
rect 14648 1309 14657 1343
rect 14657 1309 14691 1343
rect 14691 1309 14700 1343
rect 14648 1300 14700 1309
rect 14924 1343 14976 1352
rect 14924 1309 14933 1343
rect 14933 1309 14967 1343
rect 14967 1309 14976 1343
rect 14924 1300 14976 1309
rect 15200 1343 15252 1352
rect 15200 1309 15209 1343
rect 15209 1309 15243 1343
rect 15243 1309 15252 1343
rect 15200 1300 15252 1309
rect 15476 1343 15528 1352
rect 15476 1309 15485 1343
rect 15485 1309 15519 1343
rect 15519 1309 15528 1343
rect 15476 1300 15528 1309
rect 16212 1300 16264 1352
rect 16580 1300 16632 1352
rect 16764 1343 16816 1352
rect 16764 1309 16773 1343
rect 16773 1309 16807 1343
rect 16807 1309 16816 1343
rect 16764 1300 16816 1309
rect 16120 1232 16172 1284
rect 16488 1232 16540 1284
rect 17684 1343 17736 1352
rect 17684 1309 17693 1343
rect 17693 1309 17727 1343
rect 17727 1309 17736 1343
rect 17684 1300 17736 1309
rect 17776 1343 17828 1352
rect 17776 1309 17785 1343
rect 17785 1309 17819 1343
rect 17819 1309 17828 1343
rect 17776 1300 17828 1309
rect 18052 1343 18104 1352
rect 18052 1309 18061 1343
rect 18061 1309 18095 1343
rect 18095 1309 18104 1343
rect 18052 1300 18104 1309
rect 18512 1343 18564 1352
rect 18512 1309 18521 1343
rect 18521 1309 18555 1343
rect 18555 1309 18564 1343
rect 18512 1300 18564 1309
rect 18788 1343 18840 1352
rect 18788 1309 18797 1343
rect 18797 1309 18831 1343
rect 18831 1309 18840 1343
rect 18788 1300 18840 1309
rect 19156 1300 19208 1352
rect 18696 1232 18748 1284
rect 17224 1207 17276 1216
rect 17224 1173 17233 1207
rect 17233 1173 17267 1207
rect 17267 1173 17276 1207
rect 17224 1164 17276 1173
rect 19984 1436 20036 1488
rect 20904 1479 20956 1488
rect 20904 1445 20913 1479
rect 20913 1445 20947 1479
rect 20947 1445 20956 1479
rect 20904 1436 20956 1445
rect 21916 1504 21968 1556
rect 22376 1504 22428 1556
rect 23940 1504 23992 1556
rect 26240 1504 26292 1556
rect 26608 1504 26660 1556
rect 27620 1504 27672 1556
rect 19340 1300 19392 1352
rect 19432 1343 19484 1352
rect 19432 1309 19441 1343
rect 19441 1309 19475 1343
rect 19475 1309 19484 1343
rect 19432 1300 19484 1309
rect 23480 1368 23532 1420
rect 23572 1368 23624 1420
rect 19984 1300 20036 1352
rect 20352 1300 20404 1352
rect 21824 1343 21876 1352
rect 21824 1309 21833 1343
rect 21833 1309 21867 1343
rect 21867 1309 21876 1343
rect 21824 1300 21876 1309
rect 22100 1300 22152 1352
rect 23204 1343 23256 1352
rect 23204 1309 23213 1343
rect 23213 1309 23247 1343
rect 23247 1309 23256 1343
rect 23204 1300 23256 1309
rect 23296 1300 23348 1352
rect 24952 1300 25004 1352
rect 26148 1368 26200 1420
rect 26608 1368 26660 1420
rect 27712 1436 27764 1488
rect 28632 1504 28684 1556
rect 29000 1436 29052 1488
rect 28080 1368 28132 1420
rect 28264 1368 28316 1420
rect 29460 1368 29512 1420
rect 31668 1504 31720 1556
rect 31024 1436 31076 1488
rect 31668 1368 31720 1420
rect 34336 1504 34388 1556
rect 34980 1436 35032 1488
rect 36912 1504 36964 1556
rect 38108 1504 38160 1556
rect 37096 1436 37148 1488
rect 39488 1479 39540 1488
rect 39488 1445 39497 1479
rect 39497 1445 39531 1479
rect 39531 1445 39540 1479
rect 39488 1436 39540 1445
rect 20720 1275 20772 1284
rect 20720 1241 20729 1275
rect 20729 1241 20763 1275
rect 20763 1241 20772 1275
rect 20720 1232 20772 1241
rect 22192 1275 22244 1284
rect 22192 1241 22201 1275
rect 22201 1241 22235 1275
rect 22235 1241 22244 1275
rect 22192 1232 22244 1241
rect 22468 1232 22520 1284
rect 22744 1232 22796 1284
rect 23940 1232 23992 1284
rect 25872 1300 25924 1352
rect 26332 1300 26384 1352
rect 27160 1300 27212 1352
rect 27988 1300 28040 1352
rect 29368 1300 29420 1352
rect 29552 1300 29604 1352
rect 30380 1300 30432 1352
rect 31760 1300 31812 1352
rect 31944 1300 31996 1352
rect 32312 1300 32364 1352
rect 19708 1207 19760 1216
rect 19708 1173 19717 1207
rect 19717 1173 19751 1207
rect 19751 1173 19760 1207
rect 19708 1164 19760 1173
rect 20076 1207 20128 1216
rect 20076 1173 20085 1207
rect 20085 1173 20119 1207
rect 20119 1173 20128 1207
rect 20076 1164 20128 1173
rect 20444 1207 20496 1216
rect 20444 1173 20453 1207
rect 20453 1173 20487 1207
rect 20487 1173 20496 1207
rect 20444 1164 20496 1173
rect 21548 1207 21600 1216
rect 21548 1173 21557 1207
rect 21557 1173 21591 1207
rect 21591 1173 21600 1207
rect 21548 1164 21600 1173
rect 23020 1207 23072 1216
rect 23020 1173 23029 1207
rect 23029 1173 23063 1207
rect 23063 1173 23072 1207
rect 23020 1164 23072 1173
rect 23112 1164 23164 1216
rect 23756 1207 23808 1216
rect 23756 1173 23765 1207
rect 23765 1173 23799 1207
rect 23799 1173 23808 1207
rect 23756 1164 23808 1173
rect 24768 1164 24820 1216
rect 25044 1164 25096 1216
rect 29276 1232 29328 1284
rect 30472 1232 30524 1284
rect 33048 1232 33100 1284
rect 35716 1368 35768 1420
rect 38384 1368 38436 1420
rect 41420 1504 41472 1556
rect 41512 1504 41564 1556
rect 44180 1504 44232 1556
rect 44272 1436 44324 1488
rect 33600 1300 33652 1352
rect 36636 1300 36688 1352
rect 37740 1300 37792 1352
rect 38200 1300 38252 1352
rect 39028 1343 39080 1352
rect 39028 1309 39037 1343
rect 39037 1309 39071 1343
rect 39071 1309 39080 1343
rect 39028 1300 39080 1309
rect 39304 1300 39356 1352
rect 40040 1300 40092 1352
rect 34152 1232 34204 1284
rect 35348 1275 35400 1284
rect 35348 1241 35357 1275
rect 35357 1241 35391 1275
rect 35391 1241 35400 1275
rect 35348 1232 35400 1241
rect 35900 1275 35952 1284
rect 35900 1241 35909 1275
rect 35909 1241 35943 1275
rect 35943 1241 35952 1275
rect 35900 1232 35952 1241
rect 36452 1275 36504 1284
rect 36452 1241 36461 1275
rect 36461 1241 36495 1275
rect 36495 1241 36504 1275
rect 36452 1232 36504 1241
rect 36544 1232 36596 1284
rect 40224 1232 40276 1284
rect 41236 1343 41288 1352
rect 41236 1309 41245 1343
rect 41245 1309 41279 1343
rect 41279 1309 41288 1343
rect 41236 1300 41288 1309
rect 41420 1300 41472 1352
rect 42248 1300 42300 1352
rect 42708 1300 42760 1352
rect 43260 1343 43312 1352
rect 43260 1309 43269 1343
rect 43269 1309 43303 1343
rect 43303 1309 43312 1343
rect 43260 1300 43312 1309
rect 43628 1343 43680 1352
rect 43628 1309 43637 1343
rect 43637 1309 43671 1343
rect 43671 1309 43680 1343
rect 43628 1300 43680 1309
rect 41328 1232 41380 1284
rect 30012 1164 30064 1216
rect 32680 1164 32732 1216
rect 34244 1164 34296 1216
rect 37372 1164 37424 1216
rect 40500 1164 40552 1216
rect 40868 1164 40920 1216
rect 41972 1164 42024 1216
rect 42432 1207 42484 1216
rect 42432 1173 42441 1207
rect 42441 1173 42475 1207
rect 42475 1173 42484 1207
rect 42432 1164 42484 1173
rect 42708 1207 42760 1216
rect 42708 1173 42717 1207
rect 42717 1173 42751 1207
rect 42751 1173 42760 1207
rect 42708 1164 42760 1173
rect 43076 1207 43128 1216
rect 43076 1173 43085 1207
rect 43085 1173 43119 1207
rect 43119 1173 43128 1207
rect 43076 1164 43128 1173
rect 43996 1343 44048 1352
rect 43996 1309 44005 1343
rect 44005 1309 44039 1343
rect 44039 1309 44048 1343
rect 43996 1300 44048 1309
rect 44088 1300 44140 1352
rect 44732 1343 44784 1352
rect 44732 1309 44741 1343
rect 44741 1309 44775 1343
rect 44775 1309 44784 1343
rect 44732 1300 44784 1309
rect 44824 1300 44876 1352
rect 45284 1300 45336 1352
rect 44456 1232 44508 1284
rect 12128 1062 12180 1114
rect 12192 1062 12244 1114
rect 12256 1062 12308 1114
rect 12320 1062 12372 1114
rect 12384 1062 12436 1114
rect 23306 1062 23358 1114
rect 23370 1062 23422 1114
rect 23434 1062 23486 1114
rect 23498 1062 23550 1114
rect 23562 1062 23614 1114
rect 34484 1062 34536 1114
rect 34548 1062 34600 1114
rect 34612 1062 34664 1114
rect 34676 1062 34728 1114
rect 34740 1062 34792 1114
rect 45662 1062 45714 1114
rect 45726 1062 45778 1114
rect 45790 1062 45842 1114
rect 45854 1062 45906 1114
rect 45918 1062 45970 1114
rect 6552 960 6604 1012
rect 4620 892 4672 944
rect 6920 892 6972 944
rect 7288 892 7340 944
rect 7932 892 7984 944
rect 8300 892 8352 944
rect 11336 892 11388 944
rect 12808 960 12860 1012
rect 13728 892 13780 944
rect 14464 892 14516 944
rect 14556 824 14608 876
rect 21088 824 21140 876
rect 23204 824 23256 876
rect 1952 688 2004 740
rect 4988 688 5040 740
rect 6920 552 6972 604
rect 6092 484 6144 536
rect 7196 688 7248 740
rect 8484 756 8536 808
rect 12624 756 12676 808
rect 12716 756 12768 808
rect 25412 756 25464 808
rect 10140 688 10192 740
rect 14740 552 14792 604
rect 7564 484 7616 536
rect 15016 484 15068 536
rect 25504 620 25556 672
rect 27804 960 27856 1012
rect 34152 960 34204 1012
rect 35348 960 35400 1012
rect 28172 892 28224 944
rect 28540 824 28592 876
rect 28816 824 28868 876
rect 39396 960 39448 1012
rect 41236 960 41288 1012
rect 43076 960 43128 1012
rect 42432 824 42484 876
rect 42708 824 42760 876
rect 28080 756 28132 808
rect 38752 756 38804 808
rect 38844 756 38896 808
rect 28356 688 28408 740
rect 39488 688 39540 740
rect 41972 688 42024 740
rect 29644 620 29696 672
rect 29828 620 29880 672
rect 17500 552 17552 604
rect 36452 552 36504 604
rect 38752 552 38804 604
rect 40868 552 40920 604
rect 22928 484 22980 536
rect 25136 484 25188 536
rect 13084 348 13136 400
rect 13452 348 13504 400
rect 20628 348 20680 400
rect 21732 416 21784 468
rect 40500 416 40552 468
rect 22008 348 22060 400
rect 30656 348 30708 400
rect 31208 348 31260 400
rect 35900 348 35952 400
rect 3516 280 3568 332
rect 10416 280 10468 332
rect 11152 280 11204 332
rect 13360 280 13412 332
rect 22284 280 22336 332
rect 4160 212 4212 264
rect 13820 212 13872 264
rect 24032 212 24084 264
rect 25504 280 25556 332
rect 29828 212 29880 264
rect 26884 144 26936 196
rect 27344 144 27396 196
rect 20628 76 20680 128
rect 11244 8 11296 60
rect 30196 8 30248 60
<< metal2 >>
rect 1398 9840 1454 10000
rect 3606 9840 3662 10000
rect 5814 9840 5870 10000
rect 8022 9840 8078 10000
rect 10230 9840 10286 10000
rect 12438 9840 12494 10000
rect 14646 9840 14702 10000
rect 16854 9840 16910 10000
rect 19062 9840 19118 10000
rect 21270 9840 21326 10000
rect 23478 9840 23534 10000
rect 25686 9840 25742 10000
rect 27894 9840 27950 10000
rect 30102 9840 30158 10000
rect 32310 9840 32366 10000
rect 34518 9840 34574 10000
rect 34624 9846 35020 9874
rect 1412 8566 1440 9840
rect 3620 8634 3648 9840
rect 5828 8634 5856 9840
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 1400 8560 1452 8566
rect 1400 8502 1452 8508
rect 6196 8498 6224 8774
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6288 8430 6316 8774
rect 8036 8634 8064 9840
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10152 8634 10180 8774
rect 10244 8634 10272 9840
rect 12452 9058 12480 9840
rect 12452 9030 12664 9058
rect 12128 8732 12436 8741
rect 12128 8730 12134 8732
rect 12190 8730 12214 8732
rect 12270 8730 12294 8732
rect 12350 8730 12374 8732
rect 12430 8730 12436 8732
rect 12190 8678 12192 8730
rect 12372 8678 12374 8730
rect 12128 8676 12134 8678
rect 12190 8676 12214 8678
rect 12270 8676 12294 8678
rect 12350 8676 12374 8678
rect 12430 8676 12436 8678
rect 12128 8667 12436 8676
rect 12636 8634 12664 9030
rect 14660 8634 14688 9840
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14936 8498 14964 8978
rect 16868 8634 16896 9840
rect 19076 8634 19104 9840
rect 21284 8634 21312 9840
rect 23492 9058 23520 9840
rect 23020 9036 23072 9042
rect 23492 9030 23704 9058
rect 23020 8978 23072 8984
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 6539 8188 6847 8197
rect 6539 8186 6545 8188
rect 6601 8186 6625 8188
rect 6681 8186 6705 8188
rect 6761 8186 6785 8188
rect 6841 8186 6847 8188
rect 6601 8134 6603 8186
rect 6783 8134 6785 8186
rect 6539 8132 6545 8134
rect 6601 8132 6625 8134
rect 6681 8132 6705 8134
rect 6761 8132 6785 8134
rect 6841 8132 6847 8134
rect 6539 8123 6847 8132
rect 12128 7644 12436 7653
rect 12128 7642 12134 7644
rect 12190 7642 12214 7644
rect 12270 7642 12294 7644
rect 12350 7642 12374 7644
rect 12430 7642 12436 7644
rect 12190 7590 12192 7642
rect 12372 7590 12374 7642
rect 12128 7588 12134 7590
rect 12190 7588 12214 7590
rect 12270 7588 12294 7590
rect 12350 7588 12374 7590
rect 12430 7588 12436 7590
rect 12128 7579 12436 7588
rect 6539 7100 6847 7109
rect 6539 7098 6545 7100
rect 6601 7098 6625 7100
rect 6681 7098 6705 7100
rect 6761 7098 6785 7100
rect 6841 7098 6847 7100
rect 6601 7046 6603 7098
rect 6783 7046 6785 7098
rect 6539 7044 6545 7046
rect 6601 7044 6625 7046
rect 6681 7044 6705 7046
rect 6761 7044 6785 7046
rect 6841 7044 6847 7046
rect 6539 7035 6847 7044
rect 12128 6556 12436 6565
rect 12128 6554 12134 6556
rect 12190 6554 12214 6556
rect 12270 6554 12294 6556
rect 12350 6554 12374 6556
rect 12430 6554 12436 6556
rect 12190 6502 12192 6554
rect 12372 6502 12374 6554
rect 12128 6500 12134 6502
rect 12190 6500 12214 6502
rect 12270 6500 12294 6502
rect 12350 6500 12374 6502
rect 12430 6500 12436 6502
rect 12128 6491 12436 6500
rect 6539 6012 6847 6021
rect 6539 6010 6545 6012
rect 6601 6010 6625 6012
rect 6681 6010 6705 6012
rect 6761 6010 6785 6012
rect 6841 6010 6847 6012
rect 6601 5958 6603 6010
rect 6783 5958 6785 6010
rect 6539 5956 6545 5958
rect 6601 5956 6625 5958
rect 6681 5956 6705 5958
rect 6761 5956 6785 5958
rect 6841 5956 6847 5958
rect 6539 5947 6847 5956
rect 12128 5468 12436 5477
rect 12128 5466 12134 5468
rect 12190 5466 12214 5468
rect 12270 5466 12294 5468
rect 12350 5466 12374 5468
rect 12430 5466 12436 5468
rect 12190 5414 12192 5466
rect 12372 5414 12374 5466
rect 12128 5412 12134 5414
rect 12190 5412 12214 5414
rect 12270 5412 12294 5414
rect 12350 5412 12374 5414
rect 12430 5412 12436 5414
rect 12128 5403 12436 5412
rect 6539 4924 6847 4933
rect 6539 4922 6545 4924
rect 6601 4922 6625 4924
rect 6681 4922 6705 4924
rect 6761 4922 6785 4924
rect 6841 4922 6847 4924
rect 6601 4870 6603 4922
rect 6783 4870 6785 4922
rect 6539 4868 6545 4870
rect 6601 4868 6625 4870
rect 6681 4868 6705 4870
rect 6761 4868 6785 4870
rect 6841 4868 6847 4870
rect 6539 4859 6847 4868
rect 3238 4584 3294 4593
rect 3238 4519 3294 4528
rect 4988 4548 5040 4554
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2792 2106 2820 4150
rect 2780 2100 2832 2106
rect 2780 2042 2832 2048
rect 664 1964 716 1970
rect 664 1906 716 1912
rect 2596 1964 2648 1970
rect 2596 1906 2648 1912
rect 2964 1964 3016 1970
rect 2964 1906 3016 1912
rect 676 160 704 1906
rect 1032 1896 1084 1902
rect 1032 1838 1084 1844
rect 1044 160 1072 1838
rect 1584 1760 1636 1766
rect 1584 1702 1636 1708
rect 1596 1562 1624 1702
rect 1584 1556 1636 1562
rect 1584 1498 1636 1504
rect 1492 1352 1544 1358
rect 1412 1312 1492 1340
rect 1412 160 1440 1312
rect 1492 1294 1544 1300
rect 1860 1352 1912 1358
rect 1860 1294 1912 1300
rect 2228 1352 2280 1358
rect 2228 1294 2280 1300
rect 662 0 718 160
rect 1030 0 1086 160
rect 1398 0 1454 160
rect 1766 82 1822 160
rect 1872 82 1900 1294
rect 1952 1216 2004 1222
rect 1952 1158 2004 1164
rect 2044 1216 2096 1222
rect 2044 1158 2096 1164
rect 1964 746 1992 1158
rect 2056 1057 2084 1158
rect 2042 1048 2098 1057
rect 2042 983 2098 992
rect 1952 740 2004 746
rect 1952 682 2004 688
rect 1766 54 1900 82
rect 2134 82 2190 160
rect 2240 82 2268 1294
rect 2134 54 2268 82
rect 2502 82 2558 160
rect 2608 82 2636 1906
rect 2502 54 2636 82
rect 2870 82 2926 160
rect 2976 82 3004 1906
rect 3252 1358 3280 4519
rect 4988 4490 5040 4496
rect 5000 2106 5028 4490
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 6539 3836 6847 3845
rect 6539 3834 6545 3836
rect 6601 3834 6625 3836
rect 6681 3834 6705 3836
rect 6761 3834 6785 3836
rect 6841 3834 6847 3836
rect 6601 3782 6603 3834
rect 6783 3782 6785 3834
rect 6539 3780 6545 3782
rect 6601 3780 6625 3782
rect 6681 3780 6705 3782
rect 6761 3780 6785 3782
rect 6841 3780 6847 3782
rect 6539 3771 6847 3780
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 4988 2100 5040 2106
rect 4988 2042 5040 2048
rect 5644 1358 5672 2858
rect 6539 2748 6847 2757
rect 6539 2746 6545 2748
rect 6601 2746 6625 2748
rect 6681 2746 6705 2748
rect 6761 2746 6785 2748
rect 6841 2746 6847 2748
rect 6601 2694 6603 2746
rect 6783 2694 6785 2746
rect 6539 2692 6545 2694
rect 6601 2692 6625 2694
rect 6681 2692 6705 2694
rect 6761 2692 6785 2694
rect 6841 2692 6847 2694
rect 6539 2683 6847 2692
rect 6539 1660 6847 1669
rect 6539 1658 6545 1660
rect 6601 1658 6625 1660
rect 6681 1658 6705 1660
rect 6761 1658 6785 1660
rect 6841 1658 6847 1660
rect 6601 1606 6603 1658
rect 6783 1606 6785 1658
rect 6539 1604 6545 1606
rect 6601 1604 6625 1606
rect 6681 1604 6705 1606
rect 6761 1604 6785 1606
rect 6841 1604 6847 1606
rect 6539 1595 6847 1604
rect 6932 1358 6960 3538
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 7286 1456 7342 1465
rect 7286 1391 7342 1400
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 3792 1352 3844 1358
rect 3792 1294 3844 1300
rect 4068 1352 4120 1358
rect 4068 1294 4120 1300
rect 4436 1352 4488 1358
rect 4436 1294 4488 1300
rect 4804 1352 4856 1358
rect 4804 1294 4856 1300
rect 5172 1352 5224 1358
rect 5172 1294 5224 1300
rect 5540 1352 5592 1358
rect 5540 1294 5592 1300
rect 5632 1352 5684 1358
rect 5632 1294 5684 1300
rect 5908 1352 5960 1358
rect 5908 1294 5960 1300
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 6920 1352 6972 1358
rect 6920 1294 6972 1300
rect 7012 1352 7064 1358
rect 7012 1294 7064 1300
rect 2870 54 3004 82
rect 3238 82 3294 160
rect 3344 82 3372 1294
rect 3516 1216 3568 1222
rect 3516 1158 3568 1164
rect 3528 338 3556 1158
rect 3516 332 3568 338
rect 3516 274 3568 280
rect 3238 54 3372 82
rect 3606 82 3662 160
rect 3804 82 3832 1294
rect 3606 54 3832 82
rect 3974 82 4030 160
rect 4080 82 4108 1294
rect 4160 1216 4212 1222
rect 4160 1158 4212 1164
rect 4172 270 4200 1158
rect 4160 264 4212 270
rect 4160 206 4212 212
rect 3974 54 4108 82
rect 4342 82 4398 160
rect 4448 82 4476 1294
rect 4620 1216 4672 1222
rect 4620 1158 4672 1164
rect 4632 950 4660 1158
rect 4620 944 4672 950
rect 4620 886 4672 892
rect 4342 54 4476 82
rect 4710 82 4766 160
rect 4816 82 4844 1294
rect 4988 1216 5040 1222
rect 4988 1158 5040 1164
rect 5000 746 5028 1158
rect 4988 740 5040 746
rect 4988 682 5040 688
rect 4710 54 4844 82
rect 5078 82 5134 160
rect 5184 82 5212 1294
rect 5078 54 5212 82
rect 5446 82 5502 160
rect 5552 82 5580 1294
rect 5446 54 5580 82
rect 5814 82 5870 160
rect 5920 82 5948 1294
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 6104 542 6132 1158
rect 6092 536 6144 542
rect 6092 478 6144 484
rect 5814 54 5948 82
rect 6182 82 6238 160
rect 6380 82 6408 1294
rect 6552 1216 6604 1222
rect 6552 1158 6604 1164
rect 6564 1018 6592 1158
rect 6552 1012 6604 1018
rect 6552 954 6604 960
rect 6182 54 6408 82
rect 6550 82 6606 160
rect 6656 82 6684 1294
rect 6920 944 6972 950
rect 6920 886 6972 892
rect 6932 610 6960 886
rect 6920 604 6972 610
rect 6920 546 6972 552
rect 6550 54 6684 82
rect 6918 82 6974 160
rect 7024 82 7052 1294
rect 7196 1216 7248 1222
rect 7196 1158 7248 1164
rect 7208 746 7236 1158
rect 7300 950 7328 1391
rect 8496 1358 8524 2994
rect 9416 2106 9444 4422
rect 12128 4380 12436 4389
rect 12128 4378 12134 4380
rect 12190 4378 12214 4380
rect 12270 4378 12294 4380
rect 12350 4378 12374 4380
rect 12430 4378 12436 4380
rect 12190 4326 12192 4378
rect 12372 4326 12374 4378
rect 12128 4324 12134 4326
rect 12190 4324 12214 4326
rect 12270 4324 12294 4326
rect 12350 4324 12374 4326
rect 12430 4324 12436 4326
rect 12128 4315 12436 4324
rect 16854 4176 16910 4185
rect 16854 4111 16910 4120
rect 10414 4040 10470 4049
rect 10414 3975 10470 3984
rect 9586 2952 9642 2961
rect 9586 2887 9642 2896
rect 9600 2106 9628 2887
rect 9404 2100 9456 2106
rect 9404 2042 9456 2048
rect 9588 2100 9640 2106
rect 9588 2042 9640 2048
rect 9678 2000 9734 2009
rect 9220 1964 9272 1970
rect 9220 1906 9272 1912
rect 9588 1964 9640 1970
rect 9678 1935 9734 1944
rect 9588 1906 9640 1912
rect 7380 1352 7432 1358
rect 7380 1294 7432 1300
rect 7748 1352 7800 1358
rect 7748 1294 7800 1300
rect 8116 1352 8168 1358
rect 8116 1294 8168 1300
rect 8484 1352 8536 1358
rect 8484 1294 8536 1300
rect 8576 1352 8628 1358
rect 8576 1294 8628 1300
rect 7288 944 7340 950
rect 7288 886 7340 892
rect 7196 740 7248 746
rect 7196 682 7248 688
rect 6918 54 7052 82
rect 7286 82 7342 160
rect 7392 82 7420 1294
rect 7564 1216 7616 1222
rect 7564 1158 7616 1164
rect 7576 542 7604 1158
rect 7564 536 7616 542
rect 7564 478 7616 484
rect 7286 54 7420 82
rect 7654 82 7710 160
rect 7760 82 7788 1294
rect 7932 1216 7984 1222
rect 7932 1158 7984 1164
rect 7944 950 7972 1158
rect 7932 944 7984 950
rect 7932 886 7984 892
rect 7654 54 7788 82
rect 8022 82 8078 160
rect 8128 82 8156 1294
rect 8392 1284 8444 1290
rect 8392 1226 8444 1232
rect 8300 1216 8352 1222
rect 8300 1158 8352 1164
rect 8312 950 8340 1158
rect 8300 944 8352 950
rect 8300 886 8352 892
rect 8404 160 8432 1226
rect 8482 1048 8538 1057
rect 8482 983 8538 992
rect 8496 814 8524 983
rect 8484 808 8536 814
rect 8484 750 8536 756
rect 8022 54 8156 82
rect 1766 0 1822 54
rect 2134 0 2190 54
rect 2502 0 2558 54
rect 2870 0 2926 54
rect 3238 0 3294 54
rect 3606 0 3662 54
rect 3974 0 4030 54
rect 4342 0 4398 54
rect 4710 0 4766 54
rect 5078 0 5134 54
rect 5446 0 5502 54
rect 5814 0 5870 54
rect 6182 0 6238 54
rect 6550 0 6606 54
rect 6918 0 6974 54
rect 7286 0 7342 54
rect 7654 0 7710 54
rect 8022 0 8078 54
rect 8390 0 8446 160
rect 8588 82 8616 1294
rect 8760 1216 8812 1222
rect 8760 1158 8812 1164
rect 8772 513 8800 1158
rect 8758 504 8814 513
rect 8758 439 8814 448
rect 8758 82 8814 160
rect 8588 54 8814 82
rect 8758 0 8814 54
rect 9126 82 9182 160
rect 9232 82 9260 1906
rect 9496 1352 9548 1358
rect 9494 1320 9496 1329
rect 9548 1320 9550 1329
rect 9494 1255 9550 1264
rect 9126 54 9260 82
rect 9494 82 9550 160
rect 9600 82 9628 1906
rect 9692 1562 9720 1935
rect 9680 1556 9732 1562
rect 9680 1498 9732 1504
rect 9956 1352 10008 1358
rect 9956 1294 10008 1300
rect 10324 1352 10376 1358
rect 10324 1294 10376 1300
rect 9494 54 9628 82
rect 9862 82 9918 160
rect 9968 82 9996 1294
rect 10140 1216 10192 1222
rect 10140 1158 10192 1164
rect 10152 746 10180 1158
rect 10140 740 10192 746
rect 10140 682 10192 688
rect 9862 54 9996 82
rect 10230 82 10286 160
rect 10336 82 10364 1294
rect 10428 338 10456 3975
rect 16210 3632 16266 3641
rect 16210 3567 16266 3576
rect 12128 3292 12436 3301
rect 12128 3290 12134 3292
rect 12190 3290 12214 3292
rect 12270 3290 12294 3292
rect 12350 3290 12374 3292
rect 12430 3290 12436 3292
rect 12190 3238 12192 3290
rect 12372 3238 12374 3290
rect 12128 3236 12134 3238
rect 12190 3236 12214 3238
rect 12270 3236 12294 3238
rect 12350 3236 12374 3238
rect 12430 3236 12436 3238
rect 12128 3227 12436 3236
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 10692 1352 10744 1358
rect 10692 1294 10744 1300
rect 11060 1352 11112 1358
rect 11060 1294 11112 1300
rect 10416 332 10468 338
rect 10416 274 10468 280
rect 10230 54 10364 82
rect 10598 82 10654 160
rect 10704 82 10732 1294
rect 10876 1216 10928 1222
rect 10876 1158 10928 1164
rect 10888 921 10916 1158
rect 10874 912 10930 921
rect 10874 847 10930 856
rect 10598 54 10732 82
rect 10966 82 11022 160
rect 11072 82 11100 1294
rect 11164 338 11192 3130
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11440 2774 11468 3062
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 11348 2746 11468 2774
rect 11244 1216 11296 1222
rect 11244 1158 11296 1164
rect 11152 332 11204 338
rect 11152 274 11204 280
rect 10966 54 11100 82
rect 11256 66 11284 1158
rect 11348 950 11376 2746
rect 13726 2544 13782 2553
rect 13726 2479 13782 2488
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12128 2204 12436 2213
rect 12128 2202 12134 2204
rect 12190 2202 12214 2204
rect 12270 2202 12294 2204
rect 12350 2202 12374 2204
rect 12430 2202 12436 2204
rect 12190 2150 12192 2202
rect 12372 2150 12374 2202
rect 12128 2148 12134 2150
rect 12190 2148 12214 2150
rect 12270 2148 12294 2150
rect 12350 2148 12374 2150
rect 12430 2148 12436 2150
rect 12128 2139 12436 2148
rect 11520 1352 11572 1358
rect 11520 1294 11572 1300
rect 11796 1352 11848 1358
rect 12164 1352 12216 1358
rect 11796 1294 11848 1300
rect 11992 1312 12164 1340
rect 11428 1284 11480 1290
rect 11428 1226 11480 1232
rect 11336 944 11388 950
rect 11336 886 11388 892
rect 11440 785 11468 1226
rect 11426 776 11482 785
rect 11426 711 11482 720
rect 11334 82 11390 160
rect 11532 82 11560 1294
rect 11244 60 11296 66
rect 9126 0 9182 54
rect 9494 0 9550 54
rect 9862 0 9918 54
rect 10230 0 10286 54
rect 10598 0 10654 54
rect 10966 0 11022 54
rect 11244 2 11296 8
rect 11334 54 11560 82
rect 11702 82 11758 160
rect 11808 82 11836 1294
rect 11888 1216 11940 1222
rect 11888 1158 11940 1164
rect 11900 377 11928 1158
rect 11886 368 11942 377
rect 11886 303 11942 312
rect 11702 54 11836 82
rect 11992 82 12020 1312
rect 12164 1294 12216 1300
rect 12532 1352 12584 1358
rect 12532 1294 12584 1300
rect 12128 1116 12436 1125
rect 12128 1114 12134 1116
rect 12190 1114 12214 1116
rect 12270 1114 12294 1116
rect 12350 1114 12374 1116
rect 12430 1114 12436 1116
rect 12190 1062 12192 1114
rect 12372 1062 12374 1114
rect 12128 1060 12134 1062
rect 12190 1060 12214 1062
rect 12270 1060 12294 1062
rect 12350 1060 12374 1062
rect 12430 1060 12436 1062
rect 12128 1051 12436 1060
rect 12070 82 12126 160
rect 11992 54 12126 82
rect 11334 0 11390 54
rect 11702 0 11758 54
rect 12070 0 12126 54
rect 12438 82 12494 160
rect 12544 82 12572 1294
rect 12636 814 12664 2246
rect 13740 2106 13768 2479
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 13728 2100 13780 2106
rect 13728 2042 13780 2048
rect 14292 1562 14320 2314
rect 14280 1556 14332 1562
rect 14280 1498 14332 1504
rect 12808 1352 12860 1358
rect 12808 1294 12860 1300
rect 12900 1352 12952 1358
rect 12900 1294 12952 1300
rect 13268 1352 13320 1358
rect 13268 1294 13320 1300
rect 13636 1352 13688 1358
rect 13636 1294 13688 1300
rect 14096 1352 14148 1358
rect 14096 1294 14148 1300
rect 14372 1352 14424 1358
rect 14372 1294 14424 1300
rect 12716 1216 12768 1222
rect 12716 1158 12768 1164
rect 12728 814 12756 1158
rect 12820 1018 12848 1294
rect 12808 1012 12860 1018
rect 12808 954 12860 960
rect 12624 808 12676 814
rect 12624 750 12676 756
rect 12716 808 12768 814
rect 12716 750 12768 756
rect 12438 54 12572 82
rect 12806 82 12862 160
rect 12912 82 12940 1294
rect 13084 400 13136 406
rect 13084 342 13136 348
rect 13096 241 13124 342
rect 13082 232 13138 241
rect 13082 167 13138 176
rect 12806 54 12940 82
rect 13174 82 13230 160
rect 13280 82 13308 1294
rect 13360 1216 13412 1222
rect 13360 1158 13412 1164
rect 13452 1216 13504 1222
rect 13452 1158 13504 1164
rect 13372 338 13400 1158
rect 13464 406 13492 1158
rect 13452 400 13504 406
rect 13452 342 13504 348
rect 13360 332 13412 338
rect 13360 274 13412 280
rect 13174 54 13308 82
rect 13542 82 13598 160
rect 13648 82 13676 1294
rect 13820 1216 13872 1222
rect 13726 1184 13782 1193
rect 13820 1158 13872 1164
rect 13726 1119 13782 1128
rect 13740 950 13768 1119
rect 13728 944 13780 950
rect 13728 886 13780 892
rect 13832 270 13860 1158
rect 13820 264 13872 270
rect 13820 206 13872 212
rect 13542 54 13676 82
rect 13910 82 13966 160
rect 14108 82 14136 1294
rect 13910 54 14136 82
rect 14278 82 14334 160
rect 14384 82 14412 1294
rect 14464 1216 14516 1222
rect 14464 1158 14516 1164
rect 14476 950 14504 1158
rect 14464 944 14516 950
rect 14464 886 14516 892
rect 14568 882 14596 2790
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 14648 1352 14700 1358
rect 14648 1294 14700 1300
rect 14556 876 14608 882
rect 14556 818 14608 824
rect 14660 160 14688 1294
rect 14752 610 14780 2382
rect 14924 1352 14976 1358
rect 14924 1294 14976 1300
rect 14740 604 14792 610
rect 14740 546 14792 552
rect 14278 54 14412 82
rect 12438 0 12494 54
rect 12806 0 12862 54
rect 13174 0 13230 54
rect 13542 0 13598 54
rect 13910 0 13966 54
rect 14278 0 14334 54
rect 14646 0 14702 160
rect 14936 82 14964 1294
rect 15028 542 15056 2450
rect 16224 2106 16252 3567
rect 16762 3496 16818 3505
rect 16762 3431 16818 3440
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 16500 2106 16528 2926
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 16488 2100 16540 2106
rect 16488 2042 16540 2048
rect 15108 1964 15160 1970
rect 15108 1906 15160 1912
rect 15476 1964 15528 1970
rect 15476 1906 15528 1912
rect 15752 1964 15804 1970
rect 15752 1906 15804 1912
rect 16028 1964 16080 1970
rect 16028 1906 16080 1912
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 15120 1562 15148 1906
rect 15488 1562 15516 1906
rect 15658 1864 15714 1873
rect 15658 1799 15714 1808
rect 15672 1766 15700 1799
rect 15660 1760 15712 1766
rect 15660 1702 15712 1708
rect 15764 1562 15792 1906
rect 16040 1562 16068 1906
rect 16316 1562 16344 1906
rect 16776 1902 16804 3431
rect 16868 1970 16896 4111
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17144 2122 17172 3470
rect 17236 2650 17264 8434
rect 17717 8188 18025 8197
rect 17717 8186 17723 8188
rect 17779 8186 17803 8188
rect 17859 8186 17883 8188
rect 17939 8186 17963 8188
rect 18019 8186 18025 8188
rect 17779 8134 17781 8186
rect 17961 8134 17963 8186
rect 17717 8132 17723 8134
rect 17779 8132 17803 8134
rect 17859 8132 17883 8134
rect 17939 8132 17963 8134
rect 18019 8132 18025 8134
rect 17717 8123 18025 8132
rect 17717 7100 18025 7109
rect 17717 7098 17723 7100
rect 17779 7098 17803 7100
rect 17859 7098 17883 7100
rect 17939 7098 17963 7100
rect 18019 7098 18025 7100
rect 17779 7046 17781 7098
rect 17961 7046 17963 7098
rect 17717 7044 17723 7046
rect 17779 7044 17803 7046
rect 17859 7044 17883 7046
rect 17939 7044 17963 7046
rect 18019 7044 18025 7046
rect 17717 7035 18025 7044
rect 17717 6012 18025 6021
rect 17717 6010 17723 6012
rect 17779 6010 17803 6012
rect 17859 6010 17883 6012
rect 17939 6010 17963 6012
rect 18019 6010 18025 6012
rect 17779 5958 17781 6010
rect 17961 5958 17963 6010
rect 17717 5956 17723 5958
rect 17779 5956 17803 5958
rect 17859 5956 17883 5958
rect 17939 5956 17963 5958
rect 18019 5956 18025 5958
rect 17717 5947 18025 5956
rect 17717 4924 18025 4933
rect 17717 4922 17723 4924
rect 17779 4922 17803 4924
rect 17859 4922 17883 4924
rect 17939 4922 17963 4924
rect 18019 4922 18025 4924
rect 17779 4870 17781 4922
rect 17961 4870 17963 4922
rect 17717 4868 17723 4870
rect 17779 4868 17803 4870
rect 17859 4868 17883 4870
rect 17939 4868 17963 4870
rect 18019 4868 18025 4870
rect 17717 4859 18025 4868
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 17717 3836 18025 3845
rect 17717 3834 17723 3836
rect 17779 3834 17803 3836
rect 17859 3834 17883 3836
rect 17939 3834 17963 3836
rect 18019 3834 18025 3836
rect 17779 3782 17781 3834
rect 17961 3782 17963 3834
rect 17717 3780 17723 3782
rect 17779 3780 17803 3782
rect 17859 3780 17883 3782
rect 17939 3780 17963 3782
rect 18019 3780 18025 3782
rect 17717 3771 18025 3780
rect 17314 3088 17370 3097
rect 17314 3023 17370 3032
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17144 2094 17264 2122
rect 16856 1964 16908 1970
rect 16856 1906 16908 1912
rect 17132 1964 17184 1970
rect 17132 1906 17184 1912
rect 16764 1896 16816 1902
rect 16764 1838 16816 1844
rect 16948 1896 17000 1902
rect 16948 1838 17000 1844
rect 15108 1556 15160 1562
rect 15108 1498 15160 1504
rect 15476 1556 15528 1562
rect 15476 1498 15528 1504
rect 15752 1556 15804 1562
rect 15752 1498 15804 1504
rect 16028 1556 16080 1562
rect 16028 1498 16080 1504
rect 16304 1556 16356 1562
rect 16304 1498 16356 1504
rect 16488 1556 16540 1562
rect 16488 1498 16540 1504
rect 15200 1352 15252 1358
rect 15200 1294 15252 1300
rect 15476 1352 15528 1358
rect 15476 1294 15528 1300
rect 16212 1352 16264 1358
rect 16212 1294 16264 1300
rect 15016 536 15068 542
rect 15016 478 15068 484
rect 15014 82 15070 160
rect 14936 54 15070 82
rect 15212 82 15240 1294
rect 15382 82 15438 160
rect 15212 54 15438 82
rect 15488 82 15516 1294
rect 16120 1284 16172 1290
rect 16120 1226 16172 1232
rect 15672 160 15792 184
rect 16132 160 16160 1226
rect 15672 156 15806 160
rect 15672 82 15700 156
rect 15488 54 15700 82
rect 15014 0 15070 54
rect 15382 0 15438 54
rect 15750 0 15806 156
rect 16118 0 16174 160
rect 16224 82 16252 1294
rect 16500 1290 16528 1498
rect 16960 1465 16988 1838
rect 17144 1562 17172 1906
rect 17132 1556 17184 1562
rect 17132 1498 17184 1504
rect 16946 1456 17002 1465
rect 16946 1391 17002 1400
rect 16580 1352 16632 1358
rect 16580 1294 16632 1300
rect 16764 1352 16816 1358
rect 16816 1312 16988 1340
rect 16764 1294 16816 1300
rect 16488 1284 16540 1290
rect 16488 1226 16540 1232
rect 16486 82 16542 160
rect 16224 54 16542 82
rect 16592 82 16620 1294
rect 16776 160 16896 184
rect 16776 156 16910 160
rect 16776 82 16804 156
rect 16592 54 16804 82
rect 16486 0 16542 54
rect 16854 0 16910 156
rect 16960 82 16988 1312
rect 17236 1222 17264 2094
rect 17328 2038 17356 3023
rect 17717 2748 18025 2757
rect 17717 2746 17723 2748
rect 17779 2746 17803 2748
rect 17859 2746 17883 2748
rect 17939 2746 17963 2748
rect 18019 2746 18025 2748
rect 17779 2694 17781 2746
rect 17961 2694 17963 2746
rect 17717 2692 17723 2694
rect 17779 2692 17803 2694
rect 17859 2692 17883 2694
rect 17939 2692 17963 2694
rect 18019 2692 18025 2694
rect 17717 2683 18025 2692
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 17592 2440 17644 2446
rect 18052 2440 18104 2446
rect 17592 2382 17644 2388
rect 17958 2408 18014 2417
rect 17512 2038 17540 2382
rect 17604 2106 17632 2382
rect 18052 2382 18104 2388
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 17958 2343 18014 2352
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17592 2100 17644 2106
rect 17592 2042 17644 2048
rect 17316 2032 17368 2038
rect 17316 1974 17368 1980
rect 17500 2032 17552 2038
rect 17500 1974 17552 1980
rect 17590 2000 17646 2009
rect 17408 1964 17460 1970
rect 17696 1970 17724 2246
rect 17590 1935 17646 1944
rect 17684 1964 17736 1970
rect 17408 1906 17460 1912
rect 17420 1562 17448 1906
rect 17500 1760 17552 1766
rect 17500 1702 17552 1708
rect 17408 1556 17460 1562
rect 17408 1498 17460 1504
rect 17224 1216 17276 1222
rect 17224 1158 17276 1164
rect 17222 1048 17278 1057
rect 17222 983 17278 992
rect 17236 649 17264 983
rect 17222 640 17278 649
rect 17512 610 17540 1702
rect 17604 1494 17632 1935
rect 17684 1906 17736 1912
rect 17972 1766 18000 2343
rect 17960 1760 18012 1766
rect 17960 1702 18012 1708
rect 17717 1660 18025 1669
rect 17717 1658 17723 1660
rect 17779 1658 17803 1660
rect 17859 1658 17883 1660
rect 17939 1658 17963 1660
rect 18019 1658 18025 1660
rect 17779 1606 17781 1658
rect 17961 1606 17963 1658
rect 17717 1604 17723 1606
rect 17779 1604 17803 1606
rect 17859 1604 17883 1606
rect 17939 1604 17963 1606
rect 18019 1604 18025 1606
rect 17717 1595 18025 1604
rect 18064 1562 18092 2382
rect 18144 1964 18196 1970
rect 18144 1906 18196 1912
rect 18512 1964 18564 1970
rect 18512 1906 18564 1912
rect 18156 1562 18184 1906
rect 18328 1896 18380 1902
rect 18328 1838 18380 1844
rect 18236 1828 18288 1834
rect 18236 1770 18288 1776
rect 18052 1556 18104 1562
rect 18052 1498 18104 1504
rect 18144 1556 18196 1562
rect 18144 1498 18196 1504
rect 18248 1494 18276 1770
rect 17592 1488 17644 1494
rect 17592 1430 17644 1436
rect 18236 1488 18288 1494
rect 18236 1430 18288 1436
rect 18340 1426 18368 1838
rect 18524 1562 18552 1906
rect 18604 1760 18656 1766
rect 18602 1728 18604 1737
rect 18656 1728 18658 1737
rect 18602 1663 18658 1672
rect 18512 1556 18564 1562
rect 18512 1498 18564 1504
rect 18328 1420 18380 1426
rect 18328 1362 18380 1368
rect 17684 1352 17736 1358
rect 17604 1312 17684 1340
rect 17222 575 17278 584
rect 17500 604 17552 610
rect 17500 546 17552 552
rect 17604 160 17632 1312
rect 17684 1294 17736 1300
rect 17776 1352 17828 1358
rect 18052 1352 18104 1358
rect 17828 1312 18000 1340
rect 17776 1294 17828 1300
rect 17972 160 18000 1312
rect 18052 1294 18104 1300
rect 18512 1352 18564 1358
rect 18512 1294 18564 1300
rect 17222 82 17278 160
rect 16960 54 17278 82
rect 17222 0 17278 54
rect 17590 0 17646 160
rect 17958 0 18014 160
rect 18064 82 18092 1294
rect 18326 82 18382 160
rect 18064 54 18382 82
rect 18524 82 18552 1294
rect 18708 1290 18736 2382
rect 18800 1970 18828 4218
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19062 2816 19118 2825
rect 19062 2751 19118 2760
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 18984 2106 19012 2382
rect 19076 2310 19104 2751
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 18972 2100 19024 2106
rect 18972 2042 19024 2048
rect 18788 1964 18840 1970
rect 18788 1906 18840 1912
rect 19064 1964 19116 1970
rect 19064 1906 19116 1912
rect 19076 1562 19104 1906
rect 19064 1556 19116 1562
rect 19064 1498 19116 1504
rect 19168 1358 19196 3334
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 19260 2310 19288 2790
rect 19628 2582 19656 8434
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19890 2952 19946 2961
rect 19890 2887 19946 2896
rect 19616 2576 19668 2582
rect 19616 2518 19668 2524
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19708 2440 19760 2446
rect 19904 2428 19932 2887
rect 19760 2400 19932 2428
rect 19708 2382 19760 2388
rect 19248 2304 19300 2310
rect 19628 2292 19656 2382
rect 19996 2378 20024 8366
rect 20536 2916 20588 2922
rect 20536 2858 20588 2864
rect 20444 2576 20496 2582
rect 20444 2518 20496 2524
rect 20076 2440 20128 2446
rect 20352 2440 20404 2446
rect 20128 2400 20352 2428
rect 20076 2382 20128 2388
rect 20352 2382 20404 2388
rect 19984 2372 20036 2378
rect 19984 2314 20036 2320
rect 19892 2304 19944 2310
rect 19628 2264 19748 2292
rect 19248 2246 19300 2252
rect 19614 2136 19670 2145
rect 19248 2100 19300 2106
rect 19614 2071 19616 2080
rect 19248 2042 19300 2048
rect 19668 2071 19670 2080
rect 19616 2042 19668 2048
rect 19260 1601 19288 2042
rect 19720 2038 19748 2264
rect 20168 2304 20220 2310
rect 19892 2246 19944 2252
rect 19996 2252 20168 2258
rect 19996 2246 20220 2252
rect 20260 2304 20312 2310
rect 20260 2246 20312 2252
rect 19708 2032 19760 2038
rect 19338 2000 19394 2009
rect 19708 1974 19760 1980
rect 19338 1935 19340 1944
rect 19392 1935 19394 1944
rect 19616 1964 19668 1970
rect 19340 1906 19392 1912
rect 19616 1906 19668 1912
rect 19340 1828 19392 1834
rect 19340 1770 19392 1776
rect 19246 1592 19302 1601
rect 19246 1527 19302 1536
rect 19352 1358 19380 1770
rect 19628 1562 19656 1906
rect 19616 1556 19668 1562
rect 19616 1498 19668 1504
rect 18788 1352 18840 1358
rect 18788 1294 18840 1300
rect 19156 1352 19208 1358
rect 19156 1294 19208 1300
rect 19340 1352 19392 1358
rect 19340 1294 19392 1300
rect 19432 1352 19484 1358
rect 19904 1340 19932 2246
rect 19996 2230 20208 2246
rect 19996 1952 20024 2230
rect 20272 2122 20300 2246
rect 20088 2106 20300 2122
rect 20076 2100 20300 2106
rect 20128 2094 20300 2100
rect 20076 2042 20128 2048
rect 20076 1964 20128 1970
rect 19996 1924 20076 1952
rect 20076 1906 20128 1912
rect 20260 1964 20312 1970
rect 20260 1906 20312 1912
rect 20272 1850 20300 1906
rect 20180 1822 20300 1850
rect 19984 1760 20036 1766
rect 19984 1702 20036 1708
rect 19996 1494 20024 1702
rect 19984 1488 20036 1494
rect 19984 1430 20036 1436
rect 19984 1352 20036 1358
rect 19904 1312 19984 1340
rect 19432 1294 19484 1300
rect 19984 1294 20036 1300
rect 18696 1284 18748 1290
rect 18696 1226 18748 1232
rect 18694 82 18750 160
rect 18524 54 18750 82
rect 18800 82 18828 1294
rect 18984 160 19104 184
rect 19444 160 19472 1294
rect 19708 1216 19760 1222
rect 19708 1158 19760 1164
rect 20076 1216 20128 1222
rect 20076 1158 20128 1164
rect 18984 156 19118 160
rect 18984 82 19012 156
rect 18800 54 19012 82
rect 18326 0 18382 54
rect 18694 0 18750 54
rect 19062 0 19118 156
rect 19430 0 19486 160
rect 19720 82 19748 1158
rect 20088 626 20116 1158
rect 20180 762 20208 1822
rect 20260 1760 20312 1766
rect 20260 1702 20312 1708
rect 20352 1760 20404 1766
rect 20352 1702 20404 1708
rect 20272 1329 20300 1702
rect 20364 1358 20392 1702
rect 20352 1352 20404 1358
rect 20258 1320 20314 1329
rect 20352 1294 20404 1300
rect 20456 1306 20484 2518
rect 20548 1902 20576 2858
rect 21652 2446 21680 8434
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 21640 2440 21692 2446
rect 21640 2382 21692 2388
rect 20628 2304 20680 2310
rect 20916 2281 20944 2382
rect 21088 2304 21140 2310
rect 20628 2246 20680 2252
rect 20902 2272 20958 2281
rect 20640 2106 20668 2246
rect 21088 2246 21140 2252
rect 20902 2207 20958 2216
rect 21100 2106 21128 2246
rect 21192 2145 21220 2382
rect 21178 2136 21234 2145
rect 20628 2100 20680 2106
rect 20628 2042 20680 2048
rect 21088 2100 21140 2106
rect 21178 2071 21234 2080
rect 21088 2042 21140 2048
rect 20626 2000 20682 2009
rect 20626 1935 20682 1944
rect 21732 1964 21784 1970
rect 20536 1896 20588 1902
rect 20536 1838 20588 1844
rect 20640 1766 20668 1935
rect 21732 1906 21784 1912
rect 20720 1828 20772 1834
rect 20720 1770 20772 1776
rect 20628 1760 20680 1766
rect 20628 1702 20680 1708
rect 20456 1278 20576 1306
rect 20732 1290 20760 1770
rect 21088 1760 21140 1766
rect 21088 1702 21140 1708
rect 21180 1760 21232 1766
rect 21180 1702 21232 1708
rect 20904 1488 20956 1494
rect 20904 1430 20956 1436
rect 20258 1255 20314 1264
rect 20444 1216 20496 1222
rect 20548 1193 20576 1278
rect 20720 1284 20772 1290
rect 20720 1226 20772 1232
rect 20444 1158 20496 1164
rect 20534 1184 20590 1193
rect 20180 734 20300 762
rect 20088 598 20208 626
rect 20180 160 20208 598
rect 20272 241 20300 734
rect 20258 232 20314 241
rect 20258 167 20314 176
rect 19798 82 19854 160
rect 19720 54 19854 82
rect 19798 0 19854 54
rect 20166 0 20222 160
rect 20456 82 20484 1158
rect 20534 1119 20590 1128
rect 20628 400 20680 406
rect 20628 342 20680 348
rect 20534 82 20590 160
rect 20640 134 20668 342
rect 20916 160 20944 1430
rect 21100 882 21128 1702
rect 21088 876 21140 882
rect 21088 818 21140 824
rect 20456 54 20590 82
rect 20628 128 20680 134
rect 20628 70 20680 76
rect 20534 0 20590 54
rect 20902 0 20958 160
rect 21192 82 21220 1702
rect 21548 1216 21600 1222
rect 21548 1158 21600 1164
rect 21270 82 21326 160
rect 21192 54 21326 82
rect 21560 82 21588 1158
rect 21744 474 21772 1906
rect 21836 1358 21864 3402
rect 22192 2576 22244 2582
rect 22192 2518 22244 2524
rect 22100 2304 22152 2310
rect 22100 2246 22152 2252
rect 22008 1964 22060 1970
rect 22008 1906 22060 1912
rect 21916 1556 21968 1562
rect 21916 1498 21968 1504
rect 21824 1352 21876 1358
rect 21824 1294 21876 1300
rect 21732 468 21784 474
rect 21732 410 21784 416
rect 21638 82 21694 160
rect 21560 54 21694 82
rect 21928 82 21956 1498
rect 22020 406 22048 1906
rect 22112 1358 22140 2246
rect 22100 1352 22152 1358
rect 22100 1294 22152 1300
rect 22204 1290 22232 2518
rect 22480 2446 22508 3538
rect 22756 2650 22784 8910
rect 23032 2650 23060 8978
rect 23306 8732 23614 8741
rect 23306 8730 23312 8732
rect 23368 8730 23392 8732
rect 23448 8730 23472 8732
rect 23528 8730 23552 8732
rect 23608 8730 23614 8732
rect 23368 8678 23370 8730
rect 23550 8678 23552 8730
rect 23306 8676 23312 8678
rect 23368 8676 23392 8678
rect 23448 8676 23472 8678
rect 23528 8676 23552 8678
rect 23608 8676 23614 8678
rect 23306 8667 23614 8676
rect 23676 8634 23704 9030
rect 23940 8900 23992 8906
rect 23940 8842 23992 8848
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23112 8560 23164 8566
rect 23112 8502 23164 8508
rect 23124 2650 23152 8502
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 23664 8356 23716 8362
rect 23664 8298 23716 8304
rect 23306 7644 23614 7653
rect 23306 7642 23312 7644
rect 23368 7642 23392 7644
rect 23448 7642 23472 7644
rect 23528 7642 23552 7644
rect 23608 7642 23614 7644
rect 23368 7590 23370 7642
rect 23550 7590 23552 7642
rect 23306 7588 23312 7590
rect 23368 7588 23392 7590
rect 23448 7588 23472 7590
rect 23528 7588 23552 7590
rect 23608 7588 23614 7590
rect 23306 7579 23614 7588
rect 23306 6556 23614 6565
rect 23306 6554 23312 6556
rect 23368 6554 23392 6556
rect 23448 6554 23472 6556
rect 23528 6554 23552 6556
rect 23608 6554 23614 6556
rect 23368 6502 23370 6554
rect 23550 6502 23552 6554
rect 23306 6500 23312 6502
rect 23368 6500 23392 6502
rect 23448 6500 23472 6502
rect 23528 6500 23552 6502
rect 23608 6500 23614 6502
rect 23306 6491 23614 6500
rect 23306 5468 23614 5477
rect 23306 5466 23312 5468
rect 23368 5466 23392 5468
rect 23448 5466 23472 5468
rect 23528 5466 23552 5468
rect 23608 5466 23614 5468
rect 23368 5414 23370 5466
rect 23550 5414 23552 5466
rect 23306 5412 23312 5414
rect 23368 5412 23392 5414
rect 23448 5412 23472 5414
rect 23528 5412 23552 5414
rect 23608 5412 23614 5414
rect 23306 5403 23614 5412
rect 23306 4380 23614 4389
rect 23306 4378 23312 4380
rect 23368 4378 23392 4380
rect 23448 4378 23472 4380
rect 23528 4378 23552 4380
rect 23608 4378 23614 4380
rect 23368 4326 23370 4378
rect 23550 4326 23552 4378
rect 23306 4324 23312 4326
rect 23368 4324 23392 4326
rect 23448 4324 23472 4326
rect 23528 4324 23552 4326
rect 23608 4324 23614 4326
rect 23306 4315 23614 4324
rect 23306 3292 23614 3301
rect 23306 3290 23312 3292
rect 23368 3290 23392 3292
rect 23448 3290 23472 3292
rect 23528 3290 23552 3292
rect 23608 3290 23614 3292
rect 23368 3238 23370 3290
rect 23550 3238 23552 3290
rect 23306 3236 23312 3238
rect 23368 3236 23392 3238
rect 23448 3236 23472 3238
rect 23528 3236 23552 3238
rect 23608 3236 23614 3238
rect 23306 3227 23614 3236
rect 23204 3052 23256 3058
rect 23204 2994 23256 3000
rect 22744 2644 22796 2650
rect 22744 2586 22796 2592
rect 23020 2644 23072 2650
rect 23020 2586 23072 2592
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 22652 2508 22704 2514
rect 22572 2468 22652 2496
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 22468 2440 22520 2446
rect 22468 2382 22520 2388
rect 22192 1284 22244 1290
rect 22192 1226 22244 1232
rect 22008 400 22060 406
rect 22008 342 22060 348
rect 22296 338 22324 2382
rect 22572 1850 22600 2468
rect 22652 2450 22704 2456
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 22744 2304 22796 2310
rect 22744 2246 22796 2252
rect 22480 1822 22600 1850
rect 22376 1760 22428 1766
rect 22376 1702 22428 1708
rect 22388 1562 22416 1702
rect 22376 1556 22428 1562
rect 22376 1498 22428 1504
rect 22480 1290 22508 1822
rect 22560 1760 22612 1766
rect 22560 1702 22612 1708
rect 22468 1284 22520 1290
rect 22468 1226 22520 1232
rect 22572 898 22600 1702
rect 22756 1290 22784 2246
rect 22940 2106 22968 2382
rect 23032 2106 23060 2382
rect 22928 2100 22980 2106
rect 22928 2042 22980 2048
rect 23020 2100 23072 2106
rect 23020 2042 23072 2048
rect 22836 1964 22888 1970
rect 22836 1906 22888 1912
rect 22928 1964 22980 1970
rect 23216 1952 23244 2994
rect 23676 2650 23704 8298
rect 23768 2650 23796 8434
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23306 2204 23614 2213
rect 23306 2202 23312 2204
rect 23368 2202 23392 2204
rect 23448 2202 23472 2204
rect 23528 2202 23552 2204
rect 23608 2202 23614 2204
rect 23368 2150 23370 2202
rect 23550 2150 23552 2202
rect 23306 2148 23312 2150
rect 23368 2148 23392 2150
rect 23448 2148 23472 2150
rect 23528 2148 23552 2150
rect 23608 2148 23614 2150
rect 23306 2139 23614 2148
rect 23768 2106 23796 2382
rect 23756 2100 23808 2106
rect 23756 2042 23808 2048
rect 23860 1970 23888 2994
rect 23952 2650 23980 8842
rect 25700 8634 25728 9840
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 25688 8628 25740 8634
rect 25688 8570 25740 8576
rect 26056 8492 26108 8498
rect 26056 8434 26108 8440
rect 25318 4040 25374 4049
rect 25318 3975 25374 3984
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 23940 2644 23992 2650
rect 23940 2586 23992 2592
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 23388 1964 23440 1970
rect 23216 1924 23388 1952
rect 22928 1906 22980 1912
rect 23388 1906 23440 1912
rect 23848 1964 23900 1970
rect 23848 1906 23900 1912
rect 22848 1465 22876 1906
rect 22834 1456 22890 1465
rect 22834 1391 22890 1400
rect 22744 1284 22796 1290
rect 22744 1226 22796 1232
rect 22388 870 22600 898
rect 22284 332 22336 338
rect 22284 274 22336 280
rect 22388 160 22416 870
rect 22940 542 22968 1906
rect 23480 1828 23532 1834
rect 23480 1770 23532 1776
rect 23296 1760 23348 1766
rect 23296 1702 23348 1708
rect 23308 1358 23336 1702
rect 23492 1426 23520 1770
rect 23572 1760 23624 1766
rect 23572 1702 23624 1708
rect 23848 1760 23900 1766
rect 23848 1702 23900 1708
rect 23584 1426 23612 1702
rect 23480 1420 23532 1426
rect 23480 1362 23532 1368
rect 23572 1420 23624 1426
rect 23572 1362 23624 1368
rect 23204 1352 23256 1358
rect 23204 1294 23256 1300
rect 23296 1352 23348 1358
rect 23296 1294 23348 1300
rect 23020 1216 23072 1222
rect 23020 1158 23072 1164
rect 23112 1216 23164 1222
rect 23112 1158 23164 1164
rect 22928 536 22980 542
rect 22928 478 22980 484
rect 22006 82 22062 160
rect 21928 54 22062 82
rect 21270 0 21326 54
rect 21638 0 21694 54
rect 22006 0 22062 54
rect 22374 0 22430 160
rect 22742 82 22798 160
rect 23032 82 23060 1158
rect 23124 160 23152 1158
rect 23216 882 23244 1294
rect 23756 1216 23808 1222
rect 23756 1158 23808 1164
rect 23306 1116 23614 1125
rect 23306 1114 23312 1116
rect 23368 1114 23392 1116
rect 23448 1114 23472 1116
rect 23528 1114 23552 1116
rect 23608 1114 23614 1116
rect 23368 1062 23370 1114
rect 23550 1062 23552 1114
rect 23306 1060 23312 1062
rect 23368 1060 23392 1062
rect 23448 1060 23472 1062
rect 23528 1060 23552 1062
rect 23608 1060 23614 1062
rect 23306 1051 23614 1060
rect 23204 876 23256 882
rect 23204 818 23256 824
rect 23492 190 23612 218
rect 23492 160 23520 190
rect 22742 54 23060 82
rect 22742 0 22798 54
rect 23110 0 23166 160
rect 23478 0 23534 160
rect 23584 82 23612 190
rect 23768 82 23796 1158
rect 23860 160 23888 1702
rect 23940 1556 23992 1562
rect 23940 1498 23992 1504
rect 23952 1290 23980 1498
rect 23940 1284 23992 1290
rect 23940 1226 23992 1232
rect 24044 270 24072 2586
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 24136 2281 24164 2450
rect 24122 2272 24178 2281
rect 24122 2207 24178 2216
rect 24504 1970 24532 3130
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24596 2106 24624 2382
rect 25044 2372 25096 2378
rect 25044 2314 25096 2320
rect 25056 2106 25084 2314
rect 25134 2136 25190 2145
rect 24584 2100 24636 2106
rect 24584 2042 24636 2048
rect 25044 2100 25096 2106
rect 25134 2071 25136 2080
rect 25044 2042 25096 2048
rect 25188 2071 25190 2080
rect 25136 2042 25188 2048
rect 25332 1970 25360 3975
rect 26068 2582 26096 8434
rect 26606 4584 26662 4593
rect 26148 4548 26200 4554
rect 26606 4519 26662 4528
rect 26148 4490 26200 4496
rect 26056 2576 26108 2582
rect 26056 2518 26108 2524
rect 25412 2100 25464 2106
rect 25412 2042 25464 2048
rect 24492 1964 24544 1970
rect 24492 1906 24544 1912
rect 25136 1964 25188 1970
rect 25136 1906 25188 1912
rect 25320 1964 25372 1970
rect 25320 1906 25372 1912
rect 24504 1414 25084 1442
rect 24032 264 24084 270
rect 24032 206 24084 212
rect 23584 54 23796 82
rect 23846 0 23902 160
rect 24214 82 24270 160
rect 24504 82 24532 1414
rect 24952 1352 25004 1358
rect 24952 1294 25004 1300
rect 24768 1216 24820 1222
rect 24768 1158 24820 1164
rect 24780 626 24808 1158
rect 24596 598 24808 626
rect 24596 160 24624 598
rect 24964 160 24992 1294
rect 25056 1222 25084 1414
rect 25044 1216 25096 1222
rect 25044 1158 25096 1164
rect 25148 542 25176 1906
rect 25320 1828 25372 1834
rect 25320 1770 25372 1776
rect 25136 536 25188 542
rect 25136 478 25188 484
rect 25332 160 25360 1770
rect 25424 814 25452 2042
rect 26160 1970 26188 4490
rect 26424 4208 26476 4214
rect 26424 4150 26476 4156
rect 26332 3120 26384 3126
rect 26332 3062 26384 3068
rect 26344 2446 26372 3062
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 26436 1970 26464 4150
rect 26620 2446 26648 4519
rect 26700 2848 26752 2854
rect 26700 2790 26752 2796
rect 26608 2440 26660 2446
rect 26608 2382 26660 2388
rect 26712 2038 26740 2790
rect 26884 2644 26936 2650
rect 26884 2586 26936 2592
rect 26896 2446 26924 2586
rect 26884 2440 26936 2446
rect 27436 2440 27488 2446
rect 26884 2382 26936 2388
rect 27356 2400 27436 2428
rect 26792 2304 26844 2310
rect 26792 2246 26844 2252
rect 27068 2304 27120 2310
rect 27120 2264 27200 2292
rect 27068 2246 27120 2252
rect 26804 2038 26832 2246
rect 26700 2032 26752 2038
rect 26700 1974 26752 1980
rect 26792 2032 26844 2038
rect 26792 1974 26844 1980
rect 26148 1964 26200 1970
rect 26148 1906 26200 1912
rect 26424 1964 26476 1970
rect 26424 1906 26476 1912
rect 26884 1828 26936 1834
rect 26884 1770 26936 1776
rect 25872 1760 25924 1766
rect 25872 1702 25924 1708
rect 26332 1760 26384 1766
rect 26332 1702 26384 1708
rect 26424 1760 26476 1766
rect 26424 1702 26476 1708
rect 25884 1358 25912 1702
rect 26240 1556 26292 1562
rect 25976 1516 26240 1544
rect 25872 1352 25924 1358
rect 25872 1294 25924 1300
rect 25686 1184 25742 1193
rect 25686 1119 25742 1128
rect 25412 808 25464 814
rect 25412 750 25464 756
rect 25504 672 25556 678
rect 25504 614 25556 620
rect 25516 338 25544 614
rect 25700 513 25728 1119
rect 25686 504 25742 513
rect 25686 439 25742 448
rect 25504 332 25556 338
rect 25504 274 25556 280
rect 24214 54 24532 82
rect 24214 0 24270 54
rect 24582 0 24638 160
rect 24950 0 25006 160
rect 25318 0 25374 160
rect 25686 82 25742 160
rect 25976 82 26004 1516
rect 26240 1498 26292 1504
rect 26148 1420 26200 1426
rect 26148 1362 26200 1368
rect 25686 54 26004 82
rect 26054 82 26110 160
rect 26160 82 26188 1362
rect 26344 1358 26372 1702
rect 26332 1352 26384 1358
rect 26332 1294 26384 1300
rect 26436 160 26464 1702
rect 26608 1556 26660 1562
rect 26608 1498 26660 1504
rect 26620 1426 26648 1498
rect 26608 1420 26660 1426
rect 26608 1362 26660 1368
rect 26896 202 26924 1770
rect 27172 1358 27200 2264
rect 27252 1760 27304 1766
rect 27252 1702 27304 1708
rect 27160 1352 27212 1358
rect 27160 1294 27212 1300
rect 27264 218 27292 1702
rect 26884 196 26936 202
rect 26054 54 26188 82
rect 25686 0 25742 54
rect 26054 0 26110 54
rect 26422 0 26478 160
rect 26790 82 26846 160
rect 26884 138 26936 144
rect 27080 190 27292 218
rect 27356 202 27384 2400
rect 27436 2382 27488 2388
rect 27540 1902 27568 8774
rect 27908 8634 27936 9840
rect 30116 8634 30144 9840
rect 32324 8634 32352 9840
rect 34532 9738 34560 9840
rect 34624 9738 34652 9846
rect 34532 9710 34652 9738
rect 34484 8732 34792 8741
rect 34484 8730 34490 8732
rect 34546 8730 34570 8732
rect 34626 8730 34650 8732
rect 34706 8730 34730 8732
rect 34786 8730 34792 8732
rect 34546 8678 34548 8730
rect 34728 8678 34730 8730
rect 34484 8676 34490 8678
rect 34546 8676 34570 8678
rect 34626 8676 34650 8678
rect 34706 8676 34730 8678
rect 34786 8676 34792 8678
rect 34484 8667 34792 8676
rect 34992 8634 35020 9846
rect 36726 9840 36782 10000
rect 38934 9840 38990 10000
rect 41142 9840 41198 10000
rect 43350 9840 43406 10000
rect 45558 9840 45614 10000
rect 36740 8634 36768 9840
rect 38948 8634 38976 9840
rect 41156 8634 41184 9840
rect 43364 8634 43392 9840
rect 45572 8634 45600 9840
rect 45662 8732 45970 8741
rect 45662 8730 45668 8732
rect 45724 8730 45748 8732
rect 45804 8730 45828 8732
rect 45884 8730 45908 8732
rect 45964 8730 45970 8732
rect 45724 8678 45726 8730
rect 45906 8678 45908 8730
rect 45662 8676 45668 8678
rect 45724 8676 45748 8678
rect 45804 8676 45828 8678
rect 45884 8676 45908 8678
rect 45964 8676 45970 8678
rect 45662 8667 45970 8676
rect 27896 8628 27948 8634
rect 27896 8570 27948 8576
rect 30104 8628 30156 8634
rect 30104 8570 30156 8576
rect 32312 8628 32364 8634
rect 32312 8570 32364 8576
rect 34980 8628 35032 8634
rect 34980 8570 35032 8576
rect 36728 8628 36780 8634
rect 36728 8570 36780 8576
rect 38936 8628 38988 8634
rect 38936 8570 38988 8576
rect 41144 8628 41196 8634
rect 41144 8570 41196 8576
rect 43352 8628 43404 8634
rect 43352 8570 43404 8576
rect 45560 8628 45612 8634
rect 45560 8570 45612 8576
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 35072 8492 35124 8498
rect 35072 8434 35124 8440
rect 37096 8492 37148 8498
rect 37096 8434 37148 8440
rect 39304 8492 39356 8498
rect 39304 8434 39356 8440
rect 41420 8492 41472 8498
rect 41420 8434 41472 8440
rect 43720 8492 43772 8498
rect 43720 8434 43772 8440
rect 45100 8492 45152 8498
rect 45100 8434 45152 8440
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 27724 2514 27752 2790
rect 28276 2650 28304 8434
rect 28895 8188 29203 8197
rect 28895 8186 28901 8188
rect 28957 8186 28981 8188
rect 29037 8186 29061 8188
rect 29117 8186 29141 8188
rect 29197 8186 29203 8188
rect 28957 8134 28959 8186
rect 29139 8134 29141 8186
rect 28895 8132 28901 8134
rect 28957 8132 28981 8134
rect 29037 8132 29061 8134
rect 29117 8132 29141 8134
rect 29197 8132 29203 8134
rect 28895 8123 29203 8132
rect 28895 7100 29203 7109
rect 28895 7098 28901 7100
rect 28957 7098 28981 7100
rect 29037 7098 29061 7100
rect 29117 7098 29141 7100
rect 29197 7098 29203 7100
rect 28957 7046 28959 7098
rect 29139 7046 29141 7098
rect 28895 7044 28901 7046
rect 28957 7044 28981 7046
rect 29037 7044 29061 7046
rect 29117 7044 29141 7046
rect 29197 7044 29203 7046
rect 28895 7035 29203 7044
rect 28895 6012 29203 6021
rect 28895 6010 28901 6012
rect 28957 6010 28981 6012
rect 29037 6010 29061 6012
rect 29117 6010 29141 6012
rect 29197 6010 29203 6012
rect 28957 5958 28959 6010
rect 29139 5958 29141 6010
rect 28895 5956 28901 5958
rect 28957 5956 28981 5958
rect 29037 5956 29061 5958
rect 29117 5956 29141 5958
rect 29197 5956 29203 5958
rect 28895 5947 29203 5956
rect 28895 4924 29203 4933
rect 28895 4922 28901 4924
rect 28957 4922 28981 4924
rect 29037 4922 29061 4924
rect 29117 4922 29141 4924
rect 29197 4922 29203 4924
rect 28957 4870 28959 4922
rect 29139 4870 29141 4922
rect 28895 4868 28901 4870
rect 28957 4868 28981 4870
rect 29037 4868 29061 4870
rect 29117 4868 29141 4870
rect 29197 4868 29203 4870
rect 28895 4859 29203 4868
rect 28895 3836 29203 3845
rect 28895 3834 28901 3836
rect 28957 3834 28981 3836
rect 29037 3834 29061 3836
rect 29117 3834 29141 3836
rect 29197 3834 29203 3836
rect 28957 3782 28959 3834
rect 29139 3782 29141 3834
rect 28895 3780 28901 3782
rect 28957 3780 28981 3782
rect 29037 3780 29061 3782
rect 29117 3780 29141 3782
rect 29197 3780 29203 3782
rect 28895 3771 29203 3780
rect 30012 2848 30064 2854
rect 30012 2790 30064 2796
rect 30104 2848 30156 2854
rect 30104 2790 30156 2796
rect 28895 2748 29203 2757
rect 28895 2746 28901 2748
rect 28957 2746 28981 2748
rect 29037 2746 29061 2748
rect 29117 2746 29141 2748
rect 29197 2746 29203 2748
rect 28957 2694 28959 2746
rect 29139 2694 29141 2746
rect 28895 2692 28901 2694
rect 28957 2692 28981 2694
rect 29037 2692 29061 2694
rect 29117 2692 29141 2694
rect 29197 2692 29203 2694
rect 28895 2683 29203 2692
rect 28264 2644 28316 2650
rect 28264 2586 28316 2592
rect 27712 2508 27764 2514
rect 27712 2450 27764 2456
rect 27620 2440 27672 2446
rect 27620 2382 27672 2388
rect 28448 2440 28500 2446
rect 28448 2382 28500 2388
rect 29828 2440 29880 2446
rect 29828 2382 29880 2388
rect 27528 1896 27580 1902
rect 27528 1838 27580 1844
rect 27632 1834 27660 2382
rect 27988 2304 28040 2310
rect 27988 2246 28040 2252
rect 28080 2304 28132 2310
rect 28080 2246 28132 2252
rect 27620 1828 27672 1834
rect 27620 1770 27672 1776
rect 27896 1828 27948 1834
rect 27896 1770 27948 1776
rect 27802 1592 27858 1601
rect 27620 1556 27672 1562
rect 27448 1516 27620 1544
rect 27344 196 27396 202
rect 27080 82 27108 190
rect 26790 54 27108 82
rect 27158 82 27214 160
rect 27344 138 27396 144
rect 27448 82 27476 1516
rect 27802 1527 27858 1536
rect 27620 1498 27672 1504
rect 27712 1488 27764 1494
rect 27540 1436 27712 1442
rect 27540 1430 27764 1436
rect 27540 1414 27752 1430
rect 27540 160 27568 1414
rect 27816 1018 27844 1527
rect 27804 1012 27856 1018
rect 27804 954 27856 960
rect 27908 160 27936 1770
rect 28000 1358 28028 2246
rect 28092 1970 28120 2246
rect 28460 2106 28488 2382
rect 28816 2372 28868 2378
rect 28816 2314 28868 2320
rect 28908 2372 28960 2378
rect 28908 2314 28960 2320
rect 28448 2100 28500 2106
rect 28448 2042 28500 2048
rect 28080 1964 28132 1970
rect 28080 1906 28132 1912
rect 28540 1964 28592 1970
rect 28540 1906 28592 1912
rect 28356 1896 28408 1902
rect 28356 1838 28408 1844
rect 28170 1728 28226 1737
rect 28170 1663 28226 1672
rect 28080 1420 28132 1426
rect 28080 1362 28132 1368
rect 27988 1352 28040 1358
rect 27988 1294 28040 1300
rect 28092 814 28120 1362
rect 28184 950 28212 1663
rect 28264 1420 28316 1426
rect 28264 1362 28316 1368
rect 28172 944 28224 950
rect 28172 886 28224 892
rect 28080 808 28132 814
rect 28080 750 28132 756
rect 28276 160 28304 1362
rect 28368 746 28396 1838
rect 28552 882 28580 1906
rect 28632 1556 28684 1562
rect 28632 1498 28684 1504
rect 28540 876 28592 882
rect 28540 818 28592 824
rect 28356 740 28408 746
rect 28356 682 28408 688
rect 28644 160 28672 1498
rect 28828 882 28856 2314
rect 28920 2281 28948 2314
rect 28906 2272 28962 2281
rect 28906 2207 28962 2216
rect 29644 1964 29696 1970
rect 29696 1924 29776 1952
rect 29644 1906 29696 1912
rect 29368 1828 29420 1834
rect 29368 1770 29420 1776
rect 29644 1828 29696 1834
rect 29644 1770 29696 1776
rect 29276 1760 29328 1766
rect 29276 1702 29328 1708
rect 28895 1660 29203 1669
rect 28895 1658 28901 1660
rect 28957 1658 28981 1660
rect 29037 1658 29061 1660
rect 29117 1658 29141 1660
rect 29197 1658 29203 1660
rect 28957 1606 28959 1658
rect 29139 1606 29141 1658
rect 28895 1604 28901 1606
rect 28957 1604 28981 1606
rect 29037 1604 29061 1606
rect 29117 1604 29141 1606
rect 29197 1604 29203 1606
rect 28895 1595 29203 1604
rect 29000 1488 29052 1494
rect 29000 1430 29052 1436
rect 28816 876 28868 882
rect 28816 818 28868 824
rect 29012 160 29040 1430
rect 29288 1290 29316 1702
rect 29380 1358 29408 1770
rect 29552 1760 29604 1766
rect 29552 1702 29604 1708
rect 29460 1420 29512 1426
rect 29460 1362 29512 1368
rect 29368 1352 29420 1358
rect 29368 1294 29420 1300
rect 29276 1284 29328 1290
rect 29276 1226 29328 1232
rect 29472 626 29500 1362
rect 29564 1358 29592 1702
rect 29552 1352 29604 1358
rect 29552 1294 29604 1300
rect 29656 678 29684 1770
rect 29380 598 29500 626
rect 29644 672 29696 678
rect 29644 614 29696 620
rect 29380 160 29408 598
rect 29748 513 29776 1924
rect 29840 785 29868 2382
rect 30024 1970 30052 2790
rect 30012 1964 30064 1970
rect 30012 1906 30064 1912
rect 30012 1216 30064 1222
rect 30012 1158 30064 1164
rect 29826 776 29882 785
rect 29826 711 29882 720
rect 29828 672 29880 678
rect 29828 614 29880 620
rect 29734 504 29790 513
rect 29734 439 29790 448
rect 29840 270 29868 614
rect 29828 264 29880 270
rect 29828 206 29880 212
rect 27158 54 27476 82
rect 26790 0 26846 54
rect 27158 0 27214 54
rect 27526 0 27582 160
rect 27894 0 27950 160
rect 28262 0 28318 160
rect 28630 0 28686 160
rect 28998 0 29054 160
rect 29366 0 29422 160
rect 29734 82 29790 160
rect 30024 82 30052 1158
rect 30116 160 30144 2790
rect 30288 2372 30340 2378
rect 30288 2314 30340 2320
rect 30196 1964 30248 1970
rect 30196 1906 30248 1912
rect 29734 54 30052 82
rect 29734 0 29790 54
rect 30102 0 30158 160
rect 30208 66 30236 1906
rect 30300 1766 30328 2314
rect 30392 2292 30420 8434
rect 32128 4480 32180 4486
rect 32128 4422 32180 4428
rect 31760 3460 31812 3466
rect 31760 3402 31812 3408
rect 31206 2952 31262 2961
rect 31206 2887 31262 2896
rect 30932 2508 30984 2514
rect 30984 2468 31064 2496
rect 30932 2450 30984 2456
rect 30748 2440 30800 2446
rect 30668 2400 30748 2428
rect 30472 2304 30524 2310
rect 30392 2264 30472 2292
rect 30472 2246 30524 2252
rect 30380 2100 30432 2106
rect 30380 2042 30432 2048
rect 30288 1760 30340 1766
rect 30288 1702 30340 1708
rect 30392 1358 30420 2042
rect 30472 1964 30524 1970
rect 30524 1924 30604 1952
rect 30472 1906 30524 1912
rect 30472 1828 30524 1834
rect 30472 1770 30524 1776
rect 30380 1352 30432 1358
rect 30380 1294 30432 1300
rect 30484 1290 30512 1770
rect 30472 1284 30524 1290
rect 30472 1226 30524 1232
rect 30576 921 30604 1924
rect 30562 912 30618 921
rect 30562 847 30618 856
rect 30668 406 30696 2400
rect 30748 2382 30800 2388
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 30852 1193 30880 2382
rect 30932 2304 30984 2310
rect 31036 2281 31064 2468
rect 30932 2246 30984 2252
rect 31022 2272 31078 2281
rect 30944 2106 30972 2246
rect 31022 2207 31078 2216
rect 30932 2100 30984 2106
rect 30932 2042 30984 2048
rect 31024 1488 31076 1494
rect 31024 1430 31076 1436
rect 30838 1184 30894 1193
rect 30838 1119 30894 1128
rect 30656 400 30708 406
rect 30656 342 30708 348
rect 31036 218 31064 1430
rect 31220 406 31248 2887
rect 31484 2644 31536 2650
rect 31484 2586 31536 2592
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 31390 2544 31446 2553
rect 31496 2514 31524 2586
rect 31390 2479 31446 2488
rect 31484 2508 31536 2514
rect 31404 2446 31432 2479
rect 31680 2496 31708 2586
rect 31772 2514 31800 3402
rect 31852 2848 31904 2854
rect 31852 2790 31904 2796
rect 31484 2450 31536 2456
rect 31588 2468 31708 2496
rect 31760 2508 31812 2514
rect 31392 2440 31444 2446
rect 31392 2382 31444 2388
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 31312 2106 31340 2246
rect 31588 2145 31616 2468
rect 31760 2450 31812 2456
rect 31760 2304 31812 2310
rect 31760 2246 31812 2252
rect 31574 2136 31630 2145
rect 31300 2100 31352 2106
rect 31574 2071 31630 2080
rect 31300 2042 31352 2048
rect 31300 1896 31352 1902
rect 31300 1838 31352 1844
rect 31208 400 31260 406
rect 31208 342 31260 348
rect 31312 218 31340 1838
rect 31668 1556 31720 1562
rect 30484 190 30604 218
rect 30484 160 30512 190
rect 30196 60 30248 66
rect 30196 2 30248 8
rect 30470 0 30526 160
rect 30576 82 30604 190
rect 30760 190 31064 218
rect 31128 190 31340 218
rect 31496 1516 31668 1544
rect 30760 82 30788 190
rect 30576 54 30788 82
rect 30838 82 30894 160
rect 31128 82 31156 190
rect 30838 54 31156 82
rect 31206 82 31262 160
rect 31496 82 31524 1516
rect 31668 1498 31720 1504
rect 31668 1420 31720 1426
rect 31668 1362 31720 1368
rect 31206 54 31524 82
rect 31574 82 31630 160
rect 31680 82 31708 1362
rect 31772 1358 31800 2246
rect 31864 1902 31892 2790
rect 31944 2576 31996 2582
rect 31944 2518 31996 2524
rect 31852 1896 31904 1902
rect 31852 1838 31904 1844
rect 31956 1358 31984 2518
rect 32036 2440 32088 2446
rect 32036 2382 32088 2388
rect 32048 2106 32076 2382
rect 32036 2100 32088 2106
rect 32036 2042 32088 2048
rect 32140 1970 32168 4422
rect 32588 2848 32640 2854
rect 32588 2790 32640 2796
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 32312 2440 32364 2446
rect 32364 2400 32444 2428
rect 32312 2382 32364 2388
rect 32128 1964 32180 1970
rect 32128 1906 32180 1912
rect 32232 1850 32260 2382
rect 32140 1822 32260 1850
rect 32416 1834 32444 2400
rect 32600 1970 32628 2790
rect 32692 2650 32720 8434
rect 34484 7644 34792 7653
rect 34484 7642 34490 7644
rect 34546 7642 34570 7644
rect 34626 7642 34650 7644
rect 34706 7642 34730 7644
rect 34786 7642 34792 7644
rect 34546 7590 34548 7642
rect 34728 7590 34730 7642
rect 34484 7588 34490 7590
rect 34546 7588 34570 7590
rect 34626 7588 34650 7590
rect 34706 7588 34730 7590
rect 34786 7588 34792 7590
rect 34484 7579 34792 7588
rect 34484 6556 34792 6565
rect 34484 6554 34490 6556
rect 34546 6554 34570 6556
rect 34626 6554 34650 6556
rect 34706 6554 34730 6556
rect 34786 6554 34792 6556
rect 34546 6502 34548 6554
rect 34728 6502 34730 6554
rect 34484 6500 34490 6502
rect 34546 6500 34570 6502
rect 34626 6500 34650 6502
rect 34706 6500 34730 6502
rect 34786 6500 34792 6502
rect 34484 6491 34792 6500
rect 34484 5468 34792 5477
rect 34484 5466 34490 5468
rect 34546 5466 34570 5468
rect 34626 5466 34650 5468
rect 34706 5466 34730 5468
rect 34786 5466 34792 5468
rect 34546 5414 34548 5466
rect 34728 5414 34730 5466
rect 34484 5412 34490 5414
rect 34546 5412 34570 5414
rect 34626 5412 34650 5414
rect 34706 5412 34730 5414
rect 34786 5412 34792 5414
rect 34484 5403 34792 5412
rect 34484 4380 34792 4389
rect 34484 4378 34490 4380
rect 34546 4378 34570 4380
rect 34626 4378 34650 4380
rect 34706 4378 34730 4380
rect 34786 4378 34792 4380
rect 34546 4326 34548 4378
rect 34728 4326 34730 4378
rect 34484 4324 34490 4326
rect 34546 4324 34570 4326
rect 34626 4324 34650 4326
rect 34706 4324 34730 4326
rect 34786 4324 34792 4326
rect 34484 4315 34792 4324
rect 34484 3292 34792 3301
rect 34484 3290 34490 3292
rect 34546 3290 34570 3292
rect 34626 3290 34650 3292
rect 34706 3290 34730 3292
rect 34786 3290 34792 3292
rect 34546 3238 34548 3290
rect 34728 3238 34730 3290
rect 34484 3236 34490 3238
rect 34546 3236 34570 3238
rect 34626 3236 34650 3238
rect 34706 3236 34730 3238
rect 34786 3236 34792 3238
rect 34484 3227 34792 3236
rect 34336 2916 34388 2922
rect 34336 2858 34388 2864
rect 32680 2644 32732 2650
rect 32680 2586 32732 2592
rect 34348 2582 34376 2858
rect 35084 2650 35112 8434
rect 37108 6914 37136 8434
rect 36924 6886 37136 6914
rect 39316 6914 39344 8434
rect 40073 8188 40381 8197
rect 40073 8186 40079 8188
rect 40135 8186 40159 8188
rect 40215 8186 40239 8188
rect 40295 8186 40319 8188
rect 40375 8186 40381 8188
rect 40135 8134 40137 8186
rect 40317 8134 40319 8186
rect 40073 8132 40079 8134
rect 40135 8132 40159 8134
rect 40215 8132 40239 8134
rect 40295 8132 40319 8134
rect 40375 8132 40381 8134
rect 40073 8123 40381 8132
rect 40073 7100 40381 7109
rect 40073 7098 40079 7100
rect 40135 7098 40159 7100
rect 40215 7098 40239 7100
rect 40295 7098 40319 7100
rect 40375 7098 40381 7100
rect 40135 7046 40137 7098
rect 40317 7046 40319 7098
rect 40073 7044 40079 7046
rect 40135 7044 40159 7046
rect 40215 7044 40239 7046
rect 40295 7044 40319 7046
rect 40375 7044 40381 7046
rect 40073 7035 40381 7044
rect 39316 6886 39528 6914
rect 36636 3528 36688 3534
rect 36636 3470 36688 3476
rect 35532 3052 35584 3058
rect 35532 2994 35584 3000
rect 35072 2644 35124 2650
rect 35072 2586 35124 2592
rect 33140 2576 33192 2582
rect 33140 2518 33192 2524
rect 34336 2576 34388 2582
rect 34336 2518 34388 2524
rect 32956 2304 33008 2310
rect 33008 2264 33088 2292
rect 32956 2246 33008 2252
rect 32588 1964 32640 1970
rect 32588 1906 32640 1912
rect 33060 1850 33088 2264
rect 33152 2038 33180 2518
rect 33232 2440 33284 2446
rect 34888 2440 34940 2446
rect 33232 2382 33284 2388
rect 34242 2408 34298 2417
rect 33244 2310 33272 2382
rect 34888 2382 34940 2388
rect 35348 2440 35400 2446
rect 35348 2382 35400 2388
rect 34242 2343 34298 2352
rect 33232 2304 33284 2310
rect 33232 2246 33284 2252
rect 34256 2038 34284 2343
rect 34334 2272 34390 2281
rect 34334 2207 34390 2216
rect 33140 2032 33192 2038
rect 33140 1974 33192 1980
rect 34244 2032 34296 2038
rect 34244 1974 34296 1980
rect 32312 1828 32364 1834
rect 31760 1352 31812 1358
rect 31760 1294 31812 1300
rect 31944 1352 31996 1358
rect 31944 1294 31996 1300
rect 32140 649 32168 1822
rect 32312 1770 32364 1776
rect 32404 1828 32456 1834
rect 32404 1770 32456 1776
rect 32588 1828 32640 1834
rect 33060 1822 33640 1850
rect 34348 1834 34376 2207
rect 34484 2204 34792 2213
rect 34484 2202 34490 2204
rect 34546 2202 34570 2204
rect 34626 2202 34650 2204
rect 34706 2202 34730 2204
rect 34786 2202 34792 2204
rect 34546 2150 34548 2202
rect 34728 2150 34730 2202
rect 34484 2148 34490 2150
rect 34546 2148 34570 2150
rect 34626 2148 34650 2150
rect 34706 2148 34730 2150
rect 34786 2148 34792 2150
rect 34484 2139 34792 2148
rect 34900 2106 34928 2382
rect 34888 2100 34940 2106
rect 34888 2042 34940 2048
rect 35360 1970 35388 2382
rect 35544 2106 35572 2994
rect 35716 2984 35768 2990
rect 35716 2926 35768 2932
rect 35532 2100 35584 2106
rect 35532 2042 35584 2048
rect 35728 2038 35756 2926
rect 35716 2032 35768 2038
rect 35716 1974 35768 1980
rect 35348 1964 35400 1970
rect 35348 1906 35400 1912
rect 32588 1770 32640 1776
rect 32324 1358 32352 1770
rect 32312 1352 32364 1358
rect 32312 1294 32364 1300
rect 32126 640 32182 649
rect 32126 575 32182 584
rect 32600 354 32628 1770
rect 33048 1760 33100 1766
rect 33048 1702 33100 1708
rect 33416 1760 33468 1766
rect 33416 1702 33468 1708
rect 33060 1408 33088 1702
rect 32968 1380 33088 1408
rect 32680 1216 32732 1222
rect 32680 1158 32732 1164
rect 32232 326 32628 354
rect 31574 54 31708 82
rect 31942 82 31998 160
rect 32232 82 32260 326
rect 32692 218 32720 1158
rect 32600 190 32720 218
rect 31942 54 32260 82
rect 32310 82 32366 160
rect 32600 82 32628 190
rect 32310 54 32628 82
rect 32678 82 32734 160
rect 32968 82 32996 1380
rect 33048 1284 33100 1290
rect 33048 1226 33100 1232
rect 33060 160 33088 1226
rect 33428 160 33456 1702
rect 33612 1358 33640 1822
rect 34336 1828 34388 1834
rect 34336 1770 34388 1776
rect 35716 1828 35768 1834
rect 35716 1770 35768 1776
rect 34888 1760 34940 1766
rect 34888 1702 34940 1708
rect 34336 1556 34388 1562
rect 34072 1516 34336 1544
rect 33600 1352 33652 1358
rect 33600 1294 33652 1300
rect 32678 54 32996 82
rect 30838 0 30894 54
rect 31206 0 31262 54
rect 31574 0 31630 54
rect 31942 0 31998 54
rect 32310 0 32366 54
rect 32678 0 32734 54
rect 33046 0 33102 160
rect 33414 0 33470 160
rect 33782 82 33838 160
rect 34072 82 34100 1516
rect 34336 1498 34388 1504
rect 34152 1284 34204 1290
rect 34152 1226 34204 1232
rect 34164 1018 34192 1226
rect 34244 1216 34296 1222
rect 34244 1158 34296 1164
rect 34152 1012 34204 1018
rect 34152 954 34204 960
rect 34256 626 34284 1158
rect 34484 1116 34792 1125
rect 34484 1114 34490 1116
rect 34546 1114 34570 1116
rect 34626 1114 34650 1116
rect 34706 1114 34730 1116
rect 34786 1114 34792 1116
rect 34546 1062 34548 1114
rect 34728 1062 34730 1114
rect 34484 1060 34490 1062
rect 34546 1060 34570 1062
rect 34626 1060 34650 1062
rect 34706 1060 34730 1062
rect 34786 1060 34792 1062
rect 34484 1051 34792 1060
rect 34900 762 34928 1702
rect 35728 1544 35756 1770
rect 36268 1760 36320 1766
rect 36268 1702 36320 1708
rect 35544 1516 35756 1544
rect 34980 1488 35032 1494
rect 34980 1430 35032 1436
rect 34164 598 34284 626
rect 34808 734 34928 762
rect 34164 160 34192 598
rect 33782 54 34100 82
rect 33782 0 33838 54
rect 34150 0 34206 160
rect 34518 82 34574 160
rect 34808 82 34836 734
rect 34992 626 35020 1430
rect 35348 1284 35400 1290
rect 35348 1226 35400 1232
rect 35360 1018 35388 1226
rect 35348 1012 35400 1018
rect 35348 954 35400 960
rect 34900 598 35020 626
rect 34900 160 34928 598
rect 34518 54 34836 82
rect 34518 0 34574 54
rect 34886 0 34942 160
rect 35254 82 35310 160
rect 35544 82 35572 1516
rect 35716 1420 35768 1426
rect 35636 1380 35716 1408
rect 35636 160 35664 1380
rect 35716 1362 35768 1368
rect 35900 1284 35952 1290
rect 35900 1226 35952 1232
rect 35912 406 35940 1226
rect 35900 400 35952 406
rect 35900 342 35952 348
rect 35254 54 35572 82
rect 35254 0 35310 54
rect 35622 0 35678 160
rect 35990 82 36046 160
rect 36280 82 36308 1702
rect 36648 1358 36676 3470
rect 36924 2650 36952 6886
rect 39394 4176 39450 4185
rect 39394 4111 39450 4120
rect 37554 3632 37610 3641
rect 37610 3590 37780 3618
rect 37554 3567 37610 3576
rect 37464 2848 37516 2854
rect 37464 2790 37516 2796
rect 36912 2644 36964 2650
rect 36912 2586 36964 2592
rect 37188 2644 37240 2650
rect 37188 2586 37240 2592
rect 37200 2446 37228 2586
rect 37476 2446 37504 2790
rect 37556 2644 37608 2650
rect 37556 2586 37608 2592
rect 37188 2440 37240 2446
rect 37188 2382 37240 2388
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 37568 2378 37596 2586
rect 37556 2372 37608 2378
rect 37556 2314 37608 2320
rect 37188 2304 37240 2310
rect 37188 2246 37240 2252
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 37200 2088 37228 2246
rect 37384 2106 37412 2246
rect 37280 2100 37332 2106
rect 37200 2060 37280 2088
rect 37280 2042 37332 2048
rect 37372 2100 37424 2106
rect 37372 2042 37424 2048
rect 37096 1896 37148 1902
rect 37148 1844 37412 1850
rect 37096 1838 37412 1844
rect 37108 1822 37412 1838
rect 37280 1760 37332 1766
rect 37280 1702 37332 1708
rect 36912 1556 36964 1562
rect 36740 1516 36912 1544
rect 36636 1352 36688 1358
rect 36542 1320 36598 1329
rect 36452 1284 36504 1290
rect 36636 1294 36688 1300
rect 36542 1255 36544 1264
rect 36452 1226 36504 1232
rect 36596 1255 36598 1264
rect 36544 1226 36596 1232
rect 36464 610 36492 1226
rect 36452 604 36504 610
rect 36452 546 36504 552
rect 36740 218 36768 1516
rect 36912 1498 36964 1504
rect 37016 1550 37136 1578
rect 36648 190 36768 218
rect 35990 54 36308 82
rect 36358 82 36414 160
rect 36648 82 36676 190
rect 36358 54 36676 82
rect 36726 82 36782 160
rect 37016 82 37044 1550
rect 37108 1494 37136 1550
rect 37096 1488 37148 1494
rect 37096 1430 37148 1436
rect 37292 1408 37320 1702
rect 37200 1380 37320 1408
rect 36726 54 37044 82
rect 37094 82 37150 160
rect 37200 82 37228 1380
rect 37384 1222 37412 1822
rect 37752 1358 37780 3590
rect 38934 3496 38990 3505
rect 38990 3454 39068 3482
rect 38934 3431 38990 3440
rect 38660 3392 38712 3398
rect 38660 3334 38712 3340
rect 38106 3088 38162 3097
rect 38162 3046 38240 3074
rect 38106 3023 38162 3032
rect 37832 2304 37884 2310
rect 37832 2246 37884 2252
rect 37844 1970 37872 2246
rect 37832 1964 37884 1970
rect 37832 1906 37884 1912
rect 38108 1964 38160 1970
rect 38108 1906 38160 1912
rect 38120 1873 38148 1906
rect 38106 1864 38162 1873
rect 38106 1799 38162 1808
rect 38108 1556 38160 1562
rect 37936 1516 38108 1544
rect 37740 1352 37792 1358
rect 37740 1294 37792 1300
rect 37372 1216 37424 1222
rect 37372 1158 37424 1164
rect 37936 354 37964 1516
rect 38108 1498 38160 1504
rect 38212 1358 38240 3046
rect 38568 2100 38620 2106
rect 38304 2060 38568 2088
rect 38200 1352 38252 1358
rect 38200 1294 38252 1300
rect 37752 326 37964 354
rect 37094 54 37228 82
rect 37462 82 37518 160
rect 37752 82 37780 326
rect 38304 218 38332 2060
rect 38568 2042 38620 2048
rect 38672 2038 38700 3334
rect 38844 2440 38896 2446
rect 38844 2382 38896 2388
rect 38660 2032 38712 2038
rect 38660 1974 38712 1980
rect 38750 2000 38806 2009
rect 38750 1935 38752 1944
rect 38804 1935 38806 1944
rect 38752 1906 38804 1912
rect 38476 1760 38528 1766
rect 38476 1702 38528 1708
rect 38384 1420 38436 1426
rect 38384 1362 38436 1368
rect 37844 190 37964 218
rect 37844 160 37872 190
rect 37462 54 37780 82
rect 35990 0 36046 54
rect 36358 0 36414 54
rect 36726 0 36782 54
rect 37094 0 37150 54
rect 37462 0 37518 54
rect 37830 0 37886 160
rect 37936 82 37964 190
rect 38120 190 38332 218
rect 38120 82 38148 190
rect 37936 54 38148 82
rect 38198 82 38254 160
rect 38396 82 38424 1362
rect 38198 54 38424 82
rect 38488 82 38516 1702
rect 38856 814 38884 2382
rect 38936 1760 38988 1766
rect 38936 1702 38988 1708
rect 38948 1465 38976 1702
rect 38934 1456 38990 1465
rect 38934 1391 38990 1400
rect 39040 1358 39068 3454
rect 39028 1352 39080 1358
rect 39304 1352 39356 1358
rect 39028 1294 39080 1300
rect 39224 1312 39304 1340
rect 38752 808 38804 814
rect 38752 750 38804 756
rect 38844 808 38896 814
rect 38844 750 38896 756
rect 38764 610 38792 750
rect 38752 604 38804 610
rect 38752 546 38804 552
rect 38566 82 38622 160
rect 38488 54 38622 82
rect 38198 0 38254 54
rect 38566 0 38622 54
rect 38934 82 38990 160
rect 39224 82 39252 1312
rect 39304 1294 39356 1300
rect 39408 1018 39436 4111
rect 39500 2650 39528 6886
rect 40073 6012 40381 6021
rect 40073 6010 40079 6012
rect 40135 6010 40159 6012
rect 40215 6010 40239 6012
rect 40295 6010 40319 6012
rect 40375 6010 40381 6012
rect 40135 5958 40137 6010
rect 40317 5958 40319 6010
rect 40073 5956 40079 5958
rect 40135 5956 40159 5958
rect 40215 5956 40239 5958
rect 40295 5956 40319 5958
rect 40375 5956 40381 5958
rect 40073 5947 40381 5956
rect 40073 4924 40381 4933
rect 40073 4922 40079 4924
rect 40135 4922 40159 4924
rect 40215 4922 40239 4924
rect 40295 4922 40319 4924
rect 40375 4922 40381 4924
rect 40135 4870 40137 4922
rect 40317 4870 40319 4922
rect 40073 4868 40079 4870
rect 40135 4868 40159 4870
rect 40215 4868 40239 4870
rect 40295 4868 40319 4870
rect 40375 4868 40381 4870
rect 40073 4859 40381 4868
rect 40073 3836 40381 3845
rect 40073 3834 40079 3836
rect 40135 3834 40159 3836
rect 40215 3834 40239 3836
rect 40295 3834 40319 3836
rect 40375 3834 40381 3836
rect 40135 3782 40137 3834
rect 40317 3782 40319 3834
rect 40073 3780 40079 3782
rect 40135 3780 40159 3782
rect 40215 3780 40239 3782
rect 40295 3780 40319 3782
rect 40375 3780 40381 3782
rect 40073 3771 40381 3780
rect 40073 2748 40381 2757
rect 40073 2746 40079 2748
rect 40135 2746 40159 2748
rect 40215 2746 40239 2748
rect 40295 2746 40319 2748
rect 40375 2746 40381 2748
rect 40135 2694 40137 2746
rect 40317 2694 40319 2746
rect 40073 2692 40079 2694
rect 40135 2692 40159 2694
rect 40215 2692 40239 2694
rect 40295 2692 40319 2694
rect 40375 2692 40381 2694
rect 40073 2683 40381 2692
rect 41432 2650 41460 8434
rect 41604 4276 41656 4282
rect 41604 4218 41656 4224
rect 39488 2644 39540 2650
rect 39488 2586 39540 2592
rect 41420 2644 41472 2650
rect 41420 2586 41472 2592
rect 39580 2576 39632 2582
rect 39632 2524 39804 2530
rect 39580 2518 39804 2524
rect 39592 2502 39804 2518
rect 39776 2446 39804 2502
rect 39672 2440 39724 2446
rect 39672 2382 39724 2388
rect 39764 2440 39816 2446
rect 39764 2382 39816 2388
rect 41512 2440 41564 2446
rect 41512 2382 41564 2388
rect 39684 2106 39712 2382
rect 41420 2372 41472 2378
rect 41420 2314 41472 2320
rect 39672 2100 39724 2106
rect 39672 2042 39724 2048
rect 40592 1964 40644 1970
rect 40420 1924 40592 1952
rect 40073 1660 40381 1669
rect 40073 1658 40079 1660
rect 40135 1658 40159 1660
rect 40215 1658 40239 1660
rect 40295 1658 40319 1660
rect 40375 1658 40381 1660
rect 40135 1606 40137 1658
rect 40317 1606 40319 1658
rect 40073 1604 40079 1606
rect 40135 1604 40159 1606
rect 40215 1604 40239 1606
rect 40295 1604 40319 1606
rect 40375 1604 40381 1606
rect 40073 1595 40381 1604
rect 39488 1488 39540 1494
rect 39488 1430 39540 1436
rect 39396 1012 39448 1018
rect 39396 954 39448 960
rect 39500 746 39528 1430
rect 40040 1352 40092 1358
rect 39592 1312 40040 1340
rect 39488 740 39540 746
rect 39488 682 39540 688
rect 38934 54 39252 82
rect 39302 82 39358 160
rect 39592 82 39620 1312
rect 40040 1294 40092 1300
rect 40224 1284 40276 1290
rect 40224 1226 40276 1232
rect 40236 218 40264 1226
rect 40420 218 40448 1924
rect 40592 1906 40644 1912
rect 40684 1964 40736 1970
rect 40684 1906 40736 1912
rect 40500 1216 40552 1222
rect 40500 1158 40552 1164
rect 40512 474 40540 1158
rect 40500 468 40552 474
rect 40500 410 40552 416
rect 39684 190 39804 218
rect 39684 160 39712 190
rect 39302 54 39620 82
rect 38934 0 38990 54
rect 39302 0 39358 54
rect 39670 0 39726 160
rect 39776 82 39804 190
rect 39960 190 40264 218
rect 40328 190 40448 218
rect 39960 82 39988 190
rect 39776 54 39988 82
rect 40038 82 40094 160
rect 40328 82 40356 190
rect 40038 54 40356 82
rect 40406 82 40462 160
rect 40696 82 40724 1906
rect 40776 1896 40828 1902
rect 40776 1838 40828 1844
rect 40788 160 40816 1838
rect 41432 1562 41460 2314
rect 41524 1562 41552 2382
rect 41616 1970 41644 4218
rect 43732 2650 43760 8434
rect 45112 2650 45140 8434
rect 45662 7644 45970 7653
rect 45662 7642 45668 7644
rect 45724 7642 45748 7644
rect 45804 7642 45828 7644
rect 45884 7642 45908 7644
rect 45964 7642 45970 7644
rect 45724 7590 45726 7642
rect 45906 7590 45908 7642
rect 45662 7588 45668 7590
rect 45724 7588 45748 7590
rect 45804 7588 45828 7590
rect 45884 7588 45908 7590
rect 45964 7588 45970 7590
rect 45662 7579 45970 7588
rect 45662 6556 45970 6565
rect 45662 6554 45668 6556
rect 45724 6554 45748 6556
rect 45804 6554 45828 6556
rect 45884 6554 45908 6556
rect 45964 6554 45970 6556
rect 45724 6502 45726 6554
rect 45906 6502 45908 6554
rect 45662 6500 45668 6502
rect 45724 6500 45748 6502
rect 45804 6500 45828 6502
rect 45884 6500 45908 6502
rect 45964 6500 45970 6502
rect 45662 6491 45970 6500
rect 45662 5468 45970 5477
rect 45662 5466 45668 5468
rect 45724 5466 45748 5468
rect 45804 5466 45828 5468
rect 45884 5466 45908 5468
rect 45964 5466 45970 5468
rect 45724 5414 45726 5466
rect 45906 5414 45908 5466
rect 45662 5412 45668 5414
rect 45724 5412 45748 5414
rect 45804 5412 45828 5414
rect 45884 5412 45908 5414
rect 45964 5412 45970 5414
rect 45662 5403 45970 5412
rect 45662 4380 45970 4389
rect 45662 4378 45668 4380
rect 45724 4378 45748 4380
rect 45804 4378 45828 4380
rect 45884 4378 45908 4380
rect 45964 4378 45970 4380
rect 45724 4326 45726 4378
rect 45906 4326 45908 4378
rect 45662 4324 45668 4326
rect 45724 4324 45748 4326
rect 45804 4324 45828 4326
rect 45884 4324 45908 4326
rect 45964 4324 45970 4326
rect 45662 4315 45970 4324
rect 45662 3292 45970 3301
rect 45662 3290 45668 3292
rect 45724 3290 45748 3292
rect 45804 3290 45828 3292
rect 45884 3290 45908 3292
rect 45964 3290 45970 3292
rect 45724 3238 45726 3290
rect 45906 3238 45908 3290
rect 45662 3236 45668 3238
rect 45724 3236 45748 3238
rect 45804 3236 45828 3238
rect 45884 3236 45908 3238
rect 45964 3236 45970 3238
rect 45662 3227 45970 3236
rect 43720 2644 43772 2650
rect 43720 2586 43772 2592
rect 45100 2644 45152 2650
rect 45100 2586 45152 2592
rect 44456 2508 44508 2514
rect 44456 2450 44508 2456
rect 41788 2440 41840 2446
rect 41788 2382 41840 2388
rect 44180 2440 44232 2446
rect 44180 2382 44232 2388
rect 41800 2106 41828 2382
rect 44192 2106 44220 2382
rect 44272 2304 44324 2310
rect 44272 2246 44324 2252
rect 41788 2100 41840 2106
rect 41788 2042 41840 2048
rect 44180 2100 44232 2106
rect 44180 2042 44232 2048
rect 41604 1964 41656 1970
rect 41604 1906 41656 1912
rect 44180 1896 44232 1902
rect 44180 1838 44232 1844
rect 41880 1828 41932 1834
rect 41880 1770 41932 1776
rect 41420 1556 41472 1562
rect 41420 1498 41472 1504
rect 41512 1556 41564 1562
rect 41512 1498 41564 1504
rect 41156 1414 41460 1442
rect 40868 1216 40920 1222
rect 40868 1158 40920 1164
rect 40880 610 40908 1158
rect 40868 604 40920 610
rect 40868 546 40920 552
rect 41156 160 41184 1414
rect 41432 1358 41460 1414
rect 41236 1352 41288 1358
rect 41236 1294 41288 1300
rect 41420 1352 41472 1358
rect 41420 1294 41472 1300
rect 41248 1018 41276 1294
rect 41328 1284 41380 1290
rect 41328 1226 41380 1232
rect 41236 1012 41288 1018
rect 41236 954 41288 960
rect 40406 54 40724 82
rect 40038 0 40094 54
rect 40406 0 40462 54
rect 40774 0 40830 160
rect 41142 0 41198 160
rect 41340 82 41368 1226
rect 41892 160 41920 1770
rect 44192 1562 44220 1838
rect 44180 1556 44232 1562
rect 44180 1498 44232 1504
rect 44284 1494 44312 2246
rect 44272 1488 44324 1494
rect 44272 1430 44324 1436
rect 42248 1352 42300 1358
rect 42708 1352 42760 1358
rect 42248 1294 42300 1300
rect 42628 1312 42708 1340
rect 41972 1216 42024 1222
rect 41972 1158 42024 1164
rect 41984 746 42012 1158
rect 41972 740 42024 746
rect 41972 682 42024 688
rect 42260 160 42288 1294
rect 42432 1216 42484 1222
rect 42432 1158 42484 1164
rect 42444 882 42472 1158
rect 42432 876 42484 882
rect 42432 818 42484 824
rect 42628 160 42656 1312
rect 42708 1294 42760 1300
rect 43260 1352 43312 1358
rect 43260 1294 43312 1300
rect 43628 1352 43680 1358
rect 43628 1294 43680 1300
rect 43996 1352 44048 1358
rect 43996 1294 44048 1300
rect 44088 1352 44140 1358
rect 44088 1294 44140 1300
rect 42708 1216 42760 1222
rect 42708 1158 42760 1164
rect 43076 1216 43128 1222
rect 43076 1158 43128 1164
rect 42720 882 42748 1158
rect 43088 1018 43116 1158
rect 43076 1012 43128 1018
rect 43076 954 43128 960
rect 42708 876 42760 882
rect 42708 818 42760 824
rect 41510 82 41566 160
rect 41340 54 41566 82
rect 41510 0 41566 54
rect 41878 0 41934 160
rect 42246 0 42302 160
rect 42614 0 42670 160
rect 42982 82 43038 160
rect 43272 82 43300 1294
rect 42982 54 43300 82
rect 43350 82 43406 160
rect 43640 82 43668 1294
rect 43350 54 43668 82
rect 43718 82 43774 160
rect 44008 82 44036 1294
rect 44100 160 44128 1294
rect 44468 1290 44496 2450
rect 44916 2440 44968 2446
rect 44916 2382 44968 2388
rect 45192 2440 45244 2446
rect 45928 2440 45980 2446
rect 45244 2400 45416 2428
rect 45192 2382 45244 2388
rect 44928 2106 44956 2382
rect 45008 2304 45060 2310
rect 45008 2246 45060 2252
rect 45284 2304 45336 2310
rect 45284 2246 45336 2252
rect 45020 2106 45048 2246
rect 45296 2106 45324 2246
rect 44916 2100 44968 2106
rect 44916 2042 44968 2048
rect 45008 2100 45060 2106
rect 45008 2042 45060 2048
rect 45284 2100 45336 2106
rect 45284 2042 45336 2048
rect 44732 1352 44784 1358
rect 44732 1294 44784 1300
rect 44824 1352 44876 1358
rect 45284 1352 45336 1358
rect 44824 1294 44876 1300
rect 45204 1312 45284 1340
rect 44456 1284 44508 1290
rect 44456 1226 44508 1232
rect 43718 54 44036 82
rect 42982 0 43038 54
rect 43350 0 43406 54
rect 43718 0 43774 54
rect 44086 0 44142 160
rect 44454 82 44510 160
rect 44744 82 44772 1294
rect 44836 160 44864 1294
rect 45204 160 45232 1312
rect 45284 1294 45336 1300
rect 44454 54 44772 82
rect 44454 0 44510 54
rect 44822 0 44878 160
rect 45190 0 45246 160
rect 45388 82 45416 2400
rect 45980 2400 46060 2428
rect 45928 2382 45980 2388
rect 45662 2204 45970 2213
rect 45662 2202 45668 2204
rect 45724 2202 45748 2204
rect 45804 2202 45828 2204
rect 45884 2202 45908 2204
rect 45964 2202 45970 2204
rect 45724 2150 45726 2202
rect 45906 2150 45908 2202
rect 45662 2148 45668 2150
rect 45724 2148 45748 2150
rect 45804 2148 45828 2150
rect 45884 2148 45908 2150
rect 45964 2148 45970 2150
rect 45662 2139 45970 2148
rect 45468 1964 45520 1970
rect 45468 1906 45520 1912
rect 45480 1442 45508 1906
rect 45480 1414 45600 1442
rect 45572 490 45600 1414
rect 45662 1116 45970 1125
rect 45662 1114 45668 1116
rect 45724 1114 45748 1116
rect 45804 1114 45828 1116
rect 45884 1114 45908 1116
rect 45964 1114 45970 1116
rect 45724 1062 45726 1114
rect 45906 1062 45908 1114
rect 45662 1060 45668 1062
rect 45724 1060 45748 1062
rect 45804 1060 45828 1062
rect 45884 1060 45908 1062
rect 45964 1060 45970 1062
rect 45662 1051 45970 1060
rect 45572 462 45692 490
rect 45558 82 45614 160
rect 45388 54 45614 82
rect 45664 82 45692 462
rect 45926 82 45982 160
rect 45664 54 45982 82
rect 46032 82 46060 2400
rect 46294 82 46350 160
rect 46032 54 46350 82
rect 45558 0 45614 54
rect 45926 0 45982 54
rect 46294 0 46350 54
<< via2 >>
rect 12134 8730 12190 8732
rect 12214 8730 12270 8732
rect 12294 8730 12350 8732
rect 12374 8730 12430 8732
rect 12134 8678 12180 8730
rect 12180 8678 12190 8730
rect 12214 8678 12244 8730
rect 12244 8678 12256 8730
rect 12256 8678 12270 8730
rect 12294 8678 12308 8730
rect 12308 8678 12320 8730
rect 12320 8678 12350 8730
rect 12374 8678 12384 8730
rect 12384 8678 12430 8730
rect 12134 8676 12190 8678
rect 12214 8676 12270 8678
rect 12294 8676 12350 8678
rect 12374 8676 12430 8678
rect 6545 8186 6601 8188
rect 6625 8186 6681 8188
rect 6705 8186 6761 8188
rect 6785 8186 6841 8188
rect 6545 8134 6591 8186
rect 6591 8134 6601 8186
rect 6625 8134 6655 8186
rect 6655 8134 6667 8186
rect 6667 8134 6681 8186
rect 6705 8134 6719 8186
rect 6719 8134 6731 8186
rect 6731 8134 6761 8186
rect 6785 8134 6795 8186
rect 6795 8134 6841 8186
rect 6545 8132 6601 8134
rect 6625 8132 6681 8134
rect 6705 8132 6761 8134
rect 6785 8132 6841 8134
rect 12134 7642 12190 7644
rect 12214 7642 12270 7644
rect 12294 7642 12350 7644
rect 12374 7642 12430 7644
rect 12134 7590 12180 7642
rect 12180 7590 12190 7642
rect 12214 7590 12244 7642
rect 12244 7590 12256 7642
rect 12256 7590 12270 7642
rect 12294 7590 12308 7642
rect 12308 7590 12320 7642
rect 12320 7590 12350 7642
rect 12374 7590 12384 7642
rect 12384 7590 12430 7642
rect 12134 7588 12190 7590
rect 12214 7588 12270 7590
rect 12294 7588 12350 7590
rect 12374 7588 12430 7590
rect 6545 7098 6601 7100
rect 6625 7098 6681 7100
rect 6705 7098 6761 7100
rect 6785 7098 6841 7100
rect 6545 7046 6591 7098
rect 6591 7046 6601 7098
rect 6625 7046 6655 7098
rect 6655 7046 6667 7098
rect 6667 7046 6681 7098
rect 6705 7046 6719 7098
rect 6719 7046 6731 7098
rect 6731 7046 6761 7098
rect 6785 7046 6795 7098
rect 6795 7046 6841 7098
rect 6545 7044 6601 7046
rect 6625 7044 6681 7046
rect 6705 7044 6761 7046
rect 6785 7044 6841 7046
rect 12134 6554 12190 6556
rect 12214 6554 12270 6556
rect 12294 6554 12350 6556
rect 12374 6554 12430 6556
rect 12134 6502 12180 6554
rect 12180 6502 12190 6554
rect 12214 6502 12244 6554
rect 12244 6502 12256 6554
rect 12256 6502 12270 6554
rect 12294 6502 12308 6554
rect 12308 6502 12320 6554
rect 12320 6502 12350 6554
rect 12374 6502 12384 6554
rect 12384 6502 12430 6554
rect 12134 6500 12190 6502
rect 12214 6500 12270 6502
rect 12294 6500 12350 6502
rect 12374 6500 12430 6502
rect 6545 6010 6601 6012
rect 6625 6010 6681 6012
rect 6705 6010 6761 6012
rect 6785 6010 6841 6012
rect 6545 5958 6591 6010
rect 6591 5958 6601 6010
rect 6625 5958 6655 6010
rect 6655 5958 6667 6010
rect 6667 5958 6681 6010
rect 6705 5958 6719 6010
rect 6719 5958 6731 6010
rect 6731 5958 6761 6010
rect 6785 5958 6795 6010
rect 6795 5958 6841 6010
rect 6545 5956 6601 5958
rect 6625 5956 6681 5958
rect 6705 5956 6761 5958
rect 6785 5956 6841 5958
rect 12134 5466 12190 5468
rect 12214 5466 12270 5468
rect 12294 5466 12350 5468
rect 12374 5466 12430 5468
rect 12134 5414 12180 5466
rect 12180 5414 12190 5466
rect 12214 5414 12244 5466
rect 12244 5414 12256 5466
rect 12256 5414 12270 5466
rect 12294 5414 12308 5466
rect 12308 5414 12320 5466
rect 12320 5414 12350 5466
rect 12374 5414 12384 5466
rect 12384 5414 12430 5466
rect 12134 5412 12190 5414
rect 12214 5412 12270 5414
rect 12294 5412 12350 5414
rect 12374 5412 12430 5414
rect 6545 4922 6601 4924
rect 6625 4922 6681 4924
rect 6705 4922 6761 4924
rect 6785 4922 6841 4924
rect 6545 4870 6591 4922
rect 6591 4870 6601 4922
rect 6625 4870 6655 4922
rect 6655 4870 6667 4922
rect 6667 4870 6681 4922
rect 6705 4870 6719 4922
rect 6719 4870 6731 4922
rect 6731 4870 6761 4922
rect 6785 4870 6795 4922
rect 6795 4870 6841 4922
rect 6545 4868 6601 4870
rect 6625 4868 6681 4870
rect 6705 4868 6761 4870
rect 6785 4868 6841 4870
rect 3238 4528 3294 4584
rect 2042 992 2098 1048
rect 6545 3834 6601 3836
rect 6625 3834 6681 3836
rect 6705 3834 6761 3836
rect 6785 3834 6841 3836
rect 6545 3782 6591 3834
rect 6591 3782 6601 3834
rect 6625 3782 6655 3834
rect 6655 3782 6667 3834
rect 6667 3782 6681 3834
rect 6705 3782 6719 3834
rect 6719 3782 6731 3834
rect 6731 3782 6761 3834
rect 6785 3782 6795 3834
rect 6795 3782 6841 3834
rect 6545 3780 6601 3782
rect 6625 3780 6681 3782
rect 6705 3780 6761 3782
rect 6785 3780 6841 3782
rect 6545 2746 6601 2748
rect 6625 2746 6681 2748
rect 6705 2746 6761 2748
rect 6785 2746 6841 2748
rect 6545 2694 6591 2746
rect 6591 2694 6601 2746
rect 6625 2694 6655 2746
rect 6655 2694 6667 2746
rect 6667 2694 6681 2746
rect 6705 2694 6719 2746
rect 6719 2694 6731 2746
rect 6731 2694 6761 2746
rect 6785 2694 6795 2746
rect 6795 2694 6841 2746
rect 6545 2692 6601 2694
rect 6625 2692 6681 2694
rect 6705 2692 6761 2694
rect 6785 2692 6841 2694
rect 6545 1658 6601 1660
rect 6625 1658 6681 1660
rect 6705 1658 6761 1660
rect 6785 1658 6841 1660
rect 6545 1606 6591 1658
rect 6591 1606 6601 1658
rect 6625 1606 6655 1658
rect 6655 1606 6667 1658
rect 6667 1606 6681 1658
rect 6705 1606 6719 1658
rect 6719 1606 6731 1658
rect 6731 1606 6761 1658
rect 6785 1606 6795 1658
rect 6795 1606 6841 1658
rect 6545 1604 6601 1606
rect 6625 1604 6681 1606
rect 6705 1604 6761 1606
rect 6785 1604 6841 1606
rect 7286 1400 7342 1456
rect 12134 4378 12190 4380
rect 12214 4378 12270 4380
rect 12294 4378 12350 4380
rect 12374 4378 12430 4380
rect 12134 4326 12180 4378
rect 12180 4326 12190 4378
rect 12214 4326 12244 4378
rect 12244 4326 12256 4378
rect 12256 4326 12270 4378
rect 12294 4326 12308 4378
rect 12308 4326 12320 4378
rect 12320 4326 12350 4378
rect 12374 4326 12384 4378
rect 12384 4326 12430 4378
rect 12134 4324 12190 4326
rect 12214 4324 12270 4326
rect 12294 4324 12350 4326
rect 12374 4324 12430 4326
rect 16854 4120 16910 4176
rect 10414 3984 10470 4040
rect 9586 2896 9642 2952
rect 9678 1944 9734 2000
rect 8482 992 8538 1048
rect 8758 448 8814 504
rect 9494 1300 9496 1320
rect 9496 1300 9548 1320
rect 9548 1300 9550 1320
rect 9494 1264 9550 1300
rect 16210 3576 16266 3632
rect 12134 3290 12190 3292
rect 12214 3290 12270 3292
rect 12294 3290 12350 3292
rect 12374 3290 12430 3292
rect 12134 3238 12180 3290
rect 12180 3238 12190 3290
rect 12214 3238 12244 3290
rect 12244 3238 12256 3290
rect 12256 3238 12270 3290
rect 12294 3238 12308 3290
rect 12308 3238 12320 3290
rect 12320 3238 12350 3290
rect 12374 3238 12384 3290
rect 12384 3238 12430 3290
rect 12134 3236 12190 3238
rect 12214 3236 12270 3238
rect 12294 3236 12350 3238
rect 12374 3236 12430 3238
rect 10874 856 10930 912
rect 13726 2488 13782 2544
rect 12134 2202 12190 2204
rect 12214 2202 12270 2204
rect 12294 2202 12350 2204
rect 12374 2202 12430 2204
rect 12134 2150 12180 2202
rect 12180 2150 12190 2202
rect 12214 2150 12244 2202
rect 12244 2150 12256 2202
rect 12256 2150 12270 2202
rect 12294 2150 12308 2202
rect 12308 2150 12320 2202
rect 12320 2150 12350 2202
rect 12374 2150 12384 2202
rect 12384 2150 12430 2202
rect 12134 2148 12190 2150
rect 12214 2148 12270 2150
rect 12294 2148 12350 2150
rect 12374 2148 12430 2150
rect 11426 720 11482 776
rect 11886 312 11942 368
rect 12134 1114 12190 1116
rect 12214 1114 12270 1116
rect 12294 1114 12350 1116
rect 12374 1114 12430 1116
rect 12134 1062 12180 1114
rect 12180 1062 12190 1114
rect 12214 1062 12244 1114
rect 12244 1062 12256 1114
rect 12256 1062 12270 1114
rect 12294 1062 12308 1114
rect 12308 1062 12320 1114
rect 12320 1062 12350 1114
rect 12374 1062 12384 1114
rect 12384 1062 12430 1114
rect 12134 1060 12190 1062
rect 12214 1060 12270 1062
rect 12294 1060 12350 1062
rect 12374 1060 12430 1062
rect 13082 176 13138 232
rect 13726 1128 13782 1184
rect 16762 3440 16818 3496
rect 15658 1808 15714 1864
rect 17723 8186 17779 8188
rect 17803 8186 17859 8188
rect 17883 8186 17939 8188
rect 17963 8186 18019 8188
rect 17723 8134 17769 8186
rect 17769 8134 17779 8186
rect 17803 8134 17833 8186
rect 17833 8134 17845 8186
rect 17845 8134 17859 8186
rect 17883 8134 17897 8186
rect 17897 8134 17909 8186
rect 17909 8134 17939 8186
rect 17963 8134 17973 8186
rect 17973 8134 18019 8186
rect 17723 8132 17779 8134
rect 17803 8132 17859 8134
rect 17883 8132 17939 8134
rect 17963 8132 18019 8134
rect 17723 7098 17779 7100
rect 17803 7098 17859 7100
rect 17883 7098 17939 7100
rect 17963 7098 18019 7100
rect 17723 7046 17769 7098
rect 17769 7046 17779 7098
rect 17803 7046 17833 7098
rect 17833 7046 17845 7098
rect 17845 7046 17859 7098
rect 17883 7046 17897 7098
rect 17897 7046 17909 7098
rect 17909 7046 17939 7098
rect 17963 7046 17973 7098
rect 17973 7046 18019 7098
rect 17723 7044 17779 7046
rect 17803 7044 17859 7046
rect 17883 7044 17939 7046
rect 17963 7044 18019 7046
rect 17723 6010 17779 6012
rect 17803 6010 17859 6012
rect 17883 6010 17939 6012
rect 17963 6010 18019 6012
rect 17723 5958 17769 6010
rect 17769 5958 17779 6010
rect 17803 5958 17833 6010
rect 17833 5958 17845 6010
rect 17845 5958 17859 6010
rect 17883 5958 17897 6010
rect 17897 5958 17909 6010
rect 17909 5958 17939 6010
rect 17963 5958 17973 6010
rect 17973 5958 18019 6010
rect 17723 5956 17779 5958
rect 17803 5956 17859 5958
rect 17883 5956 17939 5958
rect 17963 5956 18019 5958
rect 17723 4922 17779 4924
rect 17803 4922 17859 4924
rect 17883 4922 17939 4924
rect 17963 4922 18019 4924
rect 17723 4870 17769 4922
rect 17769 4870 17779 4922
rect 17803 4870 17833 4922
rect 17833 4870 17845 4922
rect 17845 4870 17859 4922
rect 17883 4870 17897 4922
rect 17897 4870 17909 4922
rect 17909 4870 17939 4922
rect 17963 4870 17973 4922
rect 17973 4870 18019 4922
rect 17723 4868 17779 4870
rect 17803 4868 17859 4870
rect 17883 4868 17939 4870
rect 17963 4868 18019 4870
rect 17723 3834 17779 3836
rect 17803 3834 17859 3836
rect 17883 3834 17939 3836
rect 17963 3834 18019 3836
rect 17723 3782 17769 3834
rect 17769 3782 17779 3834
rect 17803 3782 17833 3834
rect 17833 3782 17845 3834
rect 17845 3782 17859 3834
rect 17883 3782 17897 3834
rect 17897 3782 17909 3834
rect 17909 3782 17939 3834
rect 17963 3782 17973 3834
rect 17973 3782 18019 3834
rect 17723 3780 17779 3782
rect 17803 3780 17859 3782
rect 17883 3780 17939 3782
rect 17963 3780 18019 3782
rect 17314 3032 17370 3088
rect 16946 1400 17002 1456
rect 17723 2746 17779 2748
rect 17803 2746 17859 2748
rect 17883 2746 17939 2748
rect 17963 2746 18019 2748
rect 17723 2694 17769 2746
rect 17769 2694 17779 2746
rect 17803 2694 17833 2746
rect 17833 2694 17845 2746
rect 17845 2694 17859 2746
rect 17883 2694 17897 2746
rect 17897 2694 17909 2746
rect 17909 2694 17939 2746
rect 17963 2694 17973 2746
rect 17973 2694 18019 2746
rect 17723 2692 17779 2694
rect 17803 2692 17859 2694
rect 17883 2692 17939 2694
rect 17963 2692 18019 2694
rect 17958 2352 18014 2408
rect 17590 1944 17646 2000
rect 17222 992 17278 1048
rect 17222 584 17278 640
rect 17723 1658 17779 1660
rect 17803 1658 17859 1660
rect 17883 1658 17939 1660
rect 17963 1658 18019 1660
rect 17723 1606 17769 1658
rect 17769 1606 17779 1658
rect 17803 1606 17833 1658
rect 17833 1606 17845 1658
rect 17845 1606 17859 1658
rect 17883 1606 17897 1658
rect 17897 1606 17909 1658
rect 17909 1606 17939 1658
rect 17963 1606 17973 1658
rect 17973 1606 18019 1658
rect 17723 1604 17779 1606
rect 17803 1604 17859 1606
rect 17883 1604 17939 1606
rect 17963 1604 18019 1606
rect 18602 1708 18604 1728
rect 18604 1708 18656 1728
rect 18656 1708 18658 1728
rect 18602 1672 18658 1708
rect 19062 2760 19118 2816
rect 19890 2896 19946 2952
rect 19614 2100 19670 2136
rect 19614 2080 19616 2100
rect 19616 2080 19668 2100
rect 19668 2080 19670 2100
rect 19338 1964 19394 2000
rect 19338 1944 19340 1964
rect 19340 1944 19392 1964
rect 19392 1944 19394 1964
rect 19246 1536 19302 1592
rect 20258 1264 20314 1320
rect 20902 2216 20958 2272
rect 21178 2080 21234 2136
rect 20626 1944 20682 2000
rect 20258 176 20314 232
rect 20534 1128 20590 1184
rect 23312 8730 23368 8732
rect 23392 8730 23448 8732
rect 23472 8730 23528 8732
rect 23552 8730 23608 8732
rect 23312 8678 23358 8730
rect 23358 8678 23368 8730
rect 23392 8678 23422 8730
rect 23422 8678 23434 8730
rect 23434 8678 23448 8730
rect 23472 8678 23486 8730
rect 23486 8678 23498 8730
rect 23498 8678 23528 8730
rect 23552 8678 23562 8730
rect 23562 8678 23608 8730
rect 23312 8676 23368 8678
rect 23392 8676 23448 8678
rect 23472 8676 23528 8678
rect 23552 8676 23608 8678
rect 23312 7642 23368 7644
rect 23392 7642 23448 7644
rect 23472 7642 23528 7644
rect 23552 7642 23608 7644
rect 23312 7590 23358 7642
rect 23358 7590 23368 7642
rect 23392 7590 23422 7642
rect 23422 7590 23434 7642
rect 23434 7590 23448 7642
rect 23472 7590 23486 7642
rect 23486 7590 23498 7642
rect 23498 7590 23528 7642
rect 23552 7590 23562 7642
rect 23562 7590 23608 7642
rect 23312 7588 23368 7590
rect 23392 7588 23448 7590
rect 23472 7588 23528 7590
rect 23552 7588 23608 7590
rect 23312 6554 23368 6556
rect 23392 6554 23448 6556
rect 23472 6554 23528 6556
rect 23552 6554 23608 6556
rect 23312 6502 23358 6554
rect 23358 6502 23368 6554
rect 23392 6502 23422 6554
rect 23422 6502 23434 6554
rect 23434 6502 23448 6554
rect 23472 6502 23486 6554
rect 23486 6502 23498 6554
rect 23498 6502 23528 6554
rect 23552 6502 23562 6554
rect 23562 6502 23608 6554
rect 23312 6500 23368 6502
rect 23392 6500 23448 6502
rect 23472 6500 23528 6502
rect 23552 6500 23608 6502
rect 23312 5466 23368 5468
rect 23392 5466 23448 5468
rect 23472 5466 23528 5468
rect 23552 5466 23608 5468
rect 23312 5414 23358 5466
rect 23358 5414 23368 5466
rect 23392 5414 23422 5466
rect 23422 5414 23434 5466
rect 23434 5414 23448 5466
rect 23472 5414 23486 5466
rect 23486 5414 23498 5466
rect 23498 5414 23528 5466
rect 23552 5414 23562 5466
rect 23562 5414 23608 5466
rect 23312 5412 23368 5414
rect 23392 5412 23448 5414
rect 23472 5412 23528 5414
rect 23552 5412 23608 5414
rect 23312 4378 23368 4380
rect 23392 4378 23448 4380
rect 23472 4378 23528 4380
rect 23552 4378 23608 4380
rect 23312 4326 23358 4378
rect 23358 4326 23368 4378
rect 23392 4326 23422 4378
rect 23422 4326 23434 4378
rect 23434 4326 23448 4378
rect 23472 4326 23486 4378
rect 23486 4326 23498 4378
rect 23498 4326 23528 4378
rect 23552 4326 23562 4378
rect 23562 4326 23608 4378
rect 23312 4324 23368 4326
rect 23392 4324 23448 4326
rect 23472 4324 23528 4326
rect 23552 4324 23608 4326
rect 23312 3290 23368 3292
rect 23392 3290 23448 3292
rect 23472 3290 23528 3292
rect 23552 3290 23608 3292
rect 23312 3238 23358 3290
rect 23358 3238 23368 3290
rect 23392 3238 23422 3290
rect 23422 3238 23434 3290
rect 23434 3238 23448 3290
rect 23472 3238 23486 3290
rect 23486 3238 23498 3290
rect 23498 3238 23528 3290
rect 23552 3238 23562 3290
rect 23562 3238 23608 3290
rect 23312 3236 23368 3238
rect 23392 3236 23448 3238
rect 23472 3236 23528 3238
rect 23552 3236 23608 3238
rect 23312 2202 23368 2204
rect 23392 2202 23448 2204
rect 23472 2202 23528 2204
rect 23552 2202 23608 2204
rect 23312 2150 23358 2202
rect 23358 2150 23368 2202
rect 23392 2150 23422 2202
rect 23422 2150 23434 2202
rect 23434 2150 23448 2202
rect 23472 2150 23486 2202
rect 23486 2150 23498 2202
rect 23498 2150 23528 2202
rect 23552 2150 23562 2202
rect 23562 2150 23608 2202
rect 23312 2148 23368 2150
rect 23392 2148 23448 2150
rect 23472 2148 23528 2150
rect 23552 2148 23608 2150
rect 25318 3984 25374 4040
rect 22834 1400 22890 1456
rect 23312 1114 23368 1116
rect 23392 1114 23448 1116
rect 23472 1114 23528 1116
rect 23552 1114 23608 1116
rect 23312 1062 23358 1114
rect 23358 1062 23368 1114
rect 23392 1062 23422 1114
rect 23422 1062 23434 1114
rect 23434 1062 23448 1114
rect 23472 1062 23486 1114
rect 23486 1062 23498 1114
rect 23498 1062 23528 1114
rect 23552 1062 23562 1114
rect 23562 1062 23608 1114
rect 23312 1060 23368 1062
rect 23392 1060 23448 1062
rect 23472 1060 23528 1062
rect 23552 1060 23608 1062
rect 24122 2216 24178 2272
rect 25134 2100 25190 2136
rect 25134 2080 25136 2100
rect 25136 2080 25188 2100
rect 25188 2080 25190 2100
rect 26606 4528 26662 4584
rect 25686 1128 25742 1184
rect 25686 448 25742 504
rect 34490 8730 34546 8732
rect 34570 8730 34626 8732
rect 34650 8730 34706 8732
rect 34730 8730 34786 8732
rect 34490 8678 34536 8730
rect 34536 8678 34546 8730
rect 34570 8678 34600 8730
rect 34600 8678 34612 8730
rect 34612 8678 34626 8730
rect 34650 8678 34664 8730
rect 34664 8678 34676 8730
rect 34676 8678 34706 8730
rect 34730 8678 34740 8730
rect 34740 8678 34786 8730
rect 34490 8676 34546 8678
rect 34570 8676 34626 8678
rect 34650 8676 34706 8678
rect 34730 8676 34786 8678
rect 45668 8730 45724 8732
rect 45748 8730 45804 8732
rect 45828 8730 45884 8732
rect 45908 8730 45964 8732
rect 45668 8678 45714 8730
rect 45714 8678 45724 8730
rect 45748 8678 45778 8730
rect 45778 8678 45790 8730
rect 45790 8678 45804 8730
rect 45828 8678 45842 8730
rect 45842 8678 45854 8730
rect 45854 8678 45884 8730
rect 45908 8678 45918 8730
rect 45918 8678 45964 8730
rect 45668 8676 45724 8678
rect 45748 8676 45804 8678
rect 45828 8676 45884 8678
rect 45908 8676 45964 8678
rect 28901 8186 28957 8188
rect 28981 8186 29037 8188
rect 29061 8186 29117 8188
rect 29141 8186 29197 8188
rect 28901 8134 28947 8186
rect 28947 8134 28957 8186
rect 28981 8134 29011 8186
rect 29011 8134 29023 8186
rect 29023 8134 29037 8186
rect 29061 8134 29075 8186
rect 29075 8134 29087 8186
rect 29087 8134 29117 8186
rect 29141 8134 29151 8186
rect 29151 8134 29197 8186
rect 28901 8132 28957 8134
rect 28981 8132 29037 8134
rect 29061 8132 29117 8134
rect 29141 8132 29197 8134
rect 28901 7098 28957 7100
rect 28981 7098 29037 7100
rect 29061 7098 29117 7100
rect 29141 7098 29197 7100
rect 28901 7046 28947 7098
rect 28947 7046 28957 7098
rect 28981 7046 29011 7098
rect 29011 7046 29023 7098
rect 29023 7046 29037 7098
rect 29061 7046 29075 7098
rect 29075 7046 29087 7098
rect 29087 7046 29117 7098
rect 29141 7046 29151 7098
rect 29151 7046 29197 7098
rect 28901 7044 28957 7046
rect 28981 7044 29037 7046
rect 29061 7044 29117 7046
rect 29141 7044 29197 7046
rect 28901 6010 28957 6012
rect 28981 6010 29037 6012
rect 29061 6010 29117 6012
rect 29141 6010 29197 6012
rect 28901 5958 28947 6010
rect 28947 5958 28957 6010
rect 28981 5958 29011 6010
rect 29011 5958 29023 6010
rect 29023 5958 29037 6010
rect 29061 5958 29075 6010
rect 29075 5958 29087 6010
rect 29087 5958 29117 6010
rect 29141 5958 29151 6010
rect 29151 5958 29197 6010
rect 28901 5956 28957 5958
rect 28981 5956 29037 5958
rect 29061 5956 29117 5958
rect 29141 5956 29197 5958
rect 28901 4922 28957 4924
rect 28981 4922 29037 4924
rect 29061 4922 29117 4924
rect 29141 4922 29197 4924
rect 28901 4870 28947 4922
rect 28947 4870 28957 4922
rect 28981 4870 29011 4922
rect 29011 4870 29023 4922
rect 29023 4870 29037 4922
rect 29061 4870 29075 4922
rect 29075 4870 29087 4922
rect 29087 4870 29117 4922
rect 29141 4870 29151 4922
rect 29151 4870 29197 4922
rect 28901 4868 28957 4870
rect 28981 4868 29037 4870
rect 29061 4868 29117 4870
rect 29141 4868 29197 4870
rect 28901 3834 28957 3836
rect 28981 3834 29037 3836
rect 29061 3834 29117 3836
rect 29141 3834 29197 3836
rect 28901 3782 28947 3834
rect 28947 3782 28957 3834
rect 28981 3782 29011 3834
rect 29011 3782 29023 3834
rect 29023 3782 29037 3834
rect 29061 3782 29075 3834
rect 29075 3782 29087 3834
rect 29087 3782 29117 3834
rect 29141 3782 29151 3834
rect 29151 3782 29197 3834
rect 28901 3780 28957 3782
rect 28981 3780 29037 3782
rect 29061 3780 29117 3782
rect 29141 3780 29197 3782
rect 28901 2746 28957 2748
rect 28981 2746 29037 2748
rect 29061 2746 29117 2748
rect 29141 2746 29197 2748
rect 28901 2694 28947 2746
rect 28947 2694 28957 2746
rect 28981 2694 29011 2746
rect 29011 2694 29023 2746
rect 29023 2694 29037 2746
rect 29061 2694 29075 2746
rect 29075 2694 29087 2746
rect 29087 2694 29117 2746
rect 29141 2694 29151 2746
rect 29151 2694 29197 2746
rect 28901 2692 28957 2694
rect 28981 2692 29037 2694
rect 29061 2692 29117 2694
rect 29141 2692 29197 2694
rect 27802 1536 27858 1592
rect 28170 1672 28226 1728
rect 28906 2216 28962 2272
rect 28901 1658 28957 1660
rect 28981 1658 29037 1660
rect 29061 1658 29117 1660
rect 29141 1658 29197 1660
rect 28901 1606 28947 1658
rect 28947 1606 28957 1658
rect 28981 1606 29011 1658
rect 29011 1606 29023 1658
rect 29023 1606 29037 1658
rect 29061 1606 29075 1658
rect 29075 1606 29087 1658
rect 29087 1606 29117 1658
rect 29141 1606 29151 1658
rect 29151 1606 29197 1658
rect 28901 1604 28957 1606
rect 28981 1604 29037 1606
rect 29061 1604 29117 1606
rect 29141 1604 29197 1606
rect 29826 720 29882 776
rect 29734 448 29790 504
rect 31206 2896 31262 2952
rect 30562 856 30618 912
rect 31022 2216 31078 2272
rect 30838 1128 30894 1184
rect 31390 2488 31446 2544
rect 31574 2080 31630 2136
rect 34490 7642 34546 7644
rect 34570 7642 34626 7644
rect 34650 7642 34706 7644
rect 34730 7642 34786 7644
rect 34490 7590 34536 7642
rect 34536 7590 34546 7642
rect 34570 7590 34600 7642
rect 34600 7590 34612 7642
rect 34612 7590 34626 7642
rect 34650 7590 34664 7642
rect 34664 7590 34676 7642
rect 34676 7590 34706 7642
rect 34730 7590 34740 7642
rect 34740 7590 34786 7642
rect 34490 7588 34546 7590
rect 34570 7588 34626 7590
rect 34650 7588 34706 7590
rect 34730 7588 34786 7590
rect 34490 6554 34546 6556
rect 34570 6554 34626 6556
rect 34650 6554 34706 6556
rect 34730 6554 34786 6556
rect 34490 6502 34536 6554
rect 34536 6502 34546 6554
rect 34570 6502 34600 6554
rect 34600 6502 34612 6554
rect 34612 6502 34626 6554
rect 34650 6502 34664 6554
rect 34664 6502 34676 6554
rect 34676 6502 34706 6554
rect 34730 6502 34740 6554
rect 34740 6502 34786 6554
rect 34490 6500 34546 6502
rect 34570 6500 34626 6502
rect 34650 6500 34706 6502
rect 34730 6500 34786 6502
rect 34490 5466 34546 5468
rect 34570 5466 34626 5468
rect 34650 5466 34706 5468
rect 34730 5466 34786 5468
rect 34490 5414 34536 5466
rect 34536 5414 34546 5466
rect 34570 5414 34600 5466
rect 34600 5414 34612 5466
rect 34612 5414 34626 5466
rect 34650 5414 34664 5466
rect 34664 5414 34676 5466
rect 34676 5414 34706 5466
rect 34730 5414 34740 5466
rect 34740 5414 34786 5466
rect 34490 5412 34546 5414
rect 34570 5412 34626 5414
rect 34650 5412 34706 5414
rect 34730 5412 34786 5414
rect 34490 4378 34546 4380
rect 34570 4378 34626 4380
rect 34650 4378 34706 4380
rect 34730 4378 34786 4380
rect 34490 4326 34536 4378
rect 34536 4326 34546 4378
rect 34570 4326 34600 4378
rect 34600 4326 34612 4378
rect 34612 4326 34626 4378
rect 34650 4326 34664 4378
rect 34664 4326 34676 4378
rect 34676 4326 34706 4378
rect 34730 4326 34740 4378
rect 34740 4326 34786 4378
rect 34490 4324 34546 4326
rect 34570 4324 34626 4326
rect 34650 4324 34706 4326
rect 34730 4324 34786 4326
rect 34490 3290 34546 3292
rect 34570 3290 34626 3292
rect 34650 3290 34706 3292
rect 34730 3290 34786 3292
rect 34490 3238 34536 3290
rect 34536 3238 34546 3290
rect 34570 3238 34600 3290
rect 34600 3238 34612 3290
rect 34612 3238 34626 3290
rect 34650 3238 34664 3290
rect 34664 3238 34676 3290
rect 34676 3238 34706 3290
rect 34730 3238 34740 3290
rect 34740 3238 34786 3290
rect 34490 3236 34546 3238
rect 34570 3236 34626 3238
rect 34650 3236 34706 3238
rect 34730 3236 34786 3238
rect 40079 8186 40135 8188
rect 40159 8186 40215 8188
rect 40239 8186 40295 8188
rect 40319 8186 40375 8188
rect 40079 8134 40125 8186
rect 40125 8134 40135 8186
rect 40159 8134 40189 8186
rect 40189 8134 40201 8186
rect 40201 8134 40215 8186
rect 40239 8134 40253 8186
rect 40253 8134 40265 8186
rect 40265 8134 40295 8186
rect 40319 8134 40329 8186
rect 40329 8134 40375 8186
rect 40079 8132 40135 8134
rect 40159 8132 40215 8134
rect 40239 8132 40295 8134
rect 40319 8132 40375 8134
rect 40079 7098 40135 7100
rect 40159 7098 40215 7100
rect 40239 7098 40295 7100
rect 40319 7098 40375 7100
rect 40079 7046 40125 7098
rect 40125 7046 40135 7098
rect 40159 7046 40189 7098
rect 40189 7046 40201 7098
rect 40201 7046 40215 7098
rect 40239 7046 40253 7098
rect 40253 7046 40265 7098
rect 40265 7046 40295 7098
rect 40319 7046 40329 7098
rect 40329 7046 40375 7098
rect 40079 7044 40135 7046
rect 40159 7044 40215 7046
rect 40239 7044 40295 7046
rect 40319 7044 40375 7046
rect 34242 2352 34298 2408
rect 34334 2216 34390 2272
rect 34490 2202 34546 2204
rect 34570 2202 34626 2204
rect 34650 2202 34706 2204
rect 34730 2202 34786 2204
rect 34490 2150 34536 2202
rect 34536 2150 34546 2202
rect 34570 2150 34600 2202
rect 34600 2150 34612 2202
rect 34612 2150 34626 2202
rect 34650 2150 34664 2202
rect 34664 2150 34676 2202
rect 34676 2150 34706 2202
rect 34730 2150 34740 2202
rect 34740 2150 34786 2202
rect 34490 2148 34546 2150
rect 34570 2148 34626 2150
rect 34650 2148 34706 2150
rect 34730 2148 34786 2150
rect 32126 584 32182 640
rect 34490 1114 34546 1116
rect 34570 1114 34626 1116
rect 34650 1114 34706 1116
rect 34730 1114 34786 1116
rect 34490 1062 34536 1114
rect 34536 1062 34546 1114
rect 34570 1062 34600 1114
rect 34600 1062 34612 1114
rect 34612 1062 34626 1114
rect 34650 1062 34664 1114
rect 34664 1062 34676 1114
rect 34676 1062 34706 1114
rect 34730 1062 34740 1114
rect 34740 1062 34786 1114
rect 34490 1060 34546 1062
rect 34570 1060 34626 1062
rect 34650 1060 34706 1062
rect 34730 1060 34786 1062
rect 39394 4120 39450 4176
rect 37554 3576 37610 3632
rect 36542 1284 36598 1320
rect 36542 1264 36544 1284
rect 36544 1264 36596 1284
rect 36596 1264 36598 1284
rect 38934 3440 38990 3496
rect 38106 3032 38162 3088
rect 38106 1808 38162 1864
rect 38750 1964 38806 2000
rect 38750 1944 38752 1964
rect 38752 1944 38804 1964
rect 38804 1944 38806 1964
rect 38934 1400 38990 1456
rect 40079 6010 40135 6012
rect 40159 6010 40215 6012
rect 40239 6010 40295 6012
rect 40319 6010 40375 6012
rect 40079 5958 40125 6010
rect 40125 5958 40135 6010
rect 40159 5958 40189 6010
rect 40189 5958 40201 6010
rect 40201 5958 40215 6010
rect 40239 5958 40253 6010
rect 40253 5958 40265 6010
rect 40265 5958 40295 6010
rect 40319 5958 40329 6010
rect 40329 5958 40375 6010
rect 40079 5956 40135 5958
rect 40159 5956 40215 5958
rect 40239 5956 40295 5958
rect 40319 5956 40375 5958
rect 40079 4922 40135 4924
rect 40159 4922 40215 4924
rect 40239 4922 40295 4924
rect 40319 4922 40375 4924
rect 40079 4870 40125 4922
rect 40125 4870 40135 4922
rect 40159 4870 40189 4922
rect 40189 4870 40201 4922
rect 40201 4870 40215 4922
rect 40239 4870 40253 4922
rect 40253 4870 40265 4922
rect 40265 4870 40295 4922
rect 40319 4870 40329 4922
rect 40329 4870 40375 4922
rect 40079 4868 40135 4870
rect 40159 4868 40215 4870
rect 40239 4868 40295 4870
rect 40319 4868 40375 4870
rect 40079 3834 40135 3836
rect 40159 3834 40215 3836
rect 40239 3834 40295 3836
rect 40319 3834 40375 3836
rect 40079 3782 40125 3834
rect 40125 3782 40135 3834
rect 40159 3782 40189 3834
rect 40189 3782 40201 3834
rect 40201 3782 40215 3834
rect 40239 3782 40253 3834
rect 40253 3782 40265 3834
rect 40265 3782 40295 3834
rect 40319 3782 40329 3834
rect 40329 3782 40375 3834
rect 40079 3780 40135 3782
rect 40159 3780 40215 3782
rect 40239 3780 40295 3782
rect 40319 3780 40375 3782
rect 40079 2746 40135 2748
rect 40159 2746 40215 2748
rect 40239 2746 40295 2748
rect 40319 2746 40375 2748
rect 40079 2694 40125 2746
rect 40125 2694 40135 2746
rect 40159 2694 40189 2746
rect 40189 2694 40201 2746
rect 40201 2694 40215 2746
rect 40239 2694 40253 2746
rect 40253 2694 40265 2746
rect 40265 2694 40295 2746
rect 40319 2694 40329 2746
rect 40329 2694 40375 2746
rect 40079 2692 40135 2694
rect 40159 2692 40215 2694
rect 40239 2692 40295 2694
rect 40319 2692 40375 2694
rect 40079 1658 40135 1660
rect 40159 1658 40215 1660
rect 40239 1658 40295 1660
rect 40319 1658 40375 1660
rect 40079 1606 40125 1658
rect 40125 1606 40135 1658
rect 40159 1606 40189 1658
rect 40189 1606 40201 1658
rect 40201 1606 40215 1658
rect 40239 1606 40253 1658
rect 40253 1606 40265 1658
rect 40265 1606 40295 1658
rect 40319 1606 40329 1658
rect 40329 1606 40375 1658
rect 40079 1604 40135 1606
rect 40159 1604 40215 1606
rect 40239 1604 40295 1606
rect 40319 1604 40375 1606
rect 45668 7642 45724 7644
rect 45748 7642 45804 7644
rect 45828 7642 45884 7644
rect 45908 7642 45964 7644
rect 45668 7590 45714 7642
rect 45714 7590 45724 7642
rect 45748 7590 45778 7642
rect 45778 7590 45790 7642
rect 45790 7590 45804 7642
rect 45828 7590 45842 7642
rect 45842 7590 45854 7642
rect 45854 7590 45884 7642
rect 45908 7590 45918 7642
rect 45918 7590 45964 7642
rect 45668 7588 45724 7590
rect 45748 7588 45804 7590
rect 45828 7588 45884 7590
rect 45908 7588 45964 7590
rect 45668 6554 45724 6556
rect 45748 6554 45804 6556
rect 45828 6554 45884 6556
rect 45908 6554 45964 6556
rect 45668 6502 45714 6554
rect 45714 6502 45724 6554
rect 45748 6502 45778 6554
rect 45778 6502 45790 6554
rect 45790 6502 45804 6554
rect 45828 6502 45842 6554
rect 45842 6502 45854 6554
rect 45854 6502 45884 6554
rect 45908 6502 45918 6554
rect 45918 6502 45964 6554
rect 45668 6500 45724 6502
rect 45748 6500 45804 6502
rect 45828 6500 45884 6502
rect 45908 6500 45964 6502
rect 45668 5466 45724 5468
rect 45748 5466 45804 5468
rect 45828 5466 45884 5468
rect 45908 5466 45964 5468
rect 45668 5414 45714 5466
rect 45714 5414 45724 5466
rect 45748 5414 45778 5466
rect 45778 5414 45790 5466
rect 45790 5414 45804 5466
rect 45828 5414 45842 5466
rect 45842 5414 45854 5466
rect 45854 5414 45884 5466
rect 45908 5414 45918 5466
rect 45918 5414 45964 5466
rect 45668 5412 45724 5414
rect 45748 5412 45804 5414
rect 45828 5412 45884 5414
rect 45908 5412 45964 5414
rect 45668 4378 45724 4380
rect 45748 4378 45804 4380
rect 45828 4378 45884 4380
rect 45908 4378 45964 4380
rect 45668 4326 45714 4378
rect 45714 4326 45724 4378
rect 45748 4326 45778 4378
rect 45778 4326 45790 4378
rect 45790 4326 45804 4378
rect 45828 4326 45842 4378
rect 45842 4326 45854 4378
rect 45854 4326 45884 4378
rect 45908 4326 45918 4378
rect 45918 4326 45964 4378
rect 45668 4324 45724 4326
rect 45748 4324 45804 4326
rect 45828 4324 45884 4326
rect 45908 4324 45964 4326
rect 45668 3290 45724 3292
rect 45748 3290 45804 3292
rect 45828 3290 45884 3292
rect 45908 3290 45964 3292
rect 45668 3238 45714 3290
rect 45714 3238 45724 3290
rect 45748 3238 45778 3290
rect 45778 3238 45790 3290
rect 45790 3238 45804 3290
rect 45828 3238 45842 3290
rect 45842 3238 45854 3290
rect 45854 3238 45884 3290
rect 45908 3238 45918 3290
rect 45918 3238 45964 3290
rect 45668 3236 45724 3238
rect 45748 3236 45804 3238
rect 45828 3236 45884 3238
rect 45908 3236 45964 3238
rect 45668 2202 45724 2204
rect 45748 2202 45804 2204
rect 45828 2202 45884 2204
rect 45908 2202 45964 2204
rect 45668 2150 45714 2202
rect 45714 2150 45724 2202
rect 45748 2150 45778 2202
rect 45778 2150 45790 2202
rect 45790 2150 45804 2202
rect 45828 2150 45842 2202
rect 45842 2150 45854 2202
rect 45854 2150 45884 2202
rect 45908 2150 45918 2202
rect 45918 2150 45964 2202
rect 45668 2148 45724 2150
rect 45748 2148 45804 2150
rect 45828 2148 45884 2150
rect 45908 2148 45964 2150
rect 45668 1114 45724 1116
rect 45748 1114 45804 1116
rect 45828 1114 45884 1116
rect 45908 1114 45964 1116
rect 45668 1062 45714 1114
rect 45714 1062 45724 1114
rect 45748 1062 45778 1114
rect 45778 1062 45790 1114
rect 45790 1062 45804 1114
rect 45828 1062 45842 1114
rect 45842 1062 45854 1114
rect 45854 1062 45884 1114
rect 45908 1062 45918 1114
rect 45918 1062 45964 1114
rect 45668 1060 45724 1062
rect 45748 1060 45804 1062
rect 45828 1060 45884 1062
rect 45908 1060 45964 1062
<< metal3 >>
rect 12124 8736 12440 8737
rect 12124 8672 12130 8736
rect 12194 8672 12210 8736
rect 12274 8672 12290 8736
rect 12354 8672 12370 8736
rect 12434 8672 12440 8736
rect 12124 8671 12440 8672
rect 23302 8736 23618 8737
rect 23302 8672 23308 8736
rect 23372 8672 23388 8736
rect 23452 8672 23468 8736
rect 23532 8672 23548 8736
rect 23612 8672 23618 8736
rect 23302 8671 23618 8672
rect 34480 8736 34796 8737
rect 34480 8672 34486 8736
rect 34550 8672 34566 8736
rect 34630 8672 34646 8736
rect 34710 8672 34726 8736
rect 34790 8672 34796 8736
rect 34480 8671 34796 8672
rect 45658 8736 45974 8737
rect 45658 8672 45664 8736
rect 45728 8672 45744 8736
rect 45808 8672 45824 8736
rect 45888 8672 45904 8736
rect 45968 8672 45974 8736
rect 45658 8671 45974 8672
rect 6535 8192 6851 8193
rect 6535 8128 6541 8192
rect 6605 8128 6621 8192
rect 6685 8128 6701 8192
rect 6765 8128 6781 8192
rect 6845 8128 6851 8192
rect 6535 8127 6851 8128
rect 17713 8192 18029 8193
rect 17713 8128 17719 8192
rect 17783 8128 17799 8192
rect 17863 8128 17879 8192
rect 17943 8128 17959 8192
rect 18023 8128 18029 8192
rect 17713 8127 18029 8128
rect 28891 8192 29207 8193
rect 28891 8128 28897 8192
rect 28961 8128 28977 8192
rect 29041 8128 29057 8192
rect 29121 8128 29137 8192
rect 29201 8128 29207 8192
rect 28891 8127 29207 8128
rect 40069 8192 40385 8193
rect 40069 8128 40075 8192
rect 40139 8128 40155 8192
rect 40219 8128 40235 8192
rect 40299 8128 40315 8192
rect 40379 8128 40385 8192
rect 40069 8127 40385 8128
rect 12124 7648 12440 7649
rect 12124 7584 12130 7648
rect 12194 7584 12210 7648
rect 12274 7584 12290 7648
rect 12354 7584 12370 7648
rect 12434 7584 12440 7648
rect 12124 7583 12440 7584
rect 23302 7648 23618 7649
rect 23302 7584 23308 7648
rect 23372 7584 23388 7648
rect 23452 7584 23468 7648
rect 23532 7584 23548 7648
rect 23612 7584 23618 7648
rect 23302 7583 23618 7584
rect 34480 7648 34796 7649
rect 34480 7584 34486 7648
rect 34550 7584 34566 7648
rect 34630 7584 34646 7648
rect 34710 7584 34726 7648
rect 34790 7584 34796 7648
rect 34480 7583 34796 7584
rect 45658 7648 45974 7649
rect 45658 7584 45664 7648
rect 45728 7584 45744 7648
rect 45808 7584 45824 7648
rect 45888 7584 45904 7648
rect 45968 7584 45974 7648
rect 45658 7583 45974 7584
rect 6535 7104 6851 7105
rect 6535 7040 6541 7104
rect 6605 7040 6621 7104
rect 6685 7040 6701 7104
rect 6765 7040 6781 7104
rect 6845 7040 6851 7104
rect 6535 7039 6851 7040
rect 17713 7104 18029 7105
rect 17713 7040 17719 7104
rect 17783 7040 17799 7104
rect 17863 7040 17879 7104
rect 17943 7040 17959 7104
rect 18023 7040 18029 7104
rect 17713 7039 18029 7040
rect 28891 7104 29207 7105
rect 28891 7040 28897 7104
rect 28961 7040 28977 7104
rect 29041 7040 29057 7104
rect 29121 7040 29137 7104
rect 29201 7040 29207 7104
rect 28891 7039 29207 7040
rect 40069 7104 40385 7105
rect 40069 7040 40075 7104
rect 40139 7040 40155 7104
rect 40219 7040 40235 7104
rect 40299 7040 40315 7104
rect 40379 7040 40385 7104
rect 40069 7039 40385 7040
rect 12124 6560 12440 6561
rect 12124 6496 12130 6560
rect 12194 6496 12210 6560
rect 12274 6496 12290 6560
rect 12354 6496 12370 6560
rect 12434 6496 12440 6560
rect 12124 6495 12440 6496
rect 23302 6560 23618 6561
rect 23302 6496 23308 6560
rect 23372 6496 23388 6560
rect 23452 6496 23468 6560
rect 23532 6496 23548 6560
rect 23612 6496 23618 6560
rect 23302 6495 23618 6496
rect 34480 6560 34796 6561
rect 34480 6496 34486 6560
rect 34550 6496 34566 6560
rect 34630 6496 34646 6560
rect 34710 6496 34726 6560
rect 34790 6496 34796 6560
rect 34480 6495 34796 6496
rect 45658 6560 45974 6561
rect 45658 6496 45664 6560
rect 45728 6496 45744 6560
rect 45808 6496 45824 6560
rect 45888 6496 45904 6560
rect 45968 6496 45974 6560
rect 45658 6495 45974 6496
rect 6535 6016 6851 6017
rect 6535 5952 6541 6016
rect 6605 5952 6621 6016
rect 6685 5952 6701 6016
rect 6765 5952 6781 6016
rect 6845 5952 6851 6016
rect 6535 5951 6851 5952
rect 17713 6016 18029 6017
rect 17713 5952 17719 6016
rect 17783 5952 17799 6016
rect 17863 5952 17879 6016
rect 17943 5952 17959 6016
rect 18023 5952 18029 6016
rect 17713 5951 18029 5952
rect 28891 6016 29207 6017
rect 28891 5952 28897 6016
rect 28961 5952 28977 6016
rect 29041 5952 29057 6016
rect 29121 5952 29137 6016
rect 29201 5952 29207 6016
rect 28891 5951 29207 5952
rect 40069 6016 40385 6017
rect 40069 5952 40075 6016
rect 40139 5952 40155 6016
rect 40219 5952 40235 6016
rect 40299 5952 40315 6016
rect 40379 5952 40385 6016
rect 40069 5951 40385 5952
rect 12124 5472 12440 5473
rect 12124 5408 12130 5472
rect 12194 5408 12210 5472
rect 12274 5408 12290 5472
rect 12354 5408 12370 5472
rect 12434 5408 12440 5472
rect 12124 5407 12440 5408
rect 23302 5472 23618 5473
rect 23302 5408 23308 5472
rect 23372 5408 23388 5472
rect 23452 5408 23468 5472
rect 23532 5408 23548 5472
rect 23612 5408 23618 5472
rect 23302 5407 23618 5408
rect 34480 5472 34796 5473
rect 34480 5408 34486 5472
rect 34550 5408 34566 5472
rect 34630 5408 34646 5472
rect 34710 5408 34726 5472
rect 34790 5408 34796 5472
rect 34480 5407 34796 5408
rect 45658 5472 45974 5473
rect 45658 5408 45664 5472
rect 45728 5408 45744 5472
rect 45808 5408 45824 5472
rect 45888 5408 45904 5472
rect 45968 5408 45974 5472
rect 45658 5407 45974 5408
rect 6535 4928 6851 4929
rect 6535 4864 6541 4928
rect 6605 4864 6621 4928
rect 6685 4864 6701 4928
rect 6765 4864 6781 4928
rect 6845 4864 6851 4928
rect 6535 4863 6851 4864
rect 17713 4928 18029 4929
rect 17713 4864 17719 4928
rect 17783 4864 17799 4928
rect 17863 4864 17879 4928
rect 17943 4864 17959 4928
rect 18023 4864 18029 4928
rect 17713 4863 18029 4864
rect 28891 4928 29207 4929
rect 28891 4864 28897 4928
rect 28961 4864 28977 4928
rect 29041 4864 29057 4928
rect 29121 4864 29137 4928
rect 29201 4864 29207 4928
rect 28891 4863 29207 4864
rect 40069 4928 40385 4929
rect 40069 4864 40075 4928
rect 40139 4864 40155 4928
rect 40219 4864 40235 4928
rect 40299 4864 40315 4928
rect 40379 4864 40385 4928
rect 40069 4863 40385 4864
rect 3233 4586 3299 4589
rect 26601 4586 26667 4589
rect 3233 4584 26667 4586
rect 3233 4528 3238 4584
rect 3294 4528 26606 4584
rect 26662 4528 26667 4584
rect 3233 4526 26667 4528
rect 3233 4523 3299 4526
rect 26601 4523 26667 4526
rect 12124 4384 12440 4385
rect 12124 4320 12130 4384
rect 12194 4320 12210 4384
rect 12274 4320 12290 4384
rect 12354 4320 12370 4384
rect 12434 4320 12440 4384
rect 12124 4319 12440 4320
rect 23302 4384 23618 4385
rect 23302 4320 23308 4384
rect 23372 4320 23388 4384
rect 23452 4320 23468 4384
rect 23532 4320 23548 4384
rect 23612 4320 23618 4384
rect 23302 4319 23618 4320
rect 34480 4384 34796 4385
rect 34480 4320 34486 4384
rect 34550 4320 34566 4384
rect 34630 4320 34646 4384
rect 34710 4320 34726 4384
rect 34790 4320 34796 4384
rect 34480 4319 34796 4320
rect 45658 4384 45974 4385
rect 45658 4320 45664 4384
rect 45728 4320 45744 4384
rect 45808 4320 45824 4384
rect 45888 4320 45904 4384
rect 45968 4320 45974 4384
rect 45658 4319 45974 4320
rect 16849 4178 16915 4181
rect 39389 4178 39455 4181
rect 16849 4176 39455 4178
rect 16849 4120 16854 4176
rect 16910 4120 39394 4176
rect 39450 4120 39455 4176
rect 16849 4118 39455 4120
rect 16849 4115 16915 4118
rect 39389 4115 39455 4118
rect 10409 4042 10475 4045
rect 25313 4042 25379 4045
rect 10409 4040 25379 4042
rect 10409 3984 10414 4040
rect 10470 3984 25318 4040
rect 25374 3984 25379 4040
rect 10409 3982 25379 3984
rect 10409 3979 10475 3982
rect 25313 3979 25379 3982
rect 6535 3840 6851 3841
rect 6535 3776 6541 3840
rect 6605 3776 6621 3840
rect 6685 3776 6701 3840
rect 6765 3776 6781 3840
rect 6845 3776 6851 3840
rect 6535 3775 6851 3776
rect 17713 3840 18029 3841
rect 17713 3776 17719 3840
rect 17783 3776 17799 3840
rect 17863 3776 17879 3840
rect 17943 3776 17959 3840
rect 18023 3776 18029 3840
rect 17713 3775 18029 3776
rect 28891 3840 29207 3841
rect 28891 3776 28897 3840
rect 28961 3776 28977 3840
rect 29041 3776 29057 3840
rect 29121 3776 29137 3840
rect 29201 3776 29207 3840
rect 28891 3775 29207 3776
rect 40069 3840 40385 3841
rect 40069 3776 40075 3840
rect 40139 3776 40155 3840
rect 40219 3776 40235 3840
rect 40299 3776 40315 3840
rect 40379 3776 40385 3840
rect 40069 3775 40385 3776
rect 16205 3634 16271 3637
rect 37549 3634 37615 3637
rect 16205 3632 37615 3634
rect 16205 3576 16210 3632
rect 16266 3576 37554 3632
rect 37610 3576 37615 3632
rect 16205 3574 37615 3576
rect 16205 3571 16271 3574
rect 37549 3571 37615 3574
rect 16757 3498 16823 3501
rect 38929 3498 38995 3501
rect 16757 3496 38995 3498
rect 16757 3440 16762 3496
rect 16818 3440 38934 3496
rect 38990 3440 38995 3496
rect 16757 3438 38995 3440
rect 16757 3435 16823 3438
rect 38929 3435 38995 3438
rect 12124 3296 12440 3297
rect 12124 3232 12130 3296
rect 12194 3232 12210 3296
rect 12274 3232 12290 3296
rect 12354 3232 12370 3296
rect 12434 3232 12440 3296
rect 12124 3231 12440 3232
rect 23302 3296 23618 3297
rect 23302 3232 23308 3296
rect 23372 3232 23388 3296
rect 23452 3232 23468 3296
rect 23532 3232 23548 3296
rect 23612 3232 23618 3296
rect 23302 3231 23618 3232
rect 34480 3296 34796 3297
rect 34480 3232 34486 3296
rect 34550 3232 34566 3296
rect 34630 3232 34646 3296
rect 34710 3232 34726 3296
rect 34790 3232 34796 3296
rect 34480 3231 34796 3232
rect 45658 3296 45974 3297
rect 45658 3232 45664 3296
rect 45728 3232 45744 3296
rect 45808 3232 45824 3296
rect 45888 3232 45904 3296
rect 45968 3232 45974 3296
rect 45658 3231 45974 3232
rect 17309 3090 17375 3093
rect 38101 3090 38167 3093
rect 17309 3088 38167 3090
rect 17309 3032 17314 3088
rect 17370 3032 38106 3088
rect 38162 3032 38167 3088
rect 17309 3030 38167 3032
rect 17309 3027 17375 3030
rect 38101 3027 38167 3030
rect 9581 2954 9647 2957
rect 19885 2954 19951 2957
rect 31201 2954 31267 2957
rect 9581 2952 19951 2954
rect 9581 2896 9586 2952
rect 9642 2896 19890 2952
rect 19946 2896 19951 2952
rect 9581 2894 19951 2896
rect 9581 2891 9647 2894
rect 19885 2891 19951 2894
rect 24166 2952 31267 2954
rect 24166 2896 31206 2952
rect 31262 2896 31267 2952
rect 24166 2894 31267 2896
rect 19057 2818 19123 2821
rect 24166 2818 24226 2894
rect 31201 2891 31267 2894
rect 19057 2816 24226 2818
rect 19057 2760 19062 2816
rect 19118 2760 24226 2816
rect 19057 2758 24226 2760
rect 19057 2755 19123 2758
rect 6535 2752 6851 2753
rect 6535 2688 6541 2752
rect 6605 2688 6621 2752
rect 6685 2688 6701 2752
rect 6765 2688 6781 2752
rect 6845 2688 6851 2752
rect 6535 2687 6851 2688
rect 17713 2752 18029 2753
rect 17713 2688 17719 2752
rect 17783 2688 17799 2752
rect 17863 2688 17879 2752
rect 17943 2688 17959 2752
rect 18023 2688 18029 2752
rect 17713 2687 18029 2688
rect 28891 2752 29207 2753
rect 28891 2688 28897 2752
rect 28961 2688 28977 2752
rect 29041 2688 29057 2752
rect 29121 2688 29137 2752
rect 29201 2688 29207 2752
rect 28891 2687 29207 2688
rect 40069 2752 40385 2753
rect 40069 2688 40075 2752
rect 40139 2688 40155 2752
rect 40219 2688 40235 2752
rect 40299 2688 40315 2752
rect 40379 2688 40385 2752
rect 40069 2687 40385 2688
rect 13721 2546 13787 2549
rect 31385 2546 31451 2549
rect 13721 2544 31451 2546
rect 13721 2488 13726 2544
rect 13782 2488 31390 2544
rect 31446 2488 31451 2544
rect 13721 2486 31451 2488
rect 13721 2483 13787 2486
rect 31385 2483 31451 2486
rect 17953 2410 18019 2413
rect 34237 2410 34303 2413
rect 17953 2408 34303 2410
rect 17953 2352 17958 2408
rect 18014 2352 34242 2408
rect 34298 2352 34303 2408
rect 17953 2350 34303 2352
rect 17953 2347 18019 2350
rect 34237 2347 34303 2350
rect 20897 2274 20963 2277
rect 16622 2272 20963 2274
rect 16622 2216 20902 2272
rect 20958 2216 20963 2272
rect 16622 2214 20963 2216
rect 12124 2208 12440 2209
rect 12124 2144 12130 2208
rect 12194 2144 12210 2208
rect 12274 2144 12290 2208
rect 12354 2144 12370 2208
rect 12434 2144 12440 2208
rect 12124 2143 12440 2144
rect 9673 2002 9739 2005
rect 16622 2002 16682 2214
rect 20897 2211 20963 2214
rect 24117 2274 24183 2277
rect 28901 2274 28967 2277
rect 24117 2272 28967 2274
rect 24117 2216 24122 2272
rect 24178 2216 28906 2272
rect 28962 2216 28967 2272
rect 24117 2214 28967 2216
rect 24117 2211 24183 2214
rect 28901 2211 28967 2214
rect 31017 2274 31083 2277
rect 34329 2274 34395 2277
rect 31017 2272 34395 2274
rect 31017 2216 31022 2272
rect 31078 2216 34334 2272
rect 34390 2216 34395 2272
rect 31017 2214 34395 2216
rect 31017 2211 31083 2214
rect 34329 2211 34395 2214
rect 23302 2208 23618 2209
rect 23302 2144 23308 2208
rect 23372 2144 23388 2208
rect 23452 2144 23468 2208
rect 23532 2144 23548 2208
rect 23612 2144 23618 2208
rect 23302 2143 23618 2144
rect 34480 2208 34796 2209
rect 34480 2144 34486 2208
rect 34550 2144 34566 2208
rect 34630 2144 34646 2208
rect 34710 2144 34726 2208
rect 34790 2144 34796 2208
rect 34480 2143 34796 2144
rect 45658 2208 45974 2209
rect 45658 2144 45664 2208
rect 45728 2144 45744 2208
rect 45808 2144 45824 2208
rect 45888 2144 45904 2208
rect 45968 2144 45974 2208
rect 45658 2143 45974 2144
rect 19609 2138 19675 2141
rect 21173 2138 21239 2141
rect 19609 2136 21239 2138
rect 19609 2080 19614 2136
rect 19670 2080 21178 2136
rect 21234 2080 21239 2136
rect 19609 2078 21239 2080
rect 19609 2075 19675 2078
rect 21173 2075 21239 2078
rect 25129 2138 25195 2141
rect 31569 2138 31635 2141
rect 25129 2136 31635 2138
rect 25129 2080 25134 2136
rect 25190 2080 31574 2136
rect 31630 2080 31635 2136
rect 25129 2078 31635 2080
rect 25129 2075 25195 2078
rect 31569 2075 31635 2078
rect 9673 2000 16682 2002
rect 9673 1944 9678 2000
rect 9734 1944 16682 2000
rect 9673 1942 16682 1944
rect 17585 2002 17651 2005
rect 19333 2002 19399 2005
rect 17585 2000 19399 2002
rect 17585 1944 17590 2000
rect 17646 1944 19338 2000
rect 19394 1944 19399 2000
rect 17585 1942 19399 1944
rect 9673 1939 9739 1942
rect 17585 1939 17651 1942
rect 19333 1939 19399 1942
rect 20621 2002 20687 2005
rect 38745 2002 38811 2005
rect 20621 2000 38811 2002
rect 20621 1944 20626 2000
rect 20682 1944 38750 2000
rect 38806 1944 38811 2000
rect 20621 1942 38811 1944
rect 20621 1939 20687 1942
rect 38745 1939 38811 1942
rect 15653 1866 15719 1869
rect 38101 1866 38167 1869
rect 15653 1864 38167 1866
rect 15653 1808 15658 1864
rect 15714 1808 38106 1864
rect 38162 1808 38167 1864
rect 15653 1806 38167 1808
rect 15653 1803 15719 1806
rect 38101 1803 38167 1806
rect 18597 1730 18663 1733
rect 28165 1730 28231 1733
rect 18597 1728 28231 1730
rect 18597 1672 18602 1728
rect 18658 1672 28170 1728
rect 28226 1672 28231 1728
rect 18597 1670 28231 1672
rect 18597 1667 18663 1670
rect 28165 1667 28231 1670
rect 6535 1664 6851 1665
rect 6535 1600 6541 1664
rect 6605 1600 6621 1664
rect 6685 1600 6701 1664
rect 6765 1600 6781 1664
rect 6845 1600 6851 1664
rect 6535 1599 6851 1600
rect 17713 1664 18029 1665
rect 17713 1600 17719 1664
rect 17783 1600 17799 1664
rect 17863 1600 17879 1664
rect 17943 1600 17959 1664
rect 18023 1600 18029 1664
rect 17713 1599 18029 1600
rect 28891 1664 29207 1665
rect 28891 1600 28897 1664
rect 28961 1600 28977 1664
rect 29041 1600 29057 1664
rect 29121 1600 29137 1664
rect 29201 1600 29207 1664
rect 28891 1599 29207 1600
rect 40069 1664 40385 1665
rect 40069 1600 40075 1664
rect 40139 1600 40155 1664
rect 40219 1600 40235 1664
rect 40299 1600 40315 1664
rect 40379 1600 40385 1664
rect 40069 1599 40385 1600
rect 19241 1594 19307 1597
rect 27797 1594 27863 1597
rect 19241 1592 27863 1594
rect 19241 1536 19246 1592
rect 19302 1536 27802 1592
rect 27858 1536 27863 1592
rect 19241 1534 27863 1536
rect 19241 1531 19307 1534
rect 27797 1531 27863 1534
rect 7281 1458 7347 1461
rect 16941 1458 17007 1461
rect 7281 1456 17007 1458
rect 7281 1400 7286 1456
rect 7342 1400 16946 1456
rect 17002 1400 17007 1456
rect 7281 1398 17007 1400
rect 7281 1395 7347 1398
rect 16941 1395 17007 1398
rect 22829 1458 22895 1461
rect 38929 1458 38995 1461
rect 22829 1456 38995 1458
rect 22829 1400 22834 1456
rect 22890 1400 38934 1456
rect 38990 1400 38995 1456
rect 22829 1398 38995 1400
rect 22829 1395 22895 1398
rect 38929 1395 38995 1398
rect 9489 1322 9555 1325
rect 20253 1322 20319 1325
rect 36537 1322 36603 1325
rect 9489 1320 13554 1322
rect 9489 1264 9494 1320
rect 9550 1264 13554 1320
rect 9489 1262 13554 1264
rect 9489 1259 9555 1262
rect 12124 1120 12440 1121
rect 12124 1056 12130 1120
rect 12194 1056 12210 1120
rect 12274 1056 12290 1120
rect 12354 1056 12370 1120
rect 12434 1056 12440 1120
rect 12124 1055 12440 1056
rect 2037 1050 2103 1053
rect 8477 1050 8543 1053
rect 2037 1048 8543 1050
rect 2037 992 2042 1048
rect 2098 992 8482 1048
rect 8538 992 8543 1048
rect 2037 990 8543 992
rect 13494 1050 13554 1262
rect 20253 1320 36603 1322
rect 20253 1264 20258 1320
rect 20314 1264 36542 1320
rect 36598 1264 36603 1320
rect 20253 1262 36603 1264
rect 20253 1259 20319 1262
rect 36537 1259 36603 1262
rect 13721 1186 13787 1189
rect 20529 1186 20595 1189
rect 13721 1184 20595 1186
rect 13721 1128 13726 1184
rect 13782 1128 20534 1184
rect 20590 1128 20595 1184
rect 13721 1126 20595 1128
rect 13721 1123 13787 1126
rect 20529 1123 20595 1126
rect 25681 1186 25747 1189
rect 30833 1186 30899 1189
rect 25681 1184 30899 1186
rect 25681 1128 25686 1184
rect 25742 1128 30838 1184
rect 30894 1128 30899 1184
rect 25681 1126 30899 1128
rect 25681 1123 25747 1126
rect 30833 1123 30899 1126
rect 23302 1120 23618 1121
rect 23302 1056 23308 1120
rect 23372 1056 23388 1120
rect 23452 1056 23468 1120
rect 23532 1056 23548 1120
rect 23612 1056 23618 1120
rect 23302 1055 23618 1056
rect 34480 1120 34796 1121
rect 34480 1056 34486 1120
rect 34550 1056 34566 1120
rect 34630 1056 34646 1120
rect 34710 1056 34726 1120
rect 34790 1056 34796 1120
rect 34480 1055 34796 1056
rect 45658 1120 45974 1121
rect 45658 1056 45664 1120
rect 45728 1056 45744 1120
rect 45808 1056 45824 1120
rect 45888 1056 45904 1120
rect 45968 1056 45974 1120
rect 45658 1055 45974 1056
rect 17217 1050 17283 1053
rect 13494 1048 17283 1050
rect 13494 992 17222 1048
rect 17278 992 17283 1048
rect 13494 990 17283 992
rect 2037 987 2103 990
rect 8477 987 8543 990
rect 17217 987 17283 990
rect 10869 914 10935 917
rect 30557 914 30623 917
rect 10869 912 30623 914
rect 10869 856 10874 912
rect 10930 856 30562 912
rect 30618 856 30623 912
rect 10869 854 30623 856
rect 10869 851 10935 854
rect 30557 851 30623 854
rect 11421 778 11487 781
rect 29821 778 29887 781
rect 11421 776 29887 778
rect 11421 720 11426 776
rect 11482 720 29826 776
rect 29882 720 29887 776
rect 11421 718 29887 720
rect 11421 715 11487 718
rect 29821 715 29887 718
rect 17217 642 17283 645
rect 32121 642 32187 645
rect 17217 640 32187 642
rect 17217 584 17222 640
rect 17278 584 32126 640
rect 32182 584 32187 640
rect 17217 582 32187 584
rect 17217 579 17283 582
rect 32121 579 32187 582
rect 8753 506 8819 509
rect 25681 506 25747 509
rect 29729 506 29795 509
rect 8753 504 25747 506
rect 8753 448 8758 504
rect 8814 448 25686 504
rect 25742 448 25747 504
rect 8753 446 25747 448
rect 8753 443 8819 446
rect 25681 443 25747 446
rect 25822 504 29795 506
rect 25822 448 29734 504
rect 29790 448 29795 504
rect 25822 446 29795 448
rect 11881 370 11947 373
rect 25822 370 25882 446
rect 29729 443 29795 446
rect 11881 368 25882 370
rect 11881 312 11886 368
rect 11942 312 25882 368
rect 11881 310 25882 312
rect 11881 307 11947 310
rect 13077 234 13143 237
rect 20253 234 20319 237
rect 13077 232 20319 234
rect 13077 176 13082 232
rect 13138 176 20258 232
rect 20314 176 20319 232
rect 13077 174 20319 176
rect 13077 171 13143 174
rect 20253 171 20319 174
<< via3 >>
rect 12130 8732 12194 8736
rect 12130 8676 12134 8732
rect 12134 8676 12190 8732
rect 12190 8676 12194 8732
rect 12130 8672 12194 8676
rect 12210 8732 12274 8736
rect 12210 8676 12214 8732
rect 12214 8676 12270 8732
rect 12270 8676 12274 8732
rect 12210 8672 12274 8676
rect 12290 8732 12354 8736
rect 12290 8676 12294 8732
rect 12294 8676 12350 8732
rect 12350 8676 12354 8732
rect 12290 8672 12354 8676
rect 12370 8732 12434 8736
rect 12370 8676 12374 8732
rect 12374 8676 12430 8732
rect 12430 8676 12434 8732
rect 12370 8672 12434 8676
rect 23308 8732 23372 8736
rect 23308 8676 23312 8732
rect 23312 8676 23368 8732
rect 23368 8676 23372 8732
rect 23308 8672 23372 8676
rect 23388 8732 23452 8736
rect 23388 8676 23392 8732
rect 23392 8676 23448 8732
rect 23448 8676 23452 8732
rect 23388 8672 23452 8676
rect 23468 8732 23532 8736
rect 23468 8676 23472 8732
rect 23472 8676 23528 8732
rect 23528 8676 23532 8732
rect 23468 8672 23532 8676
rect 23548 8732 23612 8736
rect 23548 8676 23552 8732
rect 23552 8676 23608 8732
rect 23608 8676 23612 8732
rect 23548 8672 23612 8676
rect 34486 8732 34550 8736
rect 34486 8676 34490 8732
rect 34490 8676 34546 8732
rect 34546 8676 34550 8732
rect 34486 8672 34550 8676
rect 34566 8732 34630 8736
rect 34566 8676 34570 8732
rect 34570 8676 34626 8732
rect 34626 8676 34630 8732
rect 34566 8672 34630 8676
rect 34646 8732 34710 8736
rect 34646 8676 34650 8732
rect 34650 8676 34706 8732
rect 34706 8676 34710 8732
rect 34646 8672 34710 8676
rect 34726 8732 34790 8736
rect 34726 8676 34730 8732
rect 34730 8676 34786 8732
rect 34786 8676 34790 8732
rect 34726 8672 34790 8676
rect 45664 8732 45728 8736
rect 45664 8676 45668 8732
rect 45668 8676 45724 8732
rect 45724 8676 45728 8732
rect 45664 8672 45728 8676
rect 45744 8732 45808 8736
rect 45744 8676 45748 8732
rect 45748 8676 45804 8732
rect 45804 8676 45808 8732
rect 45744 8672 45808 8676
rect 45824 8732 45888 8736
rect 45824 8676 45828 8732
rect 45828 8676 45884 8732
rect 45884 8676 45888 8732
rect 45824 8672 45888 8676
rect 45904 8732 45968 8736
rect 45904 8676 45908 8732
rect 45908 8676 45964 8732
rect 45964 8676 45968 8732
rect 45904 8672 45968 8676
rect 6541 8188 6605 8192
rect 6541 8132 6545 8188
rect 6545 8132 6601 8188
rect 6601 8132 6605 8188
rect 6541 8128 6605 8132
rect 6621 8188 6685 8192
rect 6621 8132 6625 8188
rect 6625 8132 6681 8188
rect 6681 8132 6685 8188
rect 6621 8128 6685 8132
rect 6701 8188 6765 8192
rect 6701 8132 6705 8188
rect 6705 8132 6761 8188
rect 6761 8132 6765 8188
rect 6701 8128 6765 8132
rect 6781 8188 6845 8192
rect 6781 8132 6785 8188
rect 6785 8132 6841 8188
rect 6841 8132 6845 8188
rect 6781 8128 6845 8132
rect 17719 8188 17783 8192
rect 17719 8132 17723 8188
rect 17723 8132 17779 8188
rect 17779 8132 17783 8188
rect 17719 8128 17783 8132
rect 17799 8188 17863 8192
rect 17799 8132 17803 8188
rect 17803 8132 17859 8188
rect 17859 8132 17863 8188
rect 17799 8128 17863 8132
rect 17879 8188 17943 8192
rect 17879 8132 17883 8188
rect 17883 8132 17939 8188
rect 17939 8132 17943 8188
rect 17879 8128 17943 8132
rect 17959 8188 18023 8192
rect 17959 8132 17963 8188
rect 17963 8132 18019 8188
rect 18019 8132 18023 8188
rect 17959 8128 18023 8132
rect 28897 8188 28961 8192
rect 28897 8132 28901 8188
rect 28901 8132 28957 8188
rect 28957 8132 28961 8188
rect 28897 8128 28961 8132
rect 28977 8188 29041 8192
rect 28977 8132 28981 8188
rect 28981 8132 29037 8188
rect 29037 8132 29041 8188
rect 28977 8128 29041 8132
rect 29057 8188 29121 8192
rect 29057 8132 29061 8188
rect 29061 8132 29117 8188
rect 29117 8132 29121 8188
rect 29057 8128 29121 8132
rect 29137 8188 29201 8192
rect 29137 8132 29141 8188
rect 29141 8132 29197 8188
rect 29197 8132 29201 8188
rect 29137 8128 29201 8132
rect 40075 8188 40139 8192
rect 40075 8132 40079 8188
rect 40079 8132 40135 8188
rect 40135 8132 40139 8188
rect 40075 8128 40139 8132
rect 40155 8188 40219 8192
rect 40155 8132 40159 8188
rect 40159 8132 40215 8188
rect 40215 8132 40219 8188
rect 40155 8128 40219 8132
rect 40235 8188 40299 8192
rect 40235 8132 40239 8188
rect 40239 8132 40295 8188
rect 40295 8132 40299 8188
rect 40235 8128 40299 8132
rect 40315 8188 40379 8192
rect 40315 8132 40319 8188
rect 40319 8132 40375 8188
rect 40375 8132 40379 8188
rect 40315 8128 40379 8132
rect 12130 7644 12194 7648
rect 12130 7588 12134 7644
rect 12134 7588 12190 7644
rect 12190 7588 12194 7644
rect 12130 7584 12194 7588
rect 12210 7644 12274 7648
rect 12210 7588 12214 7644
rect 12214 7588 12270 7644
rect 12270 7588 12274 7644
rect 12210 7584 12274 7588
rect 12290 7644 12354 7648
rect 12290 7588 12294 7644
rect 12294 7588 12350 7644
rect 12350 7588 12354 7644
rect 12290 7584 12354 7588
rect 12370 7644 12434 7648
rect 12370 7588 12374 7644
rect 12374 7588 12430 7644
rect 12430 7588 12434 7644
rect 12370 7584 12434 7588
rect 23308 7644 23372 7648
rect 23308 7588 23312 7644
rect 23312 7588 23368 7644
rect 23368 7588 23372 7644
rect 23308 7584 23372 7588
rect 23388 7644 23452 7648
rect 23388 7588 23392 7644
rect 23392 7588 23448 7644
rect 23448 7588 23452 7644
rect 23388 7584 23452 7588
rect 23468 7644 23532 7648
rect 23468 7588 23472 7644
rect 23472 7588 23528 7644
rect 23528 7588 23532 7644
rect 23468 7584 23532 7588
rect 23548 7644 23612 7648
rect 23548 7588 23552 7644
rect 23552 7588 23608 7644
rect 23608 7588 23612 7644
rect 23548 7584 23612 7588
rect 34486 7644 34550 7648
rect 34486 7588 34490 7644
rect 34490 7588 34546 7644
rect 34546 7588 34550 7644
rect 34486 7584 34550 7588
rect 34566 7644 34630 7648
rect 34566 7588 34570 7644
rect 34570 7588 34626 7644
rect 34626 7588 34630 7644
rect 34566 7584 34630 7588
rect 34646 7644 34710 7648
rect 34646 7588 34650 7644
rect 34650 7588 34706 7644
rect 34706 7588 34710 7644
rect 34646 7584 34710 7588
rect 34726 7644 34790 7648
rect 34726 7588 34730 7644
rect 34730 7588 34786 7644
rect 34786 7588 34790 7644
rect 34726 7584 34790 7588
rect 45664 7644 45728 7648
rect 45664 7588 45668 7644
rect 45668 7588 45724 7644
rect 45724 7588 45728 7644
rect 45664 7584 45728 7588
rect 45744 7644 45808 7648
rect 45744 7588 45748 7644
rect 45748 7588 45804 7644
rect 45804 7588 45808 7644
rect 45744 7584 45808 7588
rect 45824 7644 45888 7648
rect 45824 7588 45828 7644
rect 45828 7588 45884 7644
rect 45884 7588 45888 7644
rect 45824 7584 45888 7588
rect 45904 7644 45968 7648
rect 45904 7588 45908 7644
rect 45908 7588 45964 7644
rect 45964 7588 45968 7644
rect 45904 7584 45968 7588
rect 6541 7100 6605 7104
rect 6541 7044 6545 7100
rect 6545 7044 6601 7100
rect 6601 7044 6605 7100
rect 6541 7040 6605 7044
rect 6621 7100 6685 7104
rect 6621 7044 6625 7100
rect 6625 7044 6681 7100
rect 6681 7044 6685 7100
rect 6621 7040 6685 7044
rect 6701 7100 6765 7104
rect 6701 7044 6705 7100
rect 6705 7044 6761 7100
rect 6761 7044 6765 7100
rect 6701 7040 6765 7044
rect 6781 7100 6845 7104
rect 6781 7044 6785 7100
rect 6785 7044 6841 7100
rect 6841 7044 6845 7100
rect 6781 7040 6845 7044
rect 17719 7100 17783 7104
rect 17719 7044 17723 7100
rect 17723 7044 17779 7100
rect 17779 7044 17783 7100
rect 17719 7040 17783 7044
rect 17799 7100 17863 7104
rect 17799 7044 17803 7100
rect 17803 7044 17859 7100
rect 17859 7044 17863 7100
rect 17799 7040 17863 7044
rect 17879 7100 17943 7104
rect 17879 7044 17883 7100
rect 17883 7044 17939 7100
rect 17939 7044 17943 7100
rect 17879 7040 17943 7044
rect 17959 7100 18023 7104
rect 17959 7044 17963 7100
rect 17963 7044 18019 7100
rect 18019 7044 18023 7100
rect 17959 7040 18023 7044
rect 28897 7100 28961 7104
rect 28897 7044 28901 7100
rect 28901 7044 28957 7100
rect 28957 7044 28961 7100
rect 28897 7040 28961 7044
rect 28977 7100 29041 7104
rect 28977 7044 28981 7100
rect 28981 7044 29037 7100
rect 29037 7044 29041 7100
rect 28977 7040 29041 7044
rect 29057 7100 29121 7104
rect 29057 7044 29061 7100
rect 29061 7044 29117 7100
rect 29117 7044 29121 7100
rect 29057 7040 29121 7044
rect 29137 7100 29201 7104
rect 29137 7044 29141 7100
rect 29141 7044 29197 7100
rect 29197 7044 29201 7100
rect 29137 7040 29201 7044
rect 40075 7100 40139 7104
rect 40075 7044 40079 7100
rect 40079 7044 40135 7100
rect 40135 7044 40139 7100
rect 40075 7040 40139 7044
rect 40155 7100 40219 7104
rect 40155 7044 40159 7100
rect 40159 7044 40215 7100
rect 40215 7044 40219 7100
rect 40155 7040 40219 7044
rect 40235 7100 40299 7104
rect 40235 7044 40239 7100
rect 40239 7044 40295 7100
rect 40295 7044 40299 7100
rect 40235 7040 40299 7044
rect 40315 7100 40379 7104
rect 40315 7044 40319 7100
rect 40319 7044 40375 7100
rect 40375 7044 40379 7100
rect 40315 7040 40379 7044
rect 12130 6556 12194 6560
rect 12130 6500 12134 6556
rect 12134 6500 12190 6556
rect 12190 6500 12194 6556
rect 12130 6496 12194 6500
rect 12210 6556 12274 6560
rect 12210 6500 12214 6556
rect 12214 6500 12270 6556
rect 12270 6500 12274 6556
rect 12210 6496 12274 6500
rect 12290 6556 12354 6560
rect 12290 6500 12294 6556
rect 12294 6500 12350 6556
rect 12350 6500 12354 6556
rect 12290 6496 12354 6500
rect 12370 6556 12434 6560
rect 12370 6500 12374 6556
rect 12374 6500 12430 6556
rect 12430 6500 12434 6556
rect 12370 6496 12434 6500
rect 23308 6556 23372 6560
rect 23308 6500 23312 6556
rect 23312 6500 23368 6556
rect 23368 6500 23372 6556
rect 23308 6496 23372 6500
rect 23388 6556 23452 6560
rect 23388 6500 23392 6556
rect 23392 6500 23448 6556
rect 23448 6500 23452 6556
rect 23388 6496 23452 6500
rect 23468 6556 23532 6560
rect 23468 6500 23472 6556
rect 23472 6500 23528 6556
rect 23528 6500 23532 6556
rect 23468 6496 23532 6500
rect 23548 6556 23612 6560
rect 23548 6500 23552 6556
rect 23552 6500 23608 6556
rect 23608 6500 23612 6556
rect 23548 6496 23612 6500
rect 34486 6556 34550 6560
rect 34486 6500 34490 6556
rect 34490 6500 34546 6556
rect 34546 6500 34550 6556
rect 34486 6496 34550 6500
rect 34566 6556 34630 6560
rect 34566 6500 34570 6556
rect 34570 6500 34626 6556
rect 34626 6500 34630 6556
rect 34566 6496 34630 6500
rect 34646 6556 34710 6560
rect 34646 6500 34650 6556
rect 34650 6500 34706 6556
rect 34706 6500 34710 6556
rect 34646 6496 34710 6500
rect 34726 6556 34790 6560
rect 34726 6500 34730 6556
rect 34730 6500 34786 6556
rect 34786 6500 34790 6556
rect 34726 6496 34790 6500
rect 45664 6556 45728 6560
rect 45664 6500 45668 6556
rect 45668 6500 45724 6556
rect 45724 6500 45728 6556
rect 45664 6496 45728 6500
rect 45744 6556 45808 6560
rect 45744 6500 45748 6556
rect 45748 6500 45804 6556
rect 45804 6500 45808 6556
rect 45744 6496 45808 6500
rect 45824 6556 45888 6560
rect 45824 6500 45828 6556
rect 45828 6500 45884 6556
rect 45884 6500 45888 6556
rect 45824 6496 45888 6500
rect 45904 6556 45968 6560
rect 45904 6500 45908 6556
rect 45908 6500 45964 6556
rect 45964 6500 45968 6556
rect 45904 6496 45968 6500
rect 6541 6012 6605 6016
rect 6541 5956 6545 6012
rect 6545 5956 6601 6012
rect 6601 5956 6605 6012
rect 6541 5952 6605 5956
rect 6621 6012 6685 6016
rect 6621 5956 6625 6012
rect 6625 5956 6681 6012
rect 6681 5956 6685 6012
rect 6621 5952 6685 5956
rect 6701 6012 6765 6016
rect 6701 5956 6705 6012
rect 6705 5956 6761 6012
rect 6761 5956 6765 6012
rect 6701 5952 6765 5956
rect 6781 6012 6845 6016
rect 6781 5956 6785 6012
rect 6785 5956 6841 6012
rect 6841 5956 6845 6012
rect 6781 5952 6845 5956
rect 17719 6012 17783 6016
rect 17719 5956 17723 6012
rect 17723 5956 17779 6012
rect 17779 5956 17783 6012
rect 17719 5952 17783 5956
rect 17799 6012 17863 6016
rect 17799 5956 17803 6012
rect 17803 5956 17859 6012
rect 17859 5956 17863 6012
rect 17799 5952 17863 5956
rect 17879 6012 17943 6016
rect 17879 5956 17883 6012
rect 17883 5956 17939 6012
rect 17939 5956 17943 6012
rect 17879 5952 17943 5956
rect 17959 6012 18023 6016
rect 17959 5956 17963 6012
rect 17963 5956 18019 6012
rect 18019 5956 18023 6012
rect 17959 5952 18023 5956
rect 28897 6012 28961 6016
rect 28897 5956 28901 6012
rect 28901 5956 28957 6012
rect 28957 5956 28961 6012
rect 28897 5952 28961 5956
rect 28977 6012 29041 6016
rect 28977 5956 28981 6012
rect 28981 5956 29037 6012
rect 29037 5956 29041 6012
rect 28977 5952 29041 5956
rect 29057 6012 29121 6016
rect 29057 5956 29061 6012
rect 29061 5956 29117 6012
rect 29117 5956 29121 6012
rect 29057 5952 29121 5956
rect 29137 6012 29201 6016
rect 29137 5956 29141 6012
rect 29141 5956 29197 6012
rect 29197 5956 29201 6012
rect 29137 5952 29201 5956
rect 40075 6012 40139 6016
rect 40075 5956 40079 6012
rect 40079 5956 40135 6012
rect 40135 5956 40139 6012
rect 40075 5952 40139 5956
rect 40155 6012 40219 6016
rect 40155 5956 40159 6012
rect 40159 5956 40215 6012
rect 40215 5956 40219 6012
rect 40155 5952 40219 5956
rect 40235 6012 40299 6016
rect 40235 5956 40239 6012
rect 40239 5956 40295 6012
rect 40295 5956 40299 6012
rect 40235 5952 40299 5956
rect 40315 6012 40379 6016
rect 40315 5956 40319 6012
rect 40319 5956 40375 6012
rect 40375 5956 40379 6012
rect 40315 5952 40379 5956
rect 12130 5468 12194 5472
rect 12130 5412 12134 5468
rect 12134 5412 12190 5468
rect 12190 5412 12194 5468
rect 12130 5408 12194 5412
rect 12210 5468 12274 5472
rect 12210 5412 12214 5468
rect 12214 5412 12270 5468
rect 12270 5412 12274 5468
rect 12210 5408 12274 5412
rect 12290 5468 12354 5472
rect 12290 5412 12294 5468
rect 12294 5412 12350 5468
rect 12350 5412 12354 5468
rect 12290 5408 12354 5412
rect 12370 5468 12434 5472
rect 12370 5412 12374 5468
rect 12374 5412 12430 5468
rect 12430 5412 12434 5468
rect 12370 5408 12434 5412
rect 23308 5468 23372 5472
rect 23308 5412 23312 5468
rect 23312 5412 23368 5468
rect 23368 5412 23372 5468
rect 23308 5408 23372 5412
rect 23388 5468 23452 5472
rect 23388 5412 23392 5468
rect 23392 5412 23448 5468
rect 23448 5412 23452 5468
rect 23388 5408 23452 5412
rect 23468 5468 23532 5472
rect 23468 5412 23472 5468
rect 23472 5412 23528 5468
rect 23528 5412 23532 5468
rect 23468 5408 23532 5412
rect 23548 5468 23612 5472
rect 23548 5412 23552 5468
rect 23552 5412 23608 5468
rect 23608 5412 23612 5468
rect 23548 5408 23612 5412
rect 34486 5468 34550 5472
rect 34486 5412 34490 5468
rect 34490 5412 34546 5468
rect 34546 5412 34550 5468
rect 34486 5408 34550 5412
rect 34566 5468 34630 5472
rect 34566 5412 34570 5468
rect 34570 5412 34626 5468
rect 34626 5412 34630 5468
rect 34566 5408 34630 5412
rect 34646 5468 34710 5472
rect 34646 5412 34650 5468
rect 34650 5412 34706 5468
rect 34706 5412 34710 5468
rect 34646 5408 34710 5412
rect 34726 5468 34790 5472
rect 34726 5412 34730 5468
rect 34730 5412 34786 5468
rect 34786 5412 34790 5468
rect 34726 5408 34790 5412
rect 45664 5468 45728 5472
rect 45664 5412 45668 5468
rect 45668 5412 45724 5468
rect 45724 5412 45728 5468
rect 45664 5408 45728 5412
rect 45744 5468 45808 5472
rect 45744 5412 45748 5468
rect 45748 5412 45804 5468
rect 45804 5412 45808 5468
rect 45744 5408 45808 5412
rect 45824 5468 45888 5472
rect 45824 5412 45828 5468
rect 45828 5412 45884 5468
rect 45884 5412 45888 5468
rect 45824 5408 45888 5412
rect 45904 5468 45968 5472
rect 45904 5412 45908 5468
rect 45908 5412 45964 5468
rect 45964 5412 45968 5468
rect 45904 5408 45968 5412
rect 6541 4924 6605 4928
rect 6541 4868 6545 4924
rect 6545 4868 6601 4924
rect 6601 4868 6605 4924
rect 6541 4864 6605 4868
rect 6621 4924 6685 4928
rect 6621 4868 6625 4924
rect 6625 4868 6681 4924
rect 6681 4868 6685 4924
rect 6621 4864 6685 4868
rect 6701 4924 6765 4928
rect 6701 4868 6705 4924
rect 6705 4868 6761 4924
rect 6761 4868 6765 4924
rect 6701 4864 6765 4868
rect 6781 4924 6845 4928
rect 6781 4868 6785 4924
rect 6785 4868 6841 4924
rect 6841 4868 6845 4924
rect 6781 4864 6845 4868
rect 17719 4924 17783 4928
rect 17719 4868 17723 4924
rect 17723 4868 17779 4924
rect 17779 4868 17783 4924
rect 17719 4864 17783 4868
rect 17799 4924 17863 4928
rect 17799 4868 17803 4924
rect 17803 4868 17859 4924
rect 17859 4868 17863 4924
rect 17799 4864 17863 4868
rect 17879 4924 17943 4928
rect 17879 4868 17883 4924
rect 17883 4868 17939 4924
rect 17939 4868 17943 4924
rect 17879 4864 17943 4868
rect 17959 4924 18023 4928
rect 17959 4868 17963 4924
rect 17963 4868 18019 4924
rect 18019 4868 18023 4924
rect 17959 4864 18023 4868
rect 28897 4924 28961 4928
rect 28897 4868 28901 4924
rect 28901 4868 28957 4924
rect 28957 4868 28961 4924
rect 28897 4864 28961 4868
rect 28977 4924 29041 4928
rect 28977 4868 28981 4924
rect 28981 4868 29037 4924
rect 29037 4868 29041 4924
rect 28977 4864 29041 4868
rect 29057 4924 29121 4928
rect 29057 4868 29061 4924
rect 29061 4868 29117 4924
rect 29117 4868 29121 4924
rect 29057 4864 29121 4868
rect 29137 4924 29201 4928
rect 29137 4868 29141 4924
rect 29141 4868 29197 4924
rect 29197 4868 29201 4924
rect 29137 4864 29201 4868
rect 40075 4924 40139 4928
rect 40075 4868 40079 4924
rect 40079 4868 40135 4924
rect 40135 4868 40139 4924
rect 40075 4864 40139 4868
rect 40155 4924 40219 4928
rect 40155 4868 40159 4924
rect 40159 4868 40215 4924
rect 40215 4868 40219 4924
rect 40155 4864 40219 4868
rect 40235 4924 40299 4928
rect 40235 4868 40239 4924
rect 40239 4868 40295 4924
rect 40295 4868 40299 4924
rect 40235 4864 40299 4868
rect 40315 4924 40379 4928
rect 40315 4868 40319 4924
rect 40319 4868 40375 4924
rect 40375 4868 40379 4924
rect 40315 4864 40379 4868
rect 12130 4380 12194 4384
rect 12130 4324 12134 4380
rect 12134 4324 12190 4380
rect 12190 4324 12194 4380
rect 12130 4320 12194 4324
rect 12210 4380 12274 4384
rect 12210 4324 12214 4380
rect 12214 4324 12270 4380
rect 12270 4324 12274 4380
rect 12210 4320 12274 4324
rect 12290 4380 12354 4384
rect 12290 4324 12294 4380
rect 12294 4324 12350 4380
rect 12350 4324 12354 4380
rect 12290 4320 12354 4324
rect 12370 4380 12434 4384
rect 12370 4324 12374 4380
rect 12374 4324 12430 4380
rect 12430 4324 12434 4380
rect 12370 4320 12434 4324
rect 23308 4380 23372 4384
rect 23308 4324 23312 4380
rect 23312 4324 23368 4380
rect 23368 4324 23372 4380
rect 23308 4320 23372 4324
rect 23388 4380 23452 4384
rect 23388 4324 23392 4380
rect 23392 4324 23448 4380
rect 23448 4324 23452 4380
rect 23388 4320 23452 4324
rect 23468 4380 23532 4384
rect 23468 4324 23472 4380
rect 23472 4324 23528 4380
rect 23528 4324 23532 4380
rect 23468 4320 23532 4324
rect 23548 4380 23612 4384
rect 23548 4324 23552 4380
rect 23552 4324 23608 4380
rect 23608 4324 23612 4380
rect 23548 4320 23612 4324
rect 34486 4380 34550 4384
rect 34486 4324 34490 4380
rect 34490 4324 34546 4380
rect 34546 4324 34550 4380
rect 34486 4320 34550 4324
rect 34566 4380 34630 4384
rect 34566 4324 34570 4380
rect 34570 4324 34626 4380
rect 34626 4324 34630 4380
rect 34566 4320 34630 4324
rect 34646 4380 34710 4384
rect 34646 4324 34650 4380
rect 34650 4324 34706 4380
rect 34706 4324 34710 4380
rect 34646 4320 34710 4324
rect 34726 4380 34790 4384
rect 34726 4324 34730 4380
rect 34730 4324 34786 4380
rect 34786 4324 34790 4380
rect 34726 4320 34790 4324
rect 45664 4380 45728 4384
rect 45664 4324 45668 4380
rect 45668 4324 45724 4380
rect 45724 4324 45728 4380
rect 45664 4320 45728 4324
rect 45744 4380 45808 4384
rect 45744 4324 45748 4380
rect 45748 4324 45804 4380
rect 45804 4324 45808 4380
rect 45744 4320 45808 4324
rect 45824 4380 45888 4384
rect 45824 4324 45828 4380
rect 45828 4324 45884 4380
rect 45884 4324 45888 4380
rect 45824 4320 45888 4324
rect 45904 4380 45968 4384
rect 45904 4324 45908 4380
rect 45908 4324 45964 4380
rect 45964 4324 45968 4380
rect 45904 4320 45968 4324
rect 6541 3836 6605 3840
rect 6541 3780 6545 3836
rect 6545 3780 6601 3836
rect 6601 3780 6605 3836
rect 6541 3776 6605 3780
rect 6621 3836 6685 3840
rect 6621 3780 6625 3836
rect 6625 3780 6681 3836
rect 6681 3780 6685 3836
rect 6621 3776 6685 3780
rect 6701 3836 6765 3840
rect 6701 3780 6705 3836
rect 6705 3780 6761 3836
rect 6761 3780 6765 3836
rect 6701 3776 6765 3780
rect 6781 3836 6845 3840
rect 6781 3780 6785 3836
rect 6785 3780 6841 3836
rect 6841 3780 6845 3836
rect 6781 3776 6845 3780
rect 17719 3836 17783 3840
rect 17719 3780 17723 3836
rect 17723 3780 17779 3836
rect 17779 3780 17783 3836
rect 17719 3776 17783 3780
rect 17799 3836 17863 3840
rect 17799 3780 17803 3836
rect 17803 3780 17859 3836
rect 17859 3780 17863 3836
rect 17799 3776 17863 3780
rect 17879 3836 17943 3840
rect 17879 3780 17883 3836
rect 17883 3780 17939 3836
rect 17939 3780 17943 3836
rect 17879 3776 17943 3780
rect 17959 3836 18023 3840
rect 17959 3780 17963 3836
rect 17963 3780 18019 3836
rect 18019 3780 18023 3836
rect 17959 3776 18023 3780
rect 28897 3836 28961 3840
rect 28897 3780 28901 3836
rect 28901 3780 28957 3836
rect 28957 3780 28961 3836
rect 28897 3776 28961 3780
rect 28977 3836 29041 3840
rect 28977 3780 28981 3836
rect 28981 3780 29037 3836
rect 29037 3780 29041 3836
rect 28977 3776 29041 3780
rect 29057 3836 29121 3840
rect 29057 3780 29061 3836
rect 29061 3780 29117 3836
rect 29117 3780 29121 3836
rect 29057 3776 29121 3780
rect 29137 3836 29201 3840
rect 29137 3780 29141 3836
rect 29141 3780 29197 3836
rect 29197 3780 29201 3836
rect 29137 3776 29201 3780
rect 40075 3836 40139 3840
rect 40075 3780 40079 3836
rect 40079 3780 40135 3836
rect 40135 3780 40139 3836
rect 40075 3776 40139 3780
rect 40155 3836 40219 3840
rect 40155 3780 40159 3836
rect 40159 3780 40215 3836
rect 40215 3780 40219 3836
rect 40155 3776 40219 3780
rect 40235 3836 40299 3840
rect 40235 3780 40239 3836
rect 40239 3780 40295 3836
rect 40295 3780 40299 3836
rect 40235 3776 40299 3780
rect 40315 3836 40379 3840
rect 40315 3780 40319 3836
rect 40319 3780 40375 3836
rect 40375 3780 40379 3836
rect 40315 3776 40379 3780
rect 12130 3292 12194 3296
rect 12130 3236 12134 3292
rect 12134 3236 12190 3292
rect 12190 3236 12194 3292
rect 12130 3232 12194 3236
rect 12210 3292 12274 3296
rect 12210 3236 12214 3292
rect 12214 3236 12270 3292
rect 12270 3236 12274 3292
rect 12210 3232 12274 3236
rect 12290 3292 12354 3296
rect 12290 3236 12294 3292
rect 12294 3236 12350 3292
rect 12350 3236 12354 3292
rect 12290 3232 12354 3236
rect 12370 3292 12434 3296
rect 12370 3236 12374 3292
rect 12374 3236 12430 3292
rect 12430 3236 12434 3292
rect 12370 3232 12434 3236
rect 23308 3292 23372 3296
rect 23308 3236 23312 3292
rect 23312 3236 23368 3292
rect 23368 3236 23372 3292
rect 23308 3232 23372 3236
rect 23388 3292 23452 3296
rect 23388 3236 23392 3292
rect 23392 3236 23448 3292
rect 23448 3236 23452 3292
rect 23388 3232 23452 3236
rect 23468 3292 23532 3296
rect 23468 3236 23472 3292
rect 23472 3236 23528 3292
rect 23528 3236 23532 3292
rect 23468 3232 23532 3236
rect 23548 3292 23612 3296
rect 23548 3236 23552 3292
rect 23552 3236 23608 3292
rect 23608 3236 23612 3292
rect 23548 3232 23612 3236
rect 34486 3292 34550 3296
rect 34486 3236 34490 3292
rect 34490 3236 34546 3292
rect 34546 3236 34550 3292
rect 34486 3232 34550 3236
rect 34566 3292 34630 3296
rect 34566 3236 34570 3292
rect 34570 3236 34626 3292
rect 34626 3236 34630 3292
rect 34566 3232 34630 3236
rect 34646 3292 34710 3296
rect 34646 3236 34650 3292
rect 34650 3236 34706 3292
rect 34706 3236 34710 3292
rect 34646 3232 34710 3236
rect 34726 3292 34790 3296
rect 34726 3236 34730 3292
rect 34730 3236 34786 3292
rect 34786 3236 34790 3292
rect 34726 3232 34790 3236
rect 45664 3292 45728 3296
rect 45664 3236 45668 3292
rect 45668 3236 45724 3292
rect 45724 3236 45728 3292
rect 45664 3232 45728 3236
rect 45744 3292 45808 3296
rect 45744 3236 45748 3292
rect 45748 3236 45804 3292
rect 45804 3236 45808 3292
rect 45744 3232 45808 3236
rect 45824 3292 45888 3296
rect 45824 3236 45828 3292
rect 45828 3236 45884 3292
rect 45884 3236 45888 3292
rect 45824 3232 45888 3236
rect 45904 3292 45968 3296
rect 45904 3236 45908 3292
rect 45908 3236 45964 3292
rect 45964 3236 45968 3292
rect 45904 3232 45968 3236
rect 6541 2748 6605 2752
rect 6541 2692 6545 2748
rect 6545 2692 6601 2748
rect 6601 2692 6605 2748
rect 6541 2688 6605 2692
rect 6621 2748 6685 2752
rect 6621 2692 6625 2748
rect 6625 2692 6681 2748
rect 6681 2692 6685 2748
rect 6621 2688 6685 2692
rect 6701 2748 6765 2752
rect 6701 2692 6705 2748
rect 6705 2692 6761 2748
rect 6761 2692 6765 2748
rect 6701 2688 6765 2692
rect 6781 2748 6845 2752
rect 6781 2692 6785 2748
rect 6785 2692 6841 2748
rect 6841 2692 6845 2748
rect 6781 2688 6845 2692
rect 17719 2748 17783 2752
rect 17719 2692 17723 2748
rect 17723 2692 17779 2748
rect 17779 2692 17783 2748
rect 17719 2688 17783 2692
rect 17799 2748 17863 2752
rect 17799 2692 17803 2748
rect 17803 2692 17859 2748
rect 17859 2692 17863 2748
rect 17799 2688 17863 2692
rect 17879 2748 17943 2752
rect 17879 2692 17883 2748
rect 17883 2692 17939 2748
rect 17939 2692 17943 2748
rect 17879 2688 17943 2692
rect 17959 2748 18023 2752
rect 17959 2692 17963 2748
rect 17963 2692 18019 2748
rect 18019 2692 18023 2748
rect 17959 2688 18023 2692
rect 28897 2748 28961 2752
rect 28897 2692 28901 2748
rect 28901 2692 28957 2748
rect 28957 2692 28961 2748
rect 28897 2688 28961 2692
rect 28977 2748 29041 2752
rect 28977 2692 28981 2748
rect 28981 2692 29037 2748
rect 29037 2692 29041 2748
rect 28977 2688 29041 2692
rect 29057 2748 29121 2752
rect 29057 2692 29061 2748
rect 29061 2692 29117 2748
rect 29117 2692 29121 2748
rect 29057 2688 29121 2692
rect 29137 2748 29201 2752
rect 29137 2692 29141 2748
rect 29141 2692 29197 2748
rect 29197 2692 29201 2748
rect 29137 2688 29201 2692
rect 40075 2748 40139 2752
rect 40075 2692 40079 2748
rect 40079 2692 40135 2748
rect 40135 2692 40139 2748
rect 40075 2688 40139 2692
rect 40155 2748 40219 2752
rect 40155 2692 40159 2748
rect 40159 2692 40215 2748
rect 40215 2692 40219 2748
rect 40155 2688 40219 2692
rect 40235 2748 40299 2752
rect 40235 2692 40239 2748
rect 40239 2692 40295 2748
rect 40295 2692 40299 2748
rect 40235 2688 40299 2692
rect 40315 2748 40379 2752
rect 40315 2692 40319 2748
rect 40319 2692 40375 2748
rect 40375 2692 40379 2748
rect 40315 2688 40379 2692
rect 12130 2204 12194 2208
rect 12130 2148 12134 2204
rect 12134 2148 12190 2204
rect 12190 2148 12194 2204
rect 12130 2144 12194 2148
rect 12210 2204 12274 2208
rect 12210 2148 12214 2204
rect 12214 2148 12270 2204
rect 12270 2148 12274 2204
rect 12210 2144 12274 2148
rect 12290 2204 12354 2208
rect 12290 2148 12294 2204
rect 12294 2148 12350 2204
rect 12350 2148 12354 2204
rect 12290 2144 12354 2148
rect 12370 2204 12434 2208
rect 12370 2148 12374 2204
rect 12374 2148 12430 2204
rect 12430 2148 12434 2204
rect 12370 2144 12434 2148
rect 23308 2204 23372 2208
rect 23308 2148 23312 2204
rect 23312 2148 23368 2204
rect 23368 2148 23372 2204
rect 23308 2144 23372 2148
rect 23388 2204 23452 2208
rect 23388 2148 23392 2204
rect 23392 2148 23448 2204
rect 23448 2148 23452 2204
rect 23388 2144 23452 2148
rect 23468 2204 23532 2208
rect 23468 2148 23472 2204
rect 23472 2148 23528 2204
rect 23528 2148 23532 2204
rect 23468 2144 23532 2148
rect 23548 2204 23612 2208
rect 23548 2148 23552 2204
rect 23552 2148 23608 2204
rect 23608 2148 23612 2204
rect 23548 2144 23612 2148
rect 34486 2204 34550 2208
rect 34486 2148 34490 2204
rect 34490 2148 34546 2204
rect 34546 2148 34550 2204
rect 34486 2144 34550 2148
rect 34566 2204 34630 2208
rect 34566 2148 34570 2204
rect 34570 2148 34626 2204
rect 34626 2148 34630 2204
rect 34566 2144 34630 2148
rect 34646 2204 34710 2208
rect 34646 2148 34650 2204
rect 34650 2148 34706 2204
rect 34706 2148 34710 2204
rect 34646 2144 34710 2148
rect 34726 2204 34790 2208
rect 34726 2148 34730 2204
rect 34730 2148 34786 2204
rect 34786 2148 34790 2204
rect 34726 2144 34790 2148
rect 45664 2204 45728 2208
rect 45664 2148 45668 2204
rect 45668 2148 45724 2204
rect 45724 2148 45728 2204
rect 45664 2144 45728 2148
rect 45744 2204 45808 2208
rect 45744 2148 45748 2204
rect 45748 2148 45804 2204
rect 45804 2148 45808 2204
rect 45744 2144 45808 2148
rect 45824 2204 45888 2208
rect 45824 2148 45828 2204
rect 45828 2148 45884 2204
rect 45884 2148 45888 2204
rect 45824 2144 45888 2148
rect 45904 2204 45968 2208
rect 45904 2148 45908 2204
rect 45908 2148 45964 2204
rect 45964 2148 45968 2204
rect 45904 2144 45968 2148
rect 6541 1660 6605 1664
rect 6541 1604 6545 1660
rect 6545 1604 6601 1660
rect 6601 1604 6605 1660
rect 6541 1600 6605 1604
rect 6621 1660 6685 1664
rect 6621 1604 6625 1660
rect 6625 1604 6681 1660
rect 6681 1604 6685 1660
rect 6621 1600 6685 1604
rect 6701 1660 6765 1664
rect 6701 1604 6705 1660
rect 6705 1604 6761 1660
rect 6761 1604 6765 1660
rect 6701 1600 6765 1604
rect 6781 1660 6845 1664
rect 6781 1604 6785 1660
rect 6785 1604 6841 1660
rect 6841 1604 6845 1660
rect 6781 1600 6845 1604
rect 17719 1660 17783 1664
rect 17719 1604 17723 1660
rect 17723 1604 17779 1660
rect 17779 1604 17783 1660
rect 17719 1600 17783 1604
rect 17799 1660 17863 1664
rect 17799 1604 17803 1660
rect 17803 1604 17859 1660
rect 17859 1604 17863 1660
rect 17799 1600 17863 1604
rect 17879 1660 17943 1664
rect 17879 1604 17883 1660
rect 17883 1604 17939 1660
rect 17939 1604 17943 1660
rect 17879 1600 17943 1604
rect 17959 1660 18023 1664
rect 17959 1604 17963 1660
rect 17963 1604 18019 1660
rect 18019 1604 18023 1660
rect 17959 1600 18023 1604
rect 28897 1660 28961 1664
rect 28897 1604 28901 1660
rect 28901 1604 28957 1660
rect 28957 1604 28961 1660
rect 28897 1600 28961 1604
rect 28977 1660 29041 1664
rect 28977 1604 28981 1660
rect 28981 1604 29037 1660
rect 29037 1604 29041 1660
rect 28977 1600 29041 1604
rect 29057 1660 29121 1664
rect 29057 1604 29061 1660
rect 29061 1604 29117 1660
rect 29117 1604 29121 1660
rect 29057 1600 29121 1604
rect 29137 1660 29201 1664
rect 29137 1604 29141 1660
rect 29141 1604 29197 1660
rect 29197 1604 29201 1660
rect 29137 1600 29201 1604
rect 40075 1660 40139 1664
rect 40075 1604 40079 1660
rect 40079 1604 40135 1660
rect 40135 1604 40139 1660
rect 40075 1600 40139 1604
rect 40155 1660 40219 1664
rect 40155 1604 40159 1660
rect 40159 1604 40215 1660
rect 40215 1604 40219 1660
rect 40155 1600 40219 1604
rect 40235 1660 40299 1664
rect 40235 1604 40239 1660
rect 40239 1604 40295 1660
rect 40295 1604 40299 1660
rect 40235 1600 40299 1604
rect 40315 1660 40379 1664
rect 40315 1604 40319 1660
rect 40319 1604 40375 1660
rect 40375 1604 40379 1660
rect 40315 1600 40379 1604
rect 12130 1116 12194 1120
rect 12130 1060 12134 1116
rect 12134 1060 12190 1116
rect 12190 1060 12194 1116
rect 12130 1056 12194 1060
rect 12210 1116 12274 1120
rect 12210 1060 12214 1116
rect 12214 1060 12270 1116
rect 12270 1060 12274 1116
rect 12210 1056 12274 1060
rect 12290 1116 12354 1120
rect 12290 1060 12294 1116
rect 12294 1060 12350 1116
rect 12350 1060 12354 1116
rect 12290 1056 12354 1060
rect 12370 1116 12434 1120
rect 12370 1060 12374 1116
rect 12374 1060 12430 1116
rect 12430 1060 12434 1116
rect 12370 1056 12434 1060
rect 23308 1116 23372 1120
rect 23308 1060 23312 1116
rect 23312 1060 23368 1116
rect 23368 1060 23372 1116
rect 23308 1056 23372 1060
rect 23388 1116 23452 1120
rect 23388 1060 23392 1116
rect 23392 1060 23448 1116
rect 23448 1060 23452 1116
rect 23388 1056 23452 1060
rect 23468 1116 23532 1120
rect 23468 1060 23472 1116
rect 23472 1060 23528 1116
rect 23528 1060 23532 1116
rect 23468 1056 23532 1060
rect 23548 1116 23612 1120
rect 23548 1060 23552 1116
rect 23552 1060 23608 1116
rect 23608 1060 23612 1116
rect 23548 1056 23612 1060
rect 34486 1116 34550 1120
rect 34486 1060 34490 1116
rect 34490 1060 34546 1116
rect 34546 1060 34550 1116
rect 34486 1056 34550 1060
rect 34566 1116 34630 1120
rect 34566 1060 34570 1116
rect 34570 1060 34626 1116
rect 34626 1060 34630 1116
rect 34566 1056 34630 1060
rect 34646 1116 34710 1120
rect 34646 1060 34650 1116
rect 34650 1060 34706 1116
rect 34706 1060 34710 1116
rect 34646 1056 34710 1060
rect 34726 1116 34790 1120
rect 34726 1060 34730 1116
rect 34730 1060 34786 1116
rect 34786 1060 34790 1116
rect 34726 1056 34790 1060
rect 45664 1116 45728 1120
rect 45664 1060 45668 1116
rect 45668 1060 45724 1116
rect 45724 1060 45728 1116
rect 45664 1056 45728 1060
rect 45744 1116 45808 1120
rect 45744 1060 45748 1116
rect 45748 1060 45804 1116
rect 45804 1060 45808 1116
rect 45744 1056 45808 1060
rect 45824 1116 45888 1120
rect 45824 1060 45828 1116
rect 45828 1060 45884 1116
rect 45884 1060 45888 1116
rect 45824 1056 45888 1060
rect 45904 1116 45968 1120
rect 45904 1060 45908 1116
rect 45908 1060 45964 1116
rect 45964 1060 45968 1116
rect 45904 1056 45968 1060
<< metal4 >>
rect 6533 8192 6853 8752
rect 6533 8128 6541 8192
rect 6605 8128 6621 8192
rect 6685 8128 6701 8192
rect 6765 8128 6781 8192
rect 6845 8128 6853 8192
rect 6533 7104 6853 8128
rect 6533 7040 6541 7104
rect 6605 7040 6621 7104
rect 6685 7040 6701 7104
rect 6765 7040 6781 7104
rect 6845 7040 6853 7104
rect 6533 6016 6853 7040
rect 6533 5952 6541 6016
rect 6605 5952 6621 6016
rect 6685 5952 6701 6016
rect 6765 5952 6781 6016
rect 6845 5952 6853 6016
rect 6533 4928 6853 5952
rect 6533 4864 6541 4928
rect 6605 4864 6621 4928
rect 6685 4864 6701 4928
rect 6765 4864 6781 4928
rect 6845 4864 6853 4928
rect 6533 3840 6853 4864
rect 6533 3776 6541 3840
rect 6605 3776 6621 3840
rect 6685 3776 6701 3840
rect 6765 3776 6781 3840
rect 6845 3776 6853 3840
rect 6533 2752 6853 3776
rect 6533 2688 6541 2752
rect 6605 2688 6621 2752
rect 6685 2688 6701 2752
rect 6765 2688 6781 2752
rect 6845 2688 6853 2752
rect 6533 1664 6853 2688
rect 6533 1600 6541 1664
rect 6605 1600 6621 1664
rect 6685 1600 6701 1664
rect 6765 1600 6781 1664
rect 6845 1600 6853 1664
rect 6533 1040 6853 1600
rect 12122 8736 12442 8752
rect 12122 8672 12130 8736
rect 12194 8672 12210 8736
rect 12274 8672 12290 8736
rect 12354 8672 12370 8736
rect 12434 8672 12442 8736
rect 12122 7648 12442 8672
rect 12122 7584 12130 7648
rect 12194 7584 12210 7648
rect 12274 7584 12290 7648
rect 12354 7584 12370 7648
rect 12434 7584 12442 7648
rect 12122 6560 12442 7584
rect 12122 6496 12130 6560
rect 12194 6496 12210 6560
rect 12274 6496 12290 6560
rect 12354 6496 12370 6560
rect 12434 6496 12442 6560
rect 12122 5472 12442 6496
rect 12122 5408 12130 5472
rect 12194 5408 12210 5472
rect 12274 5408 12290 5472
rect 12354 5408 12370 5472
rect 12434 5408 12442 5472
rect 12122 4384 12442 5408
rect 12122 4320 12130 4384
rect 12194 4320 12210 4384
rect 12274 4320 12290 4384
rect 12354 4320 12370 4384
rect 12434 4320 12442 4384
rect 12122 3296 12442 4320
rect 12122 3232 12130 3296
rect 12194 3232 12210 3296
rect 12274 3232 12290 3296
rect 12354 3232 12370 3296
rect 12434 3232 12442 3296
rect 12122 2208 12442 3232
rect 12122 2144 12130 2208
rect 12194 2144 12210 2208
rect 12274 2144 12290 2208
rect 12354 2144 12370 2208
rect 12434 2144 12442 2208
rect 12122 1120 12442 2144
rect 12122 1056 12130 1120
rect 12194 1056 12210 1120
rect 12274 1056 12290 1120
rect 12354 1056 12370 1120
rect 12434 1056 12442 1120
rect 12122 1040 12442 1056
rect 17711 8192 18031 8752
rect 17711 8128 17719 8192
rect 17783 8128 17799 8192
rect 17863 8128 17879 8192
rect 17943 8128 17959 8192
rect 18023 8128 18031 8192
rect 17711 7104 18031 8128
rect 17711 7040 17719 7104
rect 17783 7040 17799 7104
rect 17863 7040 17879 7104
rect 17943 7040 17959 7104
rect 18023 7040 18031 7104
rect 17711 6016 18031 7040
rect 17711 5952 17719 6016
rect 17783 5952 17799 6016
rect 17863 5952 17879 6016
rect 17943 5952 17959 6016
rect 18023 5952 18031 6016
rect 17711 4928 18031 5952
rect 17711 4864 17719 4928
rect 17783 4864 17799 4928
rect 17863 4864 17879 4928
rect 17943 4864 17959 4928
rect 18023 4864 18031 4928
rect 17711 3840 18031 4864
rect 17711 3776 17719 3840
rect 17783 3776 17799 3840
rect 17863 3776 17879 3840
rect 17943 3776 17959 3840
rect 18023 3776 18031 3840
rect 17711 2752 18031 3776
rect 17711 2688 17719 2752
rect 17783 2688 17799 2752
rect 17863 2688 17879 2752
rect 17943 2688 17959 2752
rect 18023 2688 18031 2752
rect 17711 1664 18031 2688
rect 17711 1600 17719 1664
rect 17783 1600 17799 1664
rect 17863 1600 17879 1664
rect 17943 1600 17959 1664
rect 18023 1600 18031 1664
rect 17711 1040 18031 1600
rect 23300 8736 23620 8752
rect 23300 8672 23308 8736
rect 23372 8672 23388 8736
rect 23452 8672 23468 8736
rect 23532 8672 23548 8736
rect 23612 8672 23620 8736
rect 23300 7648 23620 8672
rect 23300 7584 23308 7648
rect 23372 7584 23388 7648
rect 23452 7584 23468 7648
rect 23532 7584 23548 7648
rect 23612 7584 23620 7648
rect 23300 6560 23620 7584
rect 23300 6496 23308 6560
rect 23372 6496 23388 6560
rect 23452 6496 23468 6560
rect 23532 6496 23548 6560
rect 23612 6496 23620 6560
rect 23300 5472 23620 6496
rect 23300 5408 23308 5472
rect 23372 5408 23388 5472
rect 23452 5408 23468 5472
rect 23532 5408 23548 5472
rect 23612 5408 23620 5472
rect 23300 4384 23620 5408
rect 23300 4320 23308 4384
rect 23372 4320 23388 4384
rect 23452 4320 23468 4384
rect 23532 4320 23548 4384
rect 23612 4320 23620 4384
rect 23300 3296 23620 4320
rect 23300 3232 23308 3296
rect 23372 3232 23388 3296
rect 23452 3232 23468 3296
rect 23532 3232 23548 3296
rect 23612 3232 23620 3296
rect 23300 2208 23620 3232
rect 23300 2144 23308 2208
rect 23372 2144 23388 2208
rect 23452 2144 23468 2208
rect 23532 2144 23548 2208
rect 23612 2144 23620 2208
rect 23300 1120 23620 2144
rect 23300 1056 23308 1120
rect 23372 1056 23388 1120
rect 23452 1056 23468 1120
rect 23532 1056 23548 1120
rect 23612 1056 23620 1120
rect 23300 1040 23620 1056
rect 28889 8192 29209 8752
rect 28889 8128 28897 8192
rect 28961 8128 28977 8192
rect 29041 8128 29057 8192
rect 29121 8128 29137 8192
rect 29201 8128 29209 8192
rect 28889 7104 29209 8128
rect 28889 7040 28897 7104
rect 28961 7040 28977 7104
rect 29041 7040 29057 7104
rect 29121 7040 29137 7104
rect 29201 7040 29209 7104
rect 28889 6016 29209 7040
rect 28889 5952 28897 6016
rect 28961 5952 28977 6016
rect 29041 5952 29057 6016
rect 29121 5952 29137 6016
rect 29201 5952 29209 6016
rect 28889 4928 29209 5952
rect 28889 4864 28897 4928
rect 28961 4864 28977 4928
rect 29041 4864 29057 4928
rect 29121 4864 29137 4928
rect 29201 4864 29209 4928
rect 28889 3840 29209 4864
rect 28889 3776 28897 3840
rect 28961 3776 28977 3840
rect 29041 3776 29057 3840
rect 29121 3776 29137 3840
rect 29201 3776 29209 3840
rect 28889 2752 29209 3776
rect 28889 2688 28897 2752
rect 28961 2688 28977 2752
rect 29041 2688 29057 2752
rect 29121 2688 29137 2752
rect 29201 2688 29209 2752
rect 28889 1664 29209 2688
rect 28889 1600 28897 1664
rect 28961 1600 28977 1664
rect 29041 1600 29057 1664
rect 29121 1600 29137 1664
rect 29201 1600 29209 1664
rect 28889 1040 29209 1600
rect 34478 8736 34798 8752
rect 34478 8672 34486 8736
rect 34550 8672 34566 8736
rect 34630 8672 34646 8736
rect 34710 8672 34726 8736
rect 34790 8672 34798 8736
rect 34478 7648 34798 8672
rect 34478 7584 34486 7648
rect 34550 7584 34566 7648
rect 34630 7584 34646 7648
rect 34710 7584 34726 7648
rect 34790 7584 34798 7648
rect 34478 6560 34798 7584
rect 34478 6496 34486 6560
rect 34550 6496 34566 6560
rect 34630 6496 34646 6560
rect 34710 6496 34726 6560
rect 34790 6496 34798 6560
rect 34478 5472 34798 6496
rect 34478 5408 34486 5472
rect 34550 5408 34566 5472
rect 34630 5408 34646 5472
rect 34710 5408 34726 5472
rect 34790 5408 34798 5472
rect 34478 4384 34798 5408
rect 34478 4320 34486 4384
rect 34550 4320 34566 4384
rect 34630 4320 34646 4384
rect 34710 4320 34726 4384
rect 34790 4320 34798 4384
rect 34478 3296 34798 4320
rect 34478 3232 34486 3296
rect 34550 3232 34566 3296
rect 34630 3232 34646 3296
rect 34710 3232 34726 3296
rect 34790 3232 34798 3296
rect 34478 2208 34798 3232
rect 34478 2144 34486 2208
rect 34550 2144 34566 2208
rect 34630 2144 34646 2208
rect 34710 2144 34726 2208
rect 34790 2144 34798 2208
rect 34478 1120 34798 2144
rect 34478 1056 34486 1120
rect 34550 1056 34566 1120
rect 34630 1056 34646 1120
rect 34710 1056 34726 1120
rect 34790 1056 34798 1120
rect 34478 1040 34798 1056
rect 40067 8192 40387 8752
rect 40067 8128 40075 8192
rect 40139 8128 40155 8192
rect 40219 8128 40235 8192
rect 40299 8128 40315 8192
rect 40379 8128 40387 8192
rect 40067 7104 40387 8128
rect 40067 7040 40075 7104
rect 40139 7040 40155 7104
rect 40219 7040 40235 7104
rect 40299 7040 40315 7104
rect 40379 7040 40387 7104
rect 40067 6016 40387 7040
rect 40067 5952 40075 6016
rect 40139 5952 40155 6016
rect 40219 5952 40235 6016
rect 40299 5952 40315 6016
rect 40379 5952 40387 6016
rect 40067 4928 40387 5952
rect 40067 4864 40075 4928
rect 40139 4864 40155 4928
rect 40219 4864 40235 4928
rect 40299 4864 40315 4928
rect 40379 4864 40387 4928
rect 40067 3840 40387 4864
rect 40067 3776 40075 3840
rect 40139 3776 40155 3840
rect 40219 3776 40235 3840
rect 40299 3776 40315 3840
rect 40379 3776 40387 3840
rect 40067 2752 40387 3776
rect 40067 2688 40075 2752
rect 40139 2688 40155 2752
rect 40219 2688 40235 2752
rect 40299 2688 40315 2752
rect 40379 2688 40387 2752
rect 40067 1664 40387 2688
rect 40067 1600 40075 1664
rect 40139 1600 40155 1664
rect 40219 1600 40235 1664
rect 40299 1600 40315 1664
rect 40379 1600 40387 1664
rect 40067 1040 40387 1600
rect 45656 8736 45976 8752
rect 45656 8672 45664 8736
rect 45728 8672 45744 8736
rect 45808 8672 45824 8736
rect 45888 8672 45904 8736
rect 45968 8672 45976 8736
rect 45656 7648 45976 8672
rect 45656 7584 45664 7648
rect 45728 7584 45744 7648
rect 45808 7584 45824 7648
rect 45888 7584 45904 7648
rect 45968 7584 45976 7648
rect 45656 6560 45976 7584
rect 45656 6496 45664 6560
rect 45728 6496 45744 6560
rect 45808 6496 45824 6560
rect 45888 6496 45904 6560
rect 45968 6496 45976 6560
rect 45656 5472 45976 6496
rect 45656 5408 45664 5472
rect 45728 5408 45744 5472
rect 45808 5408 45824 5472
rect 45888 5408 45904 5472
rect 45968 5408 45976 5472
rect 45656 4384 45976 5408
rect 45656 4320 45664 4384
rect 45728 4320 45744 4384
rect 45808 4320 45824 4384
rect 45888 4320 45904 4384
rect 45968 4320 45976 4384
rect 45656 3296 45976 4320
rect 45656 3232 45664 3296
rect 45728 3232 45744 3296
rect 45808 3232 45824 3296
rect 45888 3232 45904 3296
rect 45968 3232 45976 3296
rect 45656 2208 45976 3232
rect 45656 2144 45664 2208
rect 45728 2144 45744 2208
rect 45808 2144 45824 2208
rect 45888 2144 45904 2208
rect 45968 2144 45976 2208
rect 45656 1120 45976 2144
rect 45656 1056 45664 1120
rect 45728 1056 45744 1120
rect 45808 1056 45824 1120
rect 45888 1056 45904 1120
rect 45968 1056 45976 1120
rect 45656 1040 45976 1056
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_7
timestamp 1688980957
transform 1 0 1748 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_11
timestamp 1688980957
transform 1 0 2116 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_22 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1688980957
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_35
timestamp 1688980957
transform 1 0 4324 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_39
timestamp 1688980957
transform 1 0 4692 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_43
timestamp 1688980957
transform 1 0 5060 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_47
timestamp 1688980957
transform 1 0 5428 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_51
timestamp 1688980957
transform 1 0 5796 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_63
timestamp 1688980957
transform 1 0 6900 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_67
timestamp 1688980957
transform 1 0 7268 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_71
timestamp 1688980957
transform 1 0 7636 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_75
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_79
timestamp 1688980957
transform 1 0 8372 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_95
timestamp 1688980957
transform 1 0 9844 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_99
timestamp 1688980957
transform 1 0 10212 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_103
timestamp 1688980957
transform 1 0 10580 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_107
timestamp 1688980957
transform 1 0 10948 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_119
timestamp 1688980957
transform 1 0 12052 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_123
timestamp 1688980957
transform 1 0 12420 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_127
timestamp 1688980957
transform 1 0 12788 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_131
timestamp 1688980957
transform 1 0 13156 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_135
timestamp 1688980957
transform 1 0 13524 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_176
timestamp 1688980957
transform 1 0 17296 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_218
timestamp 1688980957
transform 1 0 21160 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_234
timestamp 1688980957
transform 1 0 22632 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_250
timestamp 1688980957
transform 1 0 24104 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_253 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_278
timestamp 1688980957
transform 1 0 26680 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_287
timestamp 1688980957
transform 1 0 27508 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_446
timestamp 1688980957
transform 1 0 42136 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_455
timestamp 1688980957
transform 1 0 42964 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_459
timestamp 1688980957
transform 1 0 43332 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_463
timestamp 1688980957
transform 1 0 43700 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_467
timestamp 1688980957
transform 1 0 44068 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_471
timestamp 1688980957
transform 1 0 44436 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_475
timestamp 1688980957
transform 1 0 44804 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_19
timestamp 1688980957
transform 1 0 2852 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3220 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_35
timestamp 1688980957
transform 1 0 4324 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_47 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_87
timestamp 1688980957
transform 1 0 9108 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_91
timestamp 1688980957
transform 1 0 9476 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_95
timestamp 1688980957
transform 1 0 9844 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_107 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10948 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_220
timestamp 1688980957
transform 1 0 21344 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_252
timestamp 1688980957
transform 1 0 24288 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_266
timestamp 1688980957
transform 1 0 25576 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_278
timestamp 1688980957
transform 1 0 26680 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_285
timestamp 1688980957
transform 1 0 27324 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_295
timestamp 1688980957
transform 1 0 28244 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_322
timestamp 1688980957
transform 1 0 30728 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_343
timestamp 1688980957
transform 1 0 32660 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_351
timestamp 1688980957
transform 1 0 33396 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_364
timestamp 1688980957
transform 1 0 34592 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_379
timestamp 1688980957
transform 1 0 35972 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_400
timestamp 1688980957
transform 1 0 37904 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_407
timestamp 1688980957
transform 1 0 38548 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_423
timestamp 1688980957
transform 1 0 40020 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_436
timestamp 1688980957
transform 1 0 41216 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_452
timestamp 1688980957
transform 1 0 42688 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_464
timestamp 1688980957
transform 1 0 43792 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_472
timestamp 1688980957
transform 1 0 44528 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_479
timestamp 1688980957
transform 1 0 45172 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_180
timestamp 1688980957
transform 1 0 17664 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_188
timestamp 1688980957
transform 1 0 18400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_192
timestamp 1688980957
transform 1 0 18768 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_205
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_213
timestamp 1688980957
transform 1 0 20700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_256
timestamp 1688980957
transform 1 0 24656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_268
timestamp 1688980957
transform 1 0 25760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_294
timestamp 1688980957
transform 1 0 28152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_298
timestamp 1688980957
transform 1 0 28520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_306
timestamp 1688980957
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_318
timestamp 1688980957
transform 1 0 30360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_325
timestamp 1688980957
transform 1 0 31004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_332
timestamp 1688980957
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_336
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_340
timestamp 1688980957
transform 1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_346
timestamp 1688980957
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_352
timestamp 1688980957
transform 1 0 33488 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_370
timestamp 1688980957
transform 1 0 35144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_382
timestamp 1688980957
transform 1 0 36248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_390
timestamp 1688980957
transform 1 0 36984 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_394
timestamp 1688980957
transform 1 0 37352 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_406
timestamp 1688980957
transform 1 0 38456 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_414
timestamp 1688980957
transform 1 0 39192 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_439
timestamp 1688980957
transform 1 0 41492 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_443
timestamp 1688980957
transform 1 0 41860 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_455
timestamp 1688980957
transform 1 0 42964 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_463
timestamp 1688980957
transform 1 0 43700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_469
timestamp 1688980957
transform 1 0 44252 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_473
timestamp 1688980957
transform 1 0 44620 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_481
timestamp 1688980957
transform 1 0 45356 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1688980957
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_477
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_473
timestamp 1688980957
transform 1 0 44620 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_481
timestamp 1688980957
transform 1 0 45356 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_469
timestamp 1688980957
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 1688980957
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_473
timestamp 1688980957
transform 1 0 44620 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_481
timestamp 1688980957
transform 1 0 45356 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 1688980957
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_477
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_473
timestamp 1688980957
transform 1 0 44620 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_481
timestamp 1688980957
transform 1 0 45356 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_469
timestamp 1688980957
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 1688980957
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_477
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_461
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_473
timestamp 1688980957
transform 1 0 44620 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_481
timestamp 1688980957
transform 1 0 45356 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_469
timestamp 1688980957
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 1688980957
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_477
timestamp 1688980957
transform 1 0 44988 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_21
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_45
timestamp 1688980957
transform 1 0 5244 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_73
timestamp 1688980957
transform 1 0 7820 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_80
timestamp 1688980957
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_97
timestamp 1688980957
transform 1 0 10028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_104
timestamp 1688980957
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_121
timestamp 1688980957
transform 1 0 12236 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_128
timestamp 1688980957
transform 1 0 12880 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_147
timestamp 1688980957
transform 1 0 14628 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_152
timestamp 1688980957
transform 1 0 15088 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_164
timestamp 1688980957
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_176
timestamp 1688980957
transform 1 0 17296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_188
timestamp 1688980957
transform 1 0 18400 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_203
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_215
timestamp 1688980957
transform 1 0 20884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_219
timestamp 1688980957
transform 1 0 21252 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_241
timestamp 1688980957
transform 1 0 23276 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_248
timestamp 1688980957
transform 1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_253
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_265
timestamp 1688980957
transform 1 0 25484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_272
timestamp 1688980957
transform 1 0 26128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_289
timestamp 1688980957
transform 1 0 27692 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_296
timestamp 1688980957
transform 1 0 28336 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_309
timestamp 1688980957
transform 1 0 29532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_313
timestamp 1688980957
transform 1 0 29900 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_320
timestamp 1688980957
transform 1 0 30544 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_332
timestamp 1688980957
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_344
timestamp 1688980957
transform 1 0 32752 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_356
timestamp 1688980957
transform 1 0 33856 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_371
timestamp 1688980957
transform 1 0 35236 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_383
timestamp 1688980957
transform 1 0 36340 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_387
timestamp 1688980957
transform 1 0 36708 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_405
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_411
timestamp 1688980957
transform 1 0 38916 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_416
timestamp 1688980957
transform 1 0 39376 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_421
timestamp 1688980957
transform 1 0 39836 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_433
timestamp 1688980957
transform 1 0 40940 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_440
timestamp 1688980957
transform 1 0 41584 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_457
timestamp 1688980957
transform 1 0 43148 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_464
timestamp 1688980957
transform 1 0 43792 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 40664 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform -1 0 43332 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform -1 0 43700 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform -1 0 44068 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform -1 0 44436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform -1 0 44804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44988 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 45264 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 45264 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform -1 0 40940 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform -1 0 40664 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform -1 0 40940 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform -1 0 41216 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform -1 0 42136 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40940 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1688980957
transform 1 0 41308 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 42688 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform -1 0 42964 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 1656 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 1472 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 1840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 5520 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 5888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 6624 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1688980957
transform 1 0 6992 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1688980957
transform 1 0 7360 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1688980957
transform 1 0 2208 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 2576 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 2944 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 3312 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 4048 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 4416 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 4784 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 8096 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 11776 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 12144 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 12512 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 13248 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 13616 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1688980957
transform 1 0 9200 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform 1 0 9568 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1688980957
transform 1 0 9936 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 10304 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1688980957
transform 1 0 10672 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1688980957
transform 1 0 11040 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform -1 0 14352 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform 1 0 17480 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform -1 0 18032 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform -1 0 18308 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform 1 0 18584 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform -1 0 14628 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform -1 0 14904 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform -1 0 15180 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1688980957
transform -1 0 15456 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1688980957
transform -1 0 15732 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1688980957
transform -1 0 16008 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1688980957
transform -1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1688980957
transform -1 0 16560 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1688980957
transform -1 0 17020 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1688980957
transform -1 0 39744 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27876 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__00_
timestamp 1688980957
transform -1 0 22448 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__01_
timestamp 1688980957
transform -1 0 23368 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__02_
timestamp 1688980957
transform -1 0 23644 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__03_
timestamp 1688980957
transform -1 0 24748 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__04_
timestamp 1688980957
transform -1 0 25576 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__05_
timestamp 1688980957
transform -1 0 26404 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__06_
timestamp 1688980957
transform -1 0 26680 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__07_
timestamp 1688980957
transform -1 0 26864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__08_
timestamp 1688980957
transform -1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__09_
timestamp 1688980957
transform -1 0 20424 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__10_
timestamp 1688980957
transform -1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__11_
timestamp 1688980957
transform -1 0 21160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__12_
timestamp 1688980957
transform -1 0 22172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__13_
timestamp 1688980957
transform -1 0 20976 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__14_
timestamp 1688980957
transform -1 0 22724 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__15_
timestamp 1688980957
transform -1 0 21712 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__16_
timestamp 1688980957
transform -1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__17_
timestamp 1688980957
transform -1 0 27692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__18_
timestamp 1688980957
transform -1 0 31004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__19_
timestamp 1688980957
transform -1 0 31648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__20_
timestamp 1688980957
transform -1 0 32384 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__21_
timestamp 1688980957
transform -1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__22_
timestamp 1688980957
transform -1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__23_
timestamp 1688980957
transform 1 0 26312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__24_
timestamp 1688980957
transform -1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__25_
timestamp 1688980957
transform -1 0 29072 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__26_
timestamp 1688980957
transform -1 0 29348 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__27_
timestamp 1688980957
transform -1 0 29624 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__28_
timestamp 1688980957
transform -1 0 29900 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__29_
timestamp 1688980957
transform -1 0 30452 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__30_
timestamp 1688980957
transform -1 0 30728 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__31_
timestamp 1688980957
transform -1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__32_
timestamp 1688980957
transform 1 0 19044 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__33_
timestamp 1688980957
transform 1 0 18492 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__34_
timestamp 1688980957
transform 1 0 15732 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__35_
timestamp 1688980957
transform 1 0 15456 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__36_
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__37_
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__38_
timestamp 1688980957
transform 1 0 19872 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__39_
timestamp 1688980957
transform 1 0 20424 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__40_
timestamp 1688980957
transform 1 0 17940 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__41_
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__42_
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__43_
timestamp 1688980957
transform 1 0 17388 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__44_
timestamp 1688980957
transform 1 0 17112 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__45_
timestamp 1688980957
transform 1 0 17020 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__46_
timestamp 1688980957
transform 1 0 16284 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__47_
timestamp 1688980957
transform 1 0 16008 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__48_
timestamp 1688980957
transform -1 0 17940 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__49_
timestamp 1688980957
transform -1 0 18492 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__50_
timestamp 1688980957
transform -1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__51_
timestamp 1688980957
transform -1 0 19596 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1688980957
transform -1 0 26128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1688980957
transform -1 0 28336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output77 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30544 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1688980957
transform -1 0 32752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform -1 0 35236 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1688980957
transform -1 0 37168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1688980957
transform -1 0 39376 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform -1 0 41584 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1688980957
transform -1 0 43792 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 44988 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1688980957
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform -1 0 8464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1688980957
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform -1 0 12880 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1688980957
transform -1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1688980957
transform -1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform -1 0 19780 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1688980957
transform -1 0 21712 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform -1 0 23920 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1688980957
transform 1 0 19504 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1688980957
transform 1 0 19872 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform 1 0 20240 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 20608 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 25208 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 24656 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1688980957
transform 1 0 25760 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform 1 0 25760 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 26128 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 26956 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1688980957
transform 1 0 26956 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1688980957
transform 1 0 27876 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1688980957
transform 1 0 20976 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1688980957
transform 1 0 21344 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 22080 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1688980957
transform 1 0 22448 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1688980957
transform 1 0 22816 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1688980957
transform 1 0 23184 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 23552 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1688980957
transform 1 0 23920 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 27692 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 30912 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 32660 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 33212 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 32844 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform 1 0 33764 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform 1 0 34040 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 28244 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1688980957
transform 1 0 28428 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform -1 0 29348 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform 1 0 29532 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 30084 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 30636 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform 1 0 31188 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 31464 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 32108 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 34684 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 38364 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 37996 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output133
timestamp 1688980957
transform 1 0 38916 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output134
timestamp 1688980957
transform 1 0 39192 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 39836 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 38640 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 33488 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform 1 0 35236 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform 1 0 35788 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 35420 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 36340 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 36616 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 37260 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 36064 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 37812 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform -1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 45816 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 45816 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 45816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 45816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 45816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 45816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 45816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 45816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 45816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 45816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 45816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 45816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 45816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 45816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 25024 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform -1 0 22172 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform -1 0 23092 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform 1 0 23644 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform -1 0 22080 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform -1 0 19872 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform -1 0 17112 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform -1 0 19044 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 22172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 24748 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 29900 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 32384 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 35144 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 37628 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 39744 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 42412 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 44620 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 44896 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_outbuf_0__0_
timestamp 1688980957
transform -1 0 24196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform -1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform -1 0 23552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform -1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform -1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform -1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform -1 0 19688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 26036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 28244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 30452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 32660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform -1 0 35144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 37076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 41584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 43976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform -1 0 44896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 44896 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 37168 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 44896 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 39302 0 39358 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 42982 0 43038 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 43350 0 43406 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 43718 0 43774 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 44086 0 44142 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 44454 0 44510 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 44822 0 44878 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 45190 0 45246 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 45558 0 45614 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 45926 0 45982 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 46294 0 46350 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 39670 0 39726 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 40038 0 40094 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 40406 0 40462 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 40774 0 40830 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 41142 0 41198 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 41510 0 41566 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 41878 0 41934 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 42246 0 42302 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 42614 0 42670 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 3606 9840 3662 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 25686 9840 25742 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 27894 9840 27950 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 30102 9840 30158 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 32310 9840 32366 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 34518 9840 34574 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 36726 9840 36782 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 38934 9840 38990 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 41142 9840 41198 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 43350 9840 43406 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 45558 9840 45614 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 5814 9840 5870 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 8022 9840 8078 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 10230 9840 10286 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 12438 9840 12494 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 14646 9840 14702 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 16854 9840 16910 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 19062 9840 19118 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 21270 9840 21326 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 23478 9840 23534 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 662 0 718 160 0 FreeSans 224 90 0 0 N1END[0]
port 40 nsew signal input
flabel metal2 s 1030 0 1086 160 0 FreeSans 224 90 0 0 N1END[1]
port 41 nsew signal input
flabel metal2 s 1398 0 1454 160 0 FreeSans 224 90 0 0 N1END[2]
port 42 nsew signal input
flabel metal2 s 1766 0 1822 160 0 FreeSans 224 90 0 0 N1END[3]
port 43 nsew signal input
flabel metal2 s 5078 0 5134 160 0 FreeSans 224 90 0 0 N2END[0]
port 44 nsew signal input
flabel metal2 s 5446 0 5502 160 0 FreeSans 224 90 0 0 N2END[1]
port 45 nsew signal input
flabel metal2 s 5814 0 5870 160 0 FreeSans 224 90 0 0 N2END[2]
port 46 nsew signal input
flabel metal2 s 6182 0 6238 160 0 FreeSans 224 90 0 0 N2END[3]
port 47 nsew signal input
flabel metal2 s 6550 0 6606 160 0 FreeSans 224 90 0 0 N2END[4]
port 48 nsew signal input
flabel metal2 s 6918 0 6974 160 0 FreeSans 224 90 0 0 N2END[5]
port 49 nsew signal input
flabel metal2 s 7286 0 7342 160 0 FreeSans 224 90 0 0 N2END[6]
port 50 nsew signal input
flabel metal2 s 7654 0 7710 160 0 FreeSans 224 90 0 0 N2END[7]
port 51 nsew signal input
flabel metal2 s 2134 0 2190 160 0 FreeSans 224 90 0 0 N2MID[0]
port 52 nsew signal input
flabel metal2 s 2502 0 2558 160 0 FreeSans 224 90 0 0 N2MID[1]
port 53 nsew signal input
flabel metal2 s 2870 0 2926 160 0 FreeSans 224 90 0 0 N2MID[2]
port 54 nsew signal input
flabel metal2 s 3238 0 3294 160 0 FreeSans 224 90 0 0 N2MID[3]
port 55 nsew signal input
flabel metal2 s 3606 0 3662 160 0 FreeSans 224 90 0 0 N2MID[4]
port 56 nsew signal input
flabel metal2 s 3974 0 4030 160 0 FreeSans 224 90 0 0 N2MID[5]
port 57 nsew signal input
flabel metal2 s 4342 0 4398 160 0 FreeSans 224 90 0 0 N2MID[6]
port 58 nsew signal input
flabel metal2 s 4710 0 4766 160 0 FreeSans 224 90 0 0 N2MID[7]
port 59 nsew signal input
flabel metal2 s 8022 0 8078 160 0 FreeSans 224 90 0 0 N4END[0]
port 60 nsew signal input
flabel metal2 s 11702 0 11758 160 0 FreeSans 224 90 0 0 N4END[10]
port 61 nsew signal input
flabel metal2 s 12070 0 12126 160 0 FreeSans 224 90 0 0 N4END[11]
port 62 nsew signal input
flabel metal2 s 12438 0 12494 160 0 FreeSans 224 90 0 0 N4END[12]
port 63 nsew signal input
flabel metal2 s 12806 0 12862 160 0 FreeSans 224 90 0 0 N4END[13]
port 64 nsew signal input
flabel metal2 s 13174 0 13230 160 0 FreeSans 224 90 0 0 N4END[14]
port 65 nsew signal input
flabel metal2 s 13542 0 13598 160 0 FreeSans 224 90 0 0 N4END[15]
port 66 nsew signal input
flabel metal2 s 8390 0 8446 160 0 FreeSans 224 90 0 0 N4END[1]
port 67 nsew signal input
flabel metal2 s 8758 0 8814 160 0 FreeSans 224 90 0 0 N4END[2]
port 68 nsew signal input
flabel metal2 s 9126 0 9182 160 0 FreeSans 224 90 0 0 N4END[3]
port 69 nsew signal input
flabel metal2 s 9494 0 9550 160 0 FreeSans 224 90 0 0 N4END[4]
port 70 nsew signal input
flabel metal2 s 9862 0 9918 160 0 FreeSans 224 90 0 0 N4END[5]
port 71 nsew signal input
flabel metal2 s 10230 0 10286 160 0 FreeSans 224 90 0 0 N4END[6]
port 72 nsew signal input
flabel metal2 s 10598 0 10654 160 0 FreeSans 224 90 0 0 N4END[7]
port 73 nsew signal input
flabel metal2 s 10966 0 11022 160 0 FreeSans 224 90 0 0 N4END[8]
port 74 nsew signal input
flabel metal2 s 11334 0 11390 160 0 FreeSans 224 90 0 0 N4END[9]
port 75 nsew signal input
flabel metal2 s 13910 0 13966 160 0 FreeSans 224 90 0 0 NN4END[0]
port 76 nsew signal input
flabel metal2 s 17590 0 17646 160 0 FreeSans 224 90 0 0 NN4END[10]
port 77 nsew signal input
flabel metal2 s 17958 0 18014 160 0 FreeSans 224 90 0 0 NN4END[11]
port 78 nsew signal input
flabel metal2 s 18326 0 18382 160 0 FreeSans 224 90 0 0 NN4END[12]
port 79 nsew signal input
flabel metal2 s 18694 0 18750 160 0 FreeSans 224 90 0 0 NN4END[13]
port 80 nsew signal input
flabel metal2 s 19062 0 19118 160 0 FreeSans 224 90 0 0 NN4END[14]
port 81 nsew signal input
flabel metal2 s 19430 0 19486 160 0 FreeSans 224 90 0 0 NN4END[15]
port 82 nsew signal input
flabel metal2 s 14278 0 14334 160 0 FreeSans 224 90 0 0 NN4END[1]
port 83 nsew signal input
flabel metal2 s 14646 0 14702 160 0 FreeSans 224 90 0 0 NN4END[2]
port 84 nsew signal input
flabel metal2 s 15014 0 15070 160 0 FreeSans 224 90 0 0 NN4END[3]
port 85 nsew signal input
flabel metal2 s 15382 0 15438 160 0 FreeSans 224 90 0 0 NN4END[4]
port 86 nsew signal input
flabel metal2 s 15750 0 15806 160 0 FreeSans 224 90 0 0 NN4END[5]
port 87 nsew signal input
flabel metal2 s 16118 0 16174 160 0 FreeSans 224 90 0 0 NN4END[6]
port 88 nsew signal input
flabel metal2 s 16486 0 16542 160 0 FreeSans 224 90 0 0 NN4END[7]
port 89 nsew signal input
flabel metal2 s 16854 0 16910 160 0 FreeSans 224 90 0 0 NN4END[8]
port 90 nsew signal input
flabel metal2 s 17222 0 17278 160 0 FreeSans 224 90 0 0 NN4END[9]
port 91 nsew signal input
flabel metal2 s 19798 0 19854 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 92 nsew signal tristate
flabel metal2 s 20166 0 20222 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 93 nsew signal tristate
flabel metal2 s 20534 0 20590 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 94 nsew signal tristate
flabel metal2 s 20902 0 20958 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 95 nsew signal tristate
flabel metal2 s 24214 0 24270 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 96 nsew signal tristate
flabel metal2 s 24582 0 24638 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 97 nsew signal tristate
flabel metal2 s 24950 0 25006 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 98 nsew signal tristate
flabel metal2 s 25318 0 25374 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 99 nsew signal tristate
flabel metal2 s 25686 0 25742 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 100 nsew signal tristate
flabel metal2 s 26054 0 26110 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 101 nsew signal tristate
flabel metal2 s 26422 0 26478 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 102 nsew signal tristate
flabel metal2 s 26790 0 26846 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 103 nsew signal tristate
flabel metal2 s 21270 0 21326 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 104 nsew signal tristate
flabel metal2 s 21638 0 21694 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 105 nsew signal tristate
flabel metal2 s 22006 0 22062 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 106 nsew signal tristate
flabel metal2 s 22374 0 22430 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 107 nsew signal tristate
flabel metal2 s 22742 0 22798 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 108 nsew signal tristate
flabel metal2 s 23110 0 23166 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 109 nsew signal tristate
flabel metal2 s 23478 0 23534 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 110 nsew signal tristate
flabel metal2 s 23846 0 23902 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 111 nsew signal tristate
flabel metal2 s 27158 0 27214 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 112 nsew signal tristate
flabel metal2 s 30838 0 30894 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 113 nsew signal tristate
flabel metal2 s 31206 0 31262 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 114 nsew signal tristate
flabel metal2 s 31574 0 31630 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 115 nsew signal tristate
flabel metal2 s 31942 0 31998 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 116 nsew signal tristate
flabel metal2 s 32310 0 32366 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 117 nsew signal tristate
flabel metal2 s 32678 0 32734 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 118 nsew signal tristate
flabel metal2 s 27526 0 27582 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 119 nsew signal tristate
flabel metal2 s 27894 0 27950 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 120 nsew signal tristate
flabel metal2 s 28262 0 28318 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 121 nsew signal tristate
flabel metal2 s 28630 0 28686 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 122 nsew signal tristate
flabel metal2 s 28998 0 29054 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 123 nsew signal tristate
flabel metal2 s 29366 0 29422 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 124 nsew signal tristate
flabel metal2 s 29734 0 29790 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 125 nsew signal tristate
flabel metal2 s 30102 0 30158 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 126 nsew signal tristate
flabel metal2 s 30470 0 30526 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 127 nsew signal tristate
flabel metal2 s 33046 0 33102 160 0 FreeSans 224 90 0 0 SS4BEG[0]
port 128 nsew signal tristate
flabel metal2 s 36726 0 36782 160 0 FreeSans 224 90 0 0 SS4BEG[10]
port 129 nsew signal tristate
flabel metal2 s 37094 0 37150 160 0 FreeSans 224 90 0 0 SS4BEG[11]
port 130 nsew signal tristate
flabel metal2 s 37462 0 37518 160 0 FreeSans 224 90 0 0 SS4BEG[12]
port 131 nsew signal tristate
flabel metal2 s 37830 0 37886 160 0 FreeSans 224 90 0 0 SS4BEG[13]
port 132 nsew signal tristate
flabel metal2 s 38198 0 38254 160 0 FreeSans 224 90 0 0 SS4BEG[14]
port 133 nsew signal tristate
flabel metal2 s 38566 0 38622 160 0 FreeSans 224 90 0 0 SS4BEG[15]
port 134 nsew signal tristate
flabel metal2 s 33414 0 33470 160 0 FreeSans 224 90 0 0 SS4BEG[1]
port 135 nsew signal tristate
flabel metal2 s 33782 0 33838 160 0 FreeSans 224 90 0 0 SS4BEG[2]
port 136 nsew signal tristate
flabel metal2 s 34150 0 34206 160 0 FreeSans 224 90 0 0 SS4BEG[3]
port 137 nsew signal tristate
flabel metal2 s 34518 0 34574 160 0 FreeSans 224 90 0 0 SS4BEG[4]
port 138 nsew signal tristate
flabel metal2 s 34886 0 34942 160 0 FreeSans 224 90 0 0 SS4BEG[5]
port 139 nsew signal tristate
flabel metal2 s 35254 0 35310 160 0 FreeSans 224 90 0 0 SS4BEG[6]
port 140 nsew signal tristate
flabel metal2 s 35622 0 35678 160 0 FreeSans 224 90 0 0 SS4BEG[7]
port 141 nsew signal tristate
flabel metal2 s 35990 0 36046 160 0 FreeSans 224 90 0 0 SS4BEG[8]
port 142 nsew signal tristate
flabel metal2 s 36358 0 36414 160 0 FreeSans 224 90 0 0 SS4BEG[9]
port 143 nsew signal tristate
flabel metal2 s 38934 0 38990 160 0 FreeSans 224 90 0 0 UserCLK
port 144 nsew signal input
flabel metal2 s 1398 9840 1454 10000 0 FreeSans 224 90 0 0 UserCLKo
port 145 nsew signal tristate
flabel metal4 s 6533 1040 6853 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 17711 1040 18031 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 28889 1040 29209 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 40067 1040 40387 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 12122 1040 12442 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 23300 1040 23620 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 34478 1040 34798 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 45656 1040 45976 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
rlabel metal1 23460 8160 23460 8160 0 vccd1
rlabel via1 23540 8704 23540 8704 0 vssd1
rlabel metal2 39475 68 39475 68 0 FrameStrobe[0]
rlabel metal2 43155 68 43155 68 0 FrameStrobe[10]
rlabel metal2 43523 68 43523 68 0 FrameStrobe[11]
rlabel metal2 43891 68 43891 68 0 FrameStrobe[12]
rlabel metal2 44114 704 44114 704 0 FrameStrobe[13]
rlabel metal2 44627 68 44627 68 0 FrameStrobe[14]
rlabel metal2 44850 704 44850 704 0 FrameStrobe[15]
rlabel metal2 45218 704 45218 704 0 FrameStrobe[16]
rlabel metal2 45402 1241 45402 1241 0 FrameStrobe[17]
rlabel metal2 45494 1683 45494 1683 0 FrameStrobe[18]
rlabel metal2 46177 68 46177 68 0 FrameStrobe[19]
rlabel metal2 39698 143 39698 143 0 FrameStrobe[1]
rlabel metal2 40211 68 40211 68 0 FrameStrobe[2]
rlabel metal2 40579 68 40579 68 0 FrameStrobe[3]
rlabel metal2 40802 976 40802 976 0 FrameStrobe[4]
rlabel metal2 41446 1377 41446 1377 0 FrameStrobe[5]
rlabel metal2 41354 663 41354 663 0 FrameStrobe[6]
rlabel metal2 41906 942 41906 942 0 FrameStrobe[7]
rlabel metal2 42274 704 42274 704 0 FrameStrobe[8]
rlabel metal2 42642 704 42642 704 0 FrameStrobe[9]
rlabel metal1 3772 8602 3772 8602 0 FrameStrobe_O[0]
rlabel metal1 25806 8602 25806 8602 0 FrameStrobe_O[10]
rlabel metal1 28014 8602 28014 8602 0 FrameStrobe_O[11]
rlabel metal2 30130 9224 30130 9224 0 FrameStrobe_O[12]
rlabel metal1 32430 8602 32430 8602 0 FrameStrobe_O[13]
rlabel metal2 34546 9785 34546 9785 0 FrameStrobe_O[14]
rlabel metal1 36846 8602 36846 8602 0 FrameStrobe_O[15]
rlabel metal1 39054 8602 39054 8602 0 FrameStrobe_O[16]
rlabel metal2 41170 9224 41170 9224 0 FrameStrobe_O[17]
rlabel metal1 43470 8602 43470 8602 0 FrameStrobe_O[18]
rlabel metal2 45586 9224 45586 9224 0 FrameStrobe_O[19]
rlabel metal1 5934 8602 5934 8602 0 FrameStrobe_O[1]
rlabel metal2 8050 9224 8050 9224 0 FrameStrobe_O[2]
rlabel metal1 10350 8602 10350 8602 0 FrameStrobe_O[3]
rlabel metal2 12466 9445 12466 9445 0 FrameStrobe_O[4]
rlabel metal1 14766 8602 14766 8602 0 FrameStrobe_O[5]
rlabel metal1 16974 8602 16974 8602 0 FrameStrobe_O[6]
rlabel metal2 19090 9224 19090 9224 0 FrameStrobe_O[7]
rlabel metal1 21390 8602 21390 8602 0 FrameStrobe_O[8]
rlabel metal2 23506 9445 23506 9445 0 FrameStrobe_O[9]
rlabel metal2 25070 2210 25070 2210 0 FrameStrobe_O_i\[0\]
rlabel metal1 26266 2380 26266 2380 0 FrameStrobe_O_i\[10\]
rlabel metal1 29210 2074 29210 2074 0 FrameStrobe_O_i\[11\]
rlabel metal2 32430 2108 32430 2108 0 FrameStrobe_O_i\[12\]
rlabel metal1 33074 2414 33074 2414 0 FrameStrobe_O_i\[13\]
rlabel metal1 35052 2074 35052 2074 0 FrameStrobe_O_i\[14\]
rlabel metal1 37536 2074 37536 2074 0 FrameStrobe_O_i\[15\]
rlabel metal1 39744 2074 39744 2074 0 FrameStrobe_O_i\[16\]
rlabel metal1 42136 2074 42136 2074 0 FrameStrobe_O_i\[17\]
rlabel metal1 44436 2074 44436 2074 0 FrameStrobe_O_i\[18\]
rlabel metal2 44942 2244 44942 2244 0 FrameStrobe_O_i\[19\]
rlabel metal1 22540 2074 22540 2074 0 FrameStrobe_O_i\[1\]
rlabel metal2 23046 2244 23046 2244 0 FrameStrobe_O_i\[2\]
rlabel metal1 23736 2074 23736 2074 0 FrameStrobe_O_i\[3\]
rlabel metal1 22264 1190 22264 1190 0 FrameStrobe_O_i\[4\]
rlabel metal1 19964 2074 19964 2074 0 FrameStrobe_O_i\[5\]
rlabel metal1 17342 2074 17342 2074 0 FrameStrobe_O_i\[6\]
rlabel metal2 18998 2244 18998 2244 0 FrameStrobe_O_i\[7\]
rlabel metal1 21850 2380 21850 2380 0 FrameStrobe_O_i\[8\]
rlabel metal1 24702 2074 24702 2074 0 FrameStrobe_O_i\[9\]
rlabel metal2 690 1010 690 1010 0 N1END[0]
rlabel metal2 1058 976 1058 976 0 N1END[1]
rlabel metal2 1426 704 1426 704 0 N1END[2]
rlabel metal2 1847 68 1847 68 0 N1END[3]
rlabel metal2 5159 68 5159 68 0 N2END[0]
rlabel metal2 5527 68 5527 68 0 N2END[1]
rlabel metal2 5895 68 5895 68 0 N2END[2]
rlabel metal2 6309 68 6309 68 0 N2END[3]
rlabel metal2 6631 68 6631 68 0 N2END[4]
rlabel metal2 6999 68 6999 68 0 N2END[5]
rlabel metal2 7367 68 7367 68 0 N2END[6]
rlabel metal2 7735 68 7735 68 0 N2END[7]
rlabel metal2 2215 68 2215 68 0 N2MID[0]
rlabel metal2 2583 68 2583 68 0 N2MID[1]
rlabel metal2 2951 68 2951 68 0 N2MID[2]
rlabel metal2 3319 68 3319 68 0 N2MID[3]
rlabel metal2 3733 68 3733 68 0 N2MID[4]
rlabel metal2 4055 68 4055 68 0 N2MID[5]
rlabel metal2 4423 68 4423 68 0 N2MID[6]
rlabel metal2 4791 68 4791 68 0 N2MID[7]
rlabel metal2 8103 68 8103 68 0 N4END[0]
rlabel metal2 11783 68 11783 68 0 N4END[10]
rlabel metal2 12045 68 12045 68 0 N4END[11]
rlabel metal2 12519 68 12519 68 0 N4END[12]
rlabel metal2 12887 68 12887 68 0 N4END[13]
rlabel metal2 13255 68 13255 68 0 N4END[14]
rlabel metal2 13623 68 13623 68 0 N4END[15]
rlabel metal2 8418 670 8418 670 0 N4END[1]
rlabel metal2 8687 68 8687 68 0 N4END[2]
rlabel metal2 9207 68 9207 68 0 N4END[3]
rlabel metal2 9575 68 9575 68 0 N4END[4]
rlabel metal2 9943 68 9943 68 0 N4END[5]
rlabel metal2 10311 68 10311 68 0 N4END[6]
rlabel metal2 10679 68 10679 68 0 N4END[7]
rlabel metal2 11047 68 11047 68 0 N4END[8]
rlabel metal2 11461 68 11461 68 0 N4END[9]
rlabel metal2 14037 68 14037 68 0 NN4END[0]
rlabel metal2 17618 704 17618 704 0 NN4END[10]
rlabel metal2 17986 704 17986 704 0 NN4END[11]
rlabel metal2 18209 68 18209 68 0 NN4END[12]
rlabel metal2 18623 68 18623 68 0 NN4END[13]
rlabel metal2 19090 126 19090 126 0 NN4END[14]
rlabel metal2 19458 704 19458 704 0 NN4END[15]
rlabel metal2 14359 68 14359 68 0 NN4END[1]
rlabel metal2 14674 704 14674 704 0 NN4END[2]
rlabel metal2 14989 68 14989 68 0 NN4END[3]
rlabel metal2 15311 68 15311 68 0 NN4END[4]
rlabel metal2 15778 126 15778 126 0 NN4END[5]
rlabel metal2 16146 670 16146 670 0 NN4END[6]
rlabel metal2 16369 68 16369 68 0 NN4END[7]
rlabel metal2 16882 126 16882 126 0 NN4END[8]
rlabel metal2 17105 68 17105 68 0 NN4END[9]
rlabel metal2 19773 68 19773 68 0 S1BEG[0]
rlabel metal2 20194 347 20194 347 0 S1BEG[1]
rlabel metal2 20509 68 20509 68 0 S1BEG[2]
rlabel metal2 20930 772 20930 772 0 S1BEG[3]
rlabel metal2 24387 68 24387 68 0 S2BEG[0]
rlabel metal2 24610 347 24610 347 0 S2BEG[1]
rlabel metal2 24978 704 24978 704 0 S2BEG[2]
rlabel metal2 25346 942 25346 942 0 S2BEG[3]
rlabel metal2 25859 68 25859 68 0 S2BEG[4]
rlabel metal2 26135 68 26135 68 0 S2BEG[5]
rlabel metal2 26450 908 26450 908 0 S2BEG[6]
rlabel metal2 26963 68 26963 68 0 S2BEG[7]
rlabel metal2 21245 68 21245 68 0 S2BEGb[0]
rlabel metal2 21613 68 21613 68 0 S2BEGb[1]
rlabel metal2 21981 68 21981 68 0 S2BEGb[2]
rlabel metal2 22402 483 22402 483 0 S2BEGb[3]
rlabel metal2 22915 68 22915 68 0 S2BEGb[4]
rlabel metal2 23138 636 23138 636 0 S2BEGb[5]
rlabel metal2 23506 143 23506 143 0 S2BEGb[6]
rlabel metal2 23874 908 23874 908 0 S2BEGb[7]
rlabel metal2 27331 68 27331 68 0 S4BEG[0]
rlabel metal2 31011 68 31011 68 0 S4BEG[10]
rlabel metal2 31379 68 31379 68 0 S4BEG[11]
rlabel metal1 33442 1462 33442 1462 0 S4BEG[12]
rlabel metal2 32115 68 32115 68 0 S4BEG[13]
rlabel metal2 32483 68 32483 68 0 S4BEG[14]
rlabel metal2 32851 68 32851 68 0 S4BEG[15]
rlabel metal2 27554 755 27554 755 0 S4BEG[1]
rlabel metal2 27922 942 27922 942 0 S4BEG[2]
rlabel metal2 28290 738 28290 738 0 S4BEG[3]
rlabel metal2 28658 806 28658 806 0 S4BEG[4]
rlabel metal2 29026 772 29026 772 0 S4BEG[5]
rlabel metal2 29394 347 29394 347 0 S4BEG[6]
rlabel metal2 29907 68 29907 68 0 S4BEG[7]
rlabel metal1 31004 2822 31004 2822 0 S4BEG[8]
rlabel metal2 30498 143 30498 143 0 S4BEG[9]
rlabel metal2 33074 670 33074 670 0 SS4BEG[0]
rlabel metal2 36899 68 36899 68 0 SS4BEG[10]
rlabel metal2 37175 68 37175 68 0 SS4BEG[11]
rlabel metal2 37635 68 37635 68 0 SS4BEG[12]
rlabel metal2 37858 143 37858 143 0 SS4BEG[13]
rlabel metal2 38325 68 38325 68 0 SS4BEG[14]
rlabel metal2 38541 68 38541 68 0 SS4BEG[15]
rlabel metal2 33442 908 33442 908 0 SS4BEG[1]
rlabel metal2 33955 68 33955 68 0 SS4BEG[2]
rlabel metal2 34178 347 34178 347 0 SS4BEG[3]
rlabel metal2 34691 68 34691 68 0 SS4BEG[4]
rlabel metal2 34914 347 34914 347 0 SS4BEG[5]
rlabel metal2 35427 68 35427 68 0 SS4BEG[6]
rlabel metal2 35650 738 35650 738 0 SS4BEG[7]
rlabel metal2 36163 68 36163 68 0 SS4BEG[8]
rlabel metal2 36531 68 36531 68 0 SS4BEG[9]
rlabel metal2 39107 68 39107 68 0 UserCLK
rlabel metal2 1426 9190 1426 9190 0 UserCLKo
rlabel metal1 38916 1190 38916 1190 0 net1
rlabel metal1 44850 1904 44850 1904 0 net10
rlabel metal1 25714 1326 25714 1326 0 net100
rlabel metal1 25806 1904 25806 1904 0 net101
rlabel metal1 26082 1326 26082 1326 0 net102
rlabel metal1 26726 1326 26726 1326 0 net103
rlabel metal1 26818 1938 26818 1938 0 net104
rlabel metal1 27922 1972 27922 1972 0 net105
rlabel metal1 21022 1972 21022 1972 0 net106
rlabel metal1 20884 1326 20884 1326 0 net107
rlabel metal2 22218 1904 22218 1904 0 net108
rlabel metal1 21114 2040 21114 2040 0 net109
rlabel metal1 45218 1938 45218 1938 0 net11
rlabel metal1 22494 1326 22494 1326 0 net110
rlabel metal2 23230 1088 23230 1088 0 net111
rlabel metal1 23230 1258 23230 1258 0 net112
rlabel metal1 23966 1904 23966 1904 0 net113
rlabel metal1 27508 1326 27508 1326 0 net114
rlabel metal1 31004 2006 31004 2006 0 net115
rlabel metal1 32292 1258 32292 1258 0 net116
rlabel metal1 32844 1326 32844 1326 0 net117
rlabel metal1 32476 2006 32476 2006 0 net118
rlabel metal1 33764 1326 33764 1326 0 net119
rlabel metal2 21758 1190 21758 1190 0 net12
rlabel metal1 34178 2040 34178 2040 0 net120
rlabel metal1 28198 1326 28198 1326 0 net121
rlabel metal1 28290 1938 28290 1938 0 net122
rlabel metal1 29302 1326 29302 1326 0 net123
rlabel metal1 29486 1258 29486 1258 0 net124
rlabel metal1 29900 1326 29900 1326 0 net125
rlabel metal1 30636 1258 30636 1258 0 net126
rlabel metal1 30866 1326 30866 1326 0 net127
rlabel metal1 31602 1870 31602 1870 0 net128
rlabel metal1 32108 1326 32108 1326 0 net129
rlabel metal2 38962 1581 38962 1581 0 net13
rlabel metal2 19274 1819 19274 1819 0 net130
rlabel metal2 38180 3060 38180 3060 0 net131
rlabel metal2 15686 1785 15686 1785 0 net132
rlabel metal2 39008 3468 39008 3468 0 net133
rlabel metal1 19136 1190 19136 1190 0 net134
rlabel metal2 20286 1513 20286 1513 0 net135
rlabel metal2 20654 1853 20654 1853 0 net136
rlabel metal1 20010 1428 20010 1428 0 net137
rlabel via2 18630 1717 18630 1717 0 net138
rlabel metal2 35926 816 35926 816 0 net139
rlabel metal1 29716 3026 29716 3026 0 net14
rlabel metal1 22678 2584 22678 2584 0 net140
rlabel metal2 17526 1156 17526 1156 0 net141
rlabel metal1 17572 1802 17572 1802 0 net142
rlabel metal2 17250 1649 17250 1649 0 net143
rlabel metal1 35972 2006 35972 2006 0 net144
rlabel metal2 37674 3604 37674 3604 0 net145
rlabel metal1 10166 8568 10166 8568 0 net146
rlabel metal1 40434 2074 40434 2074 0 net15
rlabel metal1 21022 1496 21022 1496 0 net16
rlabel metal1 40342 986 40342 986 0 net17
rlabel metal2 41630 3094 41630 3094 0 net18
rlabel metal1 42458 748 42458 748 0 net19
rlabel metal2 28842 1598 28842 1598 0 net2
rlabel metal1 42734 680 42734 680 0 net20
rlabel metal2 1610 1632 1610 1632 0 net21
rlabel metal1 1886 2040 1886 2040 0 net22
rlabel metal1 1978 646 1978 646 0 net23
rlabel metal2 12650 1530 12650 1530 0 net24
rlabel metal1 21022 1870 21022 1870 0 net25
rlabel metal1 14720 3570 14720 3570 0 net26
rlabel metal2 13110 289 13110 289 0 net27
rlabel metal2 13754 1037 13754 1037 0 net28
rlabel metal3 16652 2108 16652 2108 0 net29
rlabel metal1 42504 1530 42504 1530 0 net3
rlabel metal2 14766 1496 14766 1496 0 net30
rlabel metal2 15042 1496 15042 1496 0 net31
rlabel metal1 19826 2346 19826 2346 0 net32
rlabel metal3 14950 4556 14950 4556 0 net33
rlabel metal1 14628 4182 14628 4182 0 net34
rlabel metal1 15594 4522 15594 4522 0 net35
rlabel metal3 17894 4012 17894 4012 0 net36
rlabel metal1 17848 3162 17848 3162 0 net37
rlabel metal1 15870 3026 15870 3026 0 net38
rlabel metal1 15410 578 15410 578 0 net39
rlabel metal1 43838 1224 43838 1224 0 net4
rlabel metal1 7130 578 7130 578 0 net40
rlabel metal2 11454 2927 11454 2927 0 net41
rlabel metal1 12466 1360 12466 1360 0 net42
rlabel metal1 14490 1224 14490 1224 0 net43
rlabel metal2 12742 986 12742 986 0 net44
rlabel metal1 13386 204 13386 204 0 net45
rlabel metal2 13478 782 13478 782 0 net46
rlabel metal2 13846 714 13846 714 0 net47
rlabel metal3 13524 1156 13524 1156 0 net48
rlabel metal2 8786 833 8786 833 0 net49
rlabel metal1 44068 1190 44068 1190 0 net5
rlabel metal2 9430 3264 9430 3264 0 net50
rlabel metal2 13754 2295 13754 2295 0 net51
rlabel metal2 10166 952 10166 952 0 net52
rlabel metal2 11454 1003 11454 1003 0 net53
rlabel metal2 10902 1037 10902 1037 0 net54
rlabel metal2 11270 612 11270 612 0 net55
rlabel metal2 11914 765 11914 765 0 net56
rlabel metal2 14306 1938 14306 1938 0 net57
rlabel metal1 17480 1530 17480 1530 0 net58
rlabel metal1 18032 1530 18032 1530 0 net59
rlabel metal1 44528 1190 44528 1190 0 net6
rlabel metal1 18492 1190 18492 1190 0 net60
rlabel metal1 18262 1530 18262 1530 0 net61
rlabel metal1 18584 1530 18584 1530 0 net62
rlabel metal1 19182 1530 19182 1530 0 net63
rlabel metal1 14582 1292 14582 1292 0 net64
rlabel metal1 18906 1360 18906 1360 0 net65
rlabel metal2 15134 1734 15134 1734 0 net66
rlabel metal1 15456 1530 15456 1530 0 net67
rlabel metal1 15732 1530 15732 1530 0 net68
rlabel metal1 16008 1530 16008 1530 0 net69
rlabel metal1 44666 1462 44666 1462 0 net7
rlabel metal1 16284 1530 16284 1530 0 net70
rlabel metal1 17066 1292 17066 1292 0 net71
rlabel metal1 17066 1530 17066 1530 0 net72
rlabel metal2 39514 1088 39514 1088 0 net73
rlabel metal2 6302 8602 6302 8602 0 net74
rlabel metal2 26082 5508 26082 5508 0 net75
rlabel metal2 28290 5542 28290 5542 0 net76
rlabel metal2 30452 2278 30452 2278 0 net77
rlabel metal2 32706 5542 32706 5542 0 net78
rlabel metal2 35098 5542 35098 5542 0 net79
rlabel metal1 44758 1530 44758 1530 0 net8
rlabel metal2 37030 6900 37030 6900 0 net80
rlabel metal2 39422 6900 39422 6900 0 net81
rlabel metal1 41538 2618 41538 2618 0 net82
rlabel metal1 43884 2618 43884 2618 0 net83
rlabel metal1 44988 2618 44988 2618 0 net84
rlabel metal1 6210 8874 6210 8874 0 net85
rlabel metal1 9430 8466 9430 8466 0 net86
rlabel metal1 10626 8398 10626 8398 0 net87
rlabel metal1 13846 8466 13846 8466 0 net88
rlabel metal1 20102 2312 20102 2312 0 net89
rlabel metal1 42642 1972 42642 1972 0 net9
rlabel metal1 17342 2618 17342 2618 0 net90
rlabel metal2 19642 5508 19642 5508 0 net91
rlabel metal1 21666 2346 21666 2346 0 net92
rlabel metal1 24104 2550 24104 2550 0 net93
rlabel metal1 19550 1292 19550 1292 0 net94
rlabel metal1 19918 1360 19918 1360 0 net95
rlabel metal1 20148 1326 20148 1326 0 net96
rlabel metal2 20746 1530 20746 1530 0 net97
rlabel metal1 24656 1258 24656 1258 0 net98
rlabel metal1 24058 1326 24058 1326 0 net99
<< properties >>
string FIXED_BBOX 0 0 47000 10000
<< end >>
