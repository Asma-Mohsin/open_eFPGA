magic
tech sky130A
magscale 1 2
timestamp 1733306927
<< nwell >>
rect 1066 7877 46866 8443
rect 1066 6789 46866 7355
rect 1066 5701 46866 6267
rect 1066 4613 46866 5179
rect 1066 3525 46866 4091
rect 1066 2437 46866 3003
rect 1066 1349 46866 1915
<< obsli1 >>
rect 1104 1071 46828 8721
<< obsm1 >>
rect 1104 620 46984 9988
<< metal2 >>
rect 1122 9840 1178 10000
rect 1490 9840 1546 10000
rect 1858 9840 1914 10000
rect 2226 9840 2282 10000
rect 2594 9840 2650 10000
rect 2962 9840 3018 10000
rect 3330 9840 3386 10000
rect 3698 9840 3754 10000
rect 4066 9840 4122 10000
rect 4434 9840 4490 10000
rect 4802 9840 4858 10000
rect 5170 9840 5226 10000
rect 5538 9840 5594 10000
rect 5906 9840 5962 10000
rect 6274 9840 6330 10000
rect 6642 9840 6698 10000
rect 7010 9840 7066 10000
rect 7378 9840 7434 10000
rect 7746 9840 7802 10000
rect 8114 9840 8170 10000
rect 8482 9840 8538 10000
rect 8850 9840 8906 10000
rect 9218 9840 9274 10000
rect 9586 9840 9642 10000
rect 9954 9840 10010 10000
rect 10322 9840 10378 10000
rect 10690 9840 10746 10000
rect 11058 9840 11114 10000
rect 11426 9840 11482 10000
rect 11794 9840 11850 10000
rect 12162 9840 12218 10000
rect 12530 9840 12586 10000
rect 12898 9840 12954 10000
rect 13266 9840 13322 10000
rect 13634 9840 13690 10000
rect 14002 9840 14058 10000
rect 14370 9840 14426 10000
rect 14738 9840 14794 10000
rect 15106 9840 15162 10000
rect 15474 9840 15530 10000
rect 15842 9840 15898 10000
rect 16210 9840 16266 10000
rect 16578 9840 16634 10000
rect 16946 9840 17002 10000
rect 17314 9840 17370 10000
rect 17682 9840 17738 10000
rect 18050 9840 18106 10000
rect 18418 9840 18474 10000
rect 18786 9840 18842 10000
rect 19154 9840 19210 10000
rect 19522 9840 19578 10000
rect 19890 9840 19946 10000
rect 20258 9840 20314 10000
rect 20626 9840 20682 10000
rect 20994 9840 21050 10000
rect 21362 9840 21418 10000
rect 21730 9840 21786 10000
rect 22098 9840 22154 10000
rect 22466 9840 22522 10000
rect 22834 9840 22890 10000
rect 23202 9840 23258 10000
rect 23570 9840 23626 10000
rect 23938 9840 23994 10000
rect 24306 9840 24362 10000
rect 24674 9840 24730 10000
rect 25042 9840 25098 10000
rect 25410 9840 25466 10000
rect 25778 9840 25834 10000
rect 26146 9840 26202 10000
rect 26514 9840 26570 10000
rect 26882 9840 26938 10000
rect 27250 9840 27306 10000
rect 27618 9840 27674 10000
rect 27986 9840 28042 10000
rect 28354 9840 28410 10000
rect 28722 9840 28778 10000
rect 29090 9840 29146 10000
rect 29458 9840 29514 10000
rect 29826 9840 29882 10000
rect 30194 9840 30250 10000
rect 30562 9840 30618 10000
rect 30930 9840 30986 10000
rect 31298 9840 31354 10000
rect 31666 9840 31722 10000
rect 32034 9840 32090 10000
rect 32402 9840 32458 10000
rect 32770 9840 32826 10000
rect 33138 9840 33194 10000
rect 33506 9840 33562 10000
rect 33874 9840 33930 10000
rect 34242 9840 34298 10000
rect 34610 9840 34666 10000
rect 34978 9840 35034 10000
rect 35346 9840 35402 10000
rect 35714 9840 35770 10000
rect 36082 9840 36138 10000
rect 36450 9840 36506 10000
rect 36818 9840 36874 10000
rect 37186 9840 37242 10000
rect 37554 9840 37610 10000
rect 37922 9840 37978 10000
rect 38290 9840 38346 10000
rect 38658 9840 38714 10000
rect 39026 9840 39082 10000
rect 39394 9840 39450 10000
rect 39762 9840 39818 10000
rect 40130 9840 40186 10000
rect 40498 9840 40554 10000
rect 40866 9840 40922 10000
rect 41234 9840 41290 10000
rect 41602 9840 41658 10000
rect 41970 9840 42026 10000
rect 42338 9840 42394 10000
rect 42706 9840 42762 10000
rect 43074 9840 43130 10000
rect 43442 9840 43498 10000
rect 43810 9840 43866 10000
rect 44178 9840 44234 10000
rect 44546 9840 44602 10000
rect 44914 9840 44970 10000
rect 45282 9840 45338 10000
rect 45650 9840 45706 10000
rect 46018 9840 46074 10000
rect 46386 9840 46442 10000
rect 46754 9840 46810 10000
rect 1858 0 1914 160
rect 4066 0 4122 160
rect 6274 0 6330 160
rect 8482 0 8538 160
rect 10690 0 10746 160
rect 12898 0 12954 160
rect 15106 0 15162 160
rect 17314 0 17370 160
rect 19522 0 19578 160
rect 21730 0 21786 160
rect 23938 0 23994 160
rect 26146 0 26202 160
rect 28354 0 28410 160
rect 30562 0 30618 160
rect 32770 0 32826 160
rect 34978 0 35034 160
rect 37186 0 37242 160
rect 39394 0 39450 160
rect 41602 0 41658 160
rect 43810 0 43866 160
rect 46018 0 46074 160
<< obsm2 >>
rect 1234 9784 1434 9994
rect 1602 9784 1802 9994
rect 1970 9784 2170 9994
rect 2338 9784 2538 9994
rect 2706 9784 2906 9994
rect 3074 9784 3274 9994
rect 3442 9784 3642 9994
rect 3810 9784 4010 9994
rect 4178 9784 4378 9994
rect 4546 9784 4746 9994
rect 4914 9784 5114 9994
rect 5282 9784 5482 9994
rect 5650 9784 5850 9994
rect 6018 9784 6218 9994
rect 6386 9784 6586 9994
rect 6754 9784 6954 9994
rect 7122 9784 7322 9994
rect 7490 9784 7690 9994
rect 7858 9784 8058 9994
rect 8226 9784 8426 9994
rect 8594 9784 8794 9994
rect 8962 9784 9162 9994
rect 9330 9784 9530 9994
rect 9698 9784 9898 9994
rect 10066 9784 10266 9994
rect 10434 9784 10634 9994
rect 10802 9784 11002 9994
rect 11170 9784 11370 9994
rect 11538 9784 11738 9994
rect 11906 9784 12106 9994
rect 12274 9784 12474 9994
rect 12642 9784 12842 9994
rect 13010 9784 13210 9994
rect 13378 9784 13578 9994
rect 13746 9784 13946 9994
rect 14114 9784 14314 9994
rect 14482 9784 14682 9994
rect 14850 9784 15050 9994
rect 15218 9784 15418 9994
rect 15586 9784 15786 9994
rect 15954 9784 16154 9994
rect 16322 9784 16522 9994
rect 16690 9784 16890 9994
rect 17058 9784 17258 9994
rect 17426 9784 17626 9994
rect 17794 9784 17994 9994
rect 18162 9784 18362 9994
rect 18530 9784 18730 9994
rect 18898 9784 19098 9994
rect 19266 9784 19466 9994
rect 19634 9784 19834 9994
rect 20002 9784 20202 9994
rect 20370 9784 20570 9994
rect 20738 9784 20938 9994
rect 21106 9784 21306 9994
rect 21474 9784 21674 9994
rect 21842 9784 22042 9994
rect 22210 9784 22410 9994
rect 22578 9784 22778 9994
rect 22946 9784 23146 9994
rect 23314 9784 23514 9994
rect 23682 9784 23882 9994
rect 24050 9784 24250 9994
rect 24418 9784 24618 9994
rect 24786 9784 24986 9994
rect 25154 9784 25354 9994
rect 25522 9784 25722 9994
rect 25890 9784 26090 9994
rect 26258 9784 26458 9994
rect 26626 9784 26826 9994
rect 26994 9784 27194 9994
rect 27362 9784 27562 9994
rect 27730 9784 27930 9994
rect 28098 9784 28298 9994
rect 28466 9784 28666 9994
rect 28834 9784 29034 9994
rect 29202 9784 29402 9994
rect 29570 9784 29770 9994
rect 29938 9784 30138 9994
rect 30306 9784 30506 9994
rect 30674 9784 30874 9994
rect 31042 9784 31242 9994
rect 31410 9784 31610 9994
rect 31778 9784 31978 9994
rect 32146 9784 32346 9994
rect 32514 9784 32714 9994
rect 32882 9784 33082 9994
rect 33250 9784 33450 9994
rect 33618 9784 33818 9994
rect 33986 9784 34186 9994
rect 34354 9784 34554 9994
rect 34722 9784 34922 9994
rect 35090 9784 35290 9994
rect 35458 9784 35658 9994
rect 35826 9784 36026 9994
rect 36194 9784 36394 9994
rect 36562 9784 36762 9994
rect 36930 9784 37130 9994
rect 37298 9784 37498 9994
rect 37666 9784 37866 9994
rect 38034 9784 38234 9994
rect 38402 9784 38602 9994
rect 38770 9784 38970 9994
rect 39138 9784 39338 9994
rect 39506 9784 39706 9994
rect 39874 9784 40074 9994
rect 40242 9784 40442 9994
rect 40610 9784 40810 9994
rect 40978 9784 41178 9994
rect 41346 9784 41546 9994
rect 41714 9784 41914 9994
rect 42082 9784 42282 9994
rect 42450 9784 42650 9994
rect 42818 9784 43018 9994
rect 43186 9784 43386 9994
rect 43554 9784 43754 9994
rect 43922 9784 44122 9994
rect 44290 9784 44490 9994
rect 44658 9784 44858 9994
rect 45026 9784 45226 9994
rect 45394 9784 45594 9994
rect 45762 9784 45962 9994
rect 46130 9784 46330 9994
rect 46498 9784 46698 9994
rect 46866 9784 46978 9994
rect 1124 216 46978 9784
rect 1124 54 1802 216
rect 1970 54 4010 216
rect 4178 54 6218 216
rect 6386 54 8426 216
rect 8594 54 10634 216
rect 10802 54 12842 216
rect 13010 54 15050 216
rect 15218 54 17258 216
rect 17426 54 19466 216
rect 19634 54 21674 216
rect 21842 54 23882 216
rect 24050 54 26090 216
rect 26258 54 28298 216
rect 28466 54 30506 216
rect 30674 54 32714 216
rect 32882 54 34922 216
rect 35090 54 37130 216
rect 37298 54 39338 216
rect 39506 54 41546 216
rect 41714 54 43754 216
rect 43922 54 45962 216
rect 46130 54 46978 216
<< obsm3 >>
rect 2313 1055 46982 9890
<< metal4 >>
rect 6659 1040 6979 8752
rect 12374 1040 12694 8752
rect 18089 1040 18409 8752
rect 23804 1040 24124 8752
rect 29519 1040 29839 8752
rect 35234 1040 35554 8752
rect 40949 1040 41269 8752
rect 46664 1040 46984 8752
<< labels >>
rlabel metal2 s 4066 0 4122 160 6 FrameStrobe[0]
port 1 nsew signal input
rlabel metal2 s 26146 0 26202 160 6 FrameStrobe[10]
port 2 nsew signal input
rlabel metal2 s 28354 0 28410 160 6 FrameStrobe[11]
port 3 nsew signal input
rlabel metal2 s 30562 0 30618 160 6 FrameStrobe[12]
port 4 nsew signal input
rlabel metal2 s 32770 0 32826 160 6 FrameStrobe[13]
port 5 nsew signal input
rlabel metal2 s 34978 0 35034 160 6 FrameStrobe[14]
port 6 nsew signal input
rlabel metal2 s 37186 0 37242 160 6 FrameStrobe[15]
port 7 nsew signal input
rlabel metal2 s 39394 0 39450 160 6 FrameStrobe[16]
port 8 nsew signal input
rlabel metal2 s 41602 0 41658 160 6 FrameStrobe[17]
port 9 nsew signal input
rlabel metal2 s 43810 0 43866 160 6 FrameStrobe[18]
port 10 nsew signal input
rlabel metal2 s 46018 0 46074 160 6 FrameStrobe[19]
port 11 nsew signal input
rlabel metal2 s 6274 0 6330 160 6 FrameStrobe[1]
port 12 nsew signal input
rlabel metal2 s 8482 0 8538 160 6 FrameStrobe[2]
port 13 nsew signal input
rlabel metal2 s 10690 0 10746 160 6 FrameStrobe[3]
port 14 nsew signal input
rlabel metal2 s 12898 0 12954 160 6 FrameStrobe[4]
port 15 nsew signal input
rlabel metal2 s 15106 0 15162 160 6 FrameStrobe[5]
port 16 nsew signal input
rlabel metal2 s 17314 0 17370 160 6 FrameStrobe[6]
port 17 nsew signal input
rlabel metal2 s 19522 0 19578 160 6 FrameStrobe[7]
port 18 nsew signal input
rlabel metal2 s 21730 0 21786 160 6 FrameStrobe[8]
port 19 nsew signal input
rlabel metal2 s 23938 0 23994 160 6 FrameStrobe[9]
port 20 nsew signal input
rlabel metal2 s 39762 9840 39818 10000 6 FrameStrobe_O[0]
port 21 nsew signal output
rlabel metal2 s 43442 9840 43498 10000 6 FrameStrobe_O[10]
port 22 nsew signal output
rlabel metal2 s 43810 9840 43866 10000 6 FrameStrobe_O[11]
port 23 nsew signal output
rlabel metal2 s 44178 9840 44234 10000 6 FrameStrobe_O[12]
port 24 nsew signal output
rlabel metal2 s 44546 9840 44602 10000 6 FrameStrobe_O[13]
port 25 nsew signal output
rlabel metal2 s 44914 9840 44970 10000 6 FrameStrobe_O[14]
port 26 nsew signal output
rlabel metal2 s 45282 9840 45338 10000 6 FrameStrobe_O[15]
port 27 nsew signal output
rlabel metal2 s 45650 9840 45706 10000 6 FrameStrobe_O[16]
port 28 nsew signal output
rlabel metal2 s 46018 9840 46074 10000 6 FrameStrobe_O[17]
port 29 nsew signal output
rlabel metal2 s 46386 9840 46442 10000 6 FrameStrobe_O[18]
port 30 nsew signal output
rlabel metal2 s 46754 9840 46810 10000 6 FrameStrobe_O[19]
port 31 nsew signal output
rlabel metal2 s 40130 9840 40186 10000 6 FrameStrobe_O[1]
port 32 nsew signal output
rlabel metal2 s 40498 9840 40554 10000 6 FrameStrobe_O[2]
port 33 nsew signal output
rlabel metal2 s 40866 9840 40922 10000 6 FrameStrobe_O[3]
port 34 nsew signal output
rlabel metal2 s 41234 9840 41290 10000 6 FrameStrobe_O[4]
port 35 nsew signal output
rlabel metal2 s 41602 9840 41658 10000 6 FrameStrobe_O[5]
port 36 nsew signal output
rlabel metal2 s 41970 9840 42026 10000 6 FrameStrobe_O[6]
port 37 nsew signal output
rlabel metal2 s 42338 9840 42394 10000 6 FrameStrobe_O[7]
port 38 nsew signal output
rlabel metal2 s 42706 9840 42762 10000 6 FrameStrobe_O[8]
port 39 nsew signal output
rlabel metal2 s 43074 9840 43130 10000 6 FrameStrobe_O[9]
port 40 nsew signal output
rlabel metal2 s 1122 9840 1178 10000 6 N1BEG[0]
port 41 nsew signal output
rlabel metal2 s 1490 9840 1546 10000 6 N1BEG[1]
port 42 nsew signal output
rlabel metal2 s 1858 9840 1914 10000 6 N1BEG[2]
port 43 nsew signal output
rlabel metal2 s 2226 9840 2282 10000 6 N1BEG[3]
port 44 nsew signal output
rlabel metal2 s 2594 9840 2650 10000 6 N2BEG[0]
port 45 nsew signal output
rlabel metal2 s 2962 9840 3018 10000 6 N2BEG[1]
port 46 nsew signal output
rlabel metal2 s 3330 9840 3386 10000 6 N2BEG[2]
port 47 nsew signal output
rlabel metal2 s 3698 9840 3754 10000 6 N2BEG[3]
port 48 nsew signal output
rlabel metal2 s 4066 9840 4122 10000 6 N2BEG[4]
port 49 nsew signal output
rlabel metal2 s 4434 9840 4490 10000 6 N2BEG[5]
port 50 nsew signal output
rlabel metal2 s 4802 9840 4858 10000 6 N2BEG[6]
port 51 nsew signal output
rlabel metal2 s 5170 9840 5226 10000 6 N2BEG[7]
port 52 nsew signal output
rlabel metal2 s 5538 9840 5594 10000 6 N2BEGb[0]
port 53 nsew signal output
rlabel metal2 s 5906 9840 5962 10000 6 N2BEGb[1]
port 54 nsew signal output
rlabel metal2 s 6274 9840 6330 10000 6 N2BEGb[2]
port 55 nsew signal output
rlabel metal2 s 6642 9840 6698 10000 6 N2BEGb[3]
port 56 nsew signal output
rlabel metal2 s 7010 9840 7066 10000 6 N2BEGb[4]
port 57 nsew signal output
rlabel metal2 s 7378 9840 7434 10000 6 N2BEGb[5]
port 58 nsew signal output
rlabel metal2 s 7746 9840 7802 10000 6 N2BEGb[6]
port 59 nsew signal output
rlabel metal2 s 8114 9840 8170 10000 6 N2BEGb[7]
port 60 nsew signal output
rlabel metal2 s 8482 9840 8538 10000 6 N4BEG[0]
port 61 nsew signal output
rlabel metal2 s 12162 9840 12218 10000 6 N4BEG[10]
port 62 nsew signal output
rlabel metal2 s 12530 9840 12586 10000 6 N4BEG[11]
port 63 nsew signal output
rlabel metal2 s 12898 9840 12954 10000 6 N4BEG[12]
port 64 nsew signal output
rlabel metal2 s 13266 9840 13322 10000 6 N4BEG[13]
port 65 nsew signal output
rlabel metal2 s 13634 9840 13690 10000 6 N4BEG[14]
port 66 nsew signal output
rlabel metal2 s 14002 9840 14058 10000 6 N4BEG[15]
port 67 nsew signal output
rlabel metal2 s 8850 9840 8906 10000 6 N4BEG[1]
port 68 nsew signal output
rlabel metal2 s 9218 9840 9274 10000 6 N4BEG[2]
port 69 nsew signal output
rlabel metal2 s 9586 9840 9642 10000 6 N4BEG[3]
port 70 nsew signal output
rlabel metal2 s 9954 9840 10010 10000 6 N4BEG[4]
port 71 nsew signal output
rlabel metal2 s 10322 9840 10378 10000 6 N4BEG[5]
port 72 nsew signal output
rlabel metal2 s 10690 9840 10746 10000 6 N4BEG[6]
port 73 nsew signal output
rlabel metal2 s 11058 9840 11114 10000 6 N4BEG[7]
port 74 nsew signal output
rlabel metal2 s 11426 9840 11482 10000 6 N4BEG[8]
port 75 nsew signal output
rlabel metal2 s 11794 9840 11850 10000 6 N4BEG[9]
port 76 nsew signal output
rlabel metal2 s 14370 9840 14426 10000 6 NN4BEG[0]
port 77 nsew signal output
rlabel metal2 s 18050 9840 18106 10000 6 NN4BEG[10]
port 78 nsew signal output
rlabel metal2 s 18418 9840 18474 10000 6 NN4BEG[11]
port 79 nsew signal output
rlabel metal2 s 18786 9840 18842 10000 6 NN4BEG[12]
port 80 nsew signal output
rlabel metal2 s 19154 9840 19210 10000 6 NN4BEG[13]
port 81 nsew signal output
rlabel metal2 s 19522 9840 19578 10000 6 NN4BEG[14]
port 82 nsew signal output
rlabel metal2 s 19890 9840 19946 10000 6 NN4BEG[15]
port 83 nsew signal output
rlabel metal2 s 14738 9840 14794 10000 6 NN4BEG[1]
port 84 nsew signal output
rlabel metal2 s 15106 9840 15162 10000 6 NN4BEG[2]
port 85 nsew signal output
rlabel metal2 s 15474 9840 15530 10000 6 NN4BEG[3]
port 86 nsew signal output
rlabel metal2 s 15842 9840 15898 10000 6 NN4BEG[4]
port 87 nsew signal output
rlabel metal2 s 16210 9840 16266 10000 6 NN4BEG[5]
port 88 nsew signal output
rlabel metal2 s 16578 9840 16634 10000 6 NN4BEG[6]
port 89 nsew signal output
rlabel metal2 s 16946 9840 17002 10000 6 NN4BEG[7]
port 90 nsew signal output
rlabel metal2 s 17314 9840 17370 10000 6 NN4BEG[8]
port 91 nsew signal output
rlabel metal2 s 17682 9840 17738 10000 6 NN4BEG[9]
port 92 nsew signal output
rlabel metal2 s 20258 9840 20314 10000 6 S1END[0]
port 93 nsew signal input
rlabel metal2 s 20626 9840 20682 10000 6 S1END[1]
port 94 nsew signal input
rlabel metal2 s 20994 9840 21050 10000 6 S1END[2]
port 95 nsew signal input
rlabel metal2 s 21362 9840 21418 10000 6 S1END[3]
port 96 nsew signal input
rlabel metal2 s 21730 9840 21786 10000 6 S2END[0]
port 97 nsew signal input
rlabel metal2 s 22098 9840 22154 10000 6 S2END[1]
port 98 nsew signal input
rlabel metal2 s 22466 9840 22522 10000 6 S2END[2]
port 99 nsew signal input
rlabel metal2 s 22834 9840 22890 10000 6 S2END[3]
port 100 nsew signal input
rlabel metal2 s 23202 9840 23258 10000 6 S2END[4]
port 101 nsew signal input
rlabel metal2 s 23570 9840 23626 10000 6 S2END[5]
port 102 nsew signal input
rlabel metal2 s 23938 9840 23994 10000 6 S2END[6]
port 103 nsew signal input
rlabel metal2 s 24306 9840 24362 10000 6 S2END[7]
port 104 nsew signal input
rlabel metal2 s 24674 9840 24730 10000 6 S2MID[0]
port 105 nsew signal input
rlabel metal2 s 25042 9840 25098 10000 6 S2MID[1]
port 106 nsew signal input
rlabel metal2 s 25410 9840 25466 10000 6 S2MID[2]
port 107 nsew signal input
rlabel metal2 s 25778 9840 25834 10000 6 S2MID[3]
port 108 nsew signal input
rlabel metal2 s 26146 9840 26202 10000 6 S2MID[4]
port 109 nsew signal input
rlabel metal2 s 26514 9840 26570 10000 6 S2MID[5]
port 110 nsew signal input
rlabel metal2 s 26882 9840 26938 10000 6 S2MID[6]
port 111 nsew signal input
rlabel metal2 s 27250 9840 27306 10000 6 S2MID[7]
port 112 nsew signal input
rlabel metal2 s 27618 9840 27674 10000 6 S4END[0]
port 113 nsew signal input
rlabel metal2 s 31298 9840 31354 10000 6 S4END[10]
port 114 nsew signal input
rlabel metal2 s 31666 9840 31722 10000 6 S4END[11]
port 115 nsew signal input
rlabel metal2 s 32034 9840 32090 10000 6 S4END[12]
port 116 nsew signal input
rlabel metal2 s 32402 9840 32458 10000 6 S4END[13]
port 117 nsew signal input
rlabel metal2 s 32770 9840 32826 10000 6 S4END[14]
port 118 nsew signal input
rlabel metal2 s 33138 9840 33194 10000 6 S4END[15]
port 119 nsew signal input
rlabel metal2 s 27986 9840 28042 10000 6 S4END[1]
port 120 nsew signal input
rlabel metal2 s 28354 9840 28410 10000 6 S4END[2]
port 121 nsew signal input
rlabel metal2 s 28722 9840 28778 10000 6 S4END[3]
port 122 nsew signal input
rlabel metal2 s 29090 9840 29146 10000 6 S4END[4]
port 123 nsew signal input
rlabel metal2 s 29458 9840 29514 10000 6 S4END[5]
port 124 nsew signal input
rlabel metal2 s 29826 9840 29882 10000 6 S4END[6]
port 125 nsew signal input
rlabel metal2 s 30194 9840 30250 10000 6 S4END[7]
port 126 nsew signal input
rlabel metal2 s 30562 9840 30618 10000 6 S4END[8]
port 127 nsew signal input
rlabel metal2 s 30930 9840 30986 10000 6 S4END[9]
port 128 nsew signal input
rlabel metal2 s 33506 9840 33562 10000 6 SS4END[0]
port 129 nsew signal input
rlabel metal2 s 37186 9840 37242 10000 6 SS4END[10]
port 130 nsew signal input
rlabel metal2 s 37554 9840 37610 10000 6 SS4END[11]
port 131 nsew signal input
rlabel metal2 s 37922 9840 37978 10000 6 SS4END[12]
port 132 nsew signal input
rlabel metal2 s 38290 9840 38346 10000 6 SS4END[13]
port 133 nsew signal input
rlabel metal2 s 38658 9840 38714 10000 6 SS4END[14]
port 134 nsew signal input
rlabel metal2 s 39026 9840 39082 10000 6 SS4END[15]
port 135 nsew signal input
rlabel metal2 s 33874 9840 33930 10000 6 SS4END[1]
port 136 nsew signal input
rlabel metal2 s 34242 9840 34298 10000 6 SS4END[2]
port 137 nsew signal input
rlabel metal2 s 34610 9840 34666 10000 6 SS4END[3]
port 138 nsew signal input
rlabel metal2 s 34978 9840 35034 10000 6 SS4END[4]
port 139 nsew signal input
rlabel metal2 s 35346 9840 35402 10000 6 SS4END[5]
port 140 nsew signal input
rlabel metal2 s 35714 9840 35770 10000 6 SS4END[6]
port 141 nsew signal input
rlabel metal2 s 36082 9840 36138 10000 6 SS4END[7]
port 142 nsew signal input
rlabel metal2 s 36450 9840 36506 10000 6 SS4END[8]
port 143 nsew signal input
rlabel metal2 s 36818 9840 36874 10000 6 SS4END[9]
port 144 nsew signal input
rlabel metal2 s 1858 0 1914 160 6 UserCLK
port 145 nsew signal input
rlabel metal2 s 39394 9840 39450 10000 6 UserCLKo
port 146 nsew signal output
rlabel metal4 s 6659 1040 6979 8752 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 18089 1040 18409 8752 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 29519 1040 29839 8752 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 40949 1040 41269 8752 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 12374 1040 12694 8752 6 vssd1
port 148 nsew ground bidirectional
rlabel metal4 s 23804 1040 24124 8752 6 vssd1
port 148 nsew ground bidirectional
rlabel metal4 s 35234 1040 35554 8752 6 vssd1
port 148 nsew ground bidirectional
rlabel metal4 s 46664 1040 46984 8752 6 vssd1
port 148 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 48000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 591154
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/S_term_single2/runs/24_12_04_10_07/results/signoff/S_term_single2.magic.gds
string GDS_START 42478
<< end >>

