magic
tech sky130A
magscale 1 2
timestamp 1733242054
<< obsli1 >>
rect 1104 1071 24840 43537
<< obsm1 >>
rect 14 348 25930 44940
<< metal2 >>
rect 202 44840 258 45000
rect 478 44840 534 45000
rect 754 44840 810 45000
rect 1030 44840 1086 45000
rect 1306 44840 1362 45000
rect 1582 44840 1638 45000
rect 1858 44840 1914 45000
rect 2134 44840 2190 45000
rect 2410 44840 2466 45000
rect 2686 44840 2742 45000
rect 2962 44840 3018 45000
rect 3238 44840 3294 45000
rect 3514 44840 3570 45000
rect 3790 44840 3846 45000
rect 4066 44840 4122 45000
rect 4342 44840 4398 45000
rect 4618 44840 4674 45000
rect 4894 44840 4950 45000
rect 5170 44840 5226 45000
rect 5446 44840 5502 45000
rect 5722 44840 5778 45000
rect 5998 44840 6054 45000
rect 6274 44840 6330 45000
rect 6550 44840 6606 45000
rect 6826 44840 6882 45000
rect 7102 44840 7158 45000
rect 7378 44840 7434 45000
rect 7654 44840 7710 45000
rect 7930 44840 7986 45000
rect 8206 44840 8262 45000
rect 8482 44840 8538 45000
rect 8758 44840 8814 45000
rect 9034 44840 9090 45000
rect 9310 44840 9366 45000
rect 9586 44840 9642 45000
rect 9862 44840 9918 45000
rect 10138 44840 10194 45000
rect 10414 44840 10470 45000
rect 10690 44840 10746 45000
rect 10966 44840 11022 45000
rect 11242 44840 11298 45000
rect 11518 44840 11574 45000
rect 11794 44840 11850 45000
rect 12070 44840 12126 45000
rect 12346 44840 12402 45000
rect 12622 44840 12678 45000
rect 12898 44840 12954 45000
rect 13174 44840 13230 45000
rect 13450 44840 13506 45000
rect 13726 44840 13782 45000
rect 14002 44840 14058 45000
rect 14278 44840 14334 45000
rect 14554 44840 14610 45000
rect 14830 44840 14886 45000
rect 15106 44840 15162 45000
rect 15382 44840 15438 45000
rect 15658 44840 15714 45000
rect 15934 44840 15990 45000
rect 16210 44840 16266 45000
rect 16486 44840 16542 45000
rect 16762 44840 16818 45000
rect 17038 44840 17094 45000
rect 17314 44840 17370 45000
rect 17590 44840 17646 45000
rect 17866 44840 17922 45000
rect 18142 44840 18198 45000
rect 18418 44840 18474 45000
rect 18694 44840 18750 45000
rect 18970 44840 19026 45000
rect 19246 44840 19302 45000
rect 19522 44840 19578 45000
rect 19798 44840 19854 45000
rect 20074 44840 20130 45000
rect 20350 44840 20406 45000
rect 20626 44840 20682 45000
rect 20902 44840 20958 45000
rect 21178 44840 21234 45000
rect 21454 44840 21510 45000
rect 21730 44840 21786 45000
rect 22006 44840 22062 45000
rect 22282 44840 22338 45000
rect 22558 44840 22614 45000
rect 22834 44840 22890 45000
rect 23110 44840 23166 45000
rect 23386 44840 23442 45000
rect 23662 44840 23718 45000
rect 23938 44840 23994 45000
rect 24214 44840 24270 45000
rect 24490 44840 24546 45000
rect 24766 44840 24822 45000
rect 25042 44840 25098 45000
rect 25318 44840 25374 45000
rect 25594 44840 25650 45000
rect 202 0 258 160
rect 478 0 534 160
rect 754 0 810 160
rect 1030 0 1086 160
rect 1306 0 1362 160
rect 1582 0 1638 160
rect 1858 0 1914 160
rect 2134 0 2190 160
rect 2410 0 2466 160
rect 2686 0 2742 160
rect 2962 0 3018 160
rect 3238 0 3294 160
rect 3514 0 3570 160
rect 3790 0 3846 160
rect 4066 0 4122 160
rect 4342 0 4398 160
rect 4618 0 4674 160
rect 4894 0 4950 160
rect 5170 0 5226 160
rect 5446 0 5502 160
rect 5722 0 5778 160
rect 5998 0 6054 160
rect 6274 0 6330 160
rect 6550 0 6606 160
rect 6826 0 6882 160
rect 7102 0 7158 160
rect 7378 0 7434 160
rect 7654 0 7710 160
rect 7930 0 7986 160
rect 8206 0 8262 160
rect 8482 0 8538 160
rect 8758 0 8814 160
rect 9034 0 9090 160
rect 9310 0 9366 160
rect 9586 0 9642 160
rect 9862 0 9918 160
rect 10138 0 10194 160
rect 10414 0 10470 160
rect 10690 0 10746 160
rect 10966 0 11022 160
rect 11242 0 11298 160
rect 11518 0 11574 160
rect 11794 0 11850 160
rect 12070 0 12126 160
rect 12346 0 12402 160
rect 12622 0 12678 160
rect 12898 0 12954 160
rect 13174 0 13230 160
rect 13450 0 13506 160
rect 13726 0 13782 160
rect 14002 0 14058 160
rect 14278 0 14334 160
rect 14554 0 14610 160
rect 14830 0 14886 160
rect 15106 0 15162 160
rect 15382 0 15438 160
rect 15658 0 15714 160
rect 15934 0 15990 160
rect 16210 0 16266 160
rect 16486 0 16542 160
rect 16762 0 16818 160
rect 17038 0 17094 160
rect 17314 0 17370 160
rect 17590 0 17646 160
rect 17866 0 17922 160
rect 18142 0 18198 160
rect 18418 0 18474 160
rect 18694 0 18750 160
rect 18970 0 19026 160
rect 19246 0 19302 160
rect 19522 0 19578 160
rect 19798 0 19854 160
rect 20074 0 20130 160
rect 20350 0 20406 160
rect 20626 0 20682 160
rect 20902 0 20958 160
rect 21178 0 21234 160
rect 21454 0 21510 160
rect 21730 0 21786 160
rect 22006 0 22062 160
rect 22282 0 22338 160
rect 22558 0 22614 160
rect 22834 0 22890 160
rect 23110 0 23166 160
rect 23386 0 23442 160
rect 23662 0 23718 160
rect 23938 0 23994 160
rect 24214 0 24270 160
rect 24490 0 24546 160
rect 24766 0 24822 160
rect 25042 0 25098 160
rect 25318 0 25374 160
rect 25594 0 25650 160
<< obsm2 >>
rect 18 44784 146 44962
rect 314 44784 422 44962
rect 590 44784 698 44962
rect 866 44784 974 44962
rect 1142 44784 1250 44962
rect 1418 44784 1526 44962
rect 1694 44784 1802 44962
rect 1970 44784 2078 44962
rect 2246 44784 2354 44962
rect 2522 44784 2630 44962
rect 2798 44784 2906 44962
rect 3074 44784 3182 44962
rect 3350 44784 3458 44962
rect 3626 44784 3734 44962
rect 3902 44784 4010 44962
rect 4178 44784 4286 44962
rect 4454 44784 4562 44962
rect 4730 44784 4838 44962
rect 5006 44784 5114 44962
rect 5282 44784 5390 44962
rect 5558 44784 5666 44962
rect 5834 44784 5942 44962
rect 6110 44784 6218 44962
rect 6386 44784 6494 44962
rect 6662 44784 6770 44962
rect 6938 44784 7046 44962
rect 7214 44784 7322 44962
rect 7490 44784 7598 44962
rect 7766 44784 7874 44962
rect 8042 44784 8150 44962
rect 8318 44784 8426 44962
rect 8594 44784 8702 44962
rect 8870 44784 8978 44962
rect 9146 44784 9254 44962
rect 9422 44784 9530 44962
rect 9698 44784 9806 44962
rect 9974 44784 10082 44962
rect 10250 44784 10358 44962
rect 10526 44784 10634 44962
rect 10802 44784 10910 44962
rect 11078 44784 11186 44962
rect 11354 44784 11462 44962
rect 11630 44784 11738 44962
rect 11906 44784 12014 44962
rect 12182 44784 12290 44962
rect 12458 44784 12566 44962
rect 12734 44784 12842 44962
rect 13010 44784 13118 44962
rect 13286 44784 13394 44962
rect 13562 44784 13670 44962
rect 13838 44784 13946 44962
rect 14114 44784 14222 44962
rect 14390 44784 14498 44962
rect 14666 44784 14774 44962
rect 14942 44784 15050 44962
rect 15218 44784 15326 44962
rect 15494 44784 15602 44962
rect 15770 44784 15878 44962
rect 16046 44784 16154 44962
rect 16322 44784 16430 44962
rect 16598 44784 16706 44962
rect 16874 44784 16982 44962
rect 17150 44784 17258 44962
rect 17426 44784 17534 44962
rect 17702 44784 17810 44962
rect 17978 44784 18086 44962
rect 18254 44784 18362 44962
rect 18530 44784 18638 44962
rect 18806 44784 18914 44962
rect 19082 44784 19190 44962
rect 19358 44784 19466 44962
rect 19634 44784 19742 44962
rect 19910 44784 20018 44962
rect 20186 44784 20294 44962
rect 20462 44784 20570 44962
rect 20738 44784 20846 44962
rect 21014 44784 21122 44962
rect 21290 44784 21398 44962
rect 21566 44784 21674 44962
rect 21842 44784 21950 44962
rect 22118 44784 22226 44962
rect 22394 44784 22502 44962
rect 22670 44784 22778 44962
rect 22946 44784 23054 44962
rect 23222 44784 23330 44962
rect 23498 44784 23606 44962
rect 23774 44784 23882 44962
rect 24050 44784 24158 44962
rect 24326 44784 24434 44962
rect 24602 44784 24710 44962
rect 24878 44784 24986 44962
rect 25154 44784 25262 44962
rect 25430 44784 25538 44962
rect 25706 44784 25924 44962
rect 18 216 25924 44784
rect 18 54 146 216
rect 314 54 422 216
rect 590 54 698 216
rect 866 54 974 216
rect 1142 54 1250 216
rect 1418 54 1526 216
rect 1694 54 1802 216
rect 1970 54 2078 216
rect 2246 54 2354 216
rect 2522 54 2630 216
rect 2798 54 2906 216
rect 3074 54 3182 216
rect 3350 54 3458 216
rect 3626 54 3734 216
rect 3902 54 4010 216
rect 4178 54 4286 216
rect 4454 54 4562 216
rect 4730 54 4838 216
rect 5006 54 5114 216
rect 5282 54 5390 216
rect 5558 54 5666 216
rect 5834 54 5942 216
rect 6110 54 6218 216
rect 6386 54 6494 216
rect 6662 54 6770 216
rect 6938 54 7046 216
rect 7214 54 7322 216
rect 7490 54 7598 216
rect 7766 54 7874 216
rect 8042 54 8150 216
rect 8318 54 8426 216
rect 8594 54 8702 216
rect 8870 54 8978 216
rect 9146 54 9254 216
rect 9422 54 9530 216
rect 9698 54 9806 216
rect 9974 54 10082 216
rect 10250 54 10358 216
rect 10526 54 10634 216
rect 10802 54 10910 216
rect 11078 54 11186 216
rect 11354 54 11462 216
rect 11630 54 11738 216
rect 11906 54 12014 216
rect 12182 54 12290 216
rect 12458 54 12566 216
rect 12734 54 12842 216
rect 13010 54 13118 216
rect 13286 54 13394 216
rect 13562 54 13670 216
rect 13838 54 13946 216
rect 14114 54 14222 216
rect 14390 54 14498 216
rect 14666 54 14774 216
rect 14942 54 15050 216
rect 15218 54 15326 216
rect 15494 54 15602 216
rect 15770 54 15878 216
rect 16046 54 16154 216
rect 16322 54 16430 216
rect 16598 54 16706 216
rect 16874 54 16982 216
rect 17150 54 17258 216
rect 17426 54 17534 216
rect 17702 54 17810 216
rect 17978 54 18086 216
rect 18254 54 18362 216
rect 18530 54 18638 216
rect 18806 54 18914 216
rect 19082 54 19190 216
rect 19358 54 19466 216
rect 19634 54 19742 216
rect 19910 54 20018 216
rect 20186 54 20294 216
rect 20462 54 20570 216
rect 20738 54 20846 216
rect 21014 54 21122 216
rect 21290 54 21398 216
rect 21566 54 21674 216
rect 21842 54 21950 216
rect 22118 54 22226 216
rect 22394 54 22502 216
rect 22670 54 22778 216
rect 22946 54 23054 216
rect 23222 54 23330 216
rect 23498 54 23606 216
rect 23774 54 23882 216
rect 24050 54 24158 216
rect 24326 54 24434 216
rect 24602 54 24710 216
rect 24878 54 24986 216
rect 25154 54 25262 216
rect 25430 54 25538 216
rect 25706 54 25924 216
<< metal3 >>
rect 25840 43800 26000 43920
rect 25840 43256 26000 43376
rect 25840 42712 26000 42832
rect 25840 42168 26000 42288
rect 25840 41624 26000 41744
rect 25840 41080 26000 41200
rect 25840 40536 26000 40656
rect 25840 39992 26000 40112
rect 0 39720 160 39840
rect 0 39448 160 39568
rect 25840 39448 26000 39568
rect 0 39176 160 39296
rect 0 38904 160 39024
rect 25840 38904 26000 39024
rect 0 38632 160 38752
rect 0 38360 160 38480
rect 25840 38360 26000 38480
rect 0 38088 160 38208
rect 0 37816 160 37936
rect 25840 37816 26000 37936
rect 0 37544 160 37664
rect 0 37272 160 37392
rect 25840 37272 26000 37392
rect 0 37000 160 37120
rect 0 36728 160 36848
rect 25840 36728 26000 36848
rect 0 36456 160 36576
rect 0 36184 160 36304
rect 25840 36184 26000 36304
rect 0 35912 160 36032
rect 0 35640 160 35760
rect 25840 35640 26000 35760
rect 0 35368 160 35488
rect 0 35096 160 35216
rect 25840 35096 26000 35216
rect 0 34824 160 34944
rect 0 34552 160 34672
rect 25840 34552 26000 34672
rect 0 34280 160 34400
rect 0 34008 160 34128
rect 25840 34008 26000 34128
rect 0 33736 160 33856
rect 0 33464 160 33584
rect 25840 33464 26000 33584
rect 0 33192 160 33312
rect 0 32920 160 33040
rect 25840 32920 26000 33040
rect 0 32648 160 32768
rect 0 32376 160 32496
rect 25840 32376 26000 32496
rect 0 32104 160 32224
rect 0 31832 160 31952
rect 25840 31832 26000 31952
rect 0 31560 160 31680
rect 0 31288 160 31408
rect 25840 31288 26000 31408
rect 0 31016 160 31136
rect 0 30744 160 30864
rect 25840 30744 26000 30864
rect 0 30472 160 30592
rect 0 30200 160 30320
rect 25840 30200 26000 30320
rect 0 29928 160 30048
rect 0 29656 160 29776
rect 25840 29656 26000 29776
rect 0 29384 160 29504
rect 0 29112 160 29232
rect 25840 29112 26000 29232
rect 0 28840 160 28960
rect 0 28568 160 28688
rect 25840 28568 26000 28688
rect 0 28296 160 28416
rect 0 28024 160 28144
rect 25840 28024 26000 28144
rect 0 27752 160 27872
rect 0 27480 160 27600
rect 25840 27480 26000 27600
rect 0 27208 160 27328
rect 0 26936 160 27056
rect 25840 26936 26000 27056
rect 0 26664 160 26784
rect 0 26392 160 26512
rect 25840 26392 26000 26512
rect 0 26120 160 26240
rect 0 25848 160 25968
rect 25840 25848 26000 25968
rect 0 25576 160 25696
rect 0 25304 160 25424
rect 25840 25304 26000 25424
rect 0 25032 160 25152
rect 0 24760 160 24880
rect 25840 24760 26000 24880
rect 0 24488 160 24608
rect 0 24216 160 24336
rect 25840 24216 26000 24336
rect 0 23944 160 24064
rect 0 23672 160 23792
rect 25840 23672 26000 23792
rect 0 23400 160 23520
rect 0 23128 160 23248
rect 25840 23128 26000 23248
rect 0 22856 160 22976
rect 0 22584 160 22704
rect 25840 22584 26000 22704
rect 0 22312 160 22432
rect 0 22040 160 22160
rect 25840 22040 26000 22160
rect 0 21768 160 21888
rect 0 21496 160 21616
rect 25840 21496 26000 21616
rect 0 21224 160 21344
rect 0 20952 160 21072
rect 25840 20952 26000 21072
rect 0 20680 160 20800
rect 0 20408 160 20528
rect 25840 20408 26000 20528
rect 0 20136 160 20256
rect 0 19864 160 19984
rect 25840 19864 26000 19984
rect 0 19592 160 19712
rect 0 19320 160 19440
rect 25840 19320 26000 19440
rect 0 19048 160 19168
rect 0 18776 160 18896
rect 25840 18776 26000 18896
rect 0 18504 160 18624
rect 0 18232 160 18352
rect 25840 18232 26000 18352
rect 0 17960 160 18080
rect 0 17688 160 17808
rect 25840 17688 26000 17808
rect 0 17416 160 17536
rect 0 17144 160 17264
rect 25840 17144 26000 17264
rect 0 16872 160 16992
rect 0 16600 160 16720
rect 25840 16600 26000 16720
rect 0 16328 160 16448
rect 0 16056 160 16176
rect 25840 16056 26000 16176
rect 0 15784 160 15904
rect 0 15512 160 15632
rect 25840 15512 26000 15632
rect 0 15240 160 15360
rect 0 14968 160 15088
rect 25840 14968 26000 15088
rect 0 14696 160 14816
rect 0 14424 160 14544
rect 25840 14424 26000 14544
rect 0 14152 160 14272
rect 0 13880 160 14000
rect 25840 13880 26000 14000
rect 0 13608 160 13728
rect 0 13336 160 13456
rect 25840 13336 26000 13456
rect 0 13064 160 13184
rect 0 12792 160 12912
rect 25840 12792 26000 12912
rect 0 12520 160 12640
rect 0 12248 160 12368
rect 25840 12248 26000 12368
rect 0 11976 160 12096
rect 0 11704 160 11824
rect 25840 11704 26000 11824
rect 0 11432 160 11552
rect 0 11160 160 11280
rect 25840 11160 26000 11280
rect 0 10888 160 11008
rect 0 10616 160 10736
rect 25840 10616 26000 10736
rect 0 10344 160 10464
rect 0 10072 160 10192
rect 25840 10072 26000 10192
rect 0 9800 160 9920
rect 0 9528 160 9648
rect 25840 9528 26000 9648
rect 0 9256 160 9376
rect 0 8984 160 9104
rect 25840 8984 26000 9104
rect 0 8712 160 8832
rect 0 8440 160 8560
rect 25840 8440 26000 8560
rect 0 8168 160 8288
rect 0 7896 160 8016
rect 25840 7896 26000 8016
rect 0 7624 160 7744
rect 0 7352 160 7472
rect 25840 7352 26000 7472
rect 0 7080 160 7200
rect 0 6808 160 6928
rect 25840 6808 26000 6928
rect 0 6536 160 6656
rect 0 6264 160 6384
rect 25840 6264 26000 6384
rect 0 5992 160 6112
rect 0 5720 160 5840
rect 25840 5720 26000 5840
rect 0 5448 160 5568
rect 0 5176 160 5296
rect 25840 5176 26000 5296
rect 25840 4632 26000 4752
rect 25840 4088 26000 4208
rect 25840 3544 26000 3664
rect 25840 3000 26000 3120
rect 25840 2456 26000 2576
rect 25840 1912 26000 2032
rect 25840 1368 26000 1488
rect 25840 824 26000 944
<< obsm3 >>
rect 13 43720 25760 43893
rect 13 43456 25840 43720
rect 13 43176 25760 43456
rect 13 42912 25840 43176
rect 13 42632 25760 42912
rect 13 42368 25840 42632
rect 13 42088 25760 42368
rect 13 41824 25840 42088
rect 13 41544 25760 41824
rect 13 41280 25840 41544
rect 13 41000 25760 41280
rect 13 40736 25840 41000
rect 13 40456 25760 40736
rect 13 40192 25840 40456
rect 13 39920 25760 40192
rect 240 39912 25760 39920
rect 240 39648 25840 39912
rect 240 39368 25760 39648
rect 240 39104 25840 39368
rect 240 38824 25760 39104
rect 240 38560 25840 38824
rect 240 38280 25760 38560
rect 240 38016 25840 38280
rect 240 37736 25760 38016
rect 240 37472 25840 37736
rect 240 37192 25760 37472
rect 240 36928 25840 37192
rect 240 36648 25760 36928
rect 240 36384 25840 36648
rect 240 36104 25760 36384
rect 240 35840 25840 36104
rect 240 35560 25760 35840
rect 240 35296 25840 35560
rect 240 35016 25760 35296
rect 240 34752 25840 35016
rect 240 34472 25760 34752
rect 240 34208 25840 34472
rect 240 33928 25760 34208
rect 240 33664 25840 33928
rect 240 33384 25760 33664
rect 240 33120 25840 33384
rect 240 32840 25760 33120
rect 240 32576 25840 32840
rect 240 32296 25760 32576
rect 240 32032 25840 32296
rect 240 31752 25760 32032
rect 240 31488 25840 31752
rect 240 31208 25760 31488
rect 240 30944 25840 31208
rect 240 30664 25760 30944
rect 240 30400 25840 30664
rect 240 30120 25760 30400
rect 240 29856 25840 30120
rect 240 29576 25760 29856
rect 240 29312 25840 29576
rect 240 29032 25760 29312
rect 240 28768 25840 29032
rect 240 28488 25760 28768
rect 240 28224 25840 28488
rect 240 27944 25760 28224
rect 240 27680 25840 27944
rect 240 27400 25760 27680
rect 240 27136 25840 27400
rect 240 26856 25760 27136
rect 240 26592 25840 26856
rect 240 26312 25760 26592
rect 240 26048 25840 26312
rect 240 25768 25760 26048
rect 240 25504 25840 25768
rect 240 25224 25760 25504
rect 240 24960 25840 25224
rect 240 24680 25760 24960
rect 240 24416 25840 24680
rect 240 24136 25760 24416
rect 240 23872 25840 24136
rect 240 23592 25760 23872
rect 240 23328 25840 23592
rect 240 23048 25760 23328
rect 240 22784 25840 23048
rect 240 22504 25760 22784
rect 240 22240 25840 22504
rect 240 21960 25760 22240
rect 240 21696 25840 21960
rect 240 21416 25760 21696
rect 240 21152 25840 21416
rect 240 20872 25760 21152
rect 240 20608 25840 20872
rect 240 20328 25760 20608
rect 240 20064 25840 20328
rect 240 19784 25760 20064
rect 240 19520 25840 19784
rect 240 19240 25760 19520
rect 240 18976 25840 19240
rect 240 18696 25760 18976
rect 240 18432 25840 18696
rect 240 18152 25760 18432
rect 240 17888 25840 18152
rect 240 17608 25760 17888
rect 240 17344 25840 17608
rect 240 17064 25760 17344
rect 240 16800 25840 17064
rect 240 16520 25760 16800
rect 240 16256 25840 16520
rect 240 15976 25760 16256
rect 240 15712 25840 15976
rect 240 15432 25760 15712
rect 240 15168 25840 15432
rect 240 14888 25760 15168
rect 240 14624 25840 14888
rect 240 14344 25760 14624
rect 240 14080 25840 14344
rect 240 13800 25760 14080
rect 240 13536 25840 13800
rect 240 13256 25760 13536
rect 240 12992 25840 13256
rect 240 12712 25760 12992
rect 240 12448 25840 12712
rect 240 12168 25760 12448
rect 240 11904 25840 12168
rect 240 11624 25760 11904
rect 240 11360 25840 11624
rect 240 11080 25760 11360
rect 240 10816 25840 11080
rect 240 10536 25760 10816
rect 240 10272 25840 10536
rect 240 9992 25760 10272
rect 240 9728 25840 9992
rect 240 9448 25760 9728
rect 240 9184 25840 9448
rect 240 8904 25760 9184
rect 240 8640 25840 8904
rect 240 8360 25760 8640
rect 240 8096 25840 8360
rect 240 7816 25760 8096
rect 240 7552 25840 7816
rect 240 7272 25760 7552
rect 240 7008 25840 7272
rect 240 6728 25760 7008
rect 240 6464 25840 6728
rect 240 6184 25760 6464
rect 240 5920 25840 6184
rect 240 5640 25760 5920
rect 240 5376 25840 5640
rect 240 5096 25760 5376
rect 13 4832 25840 5096
rect 13 4552 25760 4832
rect 13 4288 25840 4552
rect 13 4008 25760 4288
rect 13 3744 25840 4008
rect 13 3464 25760 3744
rect 13 3200 25840 3464
rect 13 2920 25760 3200
rect 13 2656 25840 2920
rect 13 2376 25760 2656
rect 13 2112 25840 2376
rect 13 1832 25760 2112
rect 13 1568 25840 1832
rect 13 1288 25760 1568
rect 13 1024 25840 1288
rect 13 744 25760 1024
rect 13 715 25840 744
<< metal4 >>
rect 3911 1040 4231 43568
rect 6878 1040 7198 43568
rect 9845 1040 10165 43568
rect 12812 1040 13132 43568
rect 15779 1040 16099 43568
rect 18746 1040 19066 43568
rect 21713 1040 22033 43568
rect 24680 1040 25000 43568
<< obsm4 >>
rect 611 960 3831 43213
rect 4311 960 6798 43213
rect 7278 960 9765 43213
rect 10245 960 12732 43213
rect 13212 960 15699 43213
rect 16179 960 18666 43213
rect 19146 960 21633 43213
rect 22113 960 24229 43213
rect 611 715 24229 960
<< labels >>
rlabel metal3 s 25840 9528 26000 9648 6 Config_accessC_bit0
port 1 nsew signal output
rlabel metal3 s 25840 10072 26000 10192 6 Config_accessC_bit1
port 2 nsew signal output
rlabel metal3 s 25840 10616 26000 10736 6 Config_accessC_bit2
port 3 nsew signal output
rlabel metal3 s 25840 11160 26000 11280 6 Config_accessC_bit3
port 4 nsew signal output
rlabel metal3 s 0 18232 160 18352 6 E1END[0]
port 5 nsew signal input
rlabel metal3 s 0 18504 160 18624 6 E1END[1]
port 6 nsew signal input
rlabel metal3 s 0 18776 160 18896 6 E1END[2]
port 7 nsew signal input
rlabel metal3 s 0 19048 160 19168 6 E1END[3]
port 8 nsew signal input
rlabel metal3 s 0 21496 160 21616 6 E2END[0]
port 9 nsew signal input
rlabel metal3 s 0 21768 160 21888 6 E2END[1]
port 10 nsew signal input
rlabel metal3 s 0 22040 160 22160 6 E2END[2]
port 11 nsew signal input
rlabel metal3 s 0 22312 160 22432 6 E2END[3]
port 12 nsew signal input
rlabel metal3 s 0 22584 160 22704 6 E2END[4]
port 13 nsew signal input
rlabel metal3 s 0 22856 160 22976 6 E2END[5]
port 14 nsew signal input
rlabel metal3 s 0 23128 160 23248 6 E2END[6]
port 15 nsew signal input
rlabel metal3 s 0 23400 160 23520 6 E2END[7]
port 16 nsew signal input
rlabel metal3 s 0 19320 160 19440 6 E2MID[0]
port 17 nsew signal input
rlabel metal3 s 0 19592 160 19712 6 E2MID[1]
port 18 nsew signal input
rlabel metal3 s 0 19864 160 19984 6 E2MID[2]
port 19 nsew signal input
rlabel metal3 s 0 20136 160 20256 6 E2MID[3]
port 20 nsew signal input
rlabel metal3 s 0 20408 160 20528 6 E2MID[4]
port 21 nsew signal input
rlabel metal3 s 0 20680 160 20800 6 E2MID[5]
port 22 nsew signal input
rlabel metal3 s 0 20952 160 21072 6 E2MID[6]
port 23 nsew signal input
rlabel metal3 s 0 21224 160 21344 6 E2MID[7]
port 24 nsew signal input
rlabel metal3 s 0 28024 160 28144 6 E6END[0]
port 25 nsew signal input
rlabel metal3 s 0 30744 160 30864 6 E6END[10]
port 26 nsew signal input
rlabel metal3 s 0 31016 160 31136 6 E6END[11]
port 27 nsew signal input
rlabel metal3 s 0 28296 160 28416 6 E6END[1]
port 28 nsew signal input
rlabel metal3 s 0 28568 160 28688 6 E6END[2]
port 29 nsew signal input
rlabel metal3 s 0 28840 160 28960 6 E6END[3]
port 30 nsew signal input
rlabel metal3 s 0 29112 160 29232 6 E6END[4]
port 31 nsew signal input
rlabel metal3 s 0 29384 160 29504 6 E6END[5]
port 32 nsew signal input
rlabel metal3 s 0 29656 160 29776 6 E6END[6]
port 33 nsew signal input
rlabel metal3 s 0 29928 160 30048 6 E6END[7]
port 34 nsew signal input
rlabel metal3 s 0 30200 160 30320 6 E6END[8]
port 35 nsew signal input
rlabel metal3 s 0 30472 160 30592 6 E6END[9]
port 36 nsew signal input
rlabel metal3 s 0 23672 160 23792 6 EE4END[0]
port 37 nsew signal input
rlabel metal3 s 0 26392 160 26512 6 EE4END[10]
port 38 nsew signal input
rlabel metal3 s 0 26664 160 26784 6 EE4END[11]
port 39 nsew signal input
rlabel metal3 s 0 26936 160 27056 6 EE4END[12]
port 40 nsew signal input
rlabel metal3 s 0 27208 160 27328 6 EE4END[13]
port 41 nsew signal input
rlabel metal3 s 0 27480 160 27600 6 EE4END[14]
port 42 nsew signal input
rlabel metal3 s 0 27752 160 27872 6 EE4END[15]
port 43 nsew signal input
rlabel metal3 s 0 23944 160 24064 6 EE4END[1]
port 44 nsew signal input
rlabel metal3 s 0 24216 160 24336 6 EE4END[2]
port 45 nsew signal input
rlabel metal3 s 0 24488 160 24608 6 EE4END[3]
port 46 nsew signal input
rlabel metal3 s 0 24760 160 24880 6 EE4END[4]
port 47 nsew signal input
rlabel metal3 s 0 25032 160 25152 6 EE4END[5]
port 48 nsew signal input
rlabel metal3 s 0 25304 160 25424 6 EE4END[6]
port 49 nsew signal input
rlabel metal3 s 0 25576 160 25696 6 EE4END[7]
port 50 nsew signal input
rlabel metal3 s 0 25848 160 25968 6 EE4END[8]
port 51 nsew signal input
rlabel metal3 s 0 26120 160 26240 6 EE4END[9]
port 52 nsew signal input
rlabel metal3 s 25840 16056 26000 16176 6 FAB2RAM_A0_O0
port 53 nsew signal output
rlabel metal3 s 25840 16600 26000 16720 6 FAB2RAM_A0_O1
port 54 nsew signal output
rlabel metal3 s 25840 17144 26000 17264 6 FAB2RAM_A0_O2
port 55 nsew signal output
rlabel metal3 s 25840 17688 26000 17808 6 FAB2RAM_A0_O3
port 56 nsew signal output
rlabel metal3 s 25840 13880 26000 14000 6 FAB2RAM_A1_O0
port 57 nsew signal output
rlabel metal3 s 25840 14424 26000 14544 6 FAB2RAM_A1_O1
port 58 nsew signal output
rlabel metal3 s 25840 14968 26000 15088 6 FAB2RAM_A1_O2
port 59 nsew signal output
rlabel metal3 s 25840 15512 26000 15632 6 FAB2RAM_A1_O3
port 60 nsew signal output
rlabel metal3 s 25840 11704 26000 11824 6 FAB2RAM_C_O0
port 61 nsew signal output
rlabel metal3 s 25840 12248 26000 12368 6 FAB2RAM_C_O1
port 62 nsew signal output
rlabel metal3 s 25840 12792 26000 12912 6 FAB2RAM_C_O2
port 63 nsew signal output
rlabel metal3 s 25840 13336 26000 13456 6 FAB2RAM_C_O3
port 64 nsew signal output
rlabel metal3 s 25840 24760 26000 24880 6 FAB2RAM_D0_O0
port 65 nsew signal output
rlabel metal3 s 25840 25304 26000 25424 6 FAB2RAM_D0_O1
port 66 nsew signal output
rlabel metal3 s 25840 25848 26000 25968 6 FAB2RAM_D0_O2
port 67 nsew signal output
rlabel metal3 s 25840 26392 26000 26512 6 FAB2RAM_D0_O3
port 68 nsew signal output
rlabel metal3 s 25840 22584 26000 22704 6 FAB2RAM_D1_O0
port 69 nsew signal output
rlabel metal3 s 25840 23128 26000 23248 6 FAB2RAM_D1_O1
port 70 nsew signal output
rlabel metal3 s 25840 23672 26000 23792 6 FAB2RAM_D1_O2
port 71 nsew signal output
rlabel metal3 s 25840 24216 26000 24336 6 FAB2RAM_D1_O3
port 72 nsew signal output
rlabel metal3 s 25840 20408 26000 20528 6 FAB2RAM_D2_O0
port 73 nsew signal output
rlabel metal3 s 25840 20952 26000 21072 6 FAB2RAM_D2_O1
port 74 nsew signal output
rlabel metal3 s 25840 21496 26000 21616 6 FAB2RAM_D2_O2
port 75 nsew signal output
rlabel metal3 s 25840 22040 26000 22160 6 FAB2RAM_D2_O3
port 76 nsew signal output
rlabel metal3 s 25840 18232 26000 18352 6 FAB2RAM_D3_O0
port 77 nsew signal output
rlabel metal3 s 25840 18776 26000 18896 6 FAB2RAM_D3_O1
port 78 nsew signal output
rlabel metal3 s 25840 19320 26000 19440 6 FAB2RAM_D3_O2
port 79 nsew signal output
rlabel metal3 s 25840 19864 26000 19984 6 FAB2RAM_D3_O3
port 80 nsew signal output
rlabel metal3 s 0 31288 160 31408 6 FrameData[0]
port 81 nsew signal input
rlabel metal3 s 0 34008 160 34128 6 FrameData[10]
port 82 nsew signal input
rlabel metal3 s 0 34280 160 34400 6 FrameData[11]
port 83 nsew signal input
rlabel metal3 s 0 34552 160 34672 6 FrameData[12]
port 84 nsew signal input
rlabel metal3 s 0 34824 160 34944 6 FrameData[13]
port 85 nsew signal input
rlabel metal3 s 0 35096 160 35216 6 FrameData[14]
port 86 nsew signal input
rlabel metal3 s 0 35368 160 35488 6 FrameData[15]
port 87 nsew signal input
rlabel metal3 s 0 35640 160 35760 6 FrameData[16]
port 88 nsew signal input
rlabel metal3 s 0 35912 160 36032 6 FrameData[17]
port 89 nsew signal input
rlabel metal3 s 0 36184 160 36304 6 FrameData[18]
port 90 nsew signal input
rlabel metal3 s 0 36456 160 36576 6 FrameData[19]
port 91 nsew signal input
rlabel metal3 s 0 31560 160 31680 6 FrameData[1]
port 92 nsew signal input
rlabel metal3 s 0 36728 160 36848 6 FrameData[20]
port 93 nsew signal input
rlabel metal3 s 0 37000 160 37120 6 FrameData[21]
port 94 nsew signal input
rlabel metal3 s 0 37272 160 37392 6 FrameData[22]
port 95 nsew signal input
rlabel metal3 s 0 37544 160 37664 6 FrameData[23]
port 96 nsew signal input
rlabel metal3 s 0 37816 160 37936 6 FrameData[24]
port 97 nsew signal input
rlabel metal3 s 0 38088 160 38208 6 FrameData[25]
port 98 nsew signal input
rlabel metal3 s 0 38360 160 38480 6 FrameData[26]
port 99 nsew signal input
rlabel metal3 s 0 38632 160 38752 6 FrameData[27]
port 100 nsew signal input
rlabel metal3 s 0 38904 160 39024 6 FrameData[28]
port 101 nsew signal input
rlabel metal3 s 0 39176 160 39296 6 FrameData[29]
port 102 nsew signal input
rlabel metal3 s 0 31832 160 31952 6 FrameData[2]
port 103 nsew signal input
rlabel metal3 s 0 39448 160 39568 6 FrameData[30]
port 104 nsew signal input
rlabel metal3 s 0 39720 160 39840 6 FrameData[31]
port 105 nsew signal input
rlabel metal3 s 0 32104 160 32224 6 FrameData[3]
port 106 nsew signal input
rlabel metal3 s 0 32376 160 32496 6 FrameData[4]
port 107 nsew signal input
rlabel metal3 s 0 32648 160 32768 6 FrameData[5]
port 108 nsew signal input
rlabel metal3 s 0 32920 160 33040 6 FrameData[6]
port 109 nsew signal input
rlabel metal3 s 0 33192 160 33312 6 FrameData[7]
port 110 nsew signal input
rlabel metal3 s 0 33464 160 33584 6 FrameData[8]
port 111 nsew signal input
rlabel metal3 s 0 33736 160 33856 6 FrameData[9]
port 112 nsew signal input
rlabel metal3 s 25840 26936 26000 27056 6 FrameData_O[0]
port 113 nsew signal output
rlabel metal3 s 25840 32376 26000 32496 6 FrameData_O[10]
port 114 nsew signal output
rlabel metal3 s 25840 32920 26000 33040 6 FrameData_O[11]
port 115 nsew signal output
rlabel metal3 s 25840 33464 26000 33584 6 FrameData_O[12]
port 116 nsew signal output
rlabel metal3 s 25840 34008 26000 34128 6 FrameData_O[13]
port 117 nsew signal output
rlabel metal3 s 25840 34552 26000 34672 6 FrameData_O[14]
port 118 nsew signal output
rlabel metal3 s 25840 35096 26000 35216 6 FrameData_O[15]
port 119 nsew signal output
rlabel metal3 s 25840 35640 26000 35760 6 FrameData_O[16]
port 120 nsew signal output
rlabel metal3 s 25840 36184 26000 36304 6 FrameData_O[17]
port 121 nsew signal output
rlabel metal3 s 25840 36728 26000 36848 6 FrameData_O[18]
port 122 nsew signal output
rlabel metal3 s 25840 37272 26000 37392 6 FrameData_O[19]
port 123 nsew signal output
rlabel metal3 s 25840 27480 26000 27600 6 FrameData_O[1]
port 124 nsew signal output
rlabel metal3 s 25840 37816 26000 37936 6 FrameData_O[20]
port 125 nsew signal output
rlabel metal3 s 25840 38360 26000 38480 6 FrameData_O[21]
port 126 nsew signal output
rlabel metal3 s 25840 38904 26000 39024 6 FrameData_O[22]
port 127 nsew signal output
rlabel metal3 s 25840 39448 26000 39568 6 FrameData_O[23]
port 128 nsew signal output
rlabel metal3 s 25840 39992 26000 40112 6 FrameData_O[24]
port 129 nsew signal output
rlabel metal3 s 25840 40536 26000 40656 6 FrameData_O[25]
port 130 nsew signal output
rlabel metal3 s 25840 41080 26000 41200 6 FrameData_O[26]
port 131 nsew signal output
rlabel metal3 s 25840 41624 26000 41744 6 FrameData_O[27]
port 132 nsew signal output
rlabel metal3 s 25840 42168 26000 42288 6 FrameData_O[28]
port 133 nsew signal output
rlabel metal3 s 25840 42712 26000 42832 6 FrameData_O[29]
port 134 nsew signal output
rlabel metal3 s 25840 28024 26000 28144 6 FrameData_O[2]
port 135 nsew signal output
rlabel metal3 s 25840 43256 26000 43376 6 FrameData_O[30]
port 136 nsew signal output
rlabel metal3 s 25840 43800 26000 43920 6 FrameData_O[31]
port 137 nsew signal output
rlabel metal3 s 25840 28568 26000 28688 6 FrameData_O[3]
port 138 nsew signal output
rlabel metal3 s 25840 29112 26000 29232 6 FrameData_O[4]
port 139 nsew signal output
rlabel metal3 s 25840 29656 26000 29776 6 FrameData_O[5]
port 140 nsew signal output
rlabel metal3 s 25840 30200 26000 30320 6 FrameData_O[6]
port 141 nsew signal output
rlabel metal3 s 25840 30744 26000 30864 6 FrameData_O[7]
port 142 nsew signal output
rlabel metal3 s 25840 31288 26000 31408 6 FrameData_O[8]
port 143 nsew signal output
rlabel metal3 s 25840 31832 26000 31952 6 FrameData_O[9]
port 144 nsew signal output
rlabel metal2 s 20350 0 20406 160 6 FrameStrobe[0]
port 145 nsew signal input
rlabel metal2 s 23110 0 23166 160 6 FrameStrobe[10]
port 146 nsew signal input
rlabel metal2 s 23386 0 23442 160 6 FrameStrobe[11]
port 147 nsew signal input
rlabel metal2 s 23662 0 23718 160 6 FrameStrobe[12]
port 148 nsew signal input
rlabel metal2 s 23938 0 23994 160 6 FrameStrobe[13]
port 149 nsew signal input
rlabel metal2 s 24214 0 24270 160 6 FrameStrobe[14]
port 150 nsew signal input
rlabel metal2 s 24490 0 24546 160 6 FrameStrobe[15]
port 151 nsew signal input
rlabel metal2 s 24766 0 24822 160 6 FrameStrobe[16]
port 152 nsew signal input
rlabel metal2 s 25042 0 25098 160 6 FrameStrobe[17]
port 153 nsew signal input
rlabel metal2 s 25318 0 25374 160 6 FrameStrobe[18]
port 154 nsew signal input
rlabel metal2 s 25594 0 25650 160 6 FrameStrobe[19]
port 155 nsew signal input
rlabel metal2 s 20626 0 20682 160 6 FrameStrobe[1]
port 156 nsew signal input
rlabel metal2 s 20902 0 20958 160 6 FrameStrobe[2]
port 157 nsew signal input
rlabel metal2 s 21178 0 21234 160 6 FrameStrobe[3]
port 158 nsew signal input
rlabel metal2 s 21454 0 21510 160 6 FrameStrobe[4]
port 159 nsew signal input
rlabel metal2 s 21730 0 21786 160 6 FrameStrobe[5]
port 160 nsew signal input
rlabel metal2 s 22006 0 22062 160 6 FrameStrobe[6]
port 161 nsew signal input
rlabel metal2 s 22282 0 22338 160 6 FrameStrobe[7]
port 162 nsew signal input
rlabel metal2 s 22558 0 22614 160 6 FrameStrobe[8]
port 163 nsew signal input
rlabel metal2 s 22834 0 22890 160 6 FrameStrobe[9]
port 164 nsew signal input
rlabel metal2 s 20350 44840 20406 45000 6 FrameStrobe_O[0]
port 165 nsew signal output
rlabel metal2 s 23110 44840 23166 45000 6 FrameStrobe_O[10]
port 166 nsew signal output
rlabel metal2 s 23386 44840 23442 45000 6 FrameStrobe_O[11]
port 167 nsew signal output
rlabel metal2 s 23662 44840 23718 45000 6 FrameStrobe_O[12]
port 168 nsew signal output
rlabel metal2 s 23938 44840 23994 45000 6 FrameStrobe_O[13]
port 169 nsew signal output
rlabel metal2 s 24214 44840 24270 45000 6 FrameStrobe_O[14]
port 170 nsew signal output
rlabel metal2 s 24490 44840 24546 45000 6 FrameStrobe_O[15]
port 171 nsew signal output
rlabel metal2 s 24766 44840 24822 45000 6 FrameStrobe_O[16]
port 172 nsew signal output
rlabel metal2 s 25042 44840 25098 45000 6 FrameStrobe_O[17]
port 173 nsew signal output
rlabel metal2 s 25318 44840 25374 45000 6 FrameStrobe_O[18]
port 174 nsew signal output
rlabel metal2 s 25594 44840 25650 45000 6 FrameStrobe_O[19]
port 175 nsew signal output
rlabel metal2 s 20626 44840 20682 45000 6 FrameStrobe_O[1]
port 176 nsew signal output
rlabel metal2 s 20902 44840 20958 45000 6 FrameStrobe_O[2]
port 177 nsew signal output
rlabel metal2 s 21178 44840 21234 45000 6 FrameStrobe_O[3]
port 178 nsew signal output
rlabel metal2 s 21454 44840 21510 45000 6 FrameStrobe_O[4]
port 179 nsew signal output
rlabel metal2 s 21730 44840 21786 45000 6 FrameStrobe_O[5]
port 180 nsew signal output
rlabel metal2 s 22006 44840 22062 45000 6 FrameStrobe_O[6]
port 181 nsew signal output
rlabel metal2 s 22282 44840 22338 45000 6 FrameStrobe_O[7]
port 182 nsew signal output
rlabel metal2 s 22558 44840 22614 45000 6 FrameStrobe_O[8]
port 183 nsew signal output
rlabel metal2 s 22834 44840 22890 45000 6 FrameStrobe_O[9]
port 184 nsew signal output
rlabel metal2 s 202 44840 258 45000 6 N1BEG[0]
port 185 nsew signal output
rlabel metal2 s 478 44840 534 45000 6 N1BEG[1]
port 186 nsew signal output
rlabel metal2 s 754 44840 810 45000 6 N1BEG[2]
port 187 nsew signal output
rlabel metal2 s 1030 44840 1086 45000 6 N1BEG[3]
port 188 nsew signal output
rlabel metal2 s 202 0 258 160 6 N1END[0]
port 189 nsew signal input
rlabel metal2 s 478 0 534 160 6 N1END[1]
port 190 nsew signal input
rlabel metal2 s 754 0 810 160 6 N1END[2]
port 191 nsew signal input
rlabel metal2 s 1030 0 1086 160 6 N1END[3]
port 192 nsew signal input
rlabel metal2 s 1306 44840 1362 45000 6 N2BEG[0]
port 193 nsew signal output
rlabel metal2 s 1582 44840 1638 45000 6 N2BEG[1]
port 194 nsew signal output
rlabel metal2 s 1858 44840 1914 45000 6 N2BEG[2]
port 195 nsew signal output
rlabel metal2 s 2134 44840 2190 45000 6 N2BEG[3]
port 196 nsew signal output
rlabel metal2 s 2410 44840 2466 45000 6 N2BEG[4]
port 197 nsew signal output
rlabel metal2 s 2686 44840 2742 45000 6 N2BEG[5]
port 198 nsew signal output
rlabel metal2 s 2962 44840 3018 45000 6 N2BEG[6]
port 199 nsew signal output
rlabel metal2 s 3238 44840 3294 45000 6 N2BEG[7]
port 200 nsew signal output
rlabel metal2 s 3514 44840 3570 45000 6 N2BEGb[0]
port 201 nsew signal output
rlabel metal2 s 3790 44840 3846 45000 6 N2BEGb[1]
port 202 nsew signal output
rlabel metal2 s 4066 44840 4122 45000 6 N2BEGb[2]
port 203 nsew signal output
rlabel metal2 s 4342 44840 4398 45000 6 N2BEGb[3]
port 204 nsew signal output
rlabel metal2 s 4618 44840 4674 45000 6 N2BEGb[4]
port 205 nsew signal output
rlabel metal2 s 4894 44840 4950 45000 6 N2BEGb[5]
port 206 nsew signal output
rlabel metal2 s 5170 44840 5226 45000 6 N2BEGb[6]
port 207 nsew signal output
rlabel metal2 s 5446 44840 5502 45000 6 N2BEGb[7]
port 208 nsew signal output
rlabel metal2 s 3514 0 3570 160 6 N2END[0]
port 209 nsew signal input
rlabel metal2 s 3790 0 3846 160 6 N2END[1]
port 210 nsew signal input
rlabel metal2 s 4066 0 4122 160 6 N2END[2]
port 211 nsew signal input
rlabel metal2 s 4342 0 4398 160 6 N2END[3]
port 212 nsew signal input
rlabel metal2 s 4618 0 4674 160 6 N2END[4]
port 213 nsew signal input
rlabel metal2 s 4894 0 4950 160 6 N2END[5]
port 214 nsew signal input
rlabel metal2 s 5170 0 5226 160 6 N2END[6]
port 215 nsew signal input
rlabel metal2 s 5446 0 5502 160 6 N2END[7]
port 216 nsew signal input
rlabel metal2 s 1306 0 1362 160 6 N2MID[0]
port 217 nsew signal input
rlabel metal2 s 1582 0 1638 160 6 N2MID[1]
port 218 nsew signal input
rlabel metal2 s 1858 0 1914 160 6 N2MID[2]
port 219 nsew signal input
rlabel metal2 s 2134 0 2190 160 6 N2MID[3]
port 220 nsew signal input
rlabel metal2 s 2410 0 2466 160 6 N2MID[4]
port 221 nsew signal input
rlabel metal2 s 2686 0 2742 160 6 N2MID[5]
port 222 nsew signal input
rlabel metal2 s 2962 0 3018 160 6 N2MID[6]
port 223 nsew signal input
rlabel metal2 s 3238 0 3294 160 6 N2MID[7]
port 224 nsew signal input
rlabel metal2 s 5722 44840 5778 45000 6 N4BEG[0]
port 225 nsew signal output
rlabel metal2 s 8482 44840 8538 45000 6 N4BEG[10]
port 226 nsew signal output
rlabel metal2 s 8758 44840 8814 45000 6 N4BEG[11]
port 227 nsew signal output
rlabel metal2 s 9034 44840 9090 45000 6 N4BEG[12]
port 228 nsew signal output
rlabel metal2 s 9310 44840 9366 45000 6 N4BEG[13]
port 229 nsew signal output
rlabel metal2 s 9586 44840 9642 45000 6 N4BEG[14]
port 230 nsew signal output
rlabel metal2 s 9862 44840 9918 45000 6 N4BEG[15]
port 231 nsew signal output
rlabel metal2 s 5998 44840 6054 45000 6 N4BEG[1]
port 232 nsew signal output
rlabel metal2 s 6274 44840 6330 45000 6 N4BEG[2]
port 233 nsew signal output
rlabel metal2 s 6550 44840 6606 45000 6 N4BEG[3]
port 234 nsew signal output
rlabel metal2 s 6826 44840 6882 45000 6 N4BEG[4]
port 235 nsew signal output
rlabel metal2 s 7102 44840 7158 45000 6 N4BEG[5]
port 236 nsew signal output
rlabel metal2 s 7378 44840 7434 45000 6 N4BEG[6]
port 237 nsew signal output
rlabel metal2 s 7654 44840 7710 45000 6 N4BEG[7]
port 238 nsew signal output
rlabel metal2 s 7930 44840 7986 45000 6 N4BEG[8]
port 239 nsew signal output
rlabel metal2 s 8206 44840 8262 45000 6 N4BEG[9]
port 240 nsew signal output
rlabel metal2 s 5722 0 5778 160 6 N4END[0]
port 241 nsew signal input
rlabel metal2 s 8482 0 8538 160 6 N4END[10]
port 242 nsew signal input
rlabel metal2 s 8758 0 8814 160 6 N4END[11]
port 243 nsew signal input
rlabel metal2 s 9034 0 9090 160 6 N4END[12]
port 244 nsew signal input
rlabel metal2 s 9310 0 9366 160 6 N4END[13]
port 245 nsew signal input
rlabel metal2 s 9586 0 9642 160 6 N4END[14]
port 246 nsew signal input
rlabel metal2 s 9862 0 9918 160 6 N4END[15]
port 247 nsew signal input
rlabel metal2 s 5998 0 6054 160 6 N4END[1]
port 248 nsew signal input
rlabel metal2 s 6274 0 6330 160 6 N4END[2]
port 249 nsew signal input
rlabel metal2 s 6550 0 6606 160 6 N4END[3]
port 250 nsew signal input
rlabel metal2 s 6826 0 6882 160 6 N4END[4]
port 251 nsew signal input
rlabel metal2 s 7102 0 7158 160 6 N4END[5]
port 252 nsew signal input
rlabel metal2 s 7378 0 7434 160 6 N4END[6]
port 253 nsew signal input
rlabel metal2 s 7654 0 7710 160 6 N4END[7]
port 254 nsew signal input
rlabel metal2 s 7930 0 7986 160 6 N4END[8]
port 255 nsew signal input
rlabel metal2 s 8206 0 8262 160 6 N4END[9]
port 256 nsew signal input
rlabel metal3 s 25840 7352 26000 7472 6 RAM2FAB_D0_I0
port 257 nsew signal input
rlabel metal3 s 25840 7896 26000 8016 6 RAM2FAB_D0_I1
port 258 nsew signal input
rlabel metal3 s 25840 8440 26000 8560 6 RAM2FAB_D0_I2
port 259 nsew signal input
rlabel metal3 s 25840 8984 26000 9104 6 RAM2FAB_D0_I3
port 260 nsew signal input
rlabel metal3 s 25840 5176 26000 5296 6 RAM2FAB_D1_I0
port 261 nsew signal input
rlabel metal3 s 25840 5720 26000 5840 6 RAM2FAB_D1_I1
port 262 nsew signal input
rlabel metal3 s 25840 6264 26000 6384 6 RAM2FAB_D1_I2
port 263 nsew signal input
rlabel metal3 s 25840 6808 26000 6928 6 RAM2FAB_D1_I3
port 264 nsew signal input
rlabel metal3 s 25840 3000 26000 3120 6 RAM2FAB_D2_I0
port 265 nsew signal input
rlabel metal3 s 25840 3544 26000 3664 6 RAM2FAB_D2_I1
port 266 nsew signal input
rlabel metal3 s 25840 4088 26000 4208 6 RAM2FAB_D2_I2
port 267 nsew signal input
rlabel metal3 s 25840 4632 26000 4752 6 RAM2FAB_D2_I3
port 268 nsew signal input
rlabel metal3 s 25840 824 26000 944 6 RAM2FAB_D3_I0
port 269 nsew signal input
rlabel metal3 s 25840 1368 26000 1488 6 RAM2FAB_D3_I1
port 270 nsew signal input
rlabel metal3 s 25840 1912 26000 2032 6 RAM2FAB_D3_I2
port 271 nsew signal input
rlabel metal3 s 25840 2456 26000 2576 6 RAM2FAB_D3_I3
port 272 nsew signal input
rlabel metal2 s 10138 0 10194 160 6 S1BEG[0]
port 273 nsew signal output
rlabel metal2 s 10414 0 10470 160 6 S1BEG[1]
port 274 nsew signal output
rlabel metal2 s 10690 0 10746 160 6 S1BEG[2]
port 275 nsew signal output
rlabel metal2 s 10966 0 11022 160 6 S1BEG[3]
port 276 nsew signal output
rlabel metal2 s 10138 44840 10194 45000 6 S1END[0]
port 277 nsew signal input
rlabel metal2 s 10414 44840 10470 45000 6 S1END[1]
port 278 nsew signal input
rlabel metal2 s 10690 44840 10746 45000 6 S1END[2]
port 279 nsew signal input
rlabel metal2 s 10966 44840 11022 45000 6 S1END[3]
port 280 nsew signal input
rlabel metal2 s 13450 0 13506 160 6 S2BEG[0]
port 281 nsew signal output
rlabel metal2 s 13726 0 13782 160 6 S2BEG[1]
port 282 nsew signal output
rlabel metal2 s 14002 0 14058 160 6 S2BEG[2]
port 283 nsew signal output
rlabel metal2 s 14278 0 14334 160 6 S2BEG[3]
port 284 nsew signal output
rlabel metal2 s 14554 0 14610 160 6 S2BEG[4]
port 285 nsew signal output
rlabel metal2 s 14830 0 14886 160 6 S2BEG[5]
port 286 nsew signal output
rlabel metal2 s 15106 0 15162 160 6 S2BEG[6]
port 287 nsew signal output
rlabel metal2 s 15382 0 15438 160 6 S2BEG[7]
port 288 nsew signal output
rlabel metal2 s 11242 0 11298 160 6 S2BEGb[0]
port 289 nsew signal output
rlabel metal2 s 11518 0 11574 160 6 S2BEGb[1]
port 290 nsew signal output
rlabel metal2 s 11794 0 11850 160 6 S2BEGb[2]
port 291 nsew signal output
rlabel metal2 s 12070 0 12126 160 6 S2BEGb[3]
port 292 nsew signal output
rlabel metal2 s 12346 0 12402 160 6 S2BEGb[4]
port 293 nsew signal output
rlabel metal2 s 12622 0 12678 160 6 S2BEGb[5]
port 294 nsew signal output
rlabel metal2 s 12898 0 12954 160 6 S2BEGb[6]
port 295 nsew signal output
rlabel metal2 s 13174 0 13230 160 6 S2BEGb[7]
port 296 nsew signal output
rlabel metal2 s 11242 44840 11298 45000 6 S2END[0]
port 297 nsew signal input
rlabel metal2 s 11518 44840 11574 45000 6 S2END[1]
port 298 nsew signal input
rlabel metal2 s 11794 44840 11850 45000 6 S2END[2]
port 299 nsew signal input
rlabel metal2 s 12070 44840 12126 45000 6 S2END[3]
port 300 nsew signal input
rlabel metal2 s 12346 44840 12402 45000 6 S2END[4]
port 301 nsew signal input
rlabel metal2 s 12622 44840 12678 45000 6 S2END[5]
port 302 nsew signal input
rlabel metal2 s 12898 44840 12954 45000 6 S2END[6]
port 303 nsew signal input
rlabel metal2 s 13174 44840 13230 45000 6 S2END[7]
port 304 nsew signal input
rlabel metal2 s 13450 44840 13506 45000 6 S2MID[0]
port 305 nsew signal input
rlabel metal2 s 13726 44840 13782 45000 6 S2MID[1]
port 306 nsew signal input
rlabel metal2 s 14002 44840 14058 45000 6 S2MID[2]
port 307 nsew signal input
rlabel metal2 s 14278 44840 14334 45000 6 S2MID[3]
port 308 nsew signal input
rlabel metal2 s 14554 44840 14610 45000 6 S2MID[4]
port 309 nsew signal input
rlabel metal2 s 14830 44840 14886 45000 6 S2MID[5]
port 310 nsew signal input
rlabel metal2 s 15106 44840 15162 45000 6 S2MID[6]
port 311 nsew signal input
rlabel metal2 s 15382 44840 15438 45000 6 S2MID[7]
port 312 nsew signal input
rlabel metal2 s 15658 0 15714 160 6 S4BEG[0]
port 313 nsew signal output
rlabel metal2 s 18418 0 18474 160 6 S4BEG[10]
port 314 nsew signal output
rlabel metal2 s 18694 0 18750 160 6 S4BEG[11]
port 315 nsew signal output
rlabel metal2 s 18970 0 19026 160 6 S4BEG[12]
port 316 nsew signal output
rlabel metal2 s 19246 0 19302 160 6 S4BEG[13]
port 317 nsew signal output
rlabel metal2 s 19522 0 19578 160 6 S4BEG[14]
port 318 nsew signal output
rlabel metal2 s 19798 0 19854 160 6 S4BEG[15]
port 319 nsew signal output
rlabel metal2 s 15934 0 15990 160 6 S4BEG[1]
port 320 nsew signal output
rlabel metal2 s 16210 0 16266 160 6 S4BEG[2]
port 321 nsew signal output
rlabel metal2 s 16486 0 16542 160 6 S4BEG[3]
port 322 nsew signal output
rlabel metal2 s 16762 0 16818 160 6 S4BEG[4]
port 323 nsew signal output
rlabel metal2 s 17038 0 17094 160 6 S4BEG[5]
port 324 nsew signal output
rlabel metal2 s 17314 0 17370 160 6 S4BEG[6]
port 325 nsew signal output
rlabel metal2 s 17590 0 17646 160 6 S4BEG[7]
port 326 nsew signal output
rlabel metal2 s 17866 0 17922 160 6 S4BEG[8]
port 327 nsew signal output
rlabel metal2 s 18142 0 18198 160 6 S4BEG[9]
port 328 nsew signal output
rlabel metal2 s 15658 44840 15714 45000 6 S4END[0]
port 329 nsew signal input
rlabel metal2 s 18418 44840 18474 45000 6 S4END[10]
port 330 nsew signal input
rlabel metal2 s 18694 44840 18750 45000 6 S4END[11]
port 331 nsew signal input
rlabel metal2 s 18970 44840 19026 45000 6 S4END[12]
port 332 nsew signal input
rlabel metal2 s 19246 44840 19302 45000 6 S4END[13]
port 333 nsew signal input
rlabel metal2 s 19522 44840 19578 45000 6 S4END[14]
port 334 nsew signal input
rlabel metal2 s 19798 44840 19854 45000 6 S4END[15]
port 335 nsew signal input
rlabel metal2 s 15934 44840 15990 45000 6 S4END[1]
port 336 nsew signal input
rlabel metal2 s 16210 44840 16266 45000 6 S4END[2]
port 337 nsew signal input
rlabel metal2 s 16486 44840 16542 45000 6 S4END[3]
port 338 nsew signal input
rlabel metal2 s 16762 44840 16818 45000 6 S4END[4]
port 339 nsew signal input
rlabel metal2 s 17038 44840 17094 45000 6 S4END[5]
port 340 nsew signal input
rlabel metal2 s 17314 44840 17370 45000 6 S4END[6]
port 341 nsew signal input
rlabel metal2 s 17590 44840 17646 45000 6 S4END[7]
port 342 nsew signal input
rlabel metal2 s 17866 44840 17922 45000 6 S4END[8]
port 343 nsew signal input
rlabel metal2 s 18142 44840 18198 45000 6 S4END[9]
port 344 nsew signal input
rlabel metal2 s 20074 0 20130 160 6 UserCLK
port 345 nsew signal input
rlabel metal2 s 20074 44840 20130 45000 6 UserCLKo
port 346 nsew signal output
rlabel metal4 s 6878 1040 7198 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 12812 1040 13132 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 18746 1040 19066 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 24680 1040 25000 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 3911 1040 4231 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal4 s 9845 1040 10165 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal4 s 15779 1040 16099 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal4 s 21713 1040 22033 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal3 s 0 5176 160 5296 6 W1BEG[0]
port 349 nsew signal output
rlabel metal3 s 0 5448 160 5568 6 W1BEG[1]
port 350 nsew signal output
rlabel metal3 s 0 5720 160 5840 6 W1BEG[2]
port 351 nsew signal output
rlabel metal3 s 0 5992 160 6112 6 W1BEG[3]
port 352 nsew signal output
rlabel metal3 s 0 6264 160 6384 6 W2BEG[0]
port 353 nsew signal output
rlabel metal3 s 0 6536 160 6656 6 W2BEG[1]
port 354 nsew signal output
rlabel metal3 s 0 6808 160 6928 6 W2BEG[2]
port 355 nsew signal output
rlabel metal3 s 0 7080 160 7200 6 W2BEG[3]
port 356 nsew signal output
rlabel metal3 s 0 7352 160 7472 6 W2BEG[4]
port 357 nsew signal output
rlabel metal3 s 0 7624 160 7744 6 W2BEG[5]
port 358 nsew signal output
rlabel metal3 s 0 7896 160 8016 6 W2BEG[6]
port 359 nsew signal output
rlabel metal3 s 0 8168 160 8288 6 W2BEG[7]
port 360 nsew signal output
rlabel metal3 s 0 8440 160 8560 6 W2BEGb[0]
port 361 nsew signal output
rlabel metal3 s 0 8712 160 8832 6 W2BEGb[1]
port 362 nsew signal output
rlabel metal3 s 0 8984 160 9104 6 W2BEGb[2]
port 363 nsew signal output
rlabel metal3 s 0 9256 160 9376 6 W2BEGb[3]
port 364 nsew signal output
rlabel metal3 s 0 9528 160 9648 6 W2BEGb[4]
port 365 nsew signal output
rlabel metal3 s 0 9800 160 9920 6 W2BEGb[5]
port 366 nsew signal output
rlabel metal3 s 0 10072 160 10192 6 W2BEGb[6]
port 367 nsew signal output
rlabel metal3 s 0 10344 160 10464 6 W2BEGb[7]
port 368 nsew signal output
rlabel metal3 s 0 14968 160 15088 6 W6BEG[0]
port 369 nsew signal output
rlabel metal3 s 0 17688 160 17808 6 W6BEG[10]
port 370 nsew signal output
rlabel metal3 s 0 17960 160 18080 6 W6BEG[11]
port 371 nsew signal output
rlabel metal3 s 0 15240 160 15360 6 W6BEG[1]
port 372 nsew signal output
rlabel metal3 s 0 15512 160 15632 6 W6BEG[2]
port 373 nsew signal output
rlabel metal3 s 0 15784 160 15904 6 W6BEG[3]
port 374 nsew signal output
rlabel metal3 s 0 16056 160 16176 6 W6BEG[4]
port 375 nsew signal output
rlabel metal3 s 0 16328 160 16448 6 W6BEG[5]
port 376 nsew signal output
rlabel metal3 s 0 16600 160 16720 6 W6BEG[6]
port 377 nsew signal output
rlabel metal3 s 0 16872 160 16992 6 W6BEG[7]
port 378 nsew signal output
rlabel metal3 s 0 17144 160 17264 6 W6BEG[8]
port 379 nsew signal output
rlabel metal3 s 0 17416 160 17536 6 W6BEG[9]
port 380 nsew signal output
rlabel metal3 s 0 10616 160 10736 6 WW4BEG[0]
port 381 nsew signal output
rlabel metal3 s 0 13336 160 13456 6 WW4BEG[10]
port 382 nsew signal output
rlabel metal3 s 0 13608 160 13728 6 WW4BEG[11]
port 383 nsew signal output
rlabel metal3 s 0 13880 160 14000 6 WW4BEG[12]
port 384 nsew signal output
rlabel metal3 s 0 14152 160 14272 6 WW4BEG[13]
port 385 nsew signal output
rlabel metal3 s 0 14424 160 14544 6 WW4BEG[14]
port 386 nsew signal output
rlabel metal3 s 0 14696 160 14816 6 WW4BEG[15]
port 387 nsew signal output
rlabel metal3 s 0 10888 160 11008 6 WW4BEG[1]
port 388 nsew signal output
rlabel metal3 s 0 11160 160 11280 6 WW4BEG[2]
port 389 nsew signal output
rlabel metal3 s 0 11432 160 11552 6 WW4BEG[3]
port 390 nsew signal output
rlabel metal3 s 0 11704 160 11824 6 WW4BEG[4]
port 391 nsew signal output
rlabel metal3 s 0 11976 160 12096 6 WW4BEG[5]
port 392 nsew signal output
rlabel metal3 s 0 12248 160 12368 6 WW4BEG[6]
port 393 nsew signal output
rlabel metal3 s 0 12520 160 12640 6 WW4BEG[7]
port 394 nsew signal output
rlabel metal3 s 0 12792 160 12912 6 WW4BEG[8]
port 395 nsew signal output
rlabel metal3 s 0 13064 160 13184 6 WW4BEG[9]
port 396 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 26000 45000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4287984
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/RAM_IO/runs/24_12_03_16_04/results/signoff/RAM_IO.magic.gds
string GDS_START 173598
<< end >>

