VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DSP
  CLASS BLOCK ;
  FOREIGN DSP ;
  ORIGIN 0.000 0.000 ;
  SIZE 225.000 BY 450.000 ;
  PIN Tile_X0Y0_E1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 319.640 225.000 320.240 ;
    END
  END Tile_X0Y0_E1BEG[0]
  PIN Tile_X0Y0_E1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 321.000 225.000 321.600 ;
    END
  END Tile_X0Y0_E1BEG[1]
  PIN Tile_X0Y0_E1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 322.360 225.000 322.960 ;
    END
  END Tile_X0Y0_E1BEG[2]
  PIN Tile_X0Y0_E1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 323.720 225.000 324.320 ;
    END
  END Tile_X0Y0_E1BEG[3]
  PIN Tile_X0Y0_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 0.800 320.240 ;
    END
  END Tile_X0Y0_E1END[0]
  PIN Tile_X0Y0_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 0.800 321.600 ;
    END
  END Tile_X0Y0_E1END[1]
  PIN Tile_X0Y0_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 0.800 322.960 ;
    END
  END Tile_X0Y0_E1END[2]
  PIN Tile_X0Y0_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 0.800 324.320 ;
    END
  END Tile_X0Y0_E1END[3]
  PIN Tile_X0Y0_E2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 325.080 225.000 325.680 ;
    END
  END Tile_X0Y0_E2BEG[0]
  PIN Tile_X0Y0_E2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 326.440 225.000 327.040 ;
    END
  END Tile_X0Y0_E2BEG[1]
  PIN Tile_X0Y0_E2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 327.800 225.000 328.400 ;
    END
  END Tile_X0Y0_E2BEG[2]
  PIN Tile_X0Y0_E2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 329.160 225.000 329.760 ;
    END
  END Tile_X0Y0_E2BEG[3]
  PIN Tile_X0Y0_E2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 330.520 225.000 331.120 ;
    END
  END Tile_X0Y0_E2BEG[4]
  PIN Tile_X0Y0_E2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 331.880 225.000 332.480 ;
    END
  END Tile_X0Y0_E2BEG[5]
  PIN Tile_X0Y0_E2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 333.240 225.000 333.840 ;
    END
  END Tile_X0Y0_E2BEG[6]
  PIN Tile_X0Y0_E2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 334.600 225.000 335.200 ;
    END
  END Tile_X0Y0_E2BEG[7]
  PIN Tile_X0Y0_E2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 335.960 225.000 336.560 ;
    END
  END Tile_X0Y0_E2BEGb[0]
  PIN Tile_X0Y0_E2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 337.320 225.000 337.920 ;
    END
  END Tile_X0Y0_E2BEGb[1]
  PIN Tile_X0Y0_E2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 338.680 225.000 339.280 ;
    END
  END Tile_X0Y0_E2BEGb[2]
  PIN Tile_X0Y0_E2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 340.040 225.000 340.640 ;
    END
  END Tile_X0Y0_E2BEGb[3]
  PIN Tile_X0Y0_E2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 341.400 225.000 342.000 ;
    END
  END Tile_X0Y0_E2BEGb[4]
  PIN Tile_X0Y0_E2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 342.760 225.000 343.360 ;
    END
  END Tile_X0Y0_E2BEGb[5]
  PIN Tile_X0Y0_E2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 344.120 225.000 344.720 ;
    END
  END Tile_X0Y0_E2BEGb[6]
  PIN Tile_X0Y0_E2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 345.480 225.000 346.080 ;
    END
  END Tile_X0Y0_E2BEGb[7]
  PIN Tile_X0Y0_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 0.800 336.560 ;
    END
  END Tile_X0Y0_E2END[0]
  PIN Tile_X0Y0_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 0.800 337.920 ;
    END
  END Tile_X0Y0_E2END[1]
  PIN Tile_X0Y0_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 0.800 339.280 ;
    END
  END Tile_X0Y0_E2END[2]
  PIN Tile_X0Y0_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 0.800 340.640 ;
    END
  END Tile_X0Y0_E2END[3]
  PIN Tile_X0Y0_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 0.800 342.000 ;
    END
  END Tile_X0Y0_E2END[4]
  PIN Tile_X0Y0_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 0.800 343.360 ;
    END
  END Tile_X0Y0_E2END[5]
  PIN Tile_X0Y0_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 0.800 344.720 ;
    END
  END Tile_X0Y0_E2END[6]
  PIN Tile_X0Y0_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 0.800 346.080 ;
    END
  END Tile_X0Y0_E2END[7]
  PIN Tile_X0Y0_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 0.800 325.680 ;
    END
  END Tile_X0Y0_E2MID[0]
  PIN Tile_X0Y0_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 0.800 327.040 ;
    END
  END Tile_X0Y0_E2MID[1]
  PIN Tile_X0Y0_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 0.800 328.400 ;
    END
  END Tile_X0Y0_E2MID[2]
  PIN Tile_X0Y0_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 0.800 329.760 ;
    END
  END Tile_X0Y0_E2MID[3]
  PIN Tile_X0Y0_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 0.800 331.120 ;
    END
  END Tile_X0Y0_E2MID[4]
  PIN Tile_X0Y0_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 0.800 332.480 ;
    END
  END Tile_X0Y0_E2MID[5]
  PIN Tile_X0Y0_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 0.800 333.840 ;
    END
  END Tile_X0Y0_E2MID[6]
  PIN Tile_X0Y0_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 0.800 335.200 ;
    END
  END Tile_X0Y0_E2MID[7]
  PIN Tile_X0Y0_E6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 368.600 225.000 369.200 ;
    END
  END Tile_X0Y0_E6BEG[0]
  PIN Tile_X0Y0_E6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 382.200 225.000 382.800 ;
    END
  END Tile_X0Y0_E6BEG[10]
  PIN Tile_X0Y0_E6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 383.560 225.000 384.160 ;
    END
  END Tile_X0Y0_E6BEG[11]
  PIN Tile_X0Y0_E6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 369.960 225.000 370.560 ;
    END
  END Tile_X0Y0_E6BEG[1]
  PIN Tile_X0Y0_E6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 371.320 225.000 371.920 ;
    END
  END Tile_X0Y0_E6BEG[2]
  PIN Tile_X0Y0_E6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 372.680 225.000 373.280 ;
    END
  END Tile_X0Y0_E6BEG[3]
  PIN Tile_X0Y0_E6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 374.040 225.000 374.640 ;
    END
  END Tile_X0Y0_E6BEG[4]
  PIN Tile_X0Y0_E6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 375.400 225.000 376.000 ;
    END
  END Tile_X0Y0_E6BEG[5]
  PIN Tile_X0Y0_E6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 376.760 225.000 377.360 ;
    END
  END Tile_X0Y0_E6BEG[6]
  PIN Tile_X0Y0_E6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 378.120 225.000 378.720 ;
    END
  END Tile_X0Y0_E6BEG[7]
  PIN Tile_X0Y0_E6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 379.480 225.000 380.080 ;
    END
  END Tile_X0Y0_E6BEG[8]
  PIN Tile_X0Y0_E6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 380.840 225.000 381.440 ;
    END
  END Tile_X0Y0_E6BEG[9]
  PIN Tile_X0Y0_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 0.800 369.200 ;
    END
  END Tile_X0Y0_E6END[0]
  PIN Tile_X0Y0_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 0.800 382.800 ;
    END
  END Tile_X0Y0_E6END[10]
  PIN Tile_X0Y0_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 0.800 384.160 ;
    END
  END Tile_X0Y0_E6END[11]
  PIN Tile_X0Y0_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 0.800 370.560 ;
    END
  END Tile_X0Y0_E6END[1]
  PIN Tile_X0Y0_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 0.800 371.920 ;
    END
  END Tile_X0Y0_E6END[2]
  PIN Tile_X0Y0_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 0.800 373.280 ;
    END
  END Tile_X0Y0_E6END[3]
  PIN Tile_X0Y0_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 0.800 374.640 ;
    END
  END Tile_X0Y0_E6END[4]
  PIN Tile_X0Y0_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 0.800 376.000 ;
    END
  END Tile_X0Y0_E6END[5]
  PIN Tile_X0Y0_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 0.800 377.360 ;
    END
  END Tile_X0Y0_E6END[6]
  PIN Tile_X0Y0_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 0.800 378.720 ;
    END
  END Tile_X0Y0_E6END[7]
  PIN Tile_X0Y0_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 0.800 380.080 ;
    END
  END Tile_X0Y0_E6END[8]
  PIN Tile_X0Y0_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 0.800 381.440 ;
    END
  END Tile_X0Y0_E6END[9]
  PIN Tile_X0Y0_EE4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 346.840 225.000 347.440 ;
    END
  END Tile_X0Y0_EE4BEG[0]
  PIN Tile_X0Y0_EE4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 360.440 225.000 361.040 ;
    END
  END Tile_X0Y0_EE4BEG[10]
  PIN Tile_X0Y0_EE4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 361.800 225.000 362.400 ;
    END
  END Tile_X0Y0_EE4BEG[11]
  PIN Tile_X0Y0_EE4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 363.160 225.000 363.760 ;
    END
  END Tile_X0Y0_EE4BEG[12]
  PIN Tile_X0Y0_EE4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 364.520 225.000 365.120 ;
    END
  END Tile_X0Y0_EE4BEG[13]
  PIN Tile_X0Y0_EE4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 365.880 225.000 366.480 ;
    END
  END Tile_X0Y0_EE4BEG[14]
  PIN Tile_X0Y0_EE4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 367.240 225.000 367.840 ;
    END
  END Tile_X0Y0_EE4BEG[15]
  PIN Tile_X0Y0_EE4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 348.200 225.000 348.800 ;
    END
  END Tile_X0Y0_EE4BEG[1]
  PIN Tile_X0Y0_EE4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 349.560 225.000 350.160 ;
    END
  END Tile_X0Y0_EE4BEG[2]
  PIN Tile_X0Y0_EE4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 350.920 225.000 351.520 ;
    END
  END Tile_X0Y0_EE4BEG[3]
  PIN Tile_X0Y0_EE4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 352.280 225.000 352.880 ;
    END
  END Tile_X0Y0_EE4BEG[4]
  PIN Tile_X0Y0_EE4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 353.640 225.000 354.240 ;
    END
  END Tile_X0Y0_EE4BEG[5]
  PIN Tile_X0Y0_EE4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 355.000 225.000 355.600 ;
    END
  END Tile_X0Y0_EE4BEG[6]
  PIN Tile_X0Y0_EE4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 356.360 225.000 356.960 ;
    END
  END Tile_X0Y0_EE4BEG[7]
  PIN Tile_X0Y0_EE4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 357.720 225.000 358.320 ;
    END
  END Tile_X0Y0_EE4BEG[8]
  PIN Tile_X0Y0_EE4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 359.080 225.000 359.680 ;
    END
  END Tile_X0Y0_EE4BEG[9]
  PIN Tile_X0Y0_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 0.800 347.440 ;
    END
  END Tile_X0Y0_EE4END[0]
  PIN Tile_X0Y0_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 0.800 361.040 ;
    END
  END Tile_X0Y0_EE4END[10]
  PIN Tile_X0Y0_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 0.800 362.400 ;
    END
  END Tile_X0Y0_EE4END[11]
  PIN Tile_X0Y0_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 0.800 363.760 ;
    END
  END Tile_X0Y0_EE4END[12]
  PIN Tile_X0Y0_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 0.800 365.120 ;
    END
  END Tile_X0Y0_EE4END[13]
  PIN Tile_X0Y0_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 0.800 366.480 ;
    END
  END Tile_X0Y0_EE4END[14]
  PIN Tile_X0Y0_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 0.800 367.840 ;
    END
  END Tile_X0Y0_EE4END[15]
  PIN Tile_X0Y0_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 0.800 348.800 ;
    END
  END Tile_X0Y0_EE4END[1]
  PIN Tile_X0Y0_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 0.800 350.160 ;
    END
  END Tile_X0Y0_EE4END[2]
  PIN Tile_X0Y0_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 0.800 351.520 ;
    END
  END Tile_X0Y0_EE4END[3]
  PIN Tile_X0Y0_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 0.800 352.880 ;
    END
  END Tile_X0Y0_EE4END[4]
  PIN Tile_X0Y0_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 0.800 354.240 ;
    END
  END Tile_X0Y0_EE4END[5]
  PIN Tile_X0Y0_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 0.800 355.600 ;
    END
  END Tile_X0Y0_EE4END[6]
  PIN Tile_X0Y0_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 0.800 356.960 ;
    END
  END Tile_X0Y0_EE4END[7]
  PIN Tile_X0Y0_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 0.800 358.320 ;
    END
  END Tile_X0Y0_EE4END[8]
  PIN Tile_X0Y0_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 0.800 359.680 ;
    END
  END Tile_X0Y0_EE4END[9]
  PIN Tile_X0Y0_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 0.800 385.520 ;
    END
  END Tile_X0Y0_FrameData[0]
  PIN Tile_X0Y0_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 0.800 399.120 ;
    END
  END Tile_X0Y0_FrameData[10]
  PIN Tile_X0Y0_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 0.800 400.480 ;
    END
  END Tile_X0Y0_FrameData[11]
  PIN Tile_X0Y0_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 0.800 401.840 ;
    END
  END Tile_X0Y0_FrameData[12]
  PIN Tile_X0Y0_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 0.800 403.200 ;
    END
  END Tile_X0Y0_FrameData[13]
  PIN Tile_X0Y0_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 0.800 404.560 ;
    END
  END Tile_X0Y0_FrameData[14]
  PIN Tile_X0Y0_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 0.800 405.920 ;
    END
  END Tile_X0Y0_FrameData[15]
  PIN Tile_X0Y0_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 0.800 407.280 ;
    END
  END Tile_X0Y0_FrameData[16]
  PIN Tile_X0Y0_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 0.800 408.640 ;
    END
  END Tile_X0Y0_FrameData[17]
  PIN Tile_X0Y0_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 0.800 410.000 ;
    END
  END Tile_X0Y0_FrameData[18]
  PIN Tile_X0Y0_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 0.800 411.360 ;
    END
  END Tile_X0Y0_FrameData[19]
  PIN Tile_X0Y0_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 0.800 386.880 ;
    END
  END Tile_X0Y0_FrameData[1]
  PIN Tile_X0Y0_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 0.800 412.720 ;
    END
  END Tile_X0Y0_FrameData[20]
  PIN Tile_X0Y0_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 0.800 414.080 ;
    END
  END Tile_X0Y0_FrameData[21]
  PIN Tile_X0Y0_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 0.800 415.440 ;
    END
  END Tile_X0Y0_FrameData[22]
  PIN Tile_X0Y0_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 0.800 416.800 ;
    END
  END Tile_X0Y0_FrameData[23]
  PIN Tile_X0Y0_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 0.800 418.160 ;
    END
  END Tile_X0Y0_FrameData[24]
  PIN Tile_X0Y0_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 0.800 419.520 ;
    END
  END Tile_X0Y0_FrameData[25]
  PIN Tile_X0Y0_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 0.800 420.880 ;
    END
  END Tile_X0Y0_FrameData[26]
  PIN Tile_X0Y0_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 0.800 422.240 ;
    END
  END Tile_X0Y0_FrameData[27]
  PIN Tile_X0Y0_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 0.800 423.600 ;
    END
  END Tile_X0Y0_FrameData[28]
  PIN Tile_X0Y0_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 0.800 424.960 ;
    END
  END Tile_X0Y0_FrameData[29]
  PIN Tile_X0Y0_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 0.800 388.240 ;
    END
  END Tile_X0Y0_FrameData[2]
  PIN Tile_X0Y0_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 0.800 426.320 ;
    END
  END Tile_X0Y0_FrameData[30]
  PIN Tile_X0Y0_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 0.800 427.680 ;
    END
  END Tile_X0Y0_FrameData[31]
  PIN Tile_X0Y0_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 0.800 389.600 ;
    END
  END Tile_X0Y0_FrameData[3]
  PIN Tile_X0Y0_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 0.800 390.960 ;
    END
  END Tile_X0Y0_FrameData[4]
  PIN Tile_X0Y0_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 0.800 392.320 ;
    END
  END Tile_X0Y0_FrameData[5]
  PIN Tile_X0Y0_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 0.800 393.680 ;
    END
  END Tile_X0Y0_FrameData[6]
  PIN Tile_X0Y0_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 0.800 395.040 ;
    END
  END Tile_X0Y0_FrameData[7]
  PIN Tile_X0Y0_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 0.800 396.400 ;
    END
  END Tile_X0Y0_FrameData[8]
  PIN Tile_X0Y0_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 0.800 397.760 ;
    END
  END Tile_X0Y0_FrameData[9]
  PIN Tile_X0Y0_FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 384.920 225.000 385.520 ;
    END
  END Tile_X0Y0_FrameData_O[0]
  PIN Tile_X0Y0_FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 398.520 225.000 399.120 ;
    END
  END Tile_X0Y0_FrameData_O[10]
  PIN Tile_X0Y0_FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 399.880 225.000 400.480 ;
    END
  END Tile_X0Y0_FrameData_O[11]
  PIN Tile_X0Y0_FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 401.240 225.000 401.840 ;
    END
  END Tile_X0Y0_FrameData_O[12]
  PIN Tile_X0Y0_FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 402.600 225.000 403.200 ;
    END
  END Tile_X0Y0_FrameData_O[13]
  PIN Tile_X0Y0_FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 403.960 225.000 404.560 ;
    END
  END Tile_X0Y0_FrameData_O[14]
  PIN Tile_X0Y0_FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 405.320 225.000 405.920 ;
    END
  END Tile_X0Y0_FrameData_O[15]
  PIN Tile_X0Y0_FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 406.680 225.000 407.280 ;
    END
  END Tile_X0Y0_FrameData_O[16]
  PIN Tile_X0Y0_FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 408.040 225.000 408.640 ;
    END
  END Tile_X0Y0_FrameData_O[17]
  PIN Tile_X0Y0_FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 409.400 225.000 410.000 ;
    END
  END Tile_X0Y0_FrameData_O[18]
  PIN Tile_X0Y0_FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 410.760 225.000 411.360 ;
    END
  END Tile_X0Y0_FrameData_O[19]
  PIN Tile_X0Y0_FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 386.280 225.000 386.880 ;
    END
  END Tile_X0Y0_FrameData_O[1]
  PIN Tile_X0Y0_FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 412.120 225.000 412.720 ;
    END
  END Tile_X0Y0_FrameData_O[20]
  PIN Tile_X0Y0_FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 413.480 225.000 414.080 ;
    END
  END Tile_X0Y0_FrameData_O[21]
  PIN Tile_X0Y0_FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 414.840 225.000 415.440 ;
    END
  END Tile_X0Y0_FrameData_O[22]
  PIN Tile_X0Y0_FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 416.200 225.000 416.800 ;
    END
  END Tile_X0Y0_FrameData_O[23]
  PIN Tile_X0Y0_FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 417.560 225.000 418.160 ;
    END
  END Tile_X0Y0_FrameData_O[24]
  PIN Tile_X0Y0_FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 418.920 225.000 419.520 ;
    END
  END Tile_X0Y0_FrameData_O[25]
  PIN Tile_X0Y0_FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 420.280 225.000 420.880 ;
    END
  END Tile_X0Y0_FrameData_O[26]
  PIN Tile_X0Y0_FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 421.640 225.000 422.240 ;
    END
  END Tile_X0Y0_FrameData_O[27]
  PIN Tile_X0Y0_FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 423.000 225.000 423.600 ;
    END
  END Tile_X0Y0_FrameData_O[28]
  PIN Tile_X0Y0_FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 424.360 225.000 424.960 ;
    END
  END Tile_X0Y0_FrameData_O[29]
  PIN Tile_X0Y0_FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 387.640 225.000 388.240 ;
    END
  END Tile_X0Y0_FrameData_O[2]
  PIN Tile_X0Y0_FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 425.720 225.000 426.320 ;
    END
  END Tile_X0Y0_FrameData_O[30]
  PIN Tile_X0Y0_FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 427.080 225.000 427.680 ;
    END
  END Tile_X0Y0_FrameData_O[31]
  PIN Tile_X0Y0_FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 389.000 225.000 389.600 ;
    END
  END Tile_X0Y0_FrameData_O[3]
  PIN Tile_X0Y0_FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 390.360 225.000 390.960 ;
    END
  END Tile_X0Y0_FrameData_O[4]
  PIN Tile_X0Y0_FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 391.720 225.000 392.320 ;
    END
  END Tile_X0Y0_FrameData_O[5]
  PIN Tile_X0Y0_FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 393.080 225.000 393.680 ;
    END
  END Tile_X0Y0_FrameData_O[6]
  PIN Tile_X0Y0_FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 394.440 225.000 395.040 ;
    END
  END Tile_X0Y0_FrameData_O[7]
  PIN Tile_X0Y0_FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 395.800 225.000 396.400 ;
    END
  END Tile_X0Y0_FrameData_O[8]
  PIN Tile_X0Y0_FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 397.160 225.000 397.760 ;
    END
  END Tile_X0Y0_FrameData_O[9]
  PIN Tile_X0Y0_FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 171.670 449.200 171.950 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[0]
  PIN Tile_X0Y0_FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 185.470 449.200 185.750 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[10]
  PIN Tile_X0Y0_FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 186.850 449.200 187.130 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[11]
  PIN Tile_X0Y0_FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 188.230 449.200 188.510 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[12]
  PIN Tile_X0Y0_FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 189.610 449.200 189.890 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[13]
  PIN Tile_X0Y0_FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 190.990 449.200 191.270 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[14]
  PIN Tile_X0Y0_FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 192.370 449.200 192.650 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[15]
  PIN Tile_X0Y0_FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 193.750 449.200 194.030 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[16]
  PIN Tile_X0Y0_FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 195.130 449.200 195.410 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[17]
  PIN Tile_X0Y0_FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 196.510 449.200 196.790 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[18]
  PIN Tile_X0Y0_FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 197.890 449.200 198.170 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[19]
  PIN Tile_X0Y0_FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 173.050 449.200 173.330 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[1]
  PIN Tile_X0Y0_FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 174.430 449.200 174.710 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[2]
  PIN Tile_X0Y0_FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 175.810 449.200 176.090 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[3]
  PIN Tile_X0Y0_FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 177.190 449.200 177.470 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[4]
  PIN Tile_X0Y0_FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 178.570 449.200 178.850 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[5]
  PIN Tile_X0Y0_FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 179.950 449.200 180.230 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[6]
  PIN Tile_X0Y0_FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 181.330 449.200 181.610 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[7]
  PIN Tile_X0Y0_FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 182.710 449.200 182.990 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[8]
  PIN Tile_X0Y0_FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 184.090 449.200 184.370 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[9]
  PIN Tile_X0Y0_N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 26.770 449.200 27.050 450.000 ;
    END
  END Tile_X0Y0_N1BEG[0]
  PIN Tile_X0Y0_N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 28.150 449.200 28.430 450.000 ;
    END
  END Tile_X0Y0_N1BEG[1]
  PIN Tile_X0Y0_N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.530 449.200 29.810 450.000 ;
    END
  END Tile_X0Y0_N1BEG[2]
  PIN Tile_X0Y0_N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 30.910 449.200 31.190 450.000 ;
    END
  END Tile_X0Y0_N1BEG[3]
  PIN Tile_X0Y0_N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 449.200 32.570 450.000 ;
    END
  END Tile_X0Y0_N2BEG[0]
  PIN Tile_X0Y0_N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 33.670 449.200 33.950 450.000 ;
    END
  END Tile_X0Y0_N2BEG[1]
  PIN Tile_X0Y0_N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.050 449.200 35.330 450.000 ;
    END
  END Tile_X0Y0_N2BEG[2]
  PIN Tile_X0Y0_N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 36.430 449.200 36.710 450.000 ;
    END
  END Tile_X0Y0_N2BEG[3]
  PIN Tile_X0Y0_N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 37.810 449.200 38.090 450.000 ;
    END
  END Tile_X0Y0_N2BEG[4]
  PIN Tile_X0Y0_N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 39.190 449.200 39.470 450.000 ;
    END
  END Tile_X0Y0_N2BEG[5]
  PIN Tile_X0Y0_N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 40.570 449.200 40.850 450.000 ;
    END
  END Tile_X0Y0_N2BEG[6]
  PIN Tile_X0Y0_N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.950 449.200 42.230 450.000 ;
    END
  END Tile_X0Y0_N2BEG[7]
  PIN Tile_X0Y0_N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 43.330 449.200 43.610 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[0]
  PIN Tile_X0Y0_N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 44.710 449.200 44.990 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[1]
  PIN Tile_X0Y0_N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 46.090 449.200 46.370 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[2]
  PIN Tile_X0Y0_N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 47.470 449.200 47.750 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[3]
  PIN Tile_X0Y0_N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.850 449.200 49.130 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[4]
  PIN Tile_X0Y0_N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 50.230 449.200 50.510 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[5]
  PIN Tile_X0Y0_N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 449.200 51.890 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[6]
  PIN Tile_X0Y0_N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 52.990 449.200 53.270 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[7]
  PIN Tile_X0Y0_N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.370 449.200 54.650 450.000 ;
    END
  END Tile_X0Y0_N4BEG[0]
  PIN Tile_X0Y0_N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 68.170 449.200 68.450 450.000 ;
    END
  END Tile_X0Y0_N4BEG[10]
  PIN Tile_X0Y0_N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 69.550 449.200 69.830 450.000 ;
    END
  END Tile_X0Y0_N4BEG[11]
  PIN Tile_X0Y0_N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.930 449.200 71.210 450.000 ;
    END
  END Tile_X0Y0_N4BEG[12]
  PIN Tile_X0Y0_N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 72.310 449.200 72.590 450.000 ;
    END
  END Tile_X0Y0_N4BEG[13]
  PIN Tile_X0Y0_N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 73.690 449.200 73.970 450.000 ;
    END
  END Tile_X0Y0_N4BEG[14]
  PIN Tile_X0Y0_N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 75.070 449.200 75.350 450.000 ;
    END
  END Tile_X0Y0_N4BEG[15]
  PIN Tile_X0Y0_N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 55.750 449.200 56.030 450.000 ;
    END
  END Tile_X0Y0_N4BEG[1]
  PIN Tile_X0Y0_N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 57.130 449.200 57.410 450.000 ;
    END
  END Tile_X0Y0_N4BEG[2]
  PIN Tile_X0Y0_N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 58.510 449.200 58.790 450.000 ;
    END
  END Tile_X0Y0_N4BEG[3]
  PIN Tile_X0Y0_N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 59.890 449.200 60.170 450.000 ;
    END
  END Tile_X0Y0_N4BEG[4]
  PIN Tile_X0Y0_N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.270 449.200 61.550 450.000 ;
    END
  END Tile_X0Y0_N4BEG[5]
  PIN Tile_X0Y0_N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 62.650 449.200 62.930 450.000 ;
    END
  END Tile_X0Y0_N4BEG[6]
  PIN Tile_X0Y0_N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.030 449.200 64.310 450.000 ;
    END
  END Tile_X0Y0_N4BEG[7]
  PIN Tile_X0Y0_N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.410 449.200 65.690 450.000 ;
    END
  END Tile_X0Y0_N4BEG[8]
  PIN Tile_X0Y0_N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 66.790 449.200 67.070 450.000 ;
    END
  END Tile_X0Y0_N4BEG[9]
  PIN Tile_X0Y0_NN4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 76.450 449.200 76.730 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[0]
  PIN Tile_X0Y0_NN4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.250 449.200 90.530 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[10]
  PIN Tile_X0Y0_NN4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 91.630 449.200 91.910 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[11]
  PIN Tile_X0Y0_NN4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.010 449.200 93.290 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[12]
  PIN Tile_X0Y0_NN4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 94.390 449.200 94.670 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[13]
  PIN Tile_X0Y0_NN4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 95.770 449.200 96.050 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[14]
  PIN Tile_X0Y0_NN4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 97.150 449.200 97.430 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[15]
  PIN Tile_X0Y0_NN4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.830 449.200 78.110 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[1]
  PIN Tile_X0Y0_NN4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 79.210 449.200 79.490 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[2]
  PIN Tile_X0Y0_NN4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 449.200 80.870 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[3]
  PIN Tile_X0Y0_NN4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 81.970 449.200 82.250 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[4]
  PIN Tile_X0Y0_NN4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.350 449.200 83.630 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[5]
  PIN Tile_X0Y0_NN4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 84.730 449.200 85.010 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[6]
  PIN Tile_X0Y0_NN4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 86.110 449.200 86.390 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[7]
  PIN Tile_X0Y0_NN4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.490 449.200 87.770 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[8]
  PIN Tile_X0Y0_NN4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 88.870 449.200 89.150 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[9]
  PIN Tile_X0Y0_S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 98.530 449.200 98.810 450.000 ;
    END
  END Tile_X0Y0_S1END[0]
  PIN Tile_X0Y0_S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 449.200 100.190 450.000 ;
    END
  END Tile_X0Y0_S1END[1]
  PIN Tile_X0Y0_S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 101.290 449.200 101.570 450.000 ;
    END
  END Tile_X0Y0_S1END[2]
  PIN Tile_X0Y0_S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 102.670 449.200 102.950 450.000 ;
    END
  END Tile_X0Y0_S1END[3]
  PIN Tile_X0Y0_S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 104.050 449.200 104.330 450.000 ;
    END
  END Tile_X0Y0_S2END[0]
  PIN Tile_X0Y0_S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 105.430 449.200 105.710 450.000 ;
    END
  END Tile_X0Y0_S2END[1]
  PIN Tile_X0Y0_S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 106.810 449.200 107.090 450.000 ;
    END
  END Tile_X0Y0_S2END[2]
  PIN Tile_X0Y0_S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 108.190 449.200 108.470 450.000 ;
    END
  END Tile_X0Y0_S2END[3]
  PIN Tile_X0Y0_S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 449.200 109.850 450.000 ;
    END
  END Tile_X0Y0_S2END[4]
  PIN Tile_X0Y0_S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 110.950 449.200 111.230 450.000 ;
    END
  END Tile_X0Y0_S2END[5]
  PIN Tile_X0Y0_S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 112.330 449.200 112.610 450.000 ;
    END
  END Tile_X0Y0_S2END[6]
  PIN Tile_X0Y0_S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 113.710 449.200 113.990 450.000 ;
    END
  END Tile_X0Y0_S2END[7]
  PIN Tile_X0Y0_S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 115.090 449.200 115.370 450.000 ;
    END
  END Tile_X0Y0_S2MID[0]
  PIN Tile_X0Y0_S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 116.470 449.200 116.750 450.000 ;
    END
  END Tile_X0Y0_S2MID[1]
  PIN Tile_X0Y0_S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 117.850 449.200 118.130 450.000 ;
    END
  END Tile_X0Y0_S2MID[2]
  PIN Tile_X0Y0_S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 449.200 119.510 450.000 ;
    END
  END Tile_X0Y0_S2MID[3]
  PIN Tile_X0Y0_S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 120.610 449.200 120.890 450.000 ;
    END
  END Tile_X0Y0_S2MID[4]
  PIN Tile_X0Y0_S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 121.990 449.200 122.270 450.000 ;
    END
  END Tile_X0Y0_S2MID[5]
  PIN Tile_X0Y0_S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 123.370 449.200 123.650 450.000 ;
    END
  END Tile_X0Y0_S2MID[6]
  PIN Tile_X0Y0_S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 124.750 449.200 125.030 450.000 ;
    END
  END Tile_X0Y0_S2MID[7]
  PIN Tile_X0Y0_S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 126.130 449.200 126.410 450.000 ;
    END
  END Tile_X0Y0_S4END[0]
  PIN Tile_X0Y0_S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 139.930 449.200 140.210 450.000 ;
    END
  END Tile_X0Y0_S4END[10]
  PIN Tile_X0Y0_S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 141.310 449.200 141.590 450.000 ;
    END
  END Tile_X0Y0_S4END[11]
  PIN Tile_X0Y0_S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 142.690 449.200 142.970 450.000 ;
    END
  END Tile_X0Y0_S4END[12]
  PIN Tile_X0Y0_S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.070 449.200 144.350 450.000 ;
    END
  END Tile_X0Y0_S4END[13]
  PIN Tile_X0Y0_S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 145.450 449.200 145.730 450.000 ;
    END
  END Tile_X0Y0_S4END[14]
  PIN Tile_X0Y0_S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 146.830 449.200 147.110 450.000 ;
    END
  END Tile_X0Y0_S4END[15]
  PIN Tile_X0Y0_S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 127.510 449.200 127.790 450.000 ;
    END
  END Tile_X0Y0_S4END[1]
  PIN Tile_X0Y0_S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 449.200 129.170 450.000 ;
    END
  END Tile_X0Y0_S4END[2]
  PIN Tile_X0Y0_S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 130.270 449.200 130.550 450.000 ;
    END
  END Tile_X0Y0_S4END[3]
  PIN Tile_X0Y0_S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 131.650 449.200 131.930 450.000 ;
    END
  END Tile_X0Y0_S4END[4]
  PIN Tile_X0Y0_S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 133.030 449.200 133.310 450.000 ;
    END
  END Tile_X0Y0_S4END[5]
  PIN Tile_X0Y0_S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 134.410 449.200 134.690 450.000 ;
    END
  END Tile_X0Y0_S4END[6]
  PIN Tile_X0Y0_S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 135.790 449.200 136.070 450.000 ;
    END
  END Tile_X0Y0_S4END[7]
  PIN Tile_X0Y0_S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 137.170 449.200 137.450 450.000 ;
    END
  END Tile_X0Y0_S4END[8]
  PIN Tile_X0Y0_S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 449.200 138.830 450.000 ;
    END
  END Tile_X0Y0_S4END[9]
  PIN Tile_X0Y0_SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 449.200 148.490 450.000 ;
    END
  END Tile_X0Y0_SS4END[0]
  PIN Tile_X0Y0_SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 162.010 449.200 162.290 450.000 ;
    END
  END Tile_X0Y0_SS4END[10]
  PIN Tile_X0Y0_SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 163.390 449.200 163.670 450.000 ;
    END
  END Tile_X0Y0_SS4END[11]
  PIN Tile_X0Y0_SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 164.770 449.200 165.050 450.000 ;
    END
  END Tile_X0Y0_SS4END[12]
  PIN Tile_X0Y0_SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 166.150 449.200 166.430 450.000 ;
    END
  END Tile_X0Y0_SS4END[13]
  PIN Tile_X0Y0_SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 449.200 167.810 450.000 ;
    END
  END Tile_X0Y0_SS4END[14]
  PIN Tile_X0Y0_SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 168.910 449.200 169.190 450.000 ;
    END
  END Tile_X0Y0_SS4END[15]
  PIN Tile_X0Y0_SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 149.590 449.200 149.870 450.000 ;
    END
  END Tile_X0Y0_SS4END[1]
  PIN Tile_X0Y0_SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 150.970 449.200 151.250 450.000 ;
    END
  END Tile_X0Y0_SS4END[2]
  PIN Tile_X0Y0_SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 152.350 449.200 152.630 450.000 ;
    END
  END Tile_X0Y0_SS4END[3]
  PIN Tile_X0Y0_SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 153.730 449.200 154.010 450.000 ;
    END
  END Tile_X0Y0_SS4END[4]
  PIN Tile_X0Y0_SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 155.110 449.200 155.390 450.000 ;
    END
  END Tile_X0Y0_SS4END[5]
  PIN Tile_X0Y0_SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 156.490 449.200 156.770 450.000 ;
    END
  END Tile_X0Y0_SS4END[6]
  PIN Tile_X0Y0_SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 157.870 449.200 158.150 450.000 ;
    END
  END Tile_X0Y0_SS4END[7]
  PIN Tile_X0Y0_SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 159.250 449.200 159.530 450.000 ;
    END
  END Tile_X0Y0_SS4END[8]
  PIN Tile_X0Y0_SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 160.630 449.200 160.910 450.000 ;
    END
  END Tile_X0Y0_SS4END[9]
  PIN Tile_X0Y0_UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 170.290 449.200 170.570 450.000 ;
    END
  END Tile_X0Y0_UserCLKo
  PIN Tile_X0Y0_W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 0.800 254.960 ;
    END
  END Tile_X0Y0_W1BEG[0]
  PIN Tile_X0Y0_W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 0.800 256.320 ;
    END
  END Tile_X0Y0_W1BEG[1]
  PIN Tile_X0Y0_W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 0.800 257.680 ;
    END
  END Tile_X0Y0_W1BEG[2]
  PIN Tile_X0Y0_W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 0.800 259.040 ;
    END
  END Tile_X0Y0_W1BEG[3]
  PIN Tile_X0Y0_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 254.360 225.000 254.960 ;
    END
  END Tile_X0Y0_W1END[0]
  PIN Tile_X0Y0_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 255.720 225.000 256.320 ;
    END
  END Tile_X0Y0_W1END[1]
  PIN Tile_X0Y0_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 257.080 225.000 257.680 ;
    END
  END Tile_X0Y0_W1END[2]
  PIN Tile_X0Y0_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 258.440 225.000 259.040 ;
    END
  END Tile_X0Y0_W1END[3]
  PIN Tile_X0Y0_W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 0.800 260.400 ;
    END
  END Tile_X0Y0_W2BEG[0]
  PIN Tile_X0Y0_W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 0.800 261.760 ;
    END
  END Tile_X0Y0_W2BEG[1]
  PIN Tile_X0Y0_W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 0.800 263.120 ;
    END
  END Tile_X0Y0_W2BEG[2]
  PIN Tile_X0Y0_W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 0.800 264.480 ;
    END
  END Tile_X0Y0_W2BEG[3]
  PIN Tile_X0Y0_W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 0.800 265.840 ;
    END
  END Tile_X0Y0_W2BEG[4]
  PIN Tile_X0Y0_W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 0.800 267.200 ;
    END
  END Tile_X0Y0_W2BEG[5]
  PIN Tile_X0Y0_W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 0.800 268.560 ;
    END
  END Tile_X0Y0_W2BEG[6]
  PIN Tile_X0Y0_W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 0.800 269.920 ;
    END
  END Tile_X0Y0_W2BEG[7]
  PIN Tile_X0Y0_W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 0.800 271.280 ;
    END
  END Tile_X0Y0_W2BEGb[0]
  PIN Tile_X0Y0_W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 0.800 272.640 ;
    END
  END Tile_X0Y0_W2BEGb[1]
  PIN Tile_X0Y0_W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 0.800 274.000 ;
    END
  END Tile_X0Y0_W2BEGb[2]
  PIN Tile_X0Y0_W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 0.800 275.360 ;
    END
  END Tile_X0Y0_W2BEGb[3]
  PIN Tile_X0Y0_W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 0.800 276.720 ;
    END
  END Tile_X0Y0_W2BEGb[4]
  PIN Tile_X0Y0_W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 0.800 278.080 ;
    END
  END Tile_X0Y0_W2BEGb[5]
  PIN Tile_X0Y0_W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 0.800 279.440 ;
    END
  END Tile_X0Y0_W2BEGb[6]
  PIN Tile_X0Y0_W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 0.800 280.800 ;
    END
  END Tile_X0Y0_W2BEGb[7]
  PIN Tile_X0Y0_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 270.680 225.000 271.280 ;
    END
  END Tile_X0Y0_W2END[0]
  PIN Tile_X0Y0_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 272.040 225.000 272.640 ;
    END
  END Tile_X0Y0_W2END[1]
  PIN Tile_X0Y0_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 273.400 225.000 274.000 ;
    END
  END Tile_X0Y0_W2END[2]
  PIN Tile_X0Y0_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 274.760 225.000 275.360 ;
    END
  END Tile_X0Y0_W2END[3]
  PIN Tile_X0Y0_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 276.120 225.000 276.720 ;
    END
  END Tile_X0Y0_W2END[4]
  PIN Tile_X0Y0_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 277.480 225.000 278.080 ;
    END
  END Tile_X0Y0_W2END[5]
  PIN Tile_X0Y0_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 278.840 225.000 279.440 ;
    END
  END Tile_X0Y0_W2END[6]
  PIN Tile_X0Y0_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 280.200 225.000 280.800 ;
    END
  END Tile_X0Y0_W2END[7]
  PIN Tile_X0Y0_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 259.800 225.000 260.400 ;
    END
  END Tile_X0Y0_W2MID[0]
  PIN Tile_X0Y0_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 261.160 225.000 261.760 ;
    END
  END Tile_X0Y0_W2MID[1]
  PIN Tile_X0Y0_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 262.520 225.000 263.120 ;
    END
  END Tile_X0Y0_W2MID[2]
  PIN Tile_X0Y0_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 263.880 225.000 264.480 ;
    END
  END Tile_X0Y0_W2MID[3]
  PIN Tile_X0Y0_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 265.240 225.000 265.840 ;
    END
  END Tile_X0Y0_W2MID[4]
  PIN Tile_X0Y0_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 266.600 225.000 267.200 ;
    END
  END Tile_X0Y0_W2MID[5]
  PIN Tile_X0Y0_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 267.960 225.000 268.560 ;
    END
  END Tile_X0Y0_W2MID[6]
  PIN Tile_X0Y0_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 269.320 225.000 269.920 ;
    END
  END Tile_X0Y0_W2MID[7]
  PIN Tile_X0Y0_W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 0.800 303.920 ;
    END
  END Tile_X0Y0_W6BEG[0]
  PIN Tile_X0Y0_W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 0.800 317.520 ;
    END
  END Tile_X0Y0_W6BEG[10]
  PIN Tile_X0Y0_W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 0.800 318.880 ;
    END
  END Tile_X0Y0_W6BEG[11]
  PIN Tile_X0Y0_W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 0.800 305.280 ;
    END
  END Tile_X0Y0_W6BEG[1]
  PIN Tile_X0Y0_W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 0.800 306.640 ;
    END
  END Tile_X0Y0_W6BEG[2]
  PIN Tile_X0Y0_W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 0.800 308.000 ;
    END
  END Tile_X0Y0_W6BEG[3]
  PIN Tile_X0Y0_W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 0.800 309.360 ;
    END
  END Tile_X0Y0_W6BEG[4]
  PIN Tile_X0Y0_W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 0.800 310.720 ;
    END
  END Tile_X0Y0_W6BEG[5]
  PIN Tile_X0Y0_W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 0.800 312.080 ;
    END
  END Tile_X0Y0_W6BEG[6]
  PIN Tile_X0Y0_W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 0.800 313.440 ;
    END
  END Tile_X0Y0_W6BEG[7]
  PIN Tile_X0Y0_W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 0.800 314.800 ;
    END
  END Tile_X0Y0_W6BEG[8]
  PIN Tile_X0Y0_W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 0.800 316.160 ;
    END
  END Tile_X0Y0_W6BEG[9]
  PIN Tile_X0Y0_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 303.320 225.000 303.920 ;
    END
  END Tile_X0Y0_W6END[0]
  PIN Tile_X0Y0_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 316.920 225.000 317.520 ;
    END
  END Tile_X0Y0_W6END[10]
  PIN Tile_X0Y0_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 318.280 225.000 318.880 ;
    END
  END Tile_X0Y0_W6END[11]
  PIN Tile_X0Y0_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 304.680 225.000 305.280 ;
    END
  END Tile_X0Y0_W6END[1]
  PIN Tile_X0Y0_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 306.040 225.000 306.640 ;
    END
  END Tile_X0Y0_W6END[2]
  PIN Tile_X0Y0_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 307.400 225.000 308.000 ;
    END
  END Tile_X0Y0_W6END[3]
  PIN Tile_X0Y0_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 308.760 225.000 309.360 ;
    END
  END Tile_X0Y0_W6END[4]
  PIN Tile_X0Y0_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 310.120 225.000 310.720 ;
    END
  END Tile_X0Y0_W6END[5]
  PIN Tile_X0Y0_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 311.480 225.000 312.080 ;
    END
  END Tile_X0Y0_W6END[6]
  PIN Tile_X0Y0_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 312.840 225.000 313.440 ;
    END
  END Tile_X0Y0_W6END[7]
  PIN Tile_X0Y0_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 314.200 225.000 314.800 ;
    END
  END Tile_X0Y0_W6END[8]
  PIN Tile_X0Y0_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 315.560 225.000 316.160 ;
    END
  END Tile_X0Y0_W6END[9]
  PIN Tile_X0Y0_WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 0.800 282.160 ;
    END
  END Tile_X0Y0_WW4BEG[0]
  PIN Tile_X0Y0_WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 0.800 295.760 ;
    END
  END Tile_X0Y0_WW4BEG[10]
  PIN Tile_X0Y0_WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 0.800 297.120 ;
    END
  END Tile_X0Y0_WW4BEG[11]
  PIN Tile_X0Y0_WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 0.800 298.480 ;
    END
  END Tile_X0Y0_WW4BEG[12]
  PIN Tile_X0Y0_WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 0.800 299.840 ;
    END
  END Tile_X0Y0_WW4BEG[13]
  PIN Tile_X0Y0_WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 0.800 301.200 ;
    END
  END Tile_X0Y0_WW4BEG[14]
  PIN Tile_X0Y0_WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 0.800 302.560 ;
    END
  END Tile_X0Y0_WW4BEG[15]
  PIN Tile_X0Y0_WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 0.800 283.520 ;
    END
  END Tile_X0Y0_WW4BEG[1]
  PIN Tile_X0Y0_WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 0.800 284.880 ;
    END
  END Tile_X0Y0_WW4BEG[2]
  PIN Tile_X0Y0_WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 0.800 286.240 ;
    END
  END Tile_X0Y0_WW4BEG[3]
  PIN Tile_X0Y0_WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 0.800 287.600 ;
    END
  END Tile_X0Y0_WW4BEG[4]
  PIN Tile_X0Y0_WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 0.800 288.960 ;
    END
  END Tile_X0Y0_WW4BEG[5]
  PIN Tile_X0Y0_WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 0.800 290.320 ;
    END
  END Tile_X0Y0_WW4BEG[6]
  PIN Tile_X0Y0_WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 0.800 291.680 ;
    END
  END Tile_X0Y0_WW4BEG[7]
  PIN Tile_X0Y0_WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 0.800 293.040 ;
    END
  END Tile_X0Y0_WW4BEG[8]
  PIN Tile_X0Y0_WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 0.800 294.400 ;
    END
  END Tile_X0Y0_WW4BEG[9]
  PIN Tile_X0Y0_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 281.560 225.000 282.160 ;
    END
  END Tile_X0Y0_WW4END[0]
  PIN Tile_X0Y0_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 295.160 225.000 295.760 ;
    END
  END Tile_X0Y0_WW4END[10]
  PIN Tile_X0Y0_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 296.520 225.000 297.120 ;
    END
  END Tile_X0Y0_WW4END[11]
  PIN Tile_X0Y0_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 297.880 225.000 298.480 ;
    END
  END Tile_X0Y0_WW4END[12]
  PIN Tile_X0Y0_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 299.240 225.000 299.840 ;
    END
  END Tile_X0Y0_WW4END[13]
  PIN Tile_X0Y0_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 300.600 225.000 301.200 ;
    END
  END Tile_X0Y0_WW4END[14]
  PIN Tile_X0Y0_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 301.960 225.000 302.560 ;
    END
  END Tile_X0Y0_WW4END[15]
  PIN Tile_X0Y0_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 282.920 225.000 283.520 ;
    END
  END Tile_X0Y0_WW4END[1]
  PIN Tile_X0Y0_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 284.280 225.000 284.880 ;
    END
  END Tile_X0Y0_WW4END[2]
  PIN Tile_X0Y0_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 285.640 225.000 286.240 ;
    END
  END Tile_X0Y0_WW4END[3]
  PIN Tile_X0Y0_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 287.000 225.000 287.600 ;
    END
  END Tile_X0Y0_WW4END[4]
  PIN Tile_X0Y0_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 288.360 225.000 288.960 ;
    END
  END Tile_X0Y0_WW4END[5]
  PIN Tile_X0Y0_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 289.720 225.000 290.320 ;
    END
  END Tile_X0Y0_WW4END[6]
  PIN Tile_X0Y0_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 291.080 225.000 291.680 ;
    END
  END Tile_X0Y0_WW4END[7]
  PIN Tile_X0Y0_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 292.440 225.000 293.040 ;
    END
  END Tile_X0Y0_WW4END[8]
  PIN Tile_X0Y0_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 293.800 225.000 294.400 ;
    END
  END Tile_X0Y0_WW4END[9]
  PIN Tile_X0Y1_E1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 89.800 225.000 90.400 ;
    END
  END Tile_X0Y1_E1BEG[0]
  PIN Tile_X0Y1_E1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 91.160 225.000 91.760 ;
    END
  END Tile_X0Y1_E1BEG[1]
  PIN Tile_X0Y1_E1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 92.520 225.000 93.120 ;
    END
  END Tile_X0Y1_E1BEG[2]
  PIN Tile_X0Y1_E1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 93.880 225.000 94.480 ;
    END
  END Tile_X0Y1_E1BEG[3]
  PIN Tile_X0Y1_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 0.800 90.400 ;
    END
  END Tile_X0Y1_E1END[0]
  PIN Tile_X0Y1_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 0.800 91.760 ;
    END
  END Tile_X0Y1_E1END[1]
  PIN Tile_X0Y1_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 0.800 93.120 ;
    END
  END Tile_X0Y1_E1END[2]
  PIN Tile_X0Y1_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 0.800 94.480 ;
    END
  END Tile_X0Y1_E1END[3]
  PIN Tile_X0Y1_E2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 95.240 225.000 95.840 ;
    END
  END Tile_X0Y1_E2BEG[0]
  PIN Tile_X0Y1_E2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 96.600 225.000 97.200 ;
    END
  END Tile_X0Y1_E2BEG[1]
  PIN Tile_X0Y1_E2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 97.960 225.000 98.560 ;
    END
  END Tile_X0Y1_E2BEG[2]
  PIN Tile_X0Y1_E2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 99.320 225.000 99.920 ;
    END
  END Tile_X0Y1_E2BEG[3]
  PIN Tile_X0Y1_E2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 100.680 225.000 101.280 ;
    END
  END Tile_X0Y1_E2BEG[4]
  PIN Tile_X0Y1_E2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 102.040 225.000 102.640 ;
    END
  END Tile_X0Y1_E2BEG[5]
  PIN Tile_X0Y1_E2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 103.400 225.000 104.000 ;
    END
  END Tile_X0Y1_E2BEG[6]
  PIN Tile_X0Y1_E2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 104.760 225.000 105.360 ;
    END
  END Tile_X0Y1_E2BEG[7]
  PIN Tile_X0Y1_E2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 106.120 225.000 106.720 ;
    END
  END Tile_X0Y1_E2BEGb[0]
  PIN Tile_X0Y1_E2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 107.480 225.000 108.080 ;
    END
  END Tile_X0Y1_E2BEGb[1]
  PIN Tile_X0Y1_E2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 108.840 225.000 109.440 ;
    END
  END Tile_X0Y1_E2BEGb[2]
  PIN Tile_X0Y1_E2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 110.200 225.000 110.800 ;
    END
  END Tile_X0Y1_E2BEGb[3]
  PIN Tile_X0Y1_E2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 111.560 225.000 112.160 ;
    END
  END Tile_X0Y1_E2BEGb[4]
  PIN Tile_X0Y1_E2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 112.920 225.000 113.520 ;
    END
  END Tile_X0Y1_E2BEGb[5]
  PIN Tile_X0Y1_E2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 114.280 225.000 114.880 ;
    END
  END Tile_X0Y1_E2BEGb[6]
  PIN Tile_X0Y1_E2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 115.640 225.000 116.240 ;
    END
  END Tile_X0Y1_E2BEGb[7]
  PIN Tile_X0Y1_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 0.800 106.720 ;
    END
  END Tile_X0Y1_E2END[0]
  PIN Tile_X0Y1_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 0.800 108.080 ;
    END
  END Tile_X0Y1_E2END[1]
  PIN Tile_X0Y1_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 0.800 109.440 ;
    END
  END Tile_X0Y1_E2END[2]
  PIN Tile_X0Y1_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 0.800 110.800 ;
    END
  END Tile_X0Y1_E2END[3]
  PIN Tile_X0Y1_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 0.800 112.160 ;
    END
  END Tile_X0Y1_E2END[4]
  PIN Tile_X0Y1_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 0.800 113.520 ;
    END
  END Tile_X0Y1_E2END[5]
  PIN Tile_X0Y1_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 0.800 114.880 ;
    END
  END Tile_X0Y1_E2END[6]
  PIN Tile_X0Y1_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 0.800 116.240 ;
    END
  END Tile_X0Y1_E2END[7]
  PIN Tile_X0Y1_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 0.800 95.840 ;
    END
  END Tile_X0Y1_E2MID[0]
  PIN Tile_X0Y1_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 0.800 97.200 ;
    END
  END Tile_X0Y1_E2MID[1]
  PIN Tile_X0Y1_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 0.800 98.560 ;
    END
  END Tile_X0Y1_E2MID[2]
  PIN Tile_X0Y1_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 0.800 99.920 ;
    END
  END Tile_X0Y1_E2MID[3]
  PIN Tile_X0Y1_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 0.800 101.280 ;
    END
  END Tile_X0Y1_E2MID[4]
  PIN Tile_X0Y1_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 0.800 102.640 ;
    END
  END Tile_X0Y1_E2MID[5]
  PIN Tile_X0Y1_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 0.800 104.000 ;
    END
  END Tile_X0Y1_E2MID[6]
  PIN Tile_X0Y1_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 0.800 105.360 ;
    END
  END Tile_X0Y1_E2MID[7]
  PIN Tile_X0Y1_E6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 138.760 225.000 139.360 ;
    END
  END Tile_X0Y1_E6BEG[0]
  PIN Tile_X0Y1_E6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 152.360 225.000 152.960 ;
    END
  END Tile_X0Y1_E6BEG[10]
  PIN Tile_X0Y1_E6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 153.720 225.000 154.320 ;
    END
  END Tile_X0Y1_E6BEG[11]
  PIN Tile_X0Y1_E6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 140.120 225.000 140.720 ;
    END
  END Tile_X0Y1_E6BEG[1]
  PIN Tile_X0Y1_E6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 141.480 225.000 142.080 ;
    END
  END Tile_X0Y1_E6BEG[2]
  PIN Tile_X0Y1_E6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 142.840 225.000 143.440 ;
    END
  END Tile_X0Y1_E6BEG[3]
  PIN Tile_X0Y1_E6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 144.200 225.000 144.800 ;
    END
  END Tile_X0Y1_E6BEG[4]
  PIN Tile_X0Y1_E6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 145.560 225.000 146.160 ;
    END
  END Tile_X0Y1_E6BEG[5]
  PIN Tile_X0Y1_E6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 146.920 225.000 147.520 ;
    END
  END Tile_X0Y1_E6BEG[6]
  PIN Tile_X0Y1_E6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 148.280 225.000 148.880 ;
    END
  END Tile_X0Y1_E6BEG[7]
  PIN Tile_X0Y1_E6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 149.640 225.000 150.240 ;
    END
  END Tile_X0Y1_E6BEG[8]
  PIN Tile_X0Y1_E6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 151.000 225.000 151.600 ;
    END
  END Tile_X0Y1_E6BEG[9]
  PIN Tile_X0Y1_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 0.800 139.360 ;
    END
  END Tile_X0Y1_E6END[0]
  PIN Tile_X0Y1_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 0.800 152.960 ;
    END
  END Tile_X0Y1_E6END[10]
  PIN Tile_X0Y1_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 0.800 154.320 ;
    END
  END Tile_X0Y1_E6END[11]
  PIN Tile_X0Y1_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 0.800 140.720 ;
    END
  END Tile_X0Y1_E6END[1]
  PIN Tile_X0Y1_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 0.800 142.080 ;
    END
  END Tile_X0Y1_E6END[2]
  PIN Tile_X0Y1_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 0.800 143.440 ;
    END
  END Tile_X0Y1_E6END[3]
  PIN Tile_X0Y1_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 0.800 144.800 ;
    END
  END Tile_X0Y1_E6END[4]
  PIN Tile_X0Y1_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 0.800 146.160 ;
    END
  END Tile_X0Y1_E6END[5]
  PIN Tile_X0Y1_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 0.800 147.520 ;
    END
  END Tile_X0Y1_E6END[6]
  PIN Tile_X0Y1_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 0.800 148.880 ;
    END
  END Tile_X0Y1_E6END[7]
  PIN Tile_X0Y1_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 0.800 150.240 ;
    END
  END Tile_X0Y1_E6END[8]
  PIN Tile_X0Y1_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 0.800 151.600 ;
    END
  END Tile_X0Y1_E6END[9]
  PIN Tile_X0Y1_EE4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 117.000 225.000 117.600 ;
    END
  END Tile_X0Y1_EE4BEG[0]
  PIN Tile_X0Y1_EE4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 130.600 225.000 131.200 ;
    END
  END Tile_X0Y1_EE4BEG[10]
  PIN Tile_X0Y1_EE4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 131.960 225.000 132.560 ;
    END
  END Tile_X0Y1_EE4BEG[11]
  PIN Tile_X0Y1_EE4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 133.320 225.000 133.920 ;
    END
  END Tile_X0Y1_EE4BEG[12]
  PIN Tile_X0Y1_EE4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 134.680 225.000 135.280 ;
    END
  END Tile_X0Y1_EE4BEG[13]
  PIN Tile_X0Y1_EE4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 136.040 225.000 136.640 ;
    END
  END Tile_X0Y1_EE4BEG[14]
  PIN Tile_X0Y1_EE4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 137.400 225.000 138.000 ;
    END
  END Tile_X0Y1_EE4BEG[15]
  PIN Tile_X0Y1_EE4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 118.360 225.000 118.960 ;
    END
  END Tile_X0Y1_EE4BEG[1]
  PIN Tile_X0Y1_EE4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 119.720 225.000 120.320 ;
    END
  END Tile_X0Y1_EE4BEG[2]
  PIN Tile_X0Y1_EE4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 121.080 225.000 121.680 ;
    END
  END Tile_X0Y1_EE4BEG[3]
  PIN Tile_X0Y1_EE4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 122.440 225.000 123.040 ;
    END
  END Tile_X0Y1_EE4BEG[4]
  PIN Tile_X0Y1_EE4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 123.800 225.000 124.400 ;
    END
  END Tile_X0Y1_EE4BEG[5]
  PIN Tile_X0Y1_EE4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 125.160 225.000 125.760 ;
    END
  END Tile_X0Y1_EE4BEG[6]
  PIN Tile_X0Y1_EE4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 126.520 225.000 127.120 ;
    END
  END Tile_X0Y1_EE4BEG[7]
  PIN Tile_X0Y1_EE4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 127.880 225.000 128.480 ;
    END
  END Tile_X0Y1_EE4BEG[8]
  PIN Tile_X0Y1_EE4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 129.240 225.000 129.840 ;
    END
  END Tile_X0Y1_EE4BEG[9]
  PIN Tile_X0Y1_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 0.800 117.600 ;
    END
  END Tile_X0Y1_EE4END[0]
  PIN Tile_X0Y1_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 0.800 131.200 ;
    END
  END Tile_X0Y1_EE4END[10]
  PIN Tile_X0Y1_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 0.800 132.560 ;
    END
  END Tile_X0Y1_EE4END[11]
  PIN Tile_X0Y1_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 0.800 133.920 ;
    END
  END Tile_X0Y1_EE4END[12]
  PIN Tile_X0Y1_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 0.800 135.280 ;
    END
  END Tile_X0Y1_EE4END[13]
  PIN Tile_X0Y1_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 0.800 136.640 ;
    END
  END Tile_X0Y1_EE4END[14]
  PIN Tile_X0Y1_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 0.800 138.000 ;
    END
  END Tile_X0Y1_EE4END[15]
  PIN Tile_X0Y1_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 0.800 118.960 ;
    END
  END Tile_X0Y1_EE4END[1]
  PIN Tile_X0Y1_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 0.800 120.320 ;
    END
  END Tile_X0Y1_EE4END[2]
  PIN Tile_X0Y1_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 0.800 121.680 ;
    END
  END Tile_X0Y1_EE4END[3]
  PIN Tile_X0Y1_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 0.800 123.040 ;
    END
  END Tile_X0Y1_EE4END[4]
  PIN Tile_X0Y1_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 0.800 124.400 ;
    END
  END Tile_X0Y1_EE4END[5]
  PIN Tile_X0Y1_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 0.800 125.760 ;
    END
  END Tile_X0Y1_EE4END[6]
  PIN Tile_X0Y1_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 0.800 127.120 ;
    END
  END Tile_X0Y1_EE4END[7]
  PIN Tile_X0Y1_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 0.800 128.480 ;
    END
  END Tile_X0Y1_EE4END[8]
  PIN Tile_X0Y1_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 0.800 129.840 ;
    END
  END Tile_X0Y1_EE4END[9]
  PIN Tile_X0Y1_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 0.800 155.680 ;
    END
  END Tile_X0Y1_FrameData[0]
  PIN Tile_X0Y1_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 0.800 169.280 ;
    END
  END Tile_X0Y1_FrameData[10]
  PIN Tile_X0Y1_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 0.800 170.640 ;
    END
  END Tile_X0Y1_FrameData[11]
  PIN Tile_X0Y1_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 0.800 172.000 ;
    END
  END Tile_X0Y1_FrameData[12]
  PIN Tile_X0Y1_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 0.800 173.360 ;
    END
  END Tile_X0Y1_FrameData[13]
  PIN Tile_X0Y1_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 0.800 174.720 ;
    END
  END Tile_X0Y1_FrameData[14]
  PIN Tile_X0Y1_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 0.800 176.080 ;
    END
  END Tile_X0Y1_FrameData[15]
  PIN Tile_X0Y1_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 0.800 177.440 ;
    END
  END Tile_X0Y1_FrameData[16]
  PIN Tile_X0Y1_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 0.800 178.800 ;
    END
  END Tile_X0Y1_FrameData[17]
  PIN Tile_X0Y1_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 0.800 180.160 ;
    END
  END Tile_X0Y1_FrameData[18]
  PIN Tile_X0Y1_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 0.800 181.520 ;
    END
  END Tile_X0Y1_FrameData[19]
  PIN Tile_X0Y1_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 0.800 157.040 ;
    END
  END Tile_X0Y1_FrameData[1]
  PIN Tile_X0Y1_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 0.800 182.880 ;
    END
  END Tile_X0Y1_FrameData[20]
  PIN Tile_X0Y1_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 0.800 184.240 ;
    END
  END Tile_X0Y1_FrameData[21]
  PIN Tile_X0Y1_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 0.800 185.600 ;
    END
  END Tile_X0Y1_FrameData[22]
  PIN Tile_X0Y1_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 0.800 186.960 ;
    END
  END Tile_X0Y1_FrameData[23]
  PIN Tile_X0Y1_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 0.800 188.320 ;
    END
  END Tile_X0Y1_FrameData[24]
  PIN Tile_X0Y1_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 0.800 189.680 ;
    END
  END Tile_X0Y1_FrameData[25]
  PIN Tile_X0Y1_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 0.800 191.040 ;
    END
  END Tile_X0Y1_FrameData[26]
  PIN Tile_X0Y1_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 0.800 192.400 ;
    END
  END Tile_X0Y1_FrameData[27]
  PIN Tile_X0Y1_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 0.800 193.760 ;
    END
  END Tile_X0Y1_FrameData[28]
  PIN Tile_X0Y1_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 0.800 195.120 ;
    END
  END Tile_X0Y1_FrameData[29]
  PIN Tile_X0Y1_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 0.800 158.400 ;
    END
  END Tile_X0Y1_FrameData[2]
  PIN Tile_X0Y1_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 0.800 196.480 ;
    END
  END Tile_X0Y1_FrameData[30]
  PIN Tile_X0Y1_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 0.800 197.840 ;
    END
  END Tile_X0Y1_FrameData[31]
  PIN Tile_X0Y1_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 0.800 159.760 ;
    END
  END Tile_X0Y1_FrameData[3]
  PIN Tile_X0Y1_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 0.800 161.120 ;
    END
  END Tile_X0Y1_FrameData[4]
  PIN Tile_X0Y1_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 0.800 162.480 ;
    END
  END Tile_X0Y1_FrameData[5]
  PIN Tile_X0Y1_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 0.800 163.840 ;
    END
  END Tile_X0Y1_FrameData[6]
  PIN Tile_X0Y1_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 0.800 165.200 ;
    END
  END Tile_X0Y1_FrameData[7]
  PIN Tile_X0Y1_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 0.800 166.560 ;
    END
  END Tile_X0Y1_FrameData[8]
  PIN Tile_X0Y1_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 0.800 167.920 ;
    END
  END Tile_X0Y1_FrameData[9]
  PIN Tile_X0Y1_FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 155.080 225.000 155.680 ;
    END
  END Tile_X0Y1_FrameData_O[0]
  PIN Tile_X0Y1_FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 168.680 225.000 169.280 ;
    END
  END Tile_X0Y1_FrameData_O[10]
  PIN Tile_X0Y1_FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 170.040 225.000 170.640 ;
    END
  END Tile_X0Y1_FrameData_O[11]
  PIN Tile_X0Y1_FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 171.400 225.000 172.000 ;
    END
  END Tile_X0Y1_FrameData_O[12]
  PIN Tile_X0Y1_FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 172.760 225.000 173.360 ;
    END
  END Tile_X0Y1_FrameData_O[13]
  PIN Tile_X0Y1_FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 174.120 225.000 174.720 ;
    END
  END Tile_X0Y1_FrameData_O[14]
  PIN Tile_X0Y1_FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 175.480 225.000 176.080 ;
    END
  END Tile_X0Y1_FrameData_O[15]
  PIN Tile_X0Y1_FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 176.840 225.000 177.440 ;
    END
  END Tile_X0Y1_FrameData_O[16]
  PIN Tile_X0Y1_FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 178.200 225.000 178.800 ;
    END
  END Tile_X0Y1_FrameData_O[17]
  PIN Tile_X0Y1_FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 179.560 225.000 180.160 ;
    END
  END Tile_X0Y1_FrameData_O[18]
  PIN Tile_X0Y1_FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 180.920 225.000 181.520 ;
    END
  END Tile_X0Y1_FrameData_O[19]
  PIN Tile_X0Y1_FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 156.440 225.000 157.040 ;
    END
  END Tile_X0Y1_FrameData_O[1]
  PIN Tile_X0Y1_FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 182.280 225.000 182.880 ;
    END
  END Tile_X0Y1_FrameData_O[20]
  PIN Tile_X0Y1_FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 183.640 225.000 184.240 ;
    END
  END Tile_X0Y1_FrameData_O[21]
  PIN Tile_X0Y1_FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 185.000 225.000 185.600 ;
    END
  END Tile_X0Y1_FrameData_O[22]
  PIN Tile_X0Y1_FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 186.360 225.000 186.960 ;
    END
  END Tile_X0Y1_FrameData_O[23]
  PIN Tile_X0Y1_FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 187.720 225.000 188.320 ;
    END
  END Tile_X0Y1_FrameData_O[24]
  PIN Tile_X0Y1_FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 189.080 225.000 189.680 ;
    END
  END Tile_X0Y1_FrameData_O[25]
  PIN Tile_X0Y1_FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 190.440 225.000 191.040 ;
    END
  END Tile_X0Y1_FrameData_O[26]
  PIN Tile_X0Y1_FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 191.800 225.000 192.400 ;
    END
  END Tile_X0Y1_FrameData_O[27]
  PIN Tile_X0Y1_FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 193.160 225.000 193.760 ;
    END
  END Tile_X0Y1_FrameData_O[28]
  PIN Tile_X0Y1_FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 194.520 225.000 195.120 ;
    END
  END Tile_X0Y1_FrameData_O[29]
  PIN Tile_X0Y1_FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 157.800 225.000 158.400 ;
    END
  END Tile_X0Y1_FrameData_O[2]
  PIN Tile_X0Y1_FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 195.880 225.000 196.480 ;
    END
  END Tile_X0Y1_FrameData_O[30]
  PIN Tile_X0Y1_FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 197.240 225.000 197.840 ;
    END
  END Tile_X0Y1_FrameData_O[31]
  PIN Tile_X0Y1_FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 159.160 225.000 159.760 ;
    END
  END Tile_X0Y1_FrameData_O[3]
  PIN Tile_X0Y1_FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 160.520 225.000 161.120 ;
    END
  END Tile_X0Y1_FrameData_O[4]
  PIN Tile_X0Y1_FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 161.880 225.000 162.480 ;
    END
  END Tile_X0Y1_FrameData_O[5]
  PIN Tile_X0Y1_FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 163.240 225.000 163.840 ;
    END
  END Tile_X0Y1_FrameData_O[6]
  PIN Tile_X0Y1_FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.200 164.600 225.000 165.200 ;
    END
  END Tile_X0Y1_FrameData_O[7]
  PIN Tile_X0Y1_FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 165.960 225.000 166.560 ;
    END
  END Tile_X0Y1_FrameData_O[8]
  PIN Tile_X0Y1_FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 167.320 225.000 167.920 ;
    END
  END Tile_X0Y1_FrameData_O[9]
  PIN Tile_X0Y1_FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[0]
  PIN Tile_X0Y1_FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[10]
  PIN Tile_X0Y1_FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[11]
  PIN Tile_X0Y1_FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[12]
  PIN Tile_X0Y1_FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[13]
  PIN Tile_X0Y1_FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[14]
  PIN Tile_X0Y1_FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[15]
  PIN Tile_X0Y1_FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[16]
  PIN Tile_X0Y1_FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[17]
  PIN Tile_X0Y1_FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[18]
  PIN Tile_X0Y1_FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[19]
  PIN Tile_X0Y1_FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[1]
  PIN Tile_X0Y1_FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[2]
  PIN Tile_X0Y1_FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[3]
  PIN Tile_X0Y1_FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[4]
  PIN Tile_X0Y1_FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[5]
  PIN Tile_X0Y1_FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[6]
  PIN Tile_X0Y1_FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[7]
  PIN Tile_X0Y1_FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[8]
  PIN Tile_X0Y1_FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 0.800 ;
    END
  END Tile_X0Y1_FrameStrobe[9]
  PIN Tile_X0Y1_N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 0.800 ;
    END
  END Tile_X0Y1_N1END[0]
  PIN Tile_X0Y1_N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 0.800 ;
    END
  END Tile_X0Y1_N1END[1]
  PIN Tile_X0Y1_N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 0.800 ;
    END
  END Tile_X0Y1_N1END[2]
  PIN Tile_X0Y1_N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 0.800 ;
    END
  END Tile_X0Y1_N1END[3]
  PIN Tile_X0Y1_N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 0.800 ;
    END
  END Tile_X0Y1_N2END[0]
  PIN Tile_X0Y1_N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 0.800 ;
    END
  END Tile_X0Y1_N2END[1]
  PIN Tile_X0Y1_N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 0.800 ;
    END
  END Tile_X0Y1_N2END[2]
  PIN Tile_X0Y1_N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 0.800 ;
    END
  END Tile_X0Y1_N2END[3]
  PIN Tile_X0Y1_N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 0.800 ;
    END
  END Tile_X0Y1_N2END[4]
  PIN Tile_X0Y1_N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 0.800 ;
    END
  END Tile_X0Y1_N2END[5]
  PIN Tile_X0Y1_N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 0.800 ;
    END
  END Tile_X0Y1_N2END[6]
  PIN Tile_X0Y1_N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 0.800 ;
    END
  END Tile_X0Y1_N2END[7]
  PIN Tile_X0Y1_N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 0.800 ;
    END
  END Tile_X0Y1_N2MID[0]
  PIN Tile_X0Y1_N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 0.800 ;
    END
  END Tile_X0Y1_N2MID[1]
  PIN Tile_X0Y1_N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 0.800 ;
    END
  END Tile_X0Y1_N2MID[2]
  PIN Tile_X0Y1_N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 0.800 ;
    END
  END Tile_X0Y1_N2MID[3]
  PIN Tile_X0Y1_N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 0.800 ;
    END
  END Tile_X0Y1_N2MID[4]
  PIN Tile_X0Y1_N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 0.800 ;
    END
  END Tile_X0Y1_N2MID[5]
  PIN Tile_X0Y1_N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 0.800 ;
    END
  END Tile_X0Y1_N2MID[6]
  PIN Tile_X0Y1_N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 0.800 ;
    END
  END Tile_X0Y1_N2MID[7]
  PIN Tile_X0Y1_N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 0.800 ;
    END
  END Tile_X0Y1_N4END[0]
  PIN Tile_X0Y1_N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 0.800 ;
    END
  END Tile_X0Y1_N4END[10]
  PIN Tile_X0Y1_N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 0.800 ;
    END
  END Tile_X0Y1_N4END[11]
  PIN Tile_X0Y1_N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 0.800 ;
    END
  END Tile_X0Y1_N4END[12]
  PIN Tile_X0Y1_N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 0.800 ;
    END
  END Tile_X0Y1_N4END[13]
  PIN Tile_X0Y1_N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 0.800 ;
    END
  END Tile_X0Y1_N4END[14]
  PIN Tile_X0Y1_N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 0.800 ;
    END
  END Tile_X0Y1_N4END[15]
  PIN Tile_X0Y1_N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 0.800 ;
    END
  END Tile_X0Y1_N4END[1]
  PIN Tile_X0Y1_N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 0.800 ;
    END
  END Tile_X0Y1_N4END[2]
  PIN Tile_X0Y1_N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 0.800 ;
    END
  END Tile_X0Y1_N4END[3]
  PIN Tile_X0Y1_N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 0.800 ;
    END
  END Tile_X0Y1_N4END[4]
  PIN Tile_X0Y1_N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 0.800 ;
    END
  END Tile_X0Y1_N4END[5]
  PIN Tile_X0Y1_N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 0.800 ;
    END
  END Tile_X0Y1_N4END[6]
  PIN Tile_X0Y1_N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 0.800 ;
    END
  END Tile_X0Y1_N4END[7]
  PIN Tile_X0Y1_N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 0.800 ;
    END
  END Tile_X0Y1_N4END[8]
  PIN Tile_X0Y1_N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 0.800 ;
    END
  END Tile_X0Y1_N4END[9]
  PIN Tile_X0Y1_NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 0.800 ;
    END
  END Tile_X0Y1_NN4END[0]
  PIN Tile_X0Y1_NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 0.800 ;
    END
  END Tile_X0Y1_NN4END[10]
  PIN Tile_X0Y1_NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 0.800 ;
    END
  END Tile_X0Y1_NN4END[11]
  PIN Tile_X0Y1_NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 0.800 ;
    END
  END Tile_X0Y1_NN4END[12]
  PIN Tile_X0Y1_NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 0.800 ;
    END
  END Tile_X0Y1_NN4END[13]
  PIN Tile_X0Y1_NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 0.800 ;
    END
  END Tile_X0Y1_NN4END[14]
  PIN Tile_X0Y1_NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 0.800 ;
    END
  END Tile_X0Y1_NN4END[15]
  PIN Tile_X0Y1_NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 0.800 ;
    END
  END Tile_X0Y1_NN4END[1]
  PIN Tile_X0Y1_NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 0.800 ;
    END
  END Tile_X0Y1_NN4END[2]
  PIN Tile_X0Y1_NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 0.800 ;
    END
  END Tile_X0Y1_NN4END[3]
  PIN Tile_X0Y1_NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 0.800 ;
    END
  END Tile_X0Y1_NN4END[4]
  PIN Tile_X0Y1_NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 0.800 ;
    END
  END Tile_X0Y1_NN4END[5]
  PIN Tile_X0Y1_NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 0.800 ;
    END
  END Tile_X0Y1_NN4END[6]
  PIN Tile_X0Y1_NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 0.800 ;
    END
  END Tile_X0Y1_NN4END[7]
  PIN Tile_X0Y1_NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 0.800 ;
    END
  END Tile_X0Y1_NN4END[8]
  PIN Tile_X0Y1_NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 0.800 ;
    END
  END Tile_X0Y1_NN4END[9]
  PIN Tile_X0Y1_S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 0.800 ;
    END
  END Tile_X0Y1_S1BEG[0]
  PIN Tile_X0Y1_S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 0.800 ;
    END
  END Tile_X0Y1_S1BEG[1]
  PIN Tile_X0Y1_S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 0.800 ;
    END
  END Tile_X0Y1_S1BEG[2]
  PIN Tile_X0Y1_S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 0.800 ;
    END
  END Tile_X0Y1_S1BEG[3]
  PIN Tile_X0Y1_S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 0.800 ;
    END
  END Tile_X0Y1_S2BEG[0]
  PIN Tile_X0Y1_S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 0.800 ;
    END
  END Tile_X0Y1_S2BEG[1]
  PIN Tile_X0Y1_S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 0.800 ;
    END
  END Tile_X0Y1_S2BEG[2]
  PIN Tile_X0Y1_S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 0.800 ;
    END
  END Tile_X0Y1_S2BEG[3]
  PIN Tile_X0Y1_S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 0.800 ;
    END
  END Tile_X0Y1_S2BEG[4]
  PIN Tile_X0Y1_S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 0.800 ;
    END
  END Tile_X0Y1_S2BEG[5]
  PIN Tile_X0Y1_S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 0.800 ;
    END
  END Tile_X0Y1_S2BEG[6]
  PIN Tile_X0Y1_S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 0.800 ;
    END
  END Tile_X0Y1_S2BEG[7]
  PIN Tile_X0Y1_S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 0.800 ;
    END
  END Tile_X0Y1_S2BEGb[0]
  PIN Tile_X0Y1_S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 0.800 ;
    END
  END Tile_X0Y1_S2BEGb[1]
  PIN Tile_X0Y1_S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 0.800 ;
    END
  END Tile_X0Y1_S2BEGb[2]
  PIN Tile_X0Y1_S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 0.800 ;
    END
  END Tile_X0Y1_S2BEGb[3]
  PIN Tile_X0Y1_S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 0.800 ;
    END
  END Tile_X0Y1_S2BEGb[4]
  PIN Tile_X0Y1_S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 0.800 ;
    END
  END Tile_X0Y1_S2BEGb[5]
  PIN Tile_X0Y1_S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 0.800 ;
    END
  END Tile_X0Y1_S2BEGb[6]
  PIN Tile_X0Y1_S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 0.800 ;
    END
  END Tile_X0Y1_S2BEGb[7]
  PIN Tile_X0Y1_S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 0.800 ;
    END
  END Tile_X0Y1_S4BEG[0]
  PIN Tile_X0Y1_S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 0.800 ;
    END
  END Tile_X0Y1_S4BEG[10]
  PIN Tile_X0Y1_S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 0.800 ;
    END
  END Tile_X0Y1_S4BEG[11]
  PIN Tile_X0Y1_S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 0.800 ;
    END
  END Tile_X0Y1_S4BEG[12]
  PIN Tile_X0Y1_S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 0.800 ;
    END
  END Tile_X0Y1_S4BEG[13]
  PIN Tile_X0Y1_S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 0.800 ;
    END
  END Tile_X0Y1_S4BEG[14]
  PIN Tile_X0Y1_S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 0.800 ;
    END
  END Tile_X0Y1_S4BEG[15]
  PIN Tile_X0Y1_S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 0.800 ;
    END
  END Tile_X0Y1_S4BEG[1]
  PIN Tile_X0Y1_S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 0.800 ;
    END
  END Tile_X0Y1_S4BEG[2]
  PIN Tile_X0Y1_S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 0.800 ;
    END
  END Tile_X0Y1_S4BEG[3]
  PIN Tile_X0Y1_S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 0.800 ;
    END
  END Tile_X0Y1_S4BEG[4]
  PIN Tile_X0Y1_S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 0.800 ;
    END
  END Tile_X0Y1_S4BEG[5]
  PIN Tile_X0Y1_S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 0.800 ;
    END
  END Tile_X0Y1_S4BEG[6]
  PIN Tile_X0Y1_S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 0.800 ;
    END
  END Tile_X0Y1_S4BEG[7]
  PIN Tile_X0Y1_S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 0.800 ;
    END
  END Tile_X0Y1_S4BEG[8]
  PIN Tile_X0Y1_S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 0.800 ;
    END
  END Tile_X0Y1_S4BEG[9]
  PIN Tile_X0Y1_SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[0]
  PIN Tile_X0Y1_SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[10]
  PIN Tile_X0Y1_SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[11]
  PIN Tile_X0Y1_SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[12]
  PIN Tile_X0Y1_SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[13]
  PIN Tile_X0Y1_SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[14]
  PIN Tile_X0Y1_SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[15]
  PIN Tile_X0Y1_SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[1]
  PIN Tile_X0Y1_SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[2]
  PIN Tile_X0Y1_SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[3]
  PIN Tile_X0Y1_SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[4]
  PIN Tile_X0Y1_SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[5]
  PIN Tile_X0Y1_SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[6]
  PIN Tile_X0Y1_SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[7]
  PIN Tile_X0Y1_SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[8]
  PIN Tile_X0Y1_SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 0.800 ;
    END
  END Tile_X0Y1_SS4BEG[9]
  PIN Tile_X0Y1_UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 0.800 ;
    END
  END Tile_X0Y1_UserCLK
  PIN Tile_X0Y1_W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 0.800 25.120 ;
    END
  END Tile_X0Y1_W1BEG[0]
  PIN Tile_X0Y1_W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 0.800 26.480 ;
    END
  END Tile_X0Y1_W1BEG[1]
  PIN Tile_X0Y1_W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 0.800 27.840 ;
    END
  END Tile_X0Y1_W1BEG[2]
  PIN Tile_X0Y1_W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 0.800 29.200 ;
    END
  END Tile_X0Y1_W1BEG[3]
  PIN Tile_X0Y1_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 24.520 225.000 25.120 ;
    END
  END Tile_X0Y1_W1END[0]
  PIN Tile_X0Y1_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 25.880 225.000 26.480 ;
    END
  END Tile_X0Y1_W1END[1]
  PIN Tile_X0Y1_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 27.240 225.000 27.840 ;
    END
  END Tile_X0Y1_W1END[2]
  PIN Tile_X0Y1_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 28.600 225.000 29.200 ;
    END
  END Tile_X0Y1_W1END[3]
  PIN Tile_X0Y1_W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 0.800 30.560 ;
    END
  END Tile_X0Y1_W2BEG[0]
  PIN Tile_X0Y1_W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 0.800 31.920 ;
    END
  END Tile_X0Y1_W2BEG[1]
  PIN Tile_X0Y1_W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 0.800 33.280 ;
    END
  END Tile_X0Y1_W2BEG[2]
  PIN Tile_X0Y1_W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 0.800 34.640 ;
    END
  END Tile_X0Y1_W2BEG[3]
  PIN Tile_X0Y1_W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 0.800 36.000 ;
    END
  END Tile_X0Y1_W2BEG[4]
  PIN Tile_X0Y1_W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 0.800 37.360 ;
    END
  END Tile_X0Y1_W2BEG[5]
  PIN Tile_X0Y1_W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 0.800 38.720 ;
    END
  END Tile_X0Y1_W2BEG[6]
  PIN Tile_X0Y1_W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 0.800 40.080 ;
    END
  END Tile_X0Y1_W2BEG[7]
  PIN Tile_X0Y1_W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 0.800 41.440 ;
    END
  END Tile_X0Y1_W2BEGb[0]
  PIN Tile_X0Y1_W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 0.800 42.800 ;
    END
  END Tile_X0Y1_W2BEGb[1]
  PIN Tile_X0Y1_W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 0.800 44.160 ;
    END
  END Tile_X0Y1_W2BEGb[2]
  PIN Tile_X0Y1_W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 0.800 45.520 ;
    END
  END Tile_X0Y1_W2BEGb[3]
  PIN Tile_X0Y1_W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 0.800 46.880 ;
    END
  END Tile_X0Y1_W2BEGb[4]
  PIN Tile_X0Y1_W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 0.800 48.240 ;
    END
  END Tile_X0Y1_W2BEGb[5]
  PIN Tile_X0Y1_W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 0.800 49.600 ;
    END
  END Tile_X0Y1_W2BEGb[6]
  PIN Tile_X0Y1_W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 0.800 50.960 ;
    END
  END Tile_X0Y1_W2BEGb[7]
  PIN Tile_X0Y1_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 40.840 225.000 41.440 ;
    END
  END Tile_X0Y1_W2END[0]
  PIN Tile_X0Y1_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 42.200 225.000 42.800 ;
    END
  END Tile_X0Y1_W2END[1]
  PIN Tile_X0Y1_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 43.560 225.000 44.160 ;
    END
  END Tile_X0Y1_W2END[2]
  PIN Tile_X0Y1_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 44.920 225.000 45.520 ;
    END
  END Tile_X0Y1_W2END[3]
  PIN Tile_X0Y1_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 46.280 225.000 46.880 ;
    END
  END Tile_X0Y1_W2END[4]
  PIN Tile_X0Y1_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 47.640 225.000 48.240 ;
    END
  END Tile_X0Y1_W2END[5]
  PIN Tile_X0Y1_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 49.000 225.000 49.600 ;
    END
  END Tile_X0Y1_W2END[6]
  PIN Tile_X0Y1_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 50.360 225.000 50.960 ;
    END
  END Tile_X0Y1_W2END[7]
  PIN Tile_X0Y1_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 29.960 225.000 30.560 ;
    END
  END Tile_X0Y1_W2MID[0]
  PIN Tile_X0Y1_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 31.320 225.000 31.920 ;
    END
  END Tile_X0Y1_W2MID[1]
  PIN Tile_X0Y1_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 32.680 225.000 33.280 ;
    END
  END Tile_X0Y1_W2MID[2]
  PIN Tile_X0Y1_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 34.040 225.000 34.640 ;
    END
  END Tile_X0Y1_W2MID[3]
  PIN Tile_X0Y1_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 35.400 225.000 36.000 ;
    END
  END Tile_X0Y1_W2MID[4]
  PIN Tile_X0Y1_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 36.760 225.000 37.360 ;
    END
  END Tile_X0Y1_W2MID[5]
  PIN Tile_X0Y1_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 38.120 225.000 38.720 ;
    END
  END Tile_X0Y1_W2MID[6]
  PIN Tile_X0Y1_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 39.480 225.000 40.080 ;
    END
  END Tile_X0Y1_W2MID[7]
  PIN Tile_X0Y1_W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 0.800 74.080 ;
    END
  END Tile_X0Y1_W6BEG[0]
  PIN Tile_X0Y1_W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 0.800 87.680 ;
    END
  END Tile_X0Y1_W6BEG[10]
  PIN Tile_X0Y1_W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 0.800 89.040 ;
    END
  END Tile_X0Y1_W6BEG[11]
  PIN Tile_X0Y1_W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 0.800 75.440 ;
    END
  END Tile_X0Y1_W6BEG[1]
  PIN Tile_X0Y1_W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 0.800 76.800 ;
    END
  END Tile_X0Y1_W6BEG[2]
  PIN Tile_X0Y1_W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 0.800 78.160 ;
    END
  END Tile_X0Y1_W6BEG[3]
  PIN Tile_X0Y1_W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 0.800 79.520 ;
    END
  END Tile_X0Y1_W6BEG[4]
  PIN Tile_X0Y1_W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 0.800 80.880 ;
    END
  END Tile_X0Y1_W6BEG[5]
  PIN Tile_X0Y1_W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 0.800 82.240 ;
    END
  END Tile_X0Y1_W6BEG[6]
  PIN Tile_X0Y1_W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 0.800 83.600 ;
    END
  END Tile_X0Y1_W6BEG[7]
  PIN Tile_X0Y1_W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 0.800 84.960 ;
    END
  END Tile_X0Y1_W6BEG[8]
  PIN Tile_X0Y1_W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 0.800 86.320 ;
    END
  END Tile_X0Y1_W6BEG[9]
  PIN Tile_X0Y1_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 73.480 225.000 74.080 ;
    END
  END Tile_X0Y1_W6END[0]
  PIN Tile_X0Y1_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 87.080 225.000 87.680 ;
    END
  END Tile_X0Y1_W6END[10]
  PIN Tile_X0Y1_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 88.440 225.000 89.040 ;
    END
  END Tile_X0Y1_W6END[11]
  PIN Tile_X0Y1_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 74.840 225.000 75.440 ;
    END
  END Tile_X0Y1_W6END[1]
  PIN Tile_X0Y1_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 76.200 225.000 76.800 ;
    END
  END Tile_X0Y1_W6END[2]
  PIN Tile_X0Y1_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 77.560 225.000 78.160 ;
    END
  END Tile_X0Y1_W6END[3]
  PIN Tile_X0Y1_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 78.920 225.000 79.520 ;
    END
  END Tile_X0Y1_W6END[4]
  PIN Tile_X0Y1_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 80.280 225.000 80.880 ;
    END
  END Tile_X0Y1_W6END[5]
  PIN Tile_X0Y1_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 81.640 225.000 82.240 ;
    END
  END Tile_X0Y1_W6END[6]
  PIN Tile_X0Y1_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 83.000 225.000 83.600 ;
    END
  END Tile_X0Y1_W6END[7]
  PIN Tile_X0Y1_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 84.360 225.000 84.960 ;
    END
  END Tile_X0Y1_W6END[8]
  PIN Tile_X0Y1_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 85.720 225.000 86.320 ;
    END
  END Tile_X0Y1_W6END[9]
  PIN Tile_X0Y1_WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 0.800 52.320 ;
    END
  END Tile_X0Y1_WW4BEG[0]
  PIN Tile_X0Y1_WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 0.800 65.920 ;
    END
  END Tile_X0Y1_WW4BEG[10]
  PIN Tile_X0Y1_WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 0.800 67.280 ;
    END
  END Tile_X0Y1_WW4BEG[11]
  PIN Tile_X0Y1_WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 0.800 68.640 ;
    END
  END Tile_X0Y1_WW4BEG[12]
  PIN Tile_X0Y1_WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 0.800 70.000 ;
    END
  END Tile_X0Y1_WW4BEG[13]
  PIN Tile_X0Y1_WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 0.800 71.360 ;
    END
  END Tile_X0Y1_WW4BEG[14]
  PIN Tile_X0Y1_WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 0.800 72.720 ;
    END
  END Tile_X0Y1_WW4BEG[15]
  PIN Tile_X0Y1_WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 0.800 53.680 ;
    END
  END Tile_X0Y1_WW4BEG[1]
  PIN Tile_X0Y1_WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 0.800 55.040 ;
    END
  END Tile_X0Y1_WW4BEG[2]
  PIN Tile_X0Y1_WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 0.800 56.400 ;
    END
  END Tile_X0Y1_WW4BEG[3]
  PIN Tile_X0Y1_WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 0.800 57.760 ;
    END
  END Tile_X0Y1_WW4BEG[4]
  PIN Tile_X0Y1_WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 0.800 59.120 ;
    END
  END Tile_X0Y1_WW4BEG[5]
  PIN Tile_X0Y1_WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 0.800 60.480 ;
    END
  END Tile_X0Y1_WW4BEG[6]
  PIN Tile_X0Y1_WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 0.800 61.840 ;
    END
  END Tile_X0Y1_WW4BEG[7]
  PIN Tile_X0Y1_WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 0.800 63.200 ;
    END
  END Tile_X0Y1_WW4BEG[8]
  PIN Tile_X0Y1_WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 0.800 64.560 ;
    END
  END Tile_X0Y1_WW4BEG[9]
  PIN Tile_X0Y1_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 51.720 225.000 52.320 ;
    END
  END Tile_X0Y1_WW4END[0]
  PIN Tile_X0Y1_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 65.320 225.000 65.920 ;
    END
  END Tile_X0Y1_WW4END[10]
  PIN Tile_X0Y1_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 66.680 225.000 67.280 ;
    END
  END Tile_X0Y1_WW4END[11]
  PIN Tile_X0Y1_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 68.040 225.000 68.640 ;
    END
  END Tile_X0Y1_WW4END[12]
  PIN Tile_X0Y1_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 69.400 225.000 70.000 ;
    END
  END Tile_X0Y1_WW4END[13]
  PIN Tile_X0Y1_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 70.760 225.000 71.360 ;
    END
  END Tile_X0Y1_WW4END[14]
  PIN Tile_X0Y1_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 72.120 225.000 72.720 ;
    END
  END Tile_X0Y1_WW4END[15]
  PIN Tile_X0Y1_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 53.080 225.000 53.680 ;
    END
  END Tile_X0Y1_WW4END[1]
  PIN Tile_X0Y1_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 54.440 225.000 55.040 ;
    END
  END Tile_X0Y1_WW4END[2]
  PIN Tile_X0Y1_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 224.200 55.800 225.000 56.400 ;
    END
  END Tile_X0Y1_WW4END[3]
  PIN Tile_X0Y1_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 57.160 225.000 57.760 ;
    END
  END Tile_X0Y1_WW4END[4]
  PIN Tile_X0Y1_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 58.520 225.000 59.120 ;
    END
  END Tile_X0Y1_WW4END[5]
  PIN Tile_X0Y1_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 59.880 225.000 60.480 ;
    END
  END Tile_X0Y1_WW4END[6]
  PIN Tile_X0Y1_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 61.240 225.000 61.840 ;
    END
  END Tile_X0Y1_WW4END[7]
  PIN Tile_X0Y1_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 62.600 225.000 63.200 ;
    END
  END Tile_X0Y1_WW4END[8]
  PIN Tile_X0Y1_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.200 63.960 225.000 64.560 ;
    END
  END Tile_X0Y1_WW4END[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 5.200 99.440 443.600 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 443.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 5.200 176.240 443.600 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 219.420 443.445 ;
      LAYER met1 ;
        RECT 0.070 1.060 223.950 446.380 ;
      LAYER met2 ;
        RECT 0.100 448.920 26.490 449.890 ;
        RECT 27.330 448.920 27.870 449.890 ;
        RECT 28.710 448.920 29.250 449.890 ;
        RECT 30.090 448.920 30.630 449.890 ;
        RECT 31.470 448.920 32.010 449.890 ;
        RECT 32.850 448.920 33.390 449.890 ;
        RECT 34.230 448.920 34.770 449.890 ;
        RECT 35.610 448.920 36.150 449.890 ;
        RECT 36.990 448.920 37.530 449.890 ;
        RECT 38.370 448.920 38.910 449.890 ;
        RECT 39.750 448.920 40.290 449.890 ;
        RECT 41.130 448.920 41.670 449.890 ;
        RECT 42.510 448.920 43.050 449.890 ;
        RECT 43.890 448.920 44.430 449.890 ;
        RECT 45.270 448.920 45.810 449.890 ;
        RECT 46.650 448.920 47.190 449.890 ;
        RECT 48.030 448.920 48.570 449.890 ;
        RECT 49.410 448.920 49.950 449.890 ;
        RECT 50.790 448.920 51.330 449.890 ;
        RECT 52.170 448.920 52.710 449.890 ;
        RECT 53.550 448.920 54.090 449.890 ;
        RECT 54.930 448.920 55.470 449.890 ;
        RECT 56.310 448.920 56.850 449.890 ;
        RECT 57.690 448.920 58.230 449.890 ;
        RECT 59.070 448.920 59.610 449.890 ;
        RECT 60.450 448.920 60.990 449.890 ;
        RECT 61.830 448.920 62.370 449.890 ;
        RECT 63.210 448.920 63.750 449.890 ;
        RECT 64.590 448.920 65.130 449.890 ;
        RECT 65.970 448.920 66.510 449.890 ;
        RECT 67.350 448.920 67.890 449.890 ;
        RECT 68.730 448.920 69.270 449.890 ;
        RECT 70.110 448.920 70.650 449.890 ;
        RECT 71.490 448.920 72.030 449.890 ;
        RECT 72.870 448.920 73.410 449.890 ;
        RECT 74.250 448.920 74.790 449.890 ;
        RECT 75.630 448.920 76.170 449.890 ;
        RECT 77.010 448.920 77.550 449.890 ;
        RECT 78.390 448.920 78.930 449.890 ;
        RECT 79.770 448.920 80.310 449.890 ;
        RECT 81.150 448.920 81.690 449.890 ;
        RECT 82.530 448.920 83.070 449.890 ;
        RECT 83.910 448.920 84.450 449.890 ;
        RECT 85.290 448.920 85.830 449.890 ;
        RECT 86.670 448.920 87.210 449.890 ;
        RECT 88.050 448.920 88.590 449.890 ;
        RECT 89.430 448.920 89.970 449.890 ;
        RECT 90.810 448.920 91.350 449.890 ;
        RECT 92.190 448.920 92.730 449.890 ;
        RECT 93.570 448.920 94.110 449.890 ;
        RECT 94.950 448.920 95.490 449.890 ;
        RECT 96.330 448.920 96.870 449.890 ;
        RECT 97.710 448.920 98.250 449.890 ;
        RECT 99.090 448.920 99.630 449.890 ;
        RECT 100.470 448.920 101.010 449.890 ;
        RECT 101.850 448.920 102.390 449.890 ;
        RECT 103.230 448.920 103.770 449.890 ;
        RECT 104.610 448.920 105.150 449.890 ;
        RECT 105.990 448.920 106.530 449.890 ;
        RECT 107.370 448.920 107.910 449.890 ;
        RECT 108.750 448.920 109.290 449.890 ;
        RECT 110.130 448.920 110.670 449.890 ;
        RECT 111.510 448.920 112.050 449.890 ;
        RECT 112.890 448.920 113.430 449.890 ;
        RECT 114.270 448.920 114.810 449.890 ;
        RECT 115.650 448.920 116.190 449.890 ;
        RECT 117.030 448.920 117.570 449.890 ;
        RECT 118.410 448.920 118.950 449.890 ;
        RECT 119.790 448.920 120.330 449.890 ;
        RECT 121.170 448.920 121.710 449.890 ;
        RECT 122.550 448.920 123.090 449.890 ;
        RECT 123.930 448.920 124.470 449.890 ;
        RECT 125.310 448.920 125.850 449.890 ;
        RECT 126.690 448.920 127.230 449.890 ;
        RECT 128.070 448.920 128.610 449.890 ;
        RECT 129.450 448.920 129.990 449.890 ;
        RECT 130.830 448.920 131.370 449.890 ;
        RECT 132.210 448.920 132.750 449.890 ;
        RECT 133.590 448.920 134.130 449.890 ;
        RECT 134.970 448.920 135.510 449.890 ;
        RECT 136.350 448.920 136.890 449.890 ;
        RECT 137.730 448.920 138.270 449.890 ;
        RECT 139.110 448.920 139.650 449.890 ;
        RECT 140.490 448.920 141.030 449.890 ;
        RECT 141.870 448.920 142.410 449.890 ;
        RECT 143.250 448.920 143.790 449.890 ;
        RECT 144.630 448.920 145.170 449.890 ;
        RECT 146.010 448.920 146.550 449.890 ;
        RECT 147.390 448.920 147.930 449.890 ;
        RECT 148.770 448.920 149.310 449.890 ;
        RECT 150.150 448.920 150.690 449.890 ;
        RECT 151.530 448.920 152.070 449.890 ;
        RECT 152.910 448.920 153.450 449.890 ;
        RECT 154.290 448.920 154.830 449.890 ;
        RECT 155.670 448.920 156.210 449.890 ;
        RECT 157.050 448.920 157.590 449.890 ;
        RECT 158.430 448.920 158.970 449.890 ;
        RECT 159.810 448.920 160.350 449.890 ;
        RECT 161.190 448.920 161.730 449.890 ;
        RECT 162.570 448.920 163.110 449.890 ;
        RECT 163.950 448.920 164.490 449.890 ;
        RECT 165.330 448.920 165.870 449.890 ;
        RECT 166.710 448.920 167.250 449.890 ;
        RECT 168.090 448.920 168.630 449.890 ;
        RECT 169.470 448.920 170.010 449.890 ;
        RECT 170.850 448.920 171.390 449.890 ;
        RECT 172.230 448.920 172.770 449.890 ;
        RECT 173.610 448.920 174.150 449.890 ;
        RECT 174.990 448.920 175.530 449.890 ;
        RECT 176.370 448.920 176.910 449.890 ;
        RECT 177.750 448.920 178.290 449.890 ;
        RECT 179.130 448.920 179.670 449.890 ;
        RECT 180.510 448.920 181.050 449.890 ;
        RECT 181.890 448.920 182.430 449.890 ;
        RECT 183.270 448.920 183.810 449.890 ;
        RECT 184.650 448.920 185.190 449.890 ;
        RECT 186.030 448.920 186.570 449.890 ;
        RECT 187.410 448.920 187.950 449.890 ;
        RECT 188.790 448.920 189.330 449.890 ;
        RECT 190.170 448.920 190.710 449.890 ;
        RECT 191.550 448.920 192.090 449.890 ;
        RECT 192.930 448.920 193.470 449.890 ;
        RECT 194.310 448.920 194.850 449.890 ;
        RECT 195.690 448.920 196.230 449.890 ;
        RECT 197.070 448.920 197.610 449.890 ;
        RECT 198.450 448.920 224.390 449.890 ;
        RECT 0.100 1.080 224.390 448.920 ;
        RECT 0.100 0.270 26.490 1.080 ;
        RECT 27.330 0.270 27.870 1.080 ;
        RECT 28.710 0.270 29.250 1.080 ;
        RECT 30.090 0.270 30.630 1.080 ;
        RECT 31.470 0.270 32.010 1.080 ;
        RECT 32.850 0.270 33.390 1.080 ;
        RECT 34.230 0.270 34.770 1.080 ;
        RECT 35.610 0.270 36.150 1.080 ;
        RECT 36.990 0.270 37.530 1.080 ;
        RECT 38.370 0.270 38.910 1.080 ;
        RECT 39.750 0.270 40.290 1.080 ;
        RECT 41.130 0.270 41.670 1.080 ;
        RECT 42.510 0.270 43.050 1.080 ;
        RECT 43.890 0.270 44.430 1.080 ;
        RECT 45.270 0.270 45.810 1.080 ;
        RECT 46.650 0.270 47.190 1.080 ;
        RECT 48.030 0.270 48.570 1.080 ;
        RECT 49.410 0.270 49.950 1.080 ;
        RECT 50.790 0.270 51.330 1.080 ;
        RECT 52.170 0.270 52.710 1.080 ;
        RECT 53.550 0.270 54.090 1.080 ;
        RECT 54.930 0.270 55.470 1.080 ;
        RECT 56.310 0.270 56.850 1.080 ;
        RECT 57.690 0.270 58.230 1.080 ;
        RECT 59.070 0.270 59.610 1.080 ;
        RECT 60.450 0.270 60.990 1.080 ;
        RECT 61.830 0.270 62.370 1.080 ;
        RECT 63.210 0.270 63.750 1.080 ;
        RECT 64.590 0.270 65.130 1.080 ;
        RECT 65.970 0.270 66.510 1.080 ;
        RECT 67.350 0.270 67.890 1.080 ;
        RECT 68.730 0.270 69.270 1.080 ;
        RECT 70.110 0.270 70.650 1.080 ;
        RECT 71.490 0.270 72.030 1.080 ;
        RECT 72.870 0.270 73.410 1.080 ;
        RECT 74.250 0.270 74.790 1.080 ;
        RECT 75.630 0.270 76.170 1.080 ;
        RECT 77.010 0.270 77.550 1.080 ;
        RECT 78.390 0.270 78.930 1.080 ;
        RECT 79.770 0.270 80.310 1.080 ;
        RECT 81.150 0.270 81.690 1.080 ;
        RECT 82.530 0.270 83.070 1.080 ;
        RECT 83.910 0.270 84.450 1.080 ;
        RECT 85.290 0.270 85.830 1.080 ;
        RECT 86.670 0.270 87.210 1.080 ;
        RECT 88.050 0.270 88.590 1.080 ;
        RECT 89.430 0.270 89.970 1.080 ;
        RECT 90.810 0.270 91.350 1.080 ;
        RECT 92.190 0.270 92.730 1.080 ;
        RECT 93.570 0.270 94.110 1.080 ;
        RECT 94.950 0.270 95.490 1.080 ;
        RECT 96.330 0.270 96.870 1.080 ;
        RECT 97.710 0.270 98.250 1.080 ;
        RECT 99.090 0.270 99.630 1.080 ;
        RECT 100.470 0.270 101.010 1.080 ;
        RECT 101.850 0.270 102.390 1.080 ;
        RECT 103.230 0.270 103.770 1.080 ;
        RECT 104.610 0.270 105.150 1.080 ;
        RECT 105.990 0.270 106.530 1.080 ;
        RECT 107.370 0.270 107.910 1.080 ;
        RECT 108.750 0.270 109.290 1.080 ;
        RECT 110.130 0.270 110.670 1.080 ;
        RECT 111.510 0.270 112.050 1.080 ;
        RECT 112.890 0.270 113.430 1.080 ;
        RECT 114.270 0.270 114.810 1.080 ;
        RECT 115.650 0.270 116.190 1.080 ;
        RECT 117.030 0.270 117.570 1.080 ;
        RECT 118.410 0.270 118.950 1.080 ;
        RECT 119.790 0.270 120.330 1.080 ;
        RECT 121.170 0.270 121.710 1.080 ;
        RECT 122.550 0.270 123.090 1.080 ;
        RECT 123.930 0.270 124.470 1.080 ;
        RECT 125.310 0.270 125.850 1.080 ;
        RECT 126.690 0.270 127.230 1.080 ;
        RECT 128.070 0.270 128.610 1.080 ;
        RECT 129.450 0.270 129.990 1.080 ;
        RECT 130.830 0.270 131.370 1.080 ;
        RECT 132.210 0.270 132.750 1.080 ;
        RECT 133.590 0.270 134.130 1.080 ;
        RECT 134.970 0.270 135.510 1.080 ;
        RECT 136.350 0.270 136.890 1.080 ;
        RECT 137.730 0.270 138.270 1.080 ;
        RECT 139.110 0.270 139.650 1.080 ;
        RECT 140.490 0.270 141.030 1.080 ;
        RECT 141.870 0.270 142.410 1.080 ;
        RECT 143.250 0.270 143.790 1.080 ;
        RECT 144.630 0.270 145.170 1.080 ;
        RECT 146.010 0.270 146.550 1.080 ;
        RECT 147.390 0.270 147.930 1.080 ;
        RECT 148.770 0.270 149.310 1.080 ;
        RECT 150.150 0.270 150.690 1.080 ;
        RECT 151.530 0.270 152.070 1.080 ;
        RECT 152.910 0.270 153.450 1.080 ;
        RECT 154.290 0.270 154.830 1.080 ;
        RECT 155.670 0.270 156.210 1.080 ;
        RECT 157.050 0.270 157.590 1.080 ;
        RECT 158.430 0.270 158.970 1.080 ;
        RECT 159.810 0.270 160.350 1.080 ;
        RECT 161.190 0.270 161.730 1.080 ;
        RECT 162.570 0.270 163.110 1.080 ;
        RECT 163.950 0.270 164.490 1.080 ;
        RECT 165.330 0.270 165.870 1.080 ;
        RECT 166.710 0.270 167.250 1.080 ;
        RECT 168.090 0.270 168.630 1.080 ;
        RECT 169.470 0.270 170.010 1.080 ;
        RECT 170.850 0.270 171.390 1.080 ;
        RECT 172.230 0.270 172.770 1.080 ;
        RECT 173.610 0.270 174.150 1.080 ;
        RECT 174.990 0.270 175.530 1.080 ;
        RECT 176.370 0.270 176.910 1.080 ;
        RECT 177.750 0.270 178.290 1.080 ;
        RECT 179.130 0.270 179.670 1.080 ;
        RECT 180.510 0.270 181.050 1.080 ;
        RECT 181.890 0.270 182.430 1.080 ;
        RECT 183.270 0.270 183.810 1.080 ;
        RECT 184.650 0.270 185.190 1.080 ;
        RECT 186.030 0.270 186.570 1.080 ;
        RECT 187.410 0.270 187.950 1.080 ;
        RECT 188.790 0.270 189.330 1.080 ;
        RECT 190.170 0.270 190.710 1.080 ;
        RECT 191.550 0.270 192.090 1.080 ;
        RECT 192.930 0.270 193.470 1.080 ;
        RECT 194.310 0.270 194.850 1.080 ;
        RECT 195.690 0.270 196.230 1.080 ;
        RECT 197.070 0.270 197.610 1.080 ;
        RECT 198.450 0.270 224.390 1.080 ;
      LAYER met3 ;
        RECT 0.800 428.080 224.415 444.545 ;
        RECT 1.200 253.960 223.800 428.080 ;
        RECT 0.800 198.240 224.415 253.960 ;
        RECT 1.200 24.120 223.800 198.240 ;
        RECT 0.800 4.255 224.415 24.120 ;
      LAYER met4 ;
        RECT 2.135 444.000 208.545 444.545 ;
        RECT 2.135 4.800 20.640 444.000 ;
        RECT 23.040 4.800 97.440 444.000 ;
        RECT 99.840 4.800 174.240 444.000 ;
        RECT 176.640 4.800 208.545 444.000 ;
        RECT 2.135 4.255 208.545 4.800 ;
  END
END DSP
END LIBRARY

