magic
tech sky130A
magscale 1 2
timestamp 1733241215
<< viali >>
rect 2513 6409 2547 6443
rect 4169 6409 4203 6443
rect 4629 6409 4663 6443
rect 6377 6409 6411 6443
rect 7205 6409 7239 6443
rect 7389 6409 7423 6443
rect 8401 6409 8435 6443
rect 8585 6409 8619 6443
rect 9413 6409 9447 6443
rect 9781 6409 9815 6443
rect 10609 6409 10643 6443
rect 10977 6409 11011 6443
rect 11989 6409 12023 6443
rect 12173 6409 12207 6443
rect 12449 6409 12483 6443
rect 13185 6409 13219 6443
rect 13369 6409 13403 6443
rect 14289 6409 14323 6443
rect 14933 6409 14967 6443
rect 15393 6409 15427 6443
rect 15761 6409 15795 6443
rect 16865 6409 16899 6443
rect 17233 6409 17267 6443
rect 17785 6409 17819 6443
rect 18153 6409 18187 6443
rect 19441 6409 19475 6443
rect 19809 6409 19843 6443
rect 20361 6409 20395 6443
rect 20821 6409 20855 6443
rect 21557 6409 21591 6443
rect 21833 6409 21867 6443
rect 22937 6409 22971 6443
rect 23489 6409 23523 6443
rect 23949 6409 23983 6443
rect 1409 6341 1443 6375
rect 5733 6341 5767 6375
rect 6101 6341 6135 6375
rect 6929 6341 6963 6375
rect 8125 6341 8159 6375
rect 9321 6341 9355 6375
rect 10517 6341 10551 6375
rect 14197 6341 14231 6375
rect 15301 6341 15335 6375
rect 16773 6341 16807 6375
rect 17693 6341 17727 6375
rect 19349 6341 19383 6375
rect 22477 6341 22511 6375
rect 23857 6341 23891 6375
rect 1777 6273 1811 6307
rect 2237 6273 2271 6307
rect 2329 6273 2363 6307
rect 3893 6273 3927 6307
rect 4537 6273 4571 6307
rect 6561 6273 6595 6307
rect 7573 6273 7607 6307
rect 8769 6273 8803 6307
rect 9965 6273 9999 6307
rect 11161 6273 11195 6307
rect 11805 6273 11839 6307
rect 12357 6273 12391 6307
rect 12633 6273 12667 6307
rect 13001 6273 13035 6307
rect 13553 6273 13587 6307
rect 14657 6273 14691 6307
rect 15117 6273 15151 6307
rect 15945 6273 15979 6307
rect 17417 6273 17451 6307
rect 18337 6273 18371 6307
rect 19993 6273 20027 6307
rect 20177 6273 20211 6307
rect 20545 6273 20579 6307
rect 21005 6273 21039 6307
rect 21373 6273 21407 6307
rect 22017 6273 22051 6307
rect 23121 6273 23155 6307
rect 23673 6273 23707 6307
rect 20729 6137 20763 6171
rect 14841 6069 14875 6103
rect 22569 6069 22603 6103
rect 6101 5865 6135 5899
rect 7389 5865 7423 5899
rect 8585 5865 8619 5899
rect 9689 5865 9723 5899
rect 10885 5865 10919 5899
rect 12265 5865 12299 5899
rect 13277 5865 13311 5899
rect 14381 5865 14415 5899
rect 15761 5865 15795 5899
rect 16957 5865 16991 5899
rect 18245 5865 18279 5899
rect 19809 5865 19843 5899
rect 24133 5865 24167 5899
rect 11805 5797 11839 5831
rect 6285 5661 6319 5695
rect 7573 5661 7607 5695
rect 8769 5661 8803 5695
rect 9873 5661 9907 5695
rect 11069 5661 11103 5695
rect 11989 5661 12023 5695
rect 12449 5661 12483 5695
rect 13461 5661 13495 5695
rect 14565 5661 14599 5695
rect 14841 5661 14875 5695
rect 15945 5661 15979 5695
rect 17141 5661 17175 5695
rect 18429 5661 18463 5695
rect 19993 5661 20027 5695
rect 23857 5593 23891 5627
rect 14657 5525 14691 5559
rect 6377 5321 6411 5355
rect 7573 5321 7607 5355
rect 8769 5321 8803 5355
rect 9873 5321 9907 5355
rect 11069 5321 11103 5355
rect 11989 5321 12023 5355
rect 12449 5321 12483 5355
rect 13461 5321 13495 5355
rect 14565 5321 14599 5355
rect 14841 5321 14875 5355
rect 15945 5321 15979 5355
rect 17141 5321 17175 5355
rect 18429 5321 18463 5355
rect 19993 5321 20027 5355
rect 24133 5321 24167 5355
rect 6561 5185 6595 5219
rect 7757 5185 7791 5219
rect 8953 5185 8987 5219
rect 10057 5185 10091 5219
rect 11253 5185 11287 5219
rect 12173 5185 12207 5219
rect 12633 5185 12667 5219
rect 13185 5185 13219 5219
rect 13645 5185 13679 5219
rect 14749 5185 14783 5219
rect 15025 5185 15059 5219
rect 16129 5185 16163 5219
rect 17325 5185 17359 5219
rect 18613 5185 18647 5219
rect 20177 5185 20211 5219
rect 24317 5185 24351 5219
rect 8493 5117 8527 5151
rect 24041 4777 24075 4811
rect 23765 4709 23799 4743
rect 23949 4573 23983 4607
rect 24225 4573 24259 4607
rect 23949 3689 23983 3723
rect 24133 3485 24167 3519
rect 24133 3145 24167 3179
rect 23489 3009 23523 3043
rect 23765 3009 23799 3043
rect 24041 3009 24075 3043
rect 24317 3009 24351 3043
rect 23305 2805 23339 2839
rect 23581 2805 23615 2839
rect 23857 2805 23891 2839
rect 1593 2601 1627 2635
rect 22569 2601 22603 2635
rect 23213 2601 23247 2635
rect 1685 2533 1719 2567
rect 6285 2533 6319 2567
rect 7205 2533 7239 2567
rect 10977 2533 11011 2567
rect 11529 2533 11563 2567
rect 16589 2533 16623 2567
rect 17141 2533 17175 2567
rect 19533 2533 19567 2567
rect 23489 2533 23523 2567
rect 23765 2533 23799 2567
rect 1409 2397 1443 2431
rect 1869 2397 1903 2431
rect 2145 2397 2179 2431
rect 2237 2397 2271 2431
rect 4905 2397 4939 2431
rect 6101 2397 6135 2431
rect 7389 2397 7423 2431
rect 9597 2397 9631 2431
rect 9873 2397 9907 2431
rect 10425 2397 10459 2431
rect 11161 2397 11195 2431
rect 11713 2397 11747 2431
rect 11989 2397 12023 2431
rect 12265 2397 12299 2431
rect 12541 2397 12575 2431
rect 12817 2397 12851 2431
rect 13277 2397 13311 2431
rect 15301 2397 15335 2431
rect 15577 2397 15611 2431
rect 15945 2397 15979 2431
rect 16497 2397 16531 2431
rect 16773 2397 16807 2431
rect 17049 2397 17083 2431
rect 17325 2397 17359 2431
rect 17601 2397 17635 2431
rect 17877 2397 17911 2431
rect 18153 2397 18187 2431
rect 18429 2397 18463 2431
rect 18705 2397 18739 2431
rect 18981 2397 19015 2431
rect 19441 2397 19475 2431
rect 19717 2397 19751 2431
rect 19993 2397 20027 2431
rect 20269 2397 20303 2431
rect 20545 2397 20579 2431
rect 20821 2397 20855 2431
rect 22385 2397 22419 2431
rect 22845 2397 22879 2431
rect 23121 2397 23155 2431
rect 23397 2397 23431 2431
rect 23673 2397 23707 2431
rect 23949 2397 23983 2431
rect 24225 2397 24259 2431
rect 1961 2261 1995 2295
rect 2421 2261 2455 2295
rect 4721 2261 4755 2295
rect 9413 2261 9447 2295
rect 9689 2261 9723 2295
rect 10241 2261 10275 2295
rect 11805 2261 11839 2295
rect 12081 2261 12115 2295
rect 12357 2261 12391 2295
rect 12633 2261 12667 2295
rect 13093 2261 13127 2295
rect 15117 2261 15151 2295
rect 15393 2261 15427 2295
rect 16129 2261 16163 2295
rect 16313 2261 16347 2295
rect 16865 2261 16899 2295
rect 17417 2261 17451 2295
rect 17693 2261 17727 2295
rect 17969 2261 18003 2295
rect 18245 2261 18279 2295
rect 18521 2261 18555 2295
rect 18797 2261 18831 2295
rect 19257 2261 19291 2295
rect 19809 2261 19843 2295
rect 20085 2261 20119 2295
rect 20361 2261 20395 2295
rect 20637 2261 20671 2295
rect 22661 2261 22695 2295
rect 22937 2261 22971 2295
rect 24041 2261 24075 2295
rect 2329 2057 2363 2091
rect 2697 2057 2731 2091
rect 7205 2057 7239 2091
rect 7573 2057 7607 2091
rect 7849 2057 7883 2091
rect 8953 2057 8987 2091
rect 9229 2057 9263 2091
rect 9505 2057 9539 2091
rect 14197 2057 14231 2091
rect 17417 2057 17451 2091
rect 17693 2057 17727 2091
rect 20913 2057 20947 2091
rect 21281 2057 21315 2091
rect 21465 2057 21499 2091
rect 21833 2057 21867 2091
rect 22293 2057 22327 2091
rect 22753 2057 22787 2091
rect 23213 2057 23247 2091
rect 10977 1989 11011 2023
rect 11989 1989 12023 2023
rect 15853 1989 15887 2023
rect 18061 1989 18095 2023
rect 18613 1989 18647 2023
rect 19717 1989 19751 2023
rect 20269 1989 20303 2023
rect 20821 1989 20855 2023
rect 1685 1921 1719 1955
rect 1777 1921 1811 1955
rect 2145 1921 2179 1955
rect 2605 1921 2639 1955
rect 2881 1921 2915 1955
rect 3157 1921 3191 1955
rect 3433 1921 3467 1955
rect 3709 1921 3743 1955
rect 3985 1921 4019 1955
rect 4261 1921 4295 1955
rect 4537 1921 4571 1955
rect 4813 1921 4847 1955
rect 5089 1921 5123 1955
rect 5365 1921 5399 1955
rect 5641 1921 5675 1955
rect 5733 1921 5767 1955
rect 6193 1921 6227 1955
rect 6653 1921 6687 1955
rect 6929 1921 6963 1955
rect 7021 1921 7055 1955
rect 7481 1921 7515 1955
rect 7757 1921 7791 1955
rect 8033 1921 8067 1955
rect 8309 1921 8343 1955
rect 8585 1921 8619 1955
rect 8861 1921 8895 1955
rect 9137 1921 9171 1955
rect 9413 1921 9447 1955
rect 9689 1921 9723 1955
rect 9965 1921 9999 1955
rect 10241 1921 10275 1955
rect 10425 1921 10459 1955
rect 11529 1921 11563 1955
rect 12633 1921 12667 1955
rect 12817 1921 12851 1955
rect 13461 1921 13495 1955
rect 13737 1921 13771 1955
rect 14105 1921 14139 1955
rect 14381 1921 14415 1955
rect 14473 1921 14507 1955
rect 14841 1921 14875 1955
rect 15393 1921 15427 1955
rect 15669 1921 15703 1955
rect 16497 1921 16531 1955
rect 16957 1921 16991 1955
rect 17601 1921 17635 1955
rect 17877 1921 17911 1955
rect 19165 1921 19199 1955
rect 21097 1921 21131 1955
rect 21649 1921 21683 1955
rect 22017 1921 22051 1955
rect 22109 1921 22143 1955
rect 22661 1921 22695 1955
rect 22937 1921 22971 1955
rect 23029 1921 23063 1955
rect 23581 1921 23615 1955
rect 23857 1921 23891 1955
rect 24133 1921 24167 1955
rect 24225 1921 24259 1955
rect 2421 1785 2455 1819
rect 2973 1785 3007 1819
rect 3801 1785 3835 1819
rect 4077 1785 4111 1819
rect 4629 1785 4663 1819
rect 4905 1785 4939 1819
rect 5917 1785 5951 1819
rect 10057 1785 10091 1819
rect 13277 1785 13311 1819
rect 15209 1785 15243 1819
rect 19441 1785 19475 1819
rect 22477 1785 22511 1819
rect 23397 1785 23431 1819
rect 23949 1785 23983 1819
rect 1501 1717 1535 1751
rect 1961 1717 1995 1751
rect 3249 1717 3283 1751
rect 3525 1717 3559 1751
rect 4353 1717 4387 1751
rect 5181 1717 5215 1751
rect 5457 1717 5491 1751
rect 6009 1717 6043 1751
rect 6469 1717 6503 1751
rect 6745 1717 6779 1751
rect 7297 1717 7331 1751
rect 8125 1717 8159 1751
rect 8401 1717 8435 1751
rect 8677 1717 8711 1751
rect 9781 1717 9815 1751
rect 10517 1717 10551 1751
rect 11069 1717 11103 1751
rect 11713 1717 11747 1751
rect 12081 1717 12115 1751
rect 12449 1717 12483 1751
rect 12909 1717 12943 1751
rect 13553 1717 13587 1751
rect 13921 1717 13955 1751
rect 14657 1717 14691 1751
rect 15025 1717 15059 1751
rect 15485 1717 15519 1751
rect 15945 1717 15979 1751
rect 16313 1717 16347 1751
rect 17049 1717 17083 1751
rect 18153 1717 18187 1751
rect 18705 1717 18739 1751
rect 19809 1717 19843 1751
rect 20361 1717 20395 1751
rect 23673 1717 23707 1751
rect 24409 1717 24443 1751
rect 2605 1513 2639 1547
rect 2881 1513 2915 1547
rect 6653 1513 6687 1547
rect 11529 1513 11563 1547
rect 14289 1513 14323 1547
rect 15393 1513 15427 1547
rect 15945 1513 15979 1547
rect 16313 1513 16347 1547
rect 16865 1513 16899 1547
rect 17417 1513 17451 1547
rect 18521 1513 18555 1547
rect 19441 1513 19475 1547
rect 21097 1513 21131 1547
rect 21465 1513 21499 1547
rect 23213 1513 23247 1547
rect 1501 1445 1535 1479
rect 3433 1445 3467 1479
rect 7205 1445 7239 1479
rect 20085 1445 20119 1479
rect 20637 1445 20671 1479
rect 11069 1377 11103 1411
rect 1685 1309 1719 1343
rect 1777 1309 1811 1343
rect 2237 1309 2271 1343
rect 2513 1309 2547 1343
rect 2789 1309 2823 1343
rect 3065 1309 3099 1343
rect 3341 1309 3375 1343
rect 3617 1309 3651 1343
rect 3985 1309 4019 1343
rect 4261 1309 4295 1343
rect 4537 1309 4571 1343
rect 4629 1309 4663 1343
rect 4905 1309 4939 1343
rect 5365 1309 5399 1343
rect 5641 1309 5675 1343
rect 5733 1309 5767 1343
rect 6009 1309 6043 1343
rect 6561 1309 6595 1343
rect 6837 1309 6871 1343
rect 7113 1309 7147 1343
rect 7389 1309 7423 1343
rect 7665 1309 7699 1343
rect 7941 1309 7975 1343
rect 8217 1309 8251 1343
rect 8493 1309 8527 1343
rect 8769 1309 8803 1343
rect 9045 1309 9079 1343
rect 9505 1309 9539 1343
rect 9597 1309 9631 1343
rect 9965 1309 9999 1343
rect 10333 1309 10367 1343
rect 11713 1309 11747 1343
rect 11805 1309 11839 1343
rect 12265 1309 12299 1343
rect 12909 1309 12943 1343
rect 13277 1309 13311 1343
rect 14657 1309 14691 1343
rect 15853 1309 15887 1343
rect 16497 1309 16531 1343
rect 16773 1309 16807 1343
rect 17877 1309 17911 1343
rect 19073 1309 19107 1343
rect 19901 1309 19935 1343
rect 21005 1309 21039 1343
rect 21649 1309 21683 1343
rect 22017 1309 22051 1343
rect 22109 1309 22143 1343
rect 22385 1309 22419 1343
rect 22661 1309 22695 1343
rect 22937 1309 22971 1343
rect 23397 1309 23431 1343
rect 23489 1309 23523 1343
rect 23765 1309 23799 1343
rect 24041 1309 24075 1343
rect 10793 1241 10827 1275
rect 14197 1241 14231 1275
rect 15301 1241 15335 1275
rect 17325 1241 17359 1275
rect 18429 1241 18463 1275
rect 19349 1241 19383 1275
rect 20453 1241 20487 1275
rect 1961 1173 1995 1207
rect 2053 1173 2087 1207
rect 2329 1173 2363 1207
rect 3157 1173 3191 1207
rect 3801 1173 3835 1207
rect 4077 1173 4111 1207
rect 4353 1173 4387 1207
rect 4813 1173 4847 1207
rect 5089 1173 5123 1207
rect 5181 1173 5215 1207
rect 5457 1173 5491 1207
rect 5917 1173 5951 1207
rect 6193 1173 6227 1207
rect 6377 1173 6411 1207
rect 6929 1173 6963 1207
rect 7481 1173 7515 1207
rect 7757 1173 7791 1207
rect 8033 1173 8067 1207
rect 8309 1173 8343 1207
rect 8585 1173 8619 1207
rect 9229 1173 9263 1207
rect 9321 1173 9355 1207
rect 9781 1173 9815 1207
rect 10149 1173 10183 1207
rect 10517 1173 10551 1207
rect 11989 1173 12023 1207
rect 12357 1173 12391 1207
rect 13093 1173 13127 1207
rect 13461 1173 13495 1207
rect 14841 1173 14875 1207
rect 17969 1173 18003 1207
rect 18889 1173 18923 1207
rect 21833 1173 21867 1207
rect 22293 1173 22327 1207
rect 22569 1173 22603 1207
rect 22845 1173 22879 1207
rect 23121 1173 23155 1207
rect 23673 1173 23707 1207
rect 23949 1173 23983 1207
rect 24225 1173 24259 1207
<< metal1 >>
rect 1104 6554 25000 6576
rect 1104 6502 6884 6554
rect 6936 6502 6948 6554
rect 7000 6502 7012 6554
rect 7064 6502 7076 6554
rect 7128 6502 7140 6554
rect 7192 6502 12818 6554
rect 12870 6502 12882 6554
rect 12934 6502 12946 6554
rect 12998 6502 13010 6554
rect 13062 6502 13074 6554
rect 13126 6502 18752 6554
rect 18804 6502 18816 6554
rect 18868 6502 18880 6554
rect 18932 6502 18944 6554
rect 18996 6502 19008 6554
rect 19060 6502 24686 6554
rect 24738 6502 24750 6554
rect 24802 6502 24814 6554
rect 24866 6502 24878 6554
rect 24930 6502 24942 6554
rect 24994 6502 25000 6554
rect 1104 6480 25000 6502
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 2501 6443 2559 6449
rect 2501 6440 2513 6443
rect 2188 6412 2513 6440
rect 2188 6400 2194 6412
rect 2501 6409 2513 6412
rect 2547 6409 2559 6443
rect 2501 6403 2559 6409
rect 3786 6400 3792 6452
rect 3844 6440 3850 6452
rect 4157 6443 4215 6449
rect 4157 6440 4169 6443
rect 3844 6412 4169 6440
rect 3844 6400 3850 6412
rect 4157 6409 4169 6412
rect 4203 6409 4215 6443
rect 4157 6403 4215 6409
rect 4614 6400 4620 6452
rect 4672 6400 4678 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 5736 6412 6377 6440
rect 1394 6332 1400 6384
rect 1452 6332 1458 6384
rect 5626 6372 5632 6384
rect 2332 6344 5632 6372
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6304 1823 6307
rect 2222 6304 2228 6316
rect 1811 6276 2228 6304
rect 1811 6273 1823 6276
rect 1765 6267 1823 6273
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 2332 6313 2360 6344
rect 5626 6332 5632 6344
rect 5684 6332 5690 6384
rect 5736 6381 5764 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 7193 6443 7251 6449
rect 7193 6409 7205 6443
rect 7239 6440 7251 6443
rect 7282 6440 7288 6452
rect 7239 6412 7288 6440
rect 7239 6409 7251 6412
rect 7193 6403 7251 6409
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 7377 6443 7435 6449
rect 7377 6409 7389 6443
rect 7423 6409 7435 6443
rect 7377 6403 7435 6409
rect 5721 6375 5779 6381
rect 5721 6341 5733 6375
rect 5767 6341 5779 6375
rect 5721 6335 5779 6341
rect 6086 6332 6092 6384
rect 6144 6332 6150 6384
rect 6917 6375 6975 6381
rect 6917 6341 6929 6375
rect 6963 6372 6975 6375
rect 7392 6372 7420 6403
rect 8386 6400 8392 6452
rect 8444 6400 8450 6452
rect 8573 6443 8631 6449
rect 8573 6409 8585 6443
rect 8619 6409 8631 6443
rect 8573 6403 8631 6409
rect 6963 6344 7420 6372
rect 8113 6375 8171 6381
rect 6963 6341 6975 6344
rect 6917 6335 6975 6341
rect 8113 6341 8125 6375
rect 8159 6372 8171 6375
rect 8588 6372 8616 6403
rect 9398 6400 9404 6452
rect 9456 6400 9462 6452
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6409 9827 6443
rect 9769 6403 9827 6409
rect 8159 6344 8616 6372
rect 9309 6375 9367 6381
rect 8159 6341 8171 6344
rect 8113 6335 8171 6341
rect 9309 6341 9321 6375
rect 9355 6372 9367 6375
rect 9784 6372 9812 6403
rect 10594 6400 10600 6452
rect 10652 6400 10658 6452
rect 10965 6443 11023 6449
rect 10965 6409 10977 6443
rect 11011 6409 11023 6443
rect 10965 6403 11023 6409
rect 9355 6344 9812 6372
rect 10505 6375 10563 6381
rect 9355 6341 9367 6344
rect 9309 6335 9367 6341
rect 10505 6341 10517 6375
rect 10551 6372 10563 6375
rect 10980 6372 11008 6403
rect 11974 6400 11980 6452
rect 12032 6400 12038 6452
rect 12161 6443 12219 6449
rect 12161 6409 12173 6443
rect 12207 6409 12219 6443
rect 12161 6403 12219 6409
rect 12437 6443 12495 6449
rect 12437 6409 12449 6443
rect 12483 6409 12495 6443
rect 12437 6403 12495 6409
rect 10551 6344 11008 6372
rect 10551 6341 10563 6344
rect 10505 6335 10563 6341
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6273 2375 6307
rect 2317 6267 2375 6273
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 3896 6100 3924 6267
rect 4540 6236 4568 6267
rect 6546 6264 6552 6316
rect 6604 6264 6610 6316
rect 7558 6264 7564 6316
rect 7616 6264 7622 6316
rect 8754 6264 8760 6316
rect 8812 6264 8818 6316
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 9732 6276 9965 6304
rect 9732 6264 9738 6276
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 11146 6264 11152 6316
rect 11204 6264 11210 6316
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6304 11851 6307
rect 12176 6304 12204 6403
rect 11839 6276 12204 6304
rect 11839 6273 11851 6276
rect 11793 6267 11851 6273
rect 12342 6264 12348 6316
rect 12400 6264 12406 6316
rect 12452 6236 12480 6403
rect 13170 6400 13176 6452
rect 13228 6400 13234 6452
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6409 13415 6443
rect 13357 6403 13415 6409
rect 12618 6264 12624 6316
rect 12676 6264 12682 6316
rect 12989 6307 13047 6313
rect 12989 6273 13001 6307
rect 13035 6304 13047 6307
rect 13372 6304 13400 6403
rect 14274 6400 14280 6452
rect 14332 6400 14338 6452
rect 14921 6443 14979 6449
rect 14921 6409 14933 6443
rect 14967 6409 14979 6443
rect 14921 6403 14979 6409
rect 14185 6375 14243 6381
rect 14185 6341 14197 6375
rect 14231 6372 14243 6375
rect 14936 6372 14964 6403
rect 15378 6400 15384 6452
rect 15436 6400 15442 6452
rect 15749 6443 15807 6449
rect 15749 6409 15761 6443
rect 15795 6409 15807 6443
rect 15749 6403 15807 6409
rect 14231 6344 14964 6372
rect 15289 6375 15347 6381
rect 14231 6341 14243 6344
rect 14185 6335 14243 6341
rect 15289 6341 15301 6375
rect 15335 6372 15347 6375
rect 15764 6372 15792 6403
rect 16850 6400 16856 6452
rect 16908 6400 16914 6452
rect 17221 6443 17279 6449
rect 17221 6409 17233 6443
rect 17267 6409 17279 6443
rect 17221 6403 17279 6409
rect 15335 6344 15792 6372
rect 16761 6375 16819 6381
rect 15335 6341 15347 6344
rect 15289 6335 15347 6341
rect 16761 6341 16773 6375
rect 16807 6372 16819 6375
rect 17236 6372 17264 6403
rect 17770 6400 17776 6452
rect 17828 6400 17834 6452
rect 18141 6443 18199 6449
rect 18141 6409 18153 6443
rect 18187 6409 18199 6443
rect 18141 6403 18199 6409
rect 16807 6344 17264 6372
rect 17681 6375 17739 6381
rect 16807 6341 16819 6344
rect 16761 6335 16819 6341
rect 17681 6341 17693 6375
rect 17727 6372 17739 6375
rect 18156 6372 18184 6403
rect 19426 6400 19432 6452
rect 19484 6400 19490 6452
rect 19797 6443 19855 6449
rect 19797 6409 19809 6443
rect 19843 6409 19855 6443
rect 19797 6403 19855 6409
rect 17727 6344 18184 6372
rect 19337 6375 19395 6381
rect 17727 6341 17739 6344
rect 17681 6335 17739 6341
rect 19337 6341 19349 6375
rect 19383 6372 19395 6375
rect 19812 6372 19840 6403
rect 20346 6400 20352 6452
rect 20404 6400 20410 6452
rect 20809 6443 20867 6449
rect 20809 6409 20821 6443
rect 20855 6409 20867 6443
rect 20809 6403 20867 6409
rect 20824 6372 20852 6403
rect 21542 6400 21548 6452
rect 21600 6400 21606 6452
rect 21821 6443 21879 6449
rect 21821 6409 21833 6443
rect 21867 6409 21879 6443
rect 22925 6443 22983 6449
rect 22925 6440 22937 6443
rect 21821 6403 21879 6409
rect 22480 6412 22937 6440
rect 19383 6344 19840 6372
rect 20180 6344 20852 6372
rect 19383 6341 19395 6344
rect 19337 6335 19395 6341
rect 13035 6276 13400 6304
rect 13035 6273 13047 6276
rect 12989 6267 13047 6273
rect 13538 6264 13544 6316
rect 13596 6264 13602 6316
rect 14642 6264 14648 6316
rect 14700 6264 14706 6316
rect 15102 6264 15108 6316
rect 15160 6264 15166 6316
rect 15654 6264 15660 6316
rect 15712 6304 15718 6316
rect 15933 6307 15991 6313
rect 15933 6304 15945 6307
rect 15712 6276 15945 6304
rect 15712 6264 15718 6276
rect 15933 6273 15945 6276
rect 15979 6273 15991 6307
rect 15933 6267 15991 6273
rect 17402 6264 17408 6316
rect 17460 6264 17466 6316
rect 18322 6264 18328 6316
rect 18380 6264 18386 6316
rect 19978 6264 19984 6316
rect 20036 6264 20042 6316
rect 20180 6313 20208 6344
rect 20165 6307 20223 6313
rect 20165 6273 20177 6307
rect 20211 6273 20223 6307
rect 20165 6267 20223 6273
rect 20530 6264 20536 6316
rect 20588 6264 20594 6316
rect 20993 6307 21051 6313
rect 20993 6273 21005 6307
rect 21039 6273 21051 6307
rect 20993 6267 21051 6273
rect 21361 6307 21419 6313
rect 21361 6273 21373 6307
rect 21407 6304 21419 6307
rect 21836 6304 21864 6403
rect 22480 6381 22508 6412
rect 22925 6409 22937 6412
rect 22971 6409 22983 6443
rect 22925 6403 22983 6409
rect 23477 6443 23535 6449
rect 23477 6409 23489 6443
rect 23523 6409 23535 6443
rect 23477 6403 23535 6409
rect 22465 6375 22523 6381
rect 22465 6341 22477 6375
rect 22511 6341 22523 6375
rect 23492 6372 23520 6403
rect 23658 6400 23664 6452
rect 23716 6440 23722 6452
rect 23937 6443 23995 6449
rect 23937 6440 23949 6443
rect 23716 6412 23949 6440
rect 23716 6400 23722 6412
rect 23937 6409 23949 6412
rect 23983 6409 23995 6443
rect 23937 6403 23995 6409
rect 23845 6375 23903 6381
rect 23845 6372 23857 6375
rect 23492 6344 23857 6372
rect 22465 6335 22523 6341
rect 23845 6341 23857 6344
rect 23891 6341 23903 6375
rect 23845 6335 23903 6341
rect 21407 6276 21864 6304
rect 22005 6307 22063 6313
rect 21407 6273 21419 6276
rect 21361 6267 21419 6273
rect 22005 6273 22017 6307
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 4540 6208 12480 6236
rect 5626 6128 5632 6180
rect 5684 6168 5690 6180
rect 20717 6171 20775 6177
rect 20717 6168 20729 6171
rect 5684 6140 20729 6168
rect 5684 6128 5690 6140
rect 20717 6137 20729 6140
rect 20763 6137 20775 6171
rect 21008 6168 21036 6267
rect 21634 6196 21640 6248
rect 21692 6236 21698 6248
rect 22020 6236 22048 6267
rect 23106 6264 23112 6316
rect 23164 6264 23170 6316
rect 23658 6264 23664 6316
rect 23716 6264 23722 6316
rect 21692 6208 22048 6236
rect 21692 6196 21698 6208
rect 24210 6168 24216 6180
rect 21008 6140 24216 6168
rect 20717 6131 20775 6137
rect 24210 6128 24216 6140
rect 24268 6128 24274 6180
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 3896 6072 14841 6100
rect 14829 6069 14841 6072
rect 14875 6069 14887 6103
rect 14829 6063 14887 6069
rect 22554 6060 22560 6112
rect 22612 6060 22618 6112
rect 1104 6010 24840 6032
rect 1104 5958 3917 6010
rect 3969 5958 3981 6010
rect 4033 5958 4045 6010
rect 4097 5958 4109 6010
rect 4161 5958 4173 6010
rect 4225 5958 9851 6010
rect 9903 5958 9915 6010
rect 9967 5958 9979 6010
rect 10031 5958 10043 6010
rect 10095 5958 10107 6010
rect 10159 5958 15785 6010
rect 15837 5958 15849 6010
rect 15901 5958 15913 6010
rect 15965 5958 15977 6010
rect 16029 5958 16041 6010
rect 16093 5958 21719 6010
rect 21771 5958 21783 6010
rect 21835 5958 21847 6010
rect 21899 5958 21911 6010
rect 21963 5958 21975 6010
rect 22027 5958 24840 6010
rect 1104 5936 24840 5958
rect 6089 5899 6147 5905
rect 6089 5865 6101 5899
rect 6135 5896 6147 5899
rect 6546 5896 6552 5908
rect 6135 5868 6552 5896
rect 6135 5865 6147 5868
rect 6089 5859 6147 5865
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 7377 5899 7435 5905
rect 7377 5865 7389 5899
rect 7423 5896 7435 5899
rect 7558 5896 7564 5908
rect 7423 5868 7564 5896
rect 7423 5865 7435 5868
rect 7377 5859 7435 5865
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 8573 5899 8631 5905
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 8754 5896 8760 5908
rect 8619 5868 8760 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 9674 5856 9680 5908
rect 9732 5856 9738 5908
rect 10873 5899 10931 5905
rect 10873 5865 10885 5899
rect 10919 5896 10931 5899
rect 11146 5896 11152 5908
rect 10919 5868 11152 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 12253 5899 12311 5905
rect 12253 5865 12265 5899
rect 12299 5896 12311 5899
rect 12342 5896 12348 5908
rect 12299 5868 12348 5896
rect 12299 5865 12311 5868
rect 12253 5859 12311 5865
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 12618 5856 12624 5908
rect 12676 5856 12682 5908
rect 13265 5899 13323 5905
rect 13265 5865 13277 5899
rect 13311 5896 13323 5899
rect 13538 5896 13544 5908
rect 13311 5868 13544 5896
rect 13311 5865 13323 5868
rect 13265 5859 13323 5865
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 14642 5896 14648 5908
rect 14415 5868 14648 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 15102 5856 15108 5908
rect 15160 5856 15166 5908
rect 15654 5856 15660 5908
rect 15712 5896 15718 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15712 5868 15761 5896
rect 15712 5856 15718 5868
rect 15749 5865 15761 5868
rect 15795 5865 15807 5899
rect 15749 5859 15807 5865
rect 16945 5899 17003 5905
rect 16945 5865 16957 5899
rect 16991 5896 17003 5899
rect 17402 5896 17408 5908
rect 16991 5868 17408 5896
rect 16991 5865 17003 5868
rect 16945 5859 17003 5865
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 18233 5899 18291 5905
rect 18233 5865 18245 5899
rect 18279 5896 18291 5899
rect 18322 5896 18328 5908
rect 18279 5868 18328 5896
rect 18279 5865 18291 5868
rect 18233 5859 18291 5865
rect 18322 5856 18328 5868
rect 18380 5856 18386 5908
rect 19797 5899 19855 5905
rect 19797 5865 19809 5899
rect 19843 5896 19855 5899
rect 20530 5896 20536 5908
rect 19843 5868 20536 5896
rect 19843 5865 19855 5868
rect 19797 5859 19855 5865
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 24121 5899 24179 5905
rect 24121 5865 24133 5899
rect 24167 5896 24179 5899
rect 24486 5896 24492 5908
rect 24167 5868 24492 5896
rect 24167 5865 24179 5868
rect 24121 5859 24179 5865
rect 24486 5856 24492 5868
rect 24544 5856 24550 5908
rect 11793 5831 11851 5837
rect 11793 5797 11805 5831
rect 11839 5828 11851 5831
rect 12636 5828 12664 5856
rect 11839 5800 12664 5828
rect 11839 5797 11851 5800
rect 11793 5791 11851 5797
rect 6270 5652 6276 5704
rect 6328 5652 6334 5704
rect 7558 5652 7564 5704
rect 7616 5652 7622 5704
rect 8754 5652 8760 5704
rect 8812 5652 8818 5704
rect 9858 5652 9864 5704
rect 9916 5652 9922 5704
rect 11054 5652 11060 5704
rect 11112 5652 11118 5704
rect 11974 5652 11980 5704
rect 12032 5652 12038 5704
rect 12434 5652 12440 5704
rect 12492 5652 12498 5704
rect 13446 5652 13452 5704
rect 13504 5652 13510 5704
rect 14550 5652 14556 5704
rect 14608 5652 14614 5704
rect 14826 5652 14832 5704
rect 14884 5652 14890 5704
rect 14645 5559 14703 5565
rect 14645 5525 14657 5559
rect 14691 5556 14703 5559
rect 15120 5556 15148 5856
rect 19978 5788 19984 5840
rect 20036 5828 20042 5840
rect 24026 5828 24032 5840
rect 20036 5800 24032 5828
rect 20036 5788 20042 5800
rect 24026 5788 24032 5800
rect 24084 5788 24090 5840
rect 15930 5652 15936 5704
rect 15988 5652 15994 5704
rect 17126 5652 17132 5704
rect 17184 5652 17190 5704
rect 18414 5652 18420 5704
rect 18472 5652 18478 5704
rect 19978 5652 19984 5704
rect 20036 5652 20042 5704
rect 23842 5584 23848 5636
rect 23900 5584 23906 5636
rect 14691 5528 15148 5556
rect 14691 5525 14703 5528
rect 14645 5519 14703 5525
rect 1104 5466 25000 5488
rect 1104 5414 6884 5466
rect 6936 5414 6948 5466
rect 7000 5414 7012 5466
rect 7064 5414 7076 5466
rect 7128 5414 7140 5466
rect 7192 5414 12818 5466
rect 12870 5414 12882 5466
rect 12934 5414 12946 5466
rect 12998 5414 13010 5466
rect 13062 5414 13074 5466
rect 13126 5414 18752 5466
rect 18804 5414 18816 5466
rect 18868 5414 18880 5466
rect 18932 5414 18944 5466
rect 18996 5414 19008 5466
rect 19060 5414 24686 5466
rect 24738 5414 24750 5466
rect 24802 5414 24814 5466
rect 24866 5414 24878 5466
rect 24930 5414 24942 5466
rect 24994 5414 25000 5466
rect 1104 5392 25000 5414
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 6328 5324 6377 5352
rect 6328 5312 6334 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 7558 5312 7564 5364
rect 7616 5312 7622 5364
rect 8754 5312 8760 5364
rect 8812 5312 8818 5364
rect 9858 5312 9864 5364
rect 9916 5312 9922 5364
rect 11054 5312 11060 5364
rect 11112 5312 11118 5364
rect 11974 5312 11980 5364
rect 12032 5312 12038 5364
rect 12434 5312 12440 5364
rect 12492 5312 12498 5364
rect 13446 5312 13452 5364
rect 13504 5312 13510 5364
rect 14550 5312 14556 5364
rect 14608 5312 14614 5364
rect 14826 5312 14832 5364
rect 14884 5312 14890 5364
rect 15930 5312 15936 5364
rect 15988 5312 15994 5364
rect 17126 5312 17132 5364
rect 17184 5312 17190 5364
rect 18414 5312 18420 5364
rect 18472 5312 18478 5364
rect 19978 5312 19984 5364
rect 20036 5312 20042 5364
rect 23842 5312 23848 5364
rect 23900 5352 23906 5364
rect 24121 5355 24179 5361
rect 24121 5352 24133 5355
rect 23900 5324 24133 5352
rect 23900 5312 23906 5324
rect 24121 5321 24133 5324
rect 24167 5321 24179 5355
rect 24121 5315 24179 5321
rect 13906 5284 13912 5296
rect 10060 5256 13912 5284
rect 6546 5176 6552 5228
rect 6604 5176 6610 5228
rect 10060 5225 10088 5256
rect 13906 5244 13912 5256
rect 13964 5244 13970 5296
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 8941 5219 8999 5225
rect 8941 5185 8953 5219
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5185 10103 5219
rect 10045 5179 10103 5185
rect 7760 5012 7788 5179
rect 8481 5151 8539 5157
rect 8481 5117 8493 5151
rect 8527 5148 8539 5151
rect 8956 5148 8984 5179
rect 11238 5176 11244 5228
rect 11296 5176 11302 5228
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5216 12219 5219
rect 12621 5219 12679 5225
rect 12207 5188 12434 5216
rect 12207 5185 12219 5188
rect 12161 5179 12219 5185
rect 9582 5148 9588 5160
rect 8527 5120 9588 5148
rect 8527 5117 8539 5120
rect 8481 5111 8539 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 12406 5080 12434 5188
rect 12621 5185 12633 5219
rect 12667 5185 12679 5219
rect 12621 5179 12679 5185
rect 13173 5219 13231 5225
rect 13173 5185 13185 5219
rect 13219 5216 13231 5219
rect 13633 5219 13691 5225
rect 13633 5216 13645 5219
rect 13219 5188 13645 5216
rect 13219 5185 13231 5188
rect 13173 5179 13231 5185
rect 13633 5185 13645 5188
rect 13679 5216 13691 5219
rect 13722 5216 13728 5228
rect 13679 5188 13728 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 12636 5148 12664 5179
rect 13722 5176 13728 5188
rect 13780 5176 13786 5228
rect 14734 5176 14740 5228
rect 14792 5176 14798 5228
rect 15010 5176 15016 5228
rect 15068 5176 15074 5228
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 17313 5219 17371 5225
rect 17313 5185 17325 5219
rect 17359 5216 17371 5219
rect 17862 5216 17868 5228
rect 17359 5188 17868 5216
rect 17359 5185 17371 5188
rect 17313 5179 17371 5185
rect 12636 5120 15976 5148
rect 13630 5080 13636 5092
rect 12406 5052 13636 5080
rect 13630 5040 13636 5052
rect 13688 5040 13694 5092
rect 12618 5012 12624 5024
rect 7760 4984 12624 5012
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 15948 5012 15976 5120
rect 16132 5080 16160 5179
rect 17862 5176 17868 5188
rect 17920 5176 17926 5228
rect 18601 5219 18659 5225
rect 18601 5185 18613 5219
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 20165 5219 20223 5225
rect 20165 5185 20177 5219
rect 20211 5216 20223 5219
rect 21450 5216 21456 5228
rect 20211 5188 21456 5216
rect 20211 5185 20223 5188
rect 20165 5179 20223 5185
rect 18616 5148 18644 5179
rect 21450 5176 21456 5188
rect 21508 5176 21514 5228
rect 24302 5176 24308 5228
rect 24360 5176 24366 5228
rect 21358 5148 21364 5160
rect 18616 5120 21364 5148
rect 21358 5108 21364 5120
rect 21416 5108 21422 5160
rect 21266 5080 21272 5092
rect 16132 5052 21272 5080
rect 21266 5040 21272 5052
rect 21324 5040 21330 5092
rect 16390 5012 16396 5024
rect 15948 4984 16396 5012
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 1104 4922 24840 4944
rect 1104 4870 3917 4922
rect 3969 4870 3981 4922
rect 4033 4870 4045 4922
rect 4097 4870 4109 4922
rect 4161 4870 4173 4922
rect 4225 4870 9851 4922
rect 9903 4870 9915 4922
rect 9967 4870 9979 4922
rect 10031 4870 10043 4922
rect 10095 4870 10107 4922
rect 10159 4870 15785 4922
rect 15837 4870 15849 4922
rect 15901 4870 15913 4922
rect 15965 4870 15977 4922
rect 16029 4870 16041 4922
rect 16093 4870 21719 4922
rect 21771 4870 21783 4922
rect 21835 4870 21847 4922
rect 21899 4870 21911 4922
rect 21963 4870 21975 4922
rect 22027 4870 24840 4922
rect 1104 4848 24840 4870
rect 6546 4768 6552 4820
rect 6604 4808 6610 4820
rect 24029 4811 24087 4817
rect 6604 4780 12434 4808
rect 6604 4768 6610 4780
rect 12406 4672 12434 4780
rect 24029 4777 24041 4811
rect 24075 4808 24087 4811
rect 24302 4808 24308 4820
rect 24075 4780 24308 4808
rect 24075 4777 24087 4780
rect 24029 4771 24087 4777
rect 24302 4768 24308 4780
rect 24360 4768 24366 4820
rect 23753 4743 23811 4749
rect 23753 4709 23765 4743
rect 23799 4709 23811 4743
rect 23753 4703 23811 4709
rect 13354 4672 13360 4684
rect 12406 4644 13360 4672
rect 13354 4632 13360 4644
rect 13412 4632 13418 4684
rect 23768 4672 23796 4703
rect 23768 4644 24256 4672
rect 23934 4564 23940 4616
rect 23992 4564 23998 4616
rect 24228 4613 24256 4644
rect 24213 4607 24271 4613
rect 24213 4573 24225 4607
rect 24259 4573 24271 4607
rect 24213 4567 24271 4573
rect 1104 4378 25000 4400
rect 1104 4326 6884 4378
rect 6936 4326 6948 4378
rect 7000 4326 7012 4378
rect 7064 4326 7076 4378
rect 7128 4326 7140 4378
rect 7192 4326 12818 4378
rect 12870 4326 12882 4378
rect 12934 4326 12946 4378
rect 12998 4326 13010 4378
rect 13062 4326 13074 4378
rect 13126 4326 18752 4378
rect 18804 4326 18816 4378
rect 18868 4326 18880 4378
rect 18932 4326 18944 4378
rect 18996 4326 19008 4378
rect 19060 4326 24686 4378
rect 24738 4326 24750 4378
rect 24802 4326 24814 4378
rect 24866 4326 24878 4378
rect 24930 4326 24942 4378
rect 24994 4326 25000 4378
rect 1104 4304 25000 4326
rect 1104 3834 24840 3856
rect 1104 3782 3917 3834
rect 3969 3782 3981 3834
rect 4033 3782 4045 3834
rect 4097 3782 4109 3834
rect 4161 3782 4173 3834
rect 4225 3782 9851 3834
rect 9903 3782 9915 3834
rect 9967 3782 9979 3834
rect 10031 3782 10043 3834
rect 10095 3782 10107 3834
rect 10159 3782 15785 3834
rect 15837 3782 15849 3834
rect 15901 3782 15913 3834
rect 15965 3782 15977 3834
rect 16029 3782 16041 3834
rect 16093 3782 21719 3834
rect 21771 3782 21783 3834
rect 21835 3782 21847 3834
rect 21899 3782 21911 3834
rect 21963 3782 21975 3834
rect 22027 3782 24840 3834
rect 1104 3760 24840 3782
rect 23658 3680 23664 3732
rect 23716 3720 23722 3732
rect 23937 3723 23995 3729
rect 23937 3720 23949 3723
rect 23716 3692 23949 3720
rect 23716 3680 23722 3692
rect 23937 3689 23949 3692
rect 23983 3689 23995 3723
rect 23937 3683 23995 3689
rect 24118 3476 24124 3528
rect 24176 3476 24182 3528
rect 23198 3340 23204 3392
rect 23256 3380 23262 3392
rect 24302 3380 24308 3392
rect 23256 3352 24308 3380
rect 23256 3340 23262 3352
rect 24302 3340 24308 3352
rect 24360 3340 24366 3392
rect 1104 3290 25000 3312
rect 1104 3238 6884 3290
rect 6936 3238 6948 3290
rect 7000 3238 7012 3290
rect 7064 3238 7076 3290
rect 7128 3238 7140 3290
rect 7192 3238 12818 3290
rect 12870 3238 12882 3290
rect 12934 3238 12946 3290
rect 12998 3238 13010 3290
rect 13062 3238 13074 3290
rect 13126 3238 18752 3290
rect 18804 3238 18816 3290
rect 18868 3238 18880 3290
rect 18932 3238 18944 3290
rect 18996 3238 19008 3290
rect 19060 3238 24686 3290
rect 24738 3238 24750 3290
rect 24802 3238 24814 3290
rect 24866 3238 24878 3290
rect 24930 3238 24942 3290
rect 24994 3238 25000 3290
rect 1104 3216 25000 3238
rect 24118 3136 24124 3188
rect 24176 3136 24182 3188
rect 25038 3108 25044 3120
rect 23492 3080 25044 3108
rect 23492 3049 23520 3080
rect 25038 3068 25044 3080
rect 25096 3068 25102 3120
rect 23477 3043 23535 3049
rect 23477 3009 23489 3043
rect 23523 3009 23535 3043
rect 23477 3003 23535 3009
rect 23753 3043 23811 3049
rect 23753 3009 23765 3043
rect 23799 3009 23811 3043
rect 23753 3003 23811 3009
rect 24029 3043 24087 3049
rect 24029 3009 24041 3043
rect 24075 3009 24087 3043
rect 24029 3003 24087 3009
rect 1578 2932 1584 2984
rect 1636 2972 1642 2984
rect 14366 2972 14372 2984
rect 1636 2944 14372 2972
rect 1636 2932 1642 2944
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 17862 2864 17868 2916
rect 17920 2904 17926 2916
rect 22646 2904 22652 2916
rect 17920 2876 22652 2904
rect 17920 2864 17926 2876
rect 22646 2864 22652 2876
rect 22704 2864 22710 2916
rect 23768 2904 23796 3003
rect 24044 2972 24072 3003
rect 24302 3000 24308 3052
rect 24360 3000 24366 3052
rect 24486 2972 24492 2984
rect 24044 2944 24492 2972
rect 24486 2932 24492 2944
rect 24544 2932 24550 2984
rect 24578 2904 24584 2916
rect 23768 2876 24584 2904
rect 24578 2864 24584 2876
rect 24636 2864 24642 2916
rect 9490 2796 9496 2848
rect 9548 2836 9554 2848
rect 12526 2836 12532 2848
rect 9548 2808 12532 2836
rect 9548 2796 9554 2808
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 13170 2796 13176 2848
rect 13228 2836 13234 2848
rect 15562 2836 15568 2848
rect 13228 2808 15568 2836
rect 13228 2796 13234 2808
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 19610 2796 19616 2848
rect 19668 2836 19674 2848
rect 20990 2836 20996 2848
rect 19668 2808 20996 2836
rect 19668 2796 19674 2808
rect 20990 2796 20996 2808
rect 21048 2796 21054 2848
rect 23014 2796 23020 2848
rect 23072 2836 23078 2848
rect 23293 2839 23351 2845
rect 23293 2836 23305 2839
rect 23072 2808 23305 2836
rect 23072 2796 23078 2808
rect 23293 2805 23305 2808
rect 23339 2805 23351 2839
rect 23293 2799 23351 2805
rect 23566 2796 23572 2848
rect 23624 2796 23630 2848
rect 23845 2839 23903 2845
rect 23845 2805 23857 2839
rect 23891 2836 23903 2839
rect 24026 2836 24032 2848
rect 23891 2808 24032 2836
rect 23891 2805 23903 2808
rect 23845 2799 23903 2805
rect 24026 2796 24032 2808
rect 24084 2796 24090 2848
rect 1104 2746 24840 2768
rect 1104 2694 3917 2746
rect 3969 2694 3981 2746
rect 4033 2694 4045 2746
rect 4097 2694 4109 2746
rect 4161 2694 4173 2746
rect 4225 2694 9851 2746
rect 9903 2694 9915 2746
rect 9967 2694 9979 2746
rect 10031 2694 10043 2746
rect 10095 2694 10107 2746
rect 10159 2694 15785 2746
rect 15837 2694 15849 2746
rect 15901 2694 15913 2746
rect 15965 2694 15977 2746
rect 16029 2694 16041 2746
rect 16093 2694 21719 2746
rect 21771 2694 21783 2746
rect 21835 2694 21847 2746
rect 21899 2694 21911 2746
rect 21963 2694 21975 2746
rect 22027 2694 24840 2746
rect 1104 2672 24840 2694
rect 1578 2592 1584 2644
rect 1636 2592 1642 2644
rect 2590 2592 2596 2644
rect 2648 2632 2654 2644
rect 9122 2632 9128 2644
rect 2648 2604 9128 2632
rect 2648 2592 2654 2604
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 9232 2604 14964 2632
rect 1673 2567 1731 2573
rect 1673 2533 1685 2567
rect 1719 2564 1731 2567
rect 5718 2564 5724 2576
rect 1719 2536 5724 2564
rect 1719 2533 1731 2536
rect 1673 2527 1731 2533
rect 5718 2524 5724 2536
rect 5776 2524 5782 2576
rect 6270 2524 6276 2576
rect 6328 2524 6334 2576
rect 7190 2524 7196 2576
rect 7248 2524 7254 2576
rect 7558 2524 7564 2576
rect 7616 2564 7622 2576
rect 9232 2564 9260 2604
rect 7616 2536 9260 2564
rect 10965 2567 11023 2573
rect 7616 2524 7622 2536
rect 10965 2533 10977 2567
rect 11011 2533 11023 2567
rect 10965 2527 11023 2533
rect 11517 2567 11575 2573
rect 11517 2533 11529 2567
rect 11563 2564 11575 2567
rect 13262 2564 13268 2576
rect 11563 2536 13268 2564
rect 11563 2533 11575 2536
rect 11517 2527 11575 2533
rect 474 2456 480 2508
rect 532 2496 538 2508
rect 532 2468 2176 2496
rect 532 2456 538 2468
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 2148 2437 2176 2468
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 9030 2496 9036 2508
rect 4120 2468 9036 2496
rect 4120 2456 4126 2468
rect 9030 2456 9036 2468
rect 9088 2456 9094 2508
rect 9490 2496 9496 2508
rect 9140 2468 9496 2496
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1360 2400 1409 2428
rect 1360 2388 1366 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1857 2431 1915 2437
rect 1857 2428 1869 2431
rect 1397 2391 1455 2397
rect 1504 2400 1869 2428
rect 198 2320 204 2372
rect 256 2360 262 2372
rect 1504 2360 1532 2400
rect 1857 2397 1869 2400
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2397 2191 2431
rect 2133 2391 2191 2397
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 2240 2360 2268 2391
rect 4890 2388 4896 2440
rect 4948 2388 4954 2440
rect 6086 2388 6092 2440
rect 6144 2388 6150 2440
rect 7374 2388 7380 2440
rect 7432 2388 7438 2440
rect 3326 2360 3332 2372
rect 256 2332 1532 2360
rect 1872 2332 2268 2360
rect 2332 2332 3332 2360
rect 256 2320 262 2332
rect 1872 2304 1900 2332
rect 1854 2252 1860 2304
rect 1912 2252 1918 2304
rect 1949 2295 2007 2301
rect 1949 2261 1961 2295
rect 1995 2292 2007 2295
rect 2332 2292 2360 2332
rect 3326 2320 3332 2332
rect 3384 2320 3390 2372
rect 6730 2360 6736 2372
rect 3436 2332 6736 2360
rect 3436 2304 3464 2332
rect 6730 2320 6736 2332
rect 6788 2320 6794 2372
rect 1995 2264 2360 2292
rect 1995 2261 2007 2264
rect 1949 2255 2007 2261
rect 2406 2252 2412 2304
rect 2464 2252 2470 2304
rect 3418 2252 3424 2304
rect 3476 2252 3482 2304
rect 4430 2252 4436 2304
rect 4488 2292 4494 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 4488 2264 4721 2292
rect 4488 2252 4494 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 5074 2252 5080 2304
rect 5132 2292 5138 2304
rect 9140 2292 9168 2468
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 10980 2496 11008 2527
rect 13262 2524 13268 2536
rect 13320 2524 13326 2576
rect 14936 2564 14964 2604
rect 15010 2592 15016 2644
rect 15068 2632 15074 2644
rect 22557 2635 22615 2641
rect 22557 2632 22569 2635
rect 15068 2604 22569 2632
rect 15068 2592 15074 2604
rect 22557 2601 22569 2604
rect 22603 2601 22615 2635
rect 22557 2595 22615 2601
rect 22646 2592 22652 2644
rect 22704 2592 22710 2644
rect 23198 2592 23204 2644
rect 23256 2592 23262 2644
rect 23400 2604 23612 2632
rect 16577 2567 16635 2573
rect 14936 2536 16068 2564
rect 10980 2468 11744 2496
rect 9306 2388 9312 2440
rect 9364 2428 9370 2440
rect 9585 2431 9643 2437
rect 9585 2428 9597 2431
rect 9364 2400 9597 2428
rect 9364 2388 9370 2400
rect 9585 2397 9597 2400
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 9858 2388 9864 2440
rect 9916 2388 9922 2440
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 9214 2320 9220 2372
rect 9272 2360 9278 2372
rect 10428 2360 10456 2391
rect 10686 2388 10692 2440
rect 10744 2428 10750 2440
rect 11716 2437 11744 2468
rect 11808 2468 12112 2496
rect 11808 2440 11836 2468
rect 11149 2431 11207 2437
rect 11149 2428 11161 2431
rect 10744 2400 11161 2428
rect 10744 2388 10750 2400
rect 11149 2397 11161 2400
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 11701 2431 11759 2437
rect 11701 2397 11713 2431
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 11790 2388 11796 2440
rect 11848 2388 11854 2440
rect 11974 2388 11980 2440
rect 12032 2388 12038 2440
rect 12084 2428 12112 2468
rect 12158 2456 12164 2508
rect 12216 2496 12222 2508
rect 12216 2468 13308 2496
rect 12216 2456 12222 2468
rect 12253 2431 12311 2437
rect 12253 2428 12265 2431
rect 12084 2400 12265 2428
rect 12253 2397 12265 2400
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 13280 2437 13308 2468
rect 14182 2456 14188 2508
rect 14240 2496 14246 2508
rect 14240 2468 15308 2496
rect 14240 2456 14246 2468
rect 15280 2437 15308 2468
rect 15488 2468 15976 2496
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12636 2400 12817 2428
rect 9272 2332 10456 2360
rect 9272 2320 9278 2332
rect 11606 2320 11612 2372
rect 11664 2360 11670 2372
rect 11664 2332 11928 2360
rect 11664 2320 11670 2332
rect 5132 2264 9168 2292
rect 5132 2252 5138 2264
rect 9398 2252 9404 2304
rect 9456 2252 9462 2304
rect 9490 2252 9496 2304
rect 9548 2292 9554 2304
rect 9677 2295 9735 2301
rect 9677 2292 9689 2295
rect 9548 2264 9689 2292
rect 9548 2252 9554 2264
rect 9677 2261 9689 2264
rect 9723 2261 9735 2295
rect 9677 2255 9735 2261
rect 10229 2295 10287 2301
rect 10229 2261 10241 2295
rect 10275 2292 10287 2295
rect 11238 2292 11244 2304
rect 10275 2264 11244 2292
rect 10275 2261 10287 2264
rect 10229 2255 10287 2261
rect 11238 2252 11244 2264
rect 11296 2252 11302 2304
rect 11790 2252 11796 2304
rect 11848 2252 11854 2304
rect 11900 2292 11928 2332
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 12636 2360 12664 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2397 13323 2431
rect 15280 2431 15347 2437
rect 15280 2400 15301 2431
rect 13265 2391 13323 2397
rect 15289 2397 15301 2400
rect 15335 2397 15347 2431
rect 15289 2391 15347 2397
rect 15378 2388 15384 2440
rect 15436 2428 15442 2440
rect 15488 2428 15516 2468
rect 15436 2400 15516 2428
rect 15436 2388 15442 2400
rect 15562 2388 15568 2440
rect 15620 2388 15626 2440
rect 15948 2437 15976 2468
rect 16040 2440 16068 2536
rect 16577 2533 16589 2567
rect 16623 2533 16635 2567
rect 16577 2527 16635 2533
rect 17129 2567 17187 2573
rect 17129 2533 17141 2567
rect 17175 2564 17187 2567
rect 19426 2564 19432 2576
rect 17175 2536 19432 2564
rect 17175 2533 17187 2536
rect 17129 2527 17187 2533
rect 16592 2496 16620 2527
rect 19426 2524 19432 2536
rect 19484 2524 19490 2576
rect 19521 2567 19579 2573
rect 19521 2533 19533 2567
rect 19567 2533 19579 2567
rect 19521 2527 19579 2533
rect 19334 2496 19340 2508
rect 16592 2468 17356 2496
rect 15933 2431 15991 2437
rect 15933 2397 15945 2431
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 16022 2388 16028 2440
rect 16080 2388 16086 2440
rect 16482 2388 16488 2440
rect 16540 2388 16546 2440
rect 16761 2431 16819 2437
rect 16761 2397 16773 2431
rect 16807 2397 16819 2431
rect 16761 2391 16819 2397
rect 12492 2332 12664 2360
rect 12492 2320 12498 2332
rect 14550 2320 14556 2372
rect 14608 2360 14614 2372
rect 16776 2360 16804 2391
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17328 2437 17356 2468
rect 18432 2468 19340 2496
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 17000 2400 17049 2428
rect 17000 2388 17006 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17313 2431 17371 2437
rect 17313 2397 17325 2431
rect 17359 2397 17371 2431
rect 17313 2391 17371 2397
rect 17586 2388 17592 2440
rect 17644 2388 17650 2440
rect 17862 2388 17868 2440
rect 17920 2388 17926 2440
rect 17954 2388 17960 2440
rect 18012 2388 18018 2440
rect 18138 2388 18144 2440
rect 18196 2388 18202 2440
rect 18432 2437 18460 2468
rect 19334 2456 19340 2468
rect 19392 2456 19398 2508
rect 19536 2496 19564 2527
rect 21358 2524 21364 2576
rect 21416 2524 21422 2576
rect 22664 2564 22692 2592
rect 23400 2564 23428 2604
rect 22664 2536 23428 2564
rect 23477 2567 23535 2573
rect 23477 2533 23489 2567
rect 23523 2533 23535 2567
rect 23584 2564 23612 2604
rect 23753 2567 23811 2573
rect 23753 2564 23765 2567
rect 23584 2536 23765 2564
rect 23477 2527 23535 2533
rect 23753 2533 23765 2536
rect 23799 2533 23811 2567
rect 23753 2527 23811 2533
rect 21376 2496 21404 2524
rect 23492 2496 23520 2527
rect 25314 2496 25320 2508
rect 19536 2468 20576 2496
rect 21376 2468 23520 2496
rect 23584 2468 25320 2496
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 18693 2431 18751 2437
rect 18693 2428 18705 2431
rect 18417 2391 18475 2397
rect 18524 2400 18705 2428
rect 17972 2360 18000 2388
rect 18524 2360 18552 2400
rect 18693 2397 18705 2400
rect 18739 2397 18751 2431
rect 18693 2391 18751 2397
rect 18966 2388 18972 2440
rect 19024 2388 19030 2440
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 19444 2360 19472 2391
rect 19702 2388 19708 2440
rect 19760 2388 19766 2440
rect 19981 2431 20039 2437
rect 19981 2397 19993 2431
rect 20027 2428 20039 2431
rect 20070 2428 20076 2440
rect 20027 2400 20076 2428
rect 20027 2397 20039 2400
rect 19981 2391 20039 2397
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 20254 2388 20260 2440
rect 20312 2388 20318 2440
rect 20548 2437 20576 2468
rect 20533 2431 20591 2437
rect 20533 2397 20545 2431
rect 20579 2397 20591 2431
rect 20533 2391 20591 2397
rect 20809 2431 20867 2437
rect 20809 2397 20821 2431
rect 20855 2397 20867 2431
rect 20809 2391 20867 2397
rect 14608 2332 16804 2360
rect 17420 2332 18000 2360
rect 18156 2332 18552 2360
rect 18708 2332 19380 2360
rect 19444 2332 20116 2360
rect 14608 2320 14614 2332
rect 12069 2295 12127 2301
rect 12069 2292 12081 2295
rect 11900 2264 12081 2292
rect 12069 2261 12081 2264
rect 12115 2261 12127 2295
rect 12069 2255 12127 2261
rect 12342 2252 12348 2304
rect 12400 2252 12406 2304
rect 12621 2295 12679 2301
rect 12621 2261 12633 2295
rect 12667 2292 12679 2295
rect 12710 2292 12716 2304
rect 12667 2264 12716 2292
rect 12667 2261 12679 2264
rect 12621 2255 12679 2261
rect 12710 2252 12716 2264
rect 12768 2252 12774 2304
rect 13081 2295 13139 2301
rect 13081 2261 13093 2295
rect 13127 2292 13139 2295
rect 13998 2292 14004 2304
rect 13127 2264 14004 2292
rect 13127 2261 13139 2264
rect 13081 2255 13139 2261
rect 13998 2252 14004 2264
rect 14056 2252 14062 2304
rect 15105 2295 15163 2301
rect 15105 2261 15117 2295
rect 15151 2292 15163 2295
rect 15286 2292 15292 2304
rect 15151 2264 15292 2292
rect 15151 2261 15163 2264
rect 15105 2255 15163 2261
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 15381 2295 15439 2301
rect 15381 2261 15393 2295
rect 15427 2292 15439 2295
rect 15470 2292 15476 2304
rect 15427 2264 15476 2292
rect 15427 2261 15439 2264
rect 15381 2255 15439 2261
rect 15470 2252 15476 2264
rect 15528 2252 15534 2304
rect 15562 2252 15568 2304
rect 15620 2292 15626 2304
rect 16117 2295 16175 2301
rect 16117 2292 16129 2295
rect 15620 2264 16129 2292
rect 15620 2252 15626 2264
rect 16117 2261 16129 2264
rect 16163 2261 16175 2295
rect 16117 2255 16175 2261
rect 16301 2295 16359 2301
rect 16301 2261 16313 2295
rect 16347 2292 16359 2295
rect 16666 2292 16672 2304
rect 16347 2264 16672 2292
rect 16347 2261 16359 2264
rect 16301 2255 16359 2261
rect 16666 2252 16672 2264
rect 16724 2252 16730 2304
rect 16850 2252 16856 2304
rect 16908 2252 16914 2304
rect 17420 2301 17448 2332
rect 18156 2304 18184 2332
rect 17405 2295 17463 2301
rect 17405 2261 17417 2295
rect 17451 2261 17463 2295
rect 17405 2255 17463 2261
rect 17681 2295 17739 2301
rect 17681 2261 17693 2295
rect 17727 2292 17739 2295
rect 17770 2292 17776 2304
rect 17727 2264 17776 2292
rect 17727 2261 17739 2264
rect 17681 2255 17739 2261
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 17957 2295 18015 2301
rect 17957 2261 17969 2295
rect 18003 2292 18015 2295
rect 18046 2292 18052 2304
rect 18003 2264 18052 2292
rect 18003 2261 18015 2264
rect 17957 2255 18015 2261
rect 18046 2252 18052 2264
rect 18104 2252 18110 2304
rect 18138 2252 18144 2304
rect 18196 2252 18202 2304
rect 18230 2252 18236 2304
rect 18288 2252 18294 2304
rect 18509 2295 18567 2301
rect 18509 2261 18521 2295
rect 18555 2292 18567 2295
rect 18708 2292 18736 2332
rect 18555 2264 18736 2292
rect 18785 2295 18843 2301
rect 18555 2261 18567 2264
rect 18509 2255 18567 2261
rect 18785 2261 18797 2295
rect 18831 2292 18843 2295
rect 19150 2292 19156 2304
rect 18831 2264 19156 2292
rect 18831 2261 18843 2264
rect 18785 2255 18843 2261
rect 19150 2252 19156 2264
rect 19208 2252 19214 2304
rect 19242 2252 19248 2304
rect 19300 2252 19306 2304
rect 19352 2292 19380 2332
rect 19702 2292 19708 2304
rect 19352 2264 19708 2292
rect 19702 2252 19708 2264
rect 19760 2252 19766 2304
rect 19797 2295 19855 2301
rect 19797 2261 19809 2295
rect 19843 2292 19855 2295
rect 19978 2292 19984 2304
rect 19843 2264 19984 2292
rect 19843 2261 19855 2264
rect 19797 2255 19855 2261
rect 19978 2252 19984 2264
rect 20036 2252 20042 2304
rect 20088 2301 20116 2332
rect 20162 2320 20168 2372
rect 20220 2360 20226 2372
rect 20824 2360 20852 2391
rect 22370 2388 22376 2440
rect 22428 2388 22434 2440
rect 22830 2388 22836 2440
rect 22888 2388 22894 2440
rect 23109 2431 23167 2437
rect 23109 2397 23121 2431
rect 23155 2428 23167 2431
rect 23290 2428 23296 2440
rect 23155 2400 23296 2428
rect 23155 2397 23167 2400
rect 23109 2391 23167 2397
rect 23290 2388 23296 2400
rect 23348 2388 23354 2440
rect 23385 2431 23443 2437
rect 23385 2397 23397 2431
rect 23431 2428 23443 2431
rect 23584 2428 23612 2468
rect 25314 2456 25320 2468
rect 25372 2456 25378 2508
rect 23431 2400 23612 2428
rect 23661 2431 23719 2437
rect 23431 2397 23443 2400
rect 23385 2391 23443 2397
rect 23661 2397 23673 2431
rect 23707 2397 23719 2431
rect 23661 2391 23719 2397
rect 23676 2360 23704 2391
rect 23750 2388 23756 2440
rect 23808 2428 23814 2440
rect 23937 2431 23995 2437
rect 23937 2428 23949 2431
rect 23808 2400 23949 2428
rect 23808 2388 23814 2400
rect 23937 2397 23949 2400
rect 23983 2397 23995 2431
rect 23937 2391 23995 2397
rect 24026 2388 24032 2440
rect 24084 2428 24090 2440
rect 24213 2431 24271 2437
rect 24213 2428 24225 2431
rect 24084 2400 24225 2428
rect 24084 2388 24090 2400
rect 24213 2397 24225 2400
rect 24259 2397 24271 2431
rect 24213 2391 24271 2397
rect 23842 2360 23848 2372
rect 20220 2332 20852 2360
rect 22940 2332 23428 2360
rect 23676 2332 23848 2360
rect 20220 2320 20226 2332
rect 20073 2295 20131 2301
rect 20073 2261 20085 2295
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 20346 2252 20352 2304
rect 20404 2252 20410 2304
rect 20622 2252 20628 2304
rect 20680 2252 20686 2304
rect 22646 2252 22652 2304
rect 22704 2252 22710 2304
rect 22940 2301 22968 2332
rect 22925 2295 22983 2301
rect 22925 2261 22937 2295
rect 22971 2261 22983 2295
rect 23400 2292 23428 2332
rect 23842 2320 23848 2332
rect 23900 2320 23906 2372
rect 23934 2292 23940 2304
rect 23400 2264 23940 2292
rect 22925 2255 22983 2261
rect 23934 2252 23940 2264
rect 23992 2252 23998 2304
rect 24026 2252 24032 2304
rect 24084 2252 24090 2304
rect 1104 2202 25000 2224
rect 1104 2150 6884 2202
rect 6936 2150 6948 2202
rect 7000 2150 7012 2202
rect 7064 2150 7076 2202
rect 7128 2150 7140 2202
rect 7192 2150 12818 2202
rect 12870 2150 12882 2202
rect 12934 2150 12946 2202
rect 12998 2150 13010 2202
rect 13062 2150 13074 2202
rect 13126 2150 18752 2202
rect 18804 2150 18816 2202
rect 18868 2150 18880 2202
rect 18932 2150 18944 2202
rect 18996 2150 19008 2202
rect 19060 2150 24686 2202
rect 24738 2150 24750 2202
rect 24802 2150 24814 2202
rect 24866 2150 24878 2202
rect 24930 2150 24942 2202
rect 24994 2150 25000 2202
rect 1104 2128 25000 2150
rect 2314 2048 2320 2100
rect 2372 2048 2378 2100
rect 2685 2091 2743 2097
rect 2685 2057 2697 2091
rect 2731 2057 2743 2091
rect 2685 2051 2743 2057
rect 2884 2060 5672 2088
rect 750 1980 756 2032
rect 808 2020 814 2032
rect 2700 2020 2728 2051
rect 2884 2020 2912 2060
rect 5442 2020 5448 2032
rect 808 1992 2636 2020
rect 2700 1992 2912 2020
rect 2976 1992 4476 2020
rect 808 1980 814 1992
rect 1673 1955 1731 1961
rect 1673 1921 1685 1955
rect 1719 1921 1731 1955
rect 1673 1915 1731 1921
rect 1688 1884 1716 1915
rect 1762 1912 1768 1964
rect 1820 1912 1826 1964
rect 2130 1912 2136 1964
rect 2188 1912 2194 1964
rect 2608 1961 2636 1992
rect 2593 1955 2651 1961
rect 2593 1921 2605 1955
rect 2639 1921 2651 1955
rect 2869 1955 2927 1961
rect 2869 1952 2881 1955
rect 2593 1915 2651 1921
rect 2746 1924 2881 1952
rect 1688 1856 2452 1884
rect 1026 1776 1032 1828
rect 1084 1816 1090 1828
rect 2424 1825 2452 1856
rect 2409 1819 2467 1825
rect 1084 1788 2360 1816
rect 1084 1776 1090 1788
rect 1486 1708 1492 1760
rect 1544 1708 1550 1760
rect 1946 1708 1952 1760
rect 2004 1708 2010 1760
rect 2332 1748 2360 1788
rect 2409 1785 2421 1819
rect 2455 1785 2467 1819
rect 2409 1779 2467 1785
rect 2746 1748 2774 1924
rect 2869 1921 2881 1924
rect 2915 1921 2927 1955
rect 2869 1915 2927 1921
rect 2976 1825 3004 1992
rect 3142 1912 3148 1964
rect 3200 1912 3206 1964
rect 3421 1955 3479 1961
rect 3421 1921 3433 1955
rect 3467 1952 3479 1955
rect 3602 1952 3608 1964
rect 3467 1924 3608 1952
rect 3467 1921 3479 1924
rect 3421 1915 3479 1921
rect 3602 1912 3608 1924
rect 3660 1912 3666 1964
rect 3694 1912 3700 1964
rect 3752 1912 3758 1964
rect 3973 1955 4031 1961
rect 3973 1921 3985 1955
rect 4019 1952 4031 1955
rect 4154 1952 4160 1964
rect 4019 1924 4160 1952
rect 4019 1921 4031 1924
rect 3973 1915 4031 1921
rect 4154 1912 4160 1924
rect 4212 1912 4218 1964
rect 4249 1955 4307 1961
rect 4249 1921 4261 1955
rect 4295 1921 4307 1955
rect 4249 1915 4307 1921
rect 3234 1844 3240 1896
rect 3292 1884 3298 1896
rect 4264 1884 4292 1915
rect 3292 1856 4292 1884
rect 4448 1884 4476 1992
rect 5092 1992 5448 2020
rect 4525 1955 4583 1961
rect 4525 1921 4537 1955
rect 4571 1952 4583 1955
rect 4706 1952 4712 1964
rect 4571 1924 4712 1952
rect 4571 1921 4583 1924
rect 4525 1915 4583 1921
rect 4706 1912 4712 1924
rect 4764 1912 4770 1964
rect 4801 1955 4859 1961
rect 4801 1921 4813 1955
rect 4847 1952 4859 1955
rect 4982 1952 4988 1964
rect 4847 1924 4988 1952
rect 4847 1921 4859 1924
rect 4801 1915 4859 1921
rect 4982 1912 4988 1924
rect 5040 1912 5046 1964
rect 5092 1961 5120 1992
rect 5442 1980 5448 1992
rect 5500 1980 5506 2032
rect 5644 2020 5672 2060
rect 5718 2048 5724 2100
rect 5776 2088 5782 2100
rect 6822 2088 6828 2100
rect 5776 2060 6828 2088
rect 5776 2048 5782 2060
rect 6822 2048 6828 2060
rect 6880 2048 6886 2100
rect 7193 2091 7251 2097
rect 7193 2057 7205 2091
rect 7239 2088 7251 2091
rect 7466 2088 7472 2100
rect 7239 2060 7472 2088
rect 7239 2057 7251 2060
rect 7193 2051 7251 2057
rect 7466 2048 7472 2060
rect 7524 2048 7530 2100
rect 7558 2048 7564 2100
rect 7616 2048 7622 2100
rect 7834 2048 7840 2100
rect 7892 2048 7898 2100
rect 8941 2091 8999 2097
rect 8941 2057 8953 2091
rect 8987 2057 8999 2091
rect 8941 2051 8999 2057
rect 5644 1992 8616 2020
rect 5077 1955 5135 1961
rect 5077 1921 5089 1955
rect 5123 1921 5135 1955
rect 5077 1915 5135 1921
rect 5353 1955 5411 1961
rect 5353 1921 5365 1955
rect 5399 1921 5411 1955
rect 5353 1915 5411 1921
rect 5629 1955 5687 1961
rect 5629 1921 5641 1955
rect 5675 1921 5687 1955
rect 5629 1915 5687 1921
rect 5721 1955 5779 1961
rect 5721 1921 5733 1955
rect 5767 1921 5779 1955
rect 5721 1915 5779 1921
rect 6181 1955 6239 1961
rect 6181 1921 6193 1955
rect 6227 1952 6239 1955
rect 6546 1952 6552 1964
rect 6227 1924 6552 1952
rect 6227 1921 6239 1924
rect 6181 1915 6239 1921
rect 5368 1884 5396 1915
rect 4448 1856 4568 1884
rect 3292 1844 3298 1856
rect 2961 1819 3019 1825
rect 2961 1785 2973 1819
rect 3007 1785 3019 1819
rect 2961 1779 3019 1785
rect 3050 1776 3056 1828
rect 3108 1816 3114 1828
rect 3789 1819 3847 1825
rect 3789 1816 3801 1819
rect 3108 1788 3801 1816
rect 3108 1776 3114 1788
rect 3789 1785 3801 1788
rect 3835 1785 3847 1819
rect 3789 1779 3847 1785
rect 4062 1776 4068 1828
rect 4120 1776 4126 1828
rect 2332 1720 2774 1748
rect 3237 1751 3295 1757
rect 3237 1717 3249 1751
rect 3283 1748 3295 1751
rect 3418 1748 3424 1760
rect 3283 1720 3424 1748
rect 3283 1717 3295 1720
rect 3237 1711 3295 1717
rect 3418 1708 3424 1720
rect 3476 1708 3482 1760
rect 3510 1708 3516 1760
rect 3568 1708 3574 1760
rect 4246 1708 4252 1760
rect 4304 1748 4310 1760
rect 4341 1751 4399 1757
rect 4341 1748 4353 1751
rect 4304 1720 4353 1748
rect 4304 1708 4310 1720
rect 4341 1717 4353 1720
rect 4387 1717 4399 1751
rect 4540 1748 4568 1856
rect 4632 1856 5396 1884
rect 4632 1825 4660 1856
rect 4617 1819 4675 1825
rect 4617 1785 4629 1819
rect 4663 1785 4675 1819
rect 4617 1779 4675 1785
rect 4893 1819 4951 1825
rect 4893 1785 4905 1819
rect 4939 1816 4951 1819
rect 5644 1816 5672 1915
rect 5736 1884 5764 1915
rect 6546 1912 6552 1924
rect 6604 1912 6610 1964
rect 6638 1912 6644 1964
rect 6696 1912 6702 1964
rect 6730 1912 6736 1964
rect 6788 1952 6794 1964
rect 6917 1955 6975 1961
rect 6917 1952 6929 1955
rect 6788 1924 6929 1952
rect 6788 1912 6794 1924
rect 6917 1921 6929 1924
rect 6963 1921 6975 1955
rect 6917 1915 6975 1921
rect 7009 1955 7067 1961
rect 7009 1921 7021 1955
rect 7055 1952 7067 1955
rect 7374 1952 7380 1964
rect 7055 1924 7380 1952
rect 7055 1921 7067 1924
rect 7009 1915 7067 1921
rect 7374 1912 7380 1924
rect 7432 1912 7438 1964
rect 7466 1912 7472 1964
rect 7524 1912 7530 1964
rect 7742 1912 7748 1964
rect 7800 1912 7806 1964
rect 8018 1912 8024 1964
rect 8076 1912 8082 1964
rect 8297 1955 8355 1961
rect 8297 1921 8309 1955
rect 8343 1952 8355 1955
rect 8478 1952 8484 1964
rect 8343 1924 8484 1952
rect 8343 1921 8355 1924
rect 8297 1915 8355 1921
rect 8478 1912 8484 1924
rect 8536 1912 8542 1964
rect 8588 1961 8616 1992
rect 8573 1955 8631 1961
rect 8573 1921 8585 1955
rect 8619 1921 8631 1955
rect 8573 1915 8631 1921
rect 8846 1912 8852 1964
rect 8904 1912 8910 1964
rect 6270 1884 6276 1896
rect 5736 1856 6276 1884
rect 6270 1844 6276 1856
rect 6328 1844 6334 1896
rect 8956 1884 8984 2051
rect 9214 2048 9220 2100
rect 9272 2048 9278 2100
rect 9493 2091 9551 2097
rect 9493 2057 9505 2091
rect 9539 2088 9551 2091
rect 10870 2088 10876 2100
rect 9539 2060 10876 2088
rect 9539 2057 9551 2060
rect 9493 2051 9551 2057
rect 10870 2048 10876 2060
rect 10928 2048 10934 2100
rect 11072 2060 13768 2088
rect 10965 2023 11023 2029
rect 10965 2020 10977 2023
rect 9232 1992 10977 2020
rect 9232 1964 9260 1992
rect 10965 1989 10977 1992
rect 11011 1989 11023 2023
rect 10965 1983 11023 1989
rect 9122 1912 9128 1964
rect 9180 1912 9186 1964
rect 9214 1912 9220 1964
rect 9272 1912 9278 1964
rect 9398 1912 9404 1964
rect 9456 1912 9462 1964
rect 9677 1955 9735 1961
rect 9677 1952 9689 1955
rect 9508 1924 9689 1952
rect 9508 1884 9536 1924
rect 9677 1921 9689 1924
rect 9723 1921 9735 1955
rect 9677 1915 9735 1921
rect 9766 1912 9772 1964
rect 9824 1952 9830 1964
rect 9953 1955 10011 1961
rect 9953 1952 9965 1955
rect 9824 1924 9965 1952
rect 9824 1912 9830 1924
rect 9953 1921 9965 1924
rect 9999 1921 10011 1955
rect 9953 1915 10011 1921
rect 10226 1912 10232 1964
rect 10284 1912 10290 1964
rect 10318 1912 10324 1964
rect 10376 1952 10382 1964
rect 10413 1955 10471 1961
rect 10413 1952 10425 1955
rect 10376 1924 10425 1952
rect 10376 1912 10382 1924
rect 10413 1921 10425 1924
rect 10459 1921 10471 1955
rect 10413 1915 10471 1921
rect 11072 1884 11100 2060
rect 11422 1980 11428 2032
rect 11480 2020 11486 2032
rect 11977 2023 12035 2029
rect 11977 2020 11989 2023
rect 11480 1992 11989 2020
rect 11480 1980 11486 1992
rect 11977 1989 11989 1992
rect 12023 1989 12035 2023
rect 11977 1983 12035 1989
rect 12710 1980 12716 2032
rect 12768 2020 12774 2032
rect 12768 1992 13492 2020
rect 12768 1980 12774 1992
rect 11330 1912 11336 1964
rect 11388 1952 11394 1964
rect 11517 1955 11575 1961
rect 11517 1952 11529 1955
rect 11388 1924 11529 1952
rect 11388 1912 11394 1924
rect 11517 1921 11529 1924
rect 11563 1921 11575 1955
rect 11517 1915 11575 1921
rect 11606 1912 11612 1964
rect 11664 1912 11670 1964
rect 12342 1912 12348 1964
rect 12400 1952 12406 1964
rect 12621 1955 12679 1961
rect 12621 1952 12633 1955
rect 12400 1924 12633 1952
rect 12400 1912 12406 1924
rect 12621 1921 12633 1924
rect 12667 1921 12679 1955
rect 12621 1915 12679 1921
rect 12802 1912 12808 1964
rect 12860 1912 12866 1964
rect 13464 1961 13492 1992
rect 13740 1961 13768 2060
rect 13998 2048 14004 2100
rect 14056 2048 14062 2100
rect 14182 2048 14188 2100
rect 14240 2048 14246 2100
rect 17405 2091 17463 2097
rect 14936 2060 15976 2088
rect 14016 2020 14044 2048
rect 14016 1992 14872 2020
rect 13449 1955 13507 1961
rect 13449 1921 13461 1955
rect 13495 1921 13507 1955
rect 13449 1915 13507 1921
rect 13725 1955 13783 1961
rect 13725 1921 13737 1955
rect 13771 1921 13783 1955
rect 13725 1915 13783 1921
rect 14090 1912 14096 1964
rect 14148 1912 14154 1964
rect 14366 1912 14372 1964
rect 14424 1912 14430 1964
rect 14844 1961 14872 1992
rect 14461 1955 14519 1961
rect 14461 1921 14473 1955
rect 14507 1921 14519 1955
rect 14461 1915 14519 1921
rect 14829 1955 14887 1961
rect 14829 1921 14841 1955
rect 14875 1921 14887 1955
rect 14829 1915 14887 1921
rect 8956 1856 9536 1884
rect 9600 1856 11100 1884
rect 11624 1884 11652 1912
rect 14476 1884 14504 1915
rect 14936 1884 14964 2060
rect 15470 1980 15476 2032
rect 15528 2020 15534 2032
rect 15841 2023 15899 2029
rect 15841 2020 15853 2023
rect 15528 1992 15853 2020
rect 15528 1980 15534 1992
rect 15841 1989 15853 1992
rect 15887 1989 15899 2023
rect 15841 1983 15899 1989
rect 15378 1912 15384 1964
rect 15436 1912 15442 1964
rect 15657 1955 15715 1961
rect 15657 1921 15669 1955
rect 15703 1952 15715 1955
rect 15948 1952 15976 2060
rect 17405 2057 17417 2091
rect 17451 2088 17463 2091
rect 17586 2088 17592 2100
rect 17451 2060 17592 2088
rect 17451 2057 17463 2060
rect 17405 2051 17463 2057
rect 17586 2048 17592 2060
rect 17644 2048 17650 2100
rect 17681 2091 17739 2097
rect 17681 2057 17693 2091
rect 17727 2088 17739 2091
rect 17862 2088 17868 2100
rect 17727 2060 17868 2088
rect 17727 2057 17739 2060
rect 17681 2051 17739 2057
rect 17862 2048 17868 2060
rect 17920 2048 17926 2100
rect 17954 2048 17960 2100
rect 18012 2088 18018 2100
rect 18012 2060 18184 2088
rect 18012 2048 18018 2060
rect 16022 1980 16028 2032
rect 16080 2020 16086 2032
rect 16080 1992 17632 2020
rect 16080 1980 16086 1992
rect 15703 1924 15976 1952
rect 15703 1921 15715 1924
rect 15657 1915 15715 1921
rect 16114 1912 16120 1964
rect 16172 1952 16178 1964
rect 17604 1961 17632 1992
rect 17770 1980 17776 2032
rect 17828 2020 17834 2032
rect 18049 2023 18107 2029
rect 18049 2020 18061 2023
rect 17828 1992 18061 2020
rect 17828 1980 17834 1992
rect 18049 1989 18061 1992
rect 18095 1989 18107 2023
rect 18049 1983 18107 1989
rect 16485 1955 16543 1961
rect 16485 1952 16497 1955
rect 16172 1924 16497 1952
rect 16172 1912 16178 1924
rect 16485 1921 16497 1924
rect 16531 1921 16543 1955
rect 16485 1915 16543 1921
rect 16945 1955 17003 1961
rect 16945 1921 16957 1955
rect 16991 1921 17003 1955
rect 16945 1915 17003 1921
rect 17589 1955 17647 1961
rect 17589 1921 17601 1955
rect 17635 1921 17647 1955
rect 17589 1915 17647 1921
rect 17865 1955 17923 1961
rect 17865 1921 17877 1955
rect 17911 1921 17923 1955
rect 18156 1952 18184 2060
rect 18230 2048 18236 2100
rect 18288 2088 18294 2100
rect 18288 2060 18644 2088
rect 18288 2048 18294 2060
rect 18616 2029 18644 2060
rect 19150 2048 19156 2100
rect 19208 2048 19214 2100
rect 19242 2048 19248 2100
rect 19300 2088 19306 2100
rect 19300 2060 20300 2088
rect 19300 2048 19306 2060
rect 18601 2023 18659 2029
rect 18601 1989 18613 2023
rect 18647 1989 18659 2023
rect 19168 2020 19196 2048
rect 20272 2029 20300 2060
rect 20346 2048 20352 2100
rect 20404 2048 20410 2100
rect 20622 2048 20628 2100
rect 20680 2088 20686 2100
rect 20680 2060 20852 2088
rect 20680 2048 20686 2060
rect 19705 2023 19763 2029
rect 19705 2020 19717 2023
rect 19168 1992 19717 2020
rect 18601 1983 18659 1989
rect 19705 1989 19717 1992
rect 19751 1989 19763 2023
rect 19705 1983 19763 1989
rect 20257 2023 20315 2029
rect 20257 1989 20269 2023
rect 20303 1989 20315 2023
rect 20257 1983 20315 1989
rect 19153 1955 19211 1961
rect 19153 1952 19165 1955
rect 18156 1924 19165 1952
rect 17865 1915 17923 1921
rect 19153 1921 19165 1924
rect 19199 1921 19211 1955
rect 19153 1915 19211 1921
rect 16960 1884 16988 1915
rect 17880 1884 17908 1915
rect 19334 1912 19340 1964
rect 19392 1912 19398 1964
rect 20364 1952 20392 2048
rect 20824 2029 20852 2060
rect 20898 2048 20904 2100
rect 20956 2048 20962 2100
rect 20990 2048 20996 2100
rect 21048 2088 21054 2100
rect 21269 2091 21327 2097
rect 21269 2088 21281 2091
rect 21048 2060 21281 2088
rect 21048 2048 21054 2060
rect 21269 2057 21281 2060
rect 21315 2057 21327 2091
rect 21269 2051 21327 2057
rect 21450 2048 21456 2100
rect 21508 2048 21514 2100
rect 21634 2048 21640 2100
rect 21692 2088 21698 2100
rect 21821 2091 21879 2097
rect 21821 2088 21833 2091
rect 21692 2060 21833 2088
rect 21692 2048 21698 2060
rect 21821 2057 21833 2060
rect 21867 2057 21879 2091
rect 21821 2051 21879 2057
rect 22278 2048 22284 2100
rect 22336 2048 22342 2100
rect 22646 2048 22652 2100
rect 22704 2048 22710 2100
rect 22741 2091 22799 2097
rect 22741 2057 22753 2091
rect 22787 2088 22799 2091
rect 23106 2088 23112 2100
rect 22787 2060 23112 2088
rect 22787 2057 22799 2060
rect 22741 2051 22799 2057
rect 23106 2048 23112 2060
rect 23164 2048 23170 2100
rect 23198 2048 23204 2100
rect 23256 2048 23262 2100
rect 23934 2088 23940 2100
rect 23308 2060 23940 2088
rect 20809 2023 20867 2029
rect 20809 1989 20821 2023
rect 20855 1989 20867 2023
rect 22664 2020 22692 2048
rect 23308 2020 23336 2060
rect 23934 2048 23940 2060
rect 23992 2048 23998 2100
rect 24026 2048 24032 2100
rect 24084 2048 24090 2100
rect 22664 1992 22968 2020
rect 20809 1983 20867 1989
rect 21085 1955 21143 1961
rect 21085 1952 21097 1955
rect 20364 1924 21097 1952
rect 21085 1921 21097 1924
rect 21131 1921 21143 1955
rect 21085 1915 21143 1921
rect 21637 1955 21695 1961
rect 21637 1921 21649 1955
rect 21683 1921 21695 1955
rect 21637 1915 21695 1921
rect 11624 1856 14504 1884
rect 14568 1856 14964 1884
rect 15212 1856 16988 1884
rect 17052 1856 17908 1884
rect 19352 1884 19380 1912
rect 19352 1856 20392 1884
rect 4939 1788 5672 1816
rect 4939 1785 4951 1788
rect 4893 1779 4951 1785
rect 5902 1776 5908 1828
rect 5960 1776 5966 1828
rect 6362 1776 6368 1828
rect 6420 1816 6426 1828
rect 6420 1788 6776 1816
rect 6420 1776 6426 1788
rect 5074 1748 5080 1760
rect 4540 1720 5080 1748
rect 4341 1711 4399 1717
rect 5074 1708 5080 1720
rect 5132 1708 5138 1760
rect 5166 1708 5172 1760
rect 5224 1708 5230 1760
rect 5445 1751 5503 1757
rect 5445 1717 5457 1751
rect 5491 1748 5503 1751
rect 5534 1748 5540 1760
rect 5491 1720 5540 1748
rect 5491 1717 5503 1720
rect 5445 1711 5503 1717
rect 5534 1708 5540 1720
rect 5592 1708 5598 1760
rect 5994 1708 6000 1760
rect 6052 1708 6058 1760
rect 6454 1708 6460 1760
rect 6512 1708 6518 1760
rect 6748 1757 6776 1788
rect 7834 1776 7840 1828
rect 7892 1816 7898 1828
rect 7892 1788 8800 1816
rect 7892 1776 7898 1788
rect 6733 1751 6791 1757
rect 6733 1717 6745 1751
rect 6779 1717 6791 1751
rect 6733 1711 6791 1717
rect 7285 1751 7343 1757
rect 7285 1717 7297 1751
rect 7331 1748 7343 1751
rect 7466 1748 7472 1760
rect 7331 1720 7472 1748
rect 7331 1717 7343 1720
rect 7285 1711 7343 1717
rect 7466 1708 7472 1720
rect 7524 1708 7530 1760
rect 8018 1708 8024 1760
rect 8076 1748 8082 1760
rect 8113 1751 8171 1757
rect 8113 1748 8125 1751
rect 8076 1720 8125 1748
rect 8076 1708 8082 1720
rect 8113 1717 8125 1720
rect 8159 1717 8171 1751
rect 8113 1711 8171 1717
rect 8202 1708 8208 1760
rect 8260 1748 8266 1760
rect 8389 1751 8447 1757
rect 8389 1748 8401 1751
rect 8260 1720 8401 1748
rect 8260 1708 8266 1720
rect 8389 1717 8401 1720
rect 8435 1717 8447 1751
rect 8389 1711 8447 1717
rect 8662 1708 8668 1760
rect 8720 1708 8726 1760
rect 8772 1748 8800 1788
rect 8938 1776 8944 1828
rect 8996 1816 9002 1828
rect 9490 1816 9496 1828
rect 8996 1788 9496 1816
rect 8996 1776 9002 1788
rect 9490 1776 9496 1788
rect 9548 1776 9554 1828
rect 9600 1748 9628 1856
rect 10045 1819 10103 1825
rect 10045 1785 10057 1819
rect 10091 1816 10103 1819
rect 10134 1816 10140 1828
rect 10091 1788 10140 1816
rect 10091 1785 10103 1788
rect 10045 1779 10103 1785
rect 10134 1776 10140 1788
rect 10192 1776 10198 1828
rect 13170 1816 13176 1828
rect 10428 1788 13176 1816
rect 8772 1720 9628 1748
rect 9769 1751 9827 1757
rect 9769 1717 9781 1751
rect 9815 1748 9827 1751
rect 10428 1748 10456 1788
rect 13170 1776 13176 1788
rect 13228 1776 13234 1828
rect 13265 1819 13323 1825
rect 13265 1785 13277 1819
rect 13311 1816 13323 1819
rect 14366 1816 14372 1828
rect 13311 1788 14372 1816
rect 13311 1785 13323 1788
rect 13265 1779 13323 1785
rect 14366 1776 14372 1788
rect 14424 1776 14430 1828
rect 9815 1720 10456 1748
rect 9815 1717 9827 1720
rect 9769 1711 9827 1717
rect 10502 1708 10508 1760
rect 10560 1708 10566 1760
rect 11054 1708 11060 1760
rect 11112 1708 11118 1760
rect 11698 1708 11704 1760
rect 11756 1708 11762 1760
rect 11790 1708 11796 1760
rect 11848 1748 11854 1760
rect 12069 1751 12127 1757
rect 12069 1748 12081 1751
rect 11848 1720 12081 1748
rect 11848 1708 11854 1720
rect 12069 1717 12081 1720
rect 12115 1717 12127 1751
rect 12069 1711 12127 1717
rect 12434 1708 12440 1760
rect 12492 1708 12498 1760
rect 12618 1708 12624 1760
rect 12676 1748 12682 1760
rect 12897 1751 12955 1757
rect 12897 1748 12909 1751
rect 12676 1720 12909 1748
rect 12676 1708 12682 1720
rect 12897 1717 12909 1720
rect 12943 1717 12955 1751
rect 12897 1711 12955 1717
rect 13538 1708 13544 1760
rect 13596 1708 13602 1760
rect 13909 1751 13967 1757
rect 13909 1717 13921 1751
rect 13955 1748 13967 1751
rect 14568 1748 14596 1856
rect 15212 1825 15240 1856
rect 15197 1819 15255 1825
rect 15197 1785 15209 1819
rect 15243 1785 15255 1819
rect 17052 1816 17080 1856
rect 15197 1779 15255 1785
rect 15304 1788 17080 1816
rect 13955 1720 14596 1748
rect 13955 1717 13967 1720
rect 13909 1711 13967 1717
rect 14642 1708 14648 1760
rect 14700 1708 14706 1760
rect 14734 1708 14740 1760
rect 14792 1748 14798 1760
rect 15013 1751 15071 1757
rect 15013 1748 15025 1751
rect 14792 1720 15025 1748
rect 14792 1708 14798 1720
rect 15013 1717 15025 1720
rect 15059 1717 15071 1751
rect 15013 1711 15071 1717
rect 15102 1708 15108 1760
rect 15160 1748 15166 1760
rect 15304 1748 15332 1788
rect 17770 1776 17776 1828
rect 17828 1816 17834 1828
rect 19429 1819 19487 1825
rect 19429 1816 19441 1819
rect 17828 1788 19441 1816
rect 17828 1776 17834 1788
rect 19429 1785 19441 1788
rect 19475 1785 19487 1819
rect 19429 1779 19487 1785
rect 19518 1776 19524 1828
rect 19576 1816 19582 1828
rect 20364 1816 20392 1856
rect 20438 1844 20444 1896
rect 20496 1884 20502 1896
rect 21652 1884 21680 1915
rect 21726 1912 21732 1964
rect 21784 1952 21790 1964
rect 22005 1955 22063 1961
rect 22005 1952 22017 1955
rect 21784 1924 22017 1952
rect 21784 1912 21790 1924
rect 22005 1921 22017 1924
rect 22051 1921 22063 1955
rect 22005 1915 22063 1921
rect 22094 1912 22100 1964
rect 22152 1912 22158 1964
rect 22940 1961 22968 1992
rect 23216 1992 23336 2020
rect 22649 1955 22707 1961
rect 22649 1921 22661 1955
rect 22695 1921 22707 1955
rect 22649 1915 22707 1921
rect 22925 1955 22983 1961
rect 22925 1921 22937 1955
rect 22971 1921 22983 1955
rect 22925 1915 22983 1921
rect 20496 1856 21680 1884
rect 22664 1884 22692 1915
rect 23014 1912 23020 1964
rect 23072 1912 23078 1964
rect 23216 1884 23244 1992
rect 23382 1980 23388 2032
rect 23440 2020 23446 2032
rect 23440 1992 23980 2020
rect 23440 1980 23446 1992
rect 23569 1955 23627 1961
rect 23569 1952 23581 1955
rect 22664 1856 23244 1884
rect 23308 1924 23581 1952
rect 20496 1844 20502 1856
rect 21450 1816 21456 1828
rect 19576 1788 19932 1816
rect 20364 1788 21456 1816
rect 19576 1776 19582 1788
rect 15160 1720 15332 1748
rect 15160 1708 15166 1720
rect 15470 1708 15476 1760
rect 15528 1708 15534 1760
rect 15654 1708 15660 1760
rect 15712 1748 15718 1760
rect 15933 1751 15991 1757
rect 15933 1748 15945 1751
rect 15712 1720 15945 1748
rect 15712 1708 15718 1720
rect 15933 1717 15945 1720
rect 15979 1717 15991 1751
rect 15933 1711 15991 1717
rect 16301 1751 16359 1757
rect 16301 1717 16313 1751
rect 16347 1748 16359 1751
rect 16574 1748 16580 1760
rect 16347 1720 16580 1748
rect 16347 1717 16359 1720
rect 16301 1711 16359 1717
rect 16574 1708 16580 1720
rect 16632 1708 16638 1760
rect 16758 1708 16764 1760
rect 16816 1748 16822 1760
rect 17037 1751 17095 1757
rect 17037 1748 17049 1751
rect 16816 1720 17049 1748
rect 16816 1708 16822 1720
rect 17037 1717 17049 1720
rect 17083 1717 17095 1751
rect 17037 1711 17095 1717
rect 17954 1708 17960 1760
rect 18012 1748 18018 1760
rect 18141 1751 18199 1757
rect 18141 1748 18153 1751
rect 18012 1720 18153 1748
rect 18012 1708 18018 1720
rect 18141 1717 18153 1720
rect 18187 1717 18199 1751
rect 18141 1711 18199 1717
rect 18230 1708 18236 1760
rect 18288 1748 18294 1760
rect 18693 1751 18751 1757
rect 18693 1748 18705 1751
rect 18288 1720 18705 1748
rect 18288 1708 18294 1720
rect 18693 1717 18705 1720
rect 18739 1717 18751 1751
rect 18693 1711 18751 1717
rect 19334 1708 19340 1760
rect 19392 1748 19398 1760
rect 19797 1751 19855 1757
rect 19797 1748 19809 1751
rect 19392 1720 19809 1748
rect 19392 1708 19398 1720
rect 19797 1717 19809 1720
rect 19843 1717 19855 1751
rect 19904 1748 19932 1788
rect 21450 1776 21456 1788
rect 21508 1776 21514 1828
rect 22465 1819 22523 1825
rect 22465 1785 22477 1819
rect 22511 1816 22523 1819
rect 23308 1816 23336 1924
rect 23569 1921 23581 1924
rect 23615 1921 23627 1955
rect 23569 1915 23627 1921
rect 23845 1955 23903 1961
rect 23845 1921 23857 1955
rect 23891 1921 23903 1955
rect 23845 1915 23903 1921
rect 23860 1884 23888 1915
rect 23400 1856 23888 1884
rect 23952 1884 23980 1992
rect 24044 1952 24072 2048
rect 24121 1955 24179 1961
rect 24121 1952 24133 1955
rect 24044 1924 24133 1952
rect 24121 1921 24133 1924
rect 24167 1921 24179 1955
rect 24121 1915 24179 1921
rect 24213 1955 24271 1961
rect 24213 1921 24225 1955
rect 24259 1921 24271 1955
rect 24213 1915 24271 1921
rect 24228 1884 24256 1915
rect 23952 1856 24256 1884
rect 23400 1825 23428 1856
rect 22511 1788 23336 1816
rect 23385 1819 23443 1825
rect 22511 1785 22523 1788
rect 22465 1779 22523 1785
rect 23385 1785 23397 1819
rect 23431 1785 23443 1819
rect 23385 1779 23443 1785
rect 23937 1819 23995 1825
rect 23937 1785 23949 1819
rect 23983 1816 23995 1819
rect 24210 1816 24216 1828
rect 23983 1788 24216 1816
rect 23983 1785 23995 1788
rect 23937 1779 23995 1785
rect 24210 1776 24216 1788
rect 24268 1776 24274 1828
rect 20349 1751 20407 1757
rect 20349 1748 20361 1751
rect 19904 1720 20361 1748
rect 19797 1711 19855 1717
rect 20349 1717 20361 1720
rect 20395 1717 20407 1751
rect 20349 1711 20407 1717
rect 22370 1708 22376 1760
rect 22428 1748 22434 1760
rect 23014 1748 23020 1760
rect 22428 1720 23020 1748
rect 22428 1708 22434 1720
rect 23014 1708 23020 1720
rect 23072 1708 23078 1760
rect 23661 1751 23719 1757
rect 23661 1717 23673 1751
rect 23707 1748 23719 1751
rect 24118 1748 24124 1760
rect 23707 1720 24124 1748
rect 23707 1717 23719 1720
rect 23661 1711 23719 1717
rect 24118 1708 24124 1720
rect 24176 1708 24182 1760
rect 24397 1751 24455 1757
rect 24397 1717 24409 1751
rect 24443 1748 24455 1751
rect 24443 1720 24900 1748
rect 24443 1717 24455 1720
rect 24397 1711 24455 1717
rect 1104 1658 24840 1680
rect 1104 1606 3917 1658
rect 3969 1606 3981 1658
rect 4033 1606 4045 1658
rect 4097 1606 4109 1658
rect 4161 1606 4173 1658
rect 4225 1606 9851 1658
rect 9903 1606 9915 1658
rect 9967 1606 9979 1658
rect 10031 1606 10043 1658
rect 10095 1606 10107 1658
rect 10159 1606 15785 1658
rect 15837 1606 15849 1658
rect 15901 1606 15913 1658
rect 15965 1606 15977 1658
rect 16029 1606 16041 1658
rect 16093 1606 21719 1658
rect 21771 1606 21783 1658
rect 21835 1606 21847 1658
rect 21899 1606 21911 1658
rect 21963 1606 21975 1658
rect 22027 1606 24840 1658
rect 1104 1584 24840 1606
rect 2590 1504 2596 1556
rect 2648 1504 2654 1556
rect 2869 1547 2927 1553
rect 2869 1513 2881 1547
rect 2915 1544 2927 1547
rect 3234 1544 3240 1556
rect 2915 1516 3240 1544
rect 2915 1513 2927 1516
rect 2869 1507 2927 1513
rect 3234 1504 3240 1516
rect 3292 1504 3298 1556
rect 4430 1544 4436 1556
rect 3344 1516 4436 1544
rect 1489 1479 1547 1485
rect 1489 1445 1501 1479
rect 1535 1476 1547 1479
rect 2958 1476 2964 1488
rect 1535 1448 2964 1476
rect 1535 1445 1547 1448
rect 1489 1439 1547 1445
rect 2958 1436 2964 1448
rect 3016 1436 3022 1488
rect 3234 1408 3240 1420
rect 2700 1380 3240 1408
rect 1486 1300 1492 1352
rect 1544 1340 1550 1352
rect 1673 1343 1731 1349
rect 1673 1340 1685 1343
rect 1544 1312 1685 1340
rect 1544 1300 1550 1312
rect 1673 1309 1685 1312
rect 1719 1309 1731 1343
rect 1673 1303 1731 1309
rect 1765 1343 1823 1349
rect 1765 1309 1777 1343
rect 1811 1309 1823 1343
rect 1765 1303 1823 1309
rect 2225 1343 2283 1349
rect 2225 1309 2237 1343
rect 2271 1309 2283 1343
rect 2225 1303 2283 1309
rect 2501 1343 2559 1349
rect 2501 1309 2513 1343
rect 2547 1340 2559 1343
rect 2700 1340 2728 1380
rect 3234 1368 3240 1380
rect 3292 1368 3298 1420
rect 2547 1312 2728 1340
rect 2547 1309 2559 1312
rect 2501 1303 2559 1309
rect 1780 1272 1808 1303
rect 2240 1272 2268 1303
rect 2774 1300 2780 1352
rect 2832 1300 2838 1352
rect 3050 1300 3056 1352
rect 3108 1300 3114 1352
rect 3344 1349 3372 1516
rect 4430 1504 4436 1516
rect 4488 1504 4494 1556
rect 5994 1504 6000 1556
rect 6052 1504 6058 1556
rect 6641 1547 6699 1553
rect 6641 1513 6653 1547
rect 6687 1544 6699 1547
rect 6687 1516 7144 1544
rect 6687 1513 6699 1516
rect 6641 1507 6699 1513
rect 3421 1479 3479 1485
rect 3421 1445 3433 1479
rect 3467 1476 3479 1479
rect 3467 1448 4384 1476
rect 3467 1445 3479 1448
rect 3421 1439 3479 1445
rect 3510 1368 3516 1420
rect 3568 1408 3574 1420
rect 3568 1380 4108 1408
rect 3568 1368 3574 1380
rect 3329 1343 3387 1349
rect 3329 1309 3341 1343
rect 3375 1309 3387 1343
rect 3329 1303 3387 1309
rect 3605 1343 3663 1349
rect 3605 1309 3617 1343
rect 3651 1340 3663 1343
rect 3878 1340 3884 1352
rect 3651 1312 3884 1340
rect 3651 1309 3663 1312
rect 3605 1303 3663 1309
rect 3878 1300 3884 1312
rect 3936 1300 3942 1352
rect 3973 1343 4031 1349
rect 3973 1309 3985 1343
rect 4019 1309 4031 1343
rect 4080 1340 4108 1380
rect 4249 1343 4307 1349
rect 4249 1340 4261 1343
rect 4080 1312 4261 1340
rect 3973 1303 4031 1309
rect 4249 1309 4261 1312
rect 4295 1309 4307 1343
rect 4356 1340 4384 1448
rect 6012 1408 6040 1504
rect 6362 1436 6368 1488
rect 6420 1436 6426 1488
rect 5736 1380 6040 1408
rect 6380 1408 6408 1436
rect 7116 1408 7144 1516
rect 7466 1504 7472 1556
rect 7524 1544 7530 1556
rect 7524 1516 9904 1544
rect 7524 1504 7530 1516
rect 7193 1479 7251 1485
rect 7193 1445 7205 1479
rect 7239 1476 7251 1479
rect 9214 1476 9220 1488
rect 7239 1448 9220 1476
rect 7239 1445 7251 1448
rect 7193 1439 7251 1445
rect 9214 1436 9220 1448
rect 9272 1436 9278 1488
rect 9876 1476 9904 1516
rect 9950 1504 9956 1556
rect 10008 1544 10014 1556
rect 11422 1544 11428 1556
rect 10008 1516 11428 1544
rect 10008 1504 10014 1516
rect 11422 1504 11428 1516
rect 11480 1504 11486 1556
rect 11517 1547 11575 1553
rect 11517 1513 11529 1547
rect 11563 1544 11575 1547
rect 12158 1544 12164 1556
rect 11563 1516 12164 1544
rect 11563 1513 11575 1516
rect 11517 1507 11575 1513
rect 12158 1504 12164 1516
rect 12216 1504 12222 1556
rect 12434 1504 12440 1556
rect 12492 1544 12498 1556
rect 13170 1544 13176 1556
rect 12492 1516 13176 1544
rect 12492 1504 12498 1516
rect 13170 1504 13176 1516
rect 13228 1504 13234 1556
rect 13814 1504 13820 1556
rect 13872 1544 13878 1556
rect 14277 1547 14335 1553
rect 14277 1544 14289 1547
rect 13872 1516 14289 1544
rect 13872 1504 13878 1516
rect 14277 1513 14289 1516
rect 14323 1513 14335 1547
rect 14277 1507 14335 1513
rect 15102 1504 15108 1556
rect 15160 1504 15166 1556
rect 15378 1504 15384 1556
rect 15436 1504 15442 1556
rect 15933 1547 15991 1553
rect 15933 1513 15945 1547
rect 15979 1513 15991 1547
rect 15933 1507 15991 1513
rect 15120 1476 15148 1504
rect 9876 1448 15148 1476
rect 15286 1436 15292 1488
rect 15344 1476 15350 1488
rect 15948 1476 15976 1507
rect 16114 1504 16120 1556
rect 16172 1504 16178 1556
rect 16206 1504 16212 1556
rect 16264 1504 16270 1556
rect 16301 1547 16359 1553
rect 16301 1513 16313 1547
rect 16347 1544 16359 1547
rect 16482 1544 16488 1556
rect 16347 1516 16488 1544
rect 16347 1513 16359 1516
rect 16301 1507 16359 1513
rect 16482 1504 16488 1516
rect 16540 1504 16546 1556
rect 16853 1547 16911 1553
rect 16853 1513 16865 1547
rect 16899 1513 16911 1547
rect 16853 1507 16911 1513
rect 17405 1547 17463 1553
rect 17405 1513 17417 1547
rect 17451 1513 17463 1547
rect 17405 1507 17463 1513
rect 15344 1448 15976 1476
rect 15344 1436 15350 1448
rect 8570 1408 8576 1420
rect 6380 1380 6592 1408
rect 7116 1380 7236 1408
rect 4525 1343 4583 1349
rect 4525 1340 4537 1343
rect 4356 1312 4537 1340
rect 4249 1303 4307 1309
rect 4525 1309 4537 1312
rect 4571 1309 4583 1343
rect 4525 1303 4583 1309
rect 4617 1343 4675 1349
rect 4617 1309 4629 1343
rect 4663 1340 4675 1343
rect 4798 1340 4804 1352
rect 4663 1312 4804 1340
rect 4663 1309 4675 1312
rect 4617 1303 4675 1309
rect 2682 1272 2688 1284
rect 1780 1244 2176 1272
rect 2240 1244 2688 1272
rect 1946 1164 1952 1216
rect 2004 1164 2010 1216
rect 2038 1164 2044 1216
rect 2096 1164 2102 1216
rect 2148 1204 2176 1244
rect 2682 1232 2688 1244
rect 2740 1232 2746 1284
rect 3988 1272 4016 1303
rect 4798 1300 4804 1312
rect 4856 1300 4862 1352
rect 4893 1343 4951 1349
rect 4893 1309 4905 1343
rect 4939 1309 4951 1343
rect 4893 1303 4951 1309
rect 4908 1272 4936 1303
rect 5166 1300 5172 1352
rect 5224 1340 5230 1352
rect 5353 1343 5411 1349
rect 5353 1340 5365 1343
rect 5224 1312 5365 1340
rect 5224 1300 5230 1312
rect 5353 1309 5365 1312
rect 5399 1309 5411 1343
rect 5353 1303 5411 1309
rect 5534 1300 5540 1352
rect 5592 1340 5598 1352
rect 5736 1349 5764 1380
rect 5629 1343 5687 1349
rect 5629 1340 5641 1343
rect 5592 1312 5641 1340
rect 5592 1300 5598 1312
rect 5629 1309 5641 1312
rect 5675 1309 5687 1343
rect 5629 1303 5687 1309
rect 5721 1343 5779 1349
rect 5721 1309 5733 1343
rect 5767 1309 5779 1343
rect 5721 1303 5779 1309
rect 5997 1343 6055 1349
rect 5997 1309 6009 1343
rect 6043 1340 6055 1343
rect 6454 1340 6460 1352
rect 6043 1312 6460 1340
rect 6043 1309 6055 1312
rect 5997 1303 6055 1309
rect 6454 1300 6460 1312
rect 6512 1300 6518 1352
rect 6564 1349 6592 1380
rect 6549 1343 6607 1349
rect 6549 1309 6561 1343
rect 6595 1309 6607 1343
rect 6549 1303 6607 1309
rect 6822 1300 6828 1352
rect 6880 1300 6886 1352
rect 7101 1343 7159 1349
rect 7101 1340 7113 1343
rect 6932 1312 7113 1340
rect 3160 1244 4016 1272
rect 4080 1244 4936 1272
rect 2222 1204 2228 1216
rect 2148 1176 2228 1204
rect 2222 1164 2228 1176
rect 2280 1164 2286 1216
rect 2314 1164 2320 1216
rect 2372 1164 2378 1216
rect 3160 1213 3188 1244
rect 3145 1207 3203 1213
rect 3145 1173 3157 1207
rect 3191 1173 3203 1207
rect 3145 1167 3203 1173
rect 3789 1207 3847 1213
rect 3789 1173 3801 1207
rect 3835 1204 3847 1207
rect 3970 1204 3976 1216
rect 3835 1176 3976 1204
rect 3835 1173 3847 1176
rect 3789 1167 3847 1173
rect 3970 1164 3976 1176
rect 4028 1164 4034 1216
rect 4080 1213 4108 1244
rect 5258 1232 5264 1284
rect 5316 1272 5322 1284
rect 6932 1272 6960 1312
rect 7101 1309 7113 1312
rect 7147 1309 7159 1343
rect 7208 1340 7236 1380
rect 8128 1380 8576 1408
rect 7377 1343 7435 1349
rect 7377 1340 7389 1343
rect 7208 1312 7389 1340
rect 7101 1303 7159 1309
rect 7377 1309 7389 1312
rect 7423 1309 7435 1343
rect 7377 1303 7435 1309
rect 7653 1343 7711 1349
rect 7653 1309 7665 1343
rect 7699 1309 7711 1343
rect 7653 1303 7711 1309
rect 7668 1272 7696 1303
rect 7834 1300 7840 1352
rect 7892 1300 7898 1352
rect 7929 1343 7987 1349
rect 7929 1309 7941 1343
rect 7975 1340 7987 1343
rect 8128 1340 8156 1380
rect 8570 1368 8576 1380
rect 8628 1368 8634 1420
rect 9416 1380 10456 1408
rect 7975 1312 8156 1340
rect 7975 1309 7987 1312
rect 7929 1303 7987 1309
rect 8202 1300 8208 1352
rect 8260 1300 8266 1352
rect 8481 1343 8539 1349
rect 8481 1309 8493 1343
rect 8527 1340 8539 1343
rect 8662 1340 8668 1352
rect 8527 1312 8668 1340
rect 8527 1309 8539 1312
rect 8481 1303 8539 1309
rect 8662 1300 8668 1312
rect 8720 1300 8726 1352
rect 8754 1300 8760 1352
rect 8812 1300 8818 1352
rect 8938 1300 8944 1352
rect 8996 1340 9002 1352
rect 9033 1343 9091 1349
rect 9033 1340 9045 1343
rect 8996 1312 9045 1340
rect 8996 1300 9002 1312
rect 9033 1309 9045 1312
rect 9079 1309 9091 1343
rect 9033 1303 9091 1309
rect 9416 1336 9444 1380
rect 9493 1343 9551 1349
rect 9493 1336 9505 1343
rect 9416 1309 9505 1336
rect 9539 1309 9551 1343
rect 9416 1308 9551 1309
rect 9493 1303 9551 1308
rect 9585 1343 9643 1349
rect 9585 1309 9597 1343
rect 9631 1309 9643 1343
rect 9585 1303 9643 1309
rect 5316 1244 6500 1272
rect 5316 1232 5322 1244
rect 4065 1207 4123 1213
rect 4065 1173 4077 1207
rect 4111 1173 4123 1207
rect 4065 1167 4123 1173
rect 4341 1207 4399 1213
rect 4341 1173 4353 1207
rect 4387 1204 4399 1207
rect 4522 1204 4528 1216
rect 4387 1176 4528 1204
rect 4387 1173 4399 1176
rect 4341 1167 4399 1173
rect 4522 1164 4528 1176
rect 4580 1164 4586 1216
rect 4706 1164 4712 1216
rect 4764 1204 4770 1216
rect 4801 1207 4859 1213
rect 4801 1204 4813 1207
rect 4764 1176 4813 1204
rect 4764 1164 4770 1176
rect 4801 1173 4813 1176
rect 4847 1173 4859 1207
rect 4801 1167 4859 1173
rect 5074 1164 5080 1216
rect 5132 1164 5138 1216
rect 5166 1164 5172 1216
rect 5224 1164 5230 1216
rect 5445 1207 5503 1213
rect 5445 1173 5457 1207
rect 5491 1204 5503 1207
rect 5810 1204 5816 1216
rect 5491 1176 5816 1204
rect 5491 1173 5503 1176
rect 5445 1167 5503 1173
rect 5810 1164 5816 1176
rect 5868 1164 5874 1216
rect 5902 1164 5908 1216
rect 5960 1164 5966 1216
rect 6178 1164 6184 1216
rect 6236 1164 6242 1216
rect 6362 1164 6368 1216
rect 6420 1164 6426 1216
rect 6472 1204 6500 1244
rect 6840 1244 6960 1272
rect 7392 1244 7696 1272
rect 6840 1204 6868 1244
rect 6472 1176 6868 1204
rect 6917 1207 6975 1213
rect 6917 1173 6929 1207
rect 6963 1204 6975 1207
rect 7392 1204 7420 1244
rect 6963 1176 7420 1204
rect 6963 1173 6975 1176
rect 6917 1167 6975 1173
rect 7466 1164 7472 1216
rect 7524 1164 7530 1216
rect 7745 1207 7803 1213
rect 7745 1173 7757 1207
rect 7791 1204 7803 1207
rect 7852 1204 7880 1300
rect 9600 1272 9628 1303
rect 9950 1300 9956 1352
rect 10008 1300 10014 1352
rect 10134 1300 10140 1352
rect 10192 1340 10198 1352
rect 10321 1343 10379 1349
rect 10321 1340 10333 1343
rect 10192 1312 10333 1340
rect 10192 1300 10198 1312
rect 10321 1309 10333 1312
rect 10367 1309 10379 1343
rect 10428 1340 10456 1380
rect 10502 1368 10508 1420
rect 10560 1408 10566 1420
rect 10686 1408 10692 1420
rect 10560 1380 10692 1408
rect 10560 1368 10566 1380
rect 10686 1368 10692 1380
rect 10744 1368 10750 1420
rect 10870 1368 10876 1420
rect 10928 1368 10934 1420
rect 11054 1368 11060 1420
rect 11112 1368 11118 1420
rect 11624 1380 11836 1408
rect 10594 1340 10600 1352
rect 10428 1312 10600 1340
rect 10321 1303 10379 1309
rect 10594 1300 10600 1312
rect 10652 1300 10658 1352
rect 10686 1272 10692 1284
rect 8036 1244 9628 1272
rect 10152 1244 10692 1272
rect 8036 1213 8064 1244
rect 7791 1176 7880 1204
rect 8021 1207 8079 1213
rect 7791 1173 7803 1176
rect 7745 1167 7803 1173
rect 8021 1173 8033 1207
rect 8067 1173 8079 1207
rect 8021 1167 8079 1173
rect 8294 1164 8300 1216
rect 8352 1164 8358 1216
rect 8573 1207 8631 1213
rect 8573 1173 8585 1207
rect 8619 1204 8631 1207
rect 9122 1204 9128 1216
rect 8619 1176 9128 1204
rect 8619 1173 8631 1176
rect 8573 1167 8631 1173
rect 9122 1164 9128 1176
rect 9180 1164 9186 1216
rect 9214 1164 9220 1216
rect 9272 1164 9278 1216
rect 9309 1207 9367 1213
rect 9309 1173 9321 1207
rect 9355 1204 9367 1207
rect 9674 1204 9680 1216
rect 9355 1176 9680 1204
rect 9355 1173 9367 1176
rect 9309 1167 9367 1173
rect 9674 1164 9680 1176
rect 9732 1164 9738 1216
rect 9769 1207 9827 1213
rect 9769 1173 9781 1207
rect 9815 1204 9827 1207
rect 10042 1204 10048 1216
rect 9815 1176 10048 1204
rect 9815 1173 9827 1176
rect 9769 1167 9827 1173
rect 10042 1164 10048 1176
rect 10100 1164 10106 1216
rect 10152 1213 10180 1244
rect 10686 1232 10692 1244
rect 10744 1232 10750 1284
rect 10778 1232 10784 1284
rect 10836 1232 10842 1284
rect 10888 1272 10916 1368
rect 11624 1352 11652 1380
rect 11606 1300 11612 1352
rect 11664 1300 11670 1352
rect 11698 1300 11704 1352
rect 11756 1300 11762 1352
rect 11808 1349 11836 1380
rect 12176 1380 12572 1408
rect 11793 1343 11851 1349
rect 11793 1309 11805 1343
rect 11839 1309 11851 1343
rect 12176 1340 12204 1380
rect 11793 1303 11851 1309
rect 11900 1312 12204 1340
rect 11900 1272 11928 1312
rect 12250 1300 12256 1352
rect 12308 1300 12314 1352
rect 12544 1340 12572 1380
rect 13630 1368 13636 1420
rect 13688 1408 13694 1420
rect 16132 1408 16160 1504
rect 16224 1476 16252 1504
rect 16868 1476 16896 1507
rect 16224 1448 16896 1476
rect 13688 1380 16160 1408
rect 13688 1368 13694 1380
rect 16298 1368 16304 1420
rect 16356 1408 16362 1420
rect 17420 1408 17448 1507
rect 17494 1504 17500 1556
rect 17552 1544 17558 1556
rect 18509 1547 18567 1553
rect 18509 1544 18521 1547
rect 17552 1516 18521 1544
rect 17552 1504 17558 1516
rect 18509 1513 18521 1516
rect 18555 1513 18567 1547
rect 19429 1547 19487 1553
rect 19429 1544 19441 1547
rect 18509 1507 18567 1513
rect 18616 1516 19441 1544
rect 18616 1476 18644 1516
rect 19429 1513 19441 1516
rect 19475 1513 19487 1547
rect 19429 1507 19487 1513
rect 19794 1504 19800 1556
rect 19852 1544 19858 1556
rect 21085 1547 21143 1553
rect 21085 1544 21097 1547
rect 19852 1516 21097 1544
rect 19852 1504 19858 1516
rect 21085 1513 21097 1516
rect 21131 1513 21143 1547
rect 21085 1507 21143 1513
rect 21450 1504 21456 1556
rect 21508 1504 21514 1556
rect 21634 1504 21640 1556
rect 21692 1544 21698 1556
rect 23201 1547 23259 1553
rect 23201 1544 23213 1547
rect 21692 1516 23213 1544
rect 21692 1504 21698 1516
rect 23201 1513 23213 1516
rect 23247 1513 23259 1547
rect 23201 1507 23259 1513
rect 23474 1504 23480 1556
rect 23532 1544 23538 1556
rect 24670 1544 24676 1556
rect 23532 1516 24676 1544
rect 23532 1504 23538 1516
rect 24670 1504 24676 1516
rect 24728 1504 24734 1556
rect 17972 1448 18644 1476
rect 16356 1380 17448 1408
rect 16356 1368 16362 1380
rect 17494 1368 17500 1420
rect 17552 1408 17558 1420
rect 17972 1408 18000 1448
rect 18690 1436 18696 1488
rect 18748 1476 18754 1488
rect 20073 1479 20131 1485
rect 20073 1476 20085 1479
rect 18748 1448 20085 1476
rect 18748 1436 18754 1448
rect 20073 1445 20085 1448
rect 20119 1445 20131 1479
rect 20073 1439 20131 1445
rect 20625 1479 20683 1485
rect 20625 1445 20637 1479
rect 20671 1445 20683 1479
rect 20625 1439 20683 1445
rect 17552 1380 18000 1408
rect 17552 1368 17558 1380
rect 18046 1368 18052 1420
rect 18104 1368 18110 1420
rect 18598 1368 18604 1420
rect 18656 1408 18662 1420
rect 20640 1408 20668 1439
rect 21266 1436 21272 1488
rect 21324 1476 21330 1488
rect 24872 1476 24900 1720
rect 21324 1448 24900 1476
rect 21324 1436 21330 1448
rect 18656 1380 20668 1408
rect 18656 1368 18662 1380
rect 21082 1368 21088 1420
rect 21140 1408 21146 1420
rect 21140 1380 22232 1408
rect 21140 1368 21146 1380
rect 12897 1343 12955 1349
rect 12897 1340 12909 1343
rect 12360 1312 12480 1340
rect 12544 1312 12909 1340
rect 12360 1272 12388 1312
rect 10888 1244 11928 1272
rect 11992 1244 12388 1272
rect 10137 1207 10195 1213
rect 10137 1173 10149 1207
rect 10183 1173 10195 1207
rect 10137 1167 10195 1173
rect 10505 1207 10563 1213
rect 10505 1173 10517 1207
rect 10551 1204 10563 1207
rect 11422 1204 11428 1216
rect 10551 1176 11428 1204
rect 10551 1173 10563 1176
rect 10505 1167 10563 1173
rect 11422 1164 11428 1176
rect 11480 1164 11486 1216
rect 11992 1213 12020 1244
rect 11977 1207 12035 1213
rect 11977 1173 11989 1207
rect 12023 1173 12035 1207
rect 11977 1167 12035 1173
rect 12342 1164 12348 1216
rect 12400 1164 12406 1216
rect 12452 1204 12480 1312
rect 12897 1309 12909 1312
rect 12943 1309 12955 1343
rect 12897 1303 12955 1309
rect 13170 1300 13176 1352
rect 13228 1300 13234 1352
rect 13262 1300 13268 1352
rect 13320 1300 13326 1352
rect 14366 1300 14372 1352
rect 14424 1300 14430 1352
rect 14642 1300 14648 1352
rect 14700 1300 14706 1352
rect 14918 1300 14924 1352
rect 14976 1340 14982 1352
rect 15378 1340 15384 1352
rect 14976 1312 15384 1340
rect 14976 1300 14982 1312
rect 15378 1300 15384 1312
rect 15436 1300 15442 1352
rect 15470 1300 15476 1352
rect 15528 1340 15534 1352
rect 15841 1343 15899 1349
rect 15841 1340 15853 1343
rect 15528 1312 15853 1340
rect 15528 1300 15534 1312
rect 15841 1309 15853 1312
rect 15887 1309 15899 1343
rect 15841 1303 15899 1309
rect 16114 1300 16120 1352
rect 16172 1340 16178 1352
rect 16485 1343 16543 1349
rect 16485 1340 16497 1343
rect 16172 1312 16497 1340
rect 16172 1300 16178 1312
rect 16485 1309 16497 1312
rect 16531 1309 16543 1343
rect 16485 1303 16543 1309
rect 16574 1300 16580 1352
rect 16632 1340 16638 1352
rect 16761 1343 16819 1349
rect 16761 1340 16773 1343
rect 16632 1312 16773 1340
rect 16632 1300 16638 1312
rect 16761 1309 16773 1312
rect 16807 1309 16819 1343
rect 16761 1303 16819 1309
rect 16850 1300 16856 1352
rect 16908 1340 16914 1352
rect 17865 1343 17923 1349
rect 17865 1340 17877 1343
rect 16908 1312 17877 1340
rect 16908 1300 16914 1312
rect 17865 1309 17877 1312
rect 17911 1309 17923 1343
rect 18064 1340 18092 1368
rect 19061 1343 19119 1349
rect 19061 1340 19073 1343
rect 18064 1312 19073 1340
rect 17865 1303 17923 1309
rect 19061 1309 19073 1312
rect 19107 1309 19119 1343
rect 19889 1343 19947 1349
rect 19889 1340 19901 1343
rect 19061 1303 19119 1309
rect 19260 1312 19901 1340
rect 13188 1272 13216 1300
rect 14185 1275 14243 1281
rect 14185 1272 14197 1275
rect 13188 1244 14197 1272
rect 14185 1241 14197 1244
rect 14231 1241 14243 1275
rect 14384 1272 14412 1300
rect 15289 1275 15347 1281
rect 15289 1272 15301 1275
rect 14384 1244 15301 1272
rect 14185 1235 14243 1241
rect 15289 1241 15301 1244
rect 15335 1241 15347 1275
rect 17313 1275 17371 1281
rect 17313 1272 17325 1275
rect 15289 1235 15347 1241
rect 15396 1244 17325 1272
rect 12710 1204 12716 1216
rect 12452 1176 12716 1204
rect 12710 1164 12716 1176
rect 12768 1164 12774 1216
rect 13078 1164 13084 1216
rect 13136 1164 13142 1216
rect 13446 1164 13452 1216
rect 13504 1164 13510 1216
rect 13998 1164 14004 1216
rect 14056 1204 14062 1216
rect 14829 1207 14887 1213
rect 14829 1204 14841 1207
rect 14056 1176 14841 1204
rect 14056 1164 14062 1176
rect 14829 1173 14841 1176
rect 14875 1173 14887 1207
rect 14829 1167 14887 1173
rect 14918 1164 14924 1216
rect 14976 1204 14982 1216
rect 15396 1204 15424 1244
rect 17313 1241 17325 1244
rect 17359 1241 17371 1275
rect 17313 1235 17371 1241
rect 17402 1232 17408 1284
rect 17460 1272 17466 1284
rect 18417 1275 18475 1281
rect 18417 1272 18429 1275
rect 17460 1244 18429 1272
rect 17460 1232 17466 1244
rect 18417 1241 18429 1244
rect 18463 1241 18475 1275
rect 18417 1235 18475 1241
rect 14976 1176 15424 1204
rect 14976 1164 14982 1176
rect 16482 1164 16488 1216
rect 16540 1204 16546 1216
rect 17957 1207 18015 1213
rect 17957 1204 17969 1207
rect 16540 1176 17969 1204
rect 16540 1164 16546 1176
rect 17957 1173 17969 1176
rect 18003 1173 18015 1207
rect 17957 1167 18015 1173
rect 18877 1207 18935 1213
rect 18877 1173 18889 1207
rect 18923 1204 18935 1207
rect 19260 1204 19288 1312
rect 19889 1309 19901 1312
rect 19935 1309 19947 1343
rect 19889 1303 19947 1309
rect 19978 1300 19984 1352
rect 20036 1340 20042 1352
rect 20993 1343 21051 1349
rect 20993 1340 21005 1343
rect 20036 1312 21005 1340
rect 20036 1300 20042 1312
rect 20993 1309 21005 1312
rect 21039 1309 21051 1343
rect 20993 1303 21051 1309
rect 21174 1300 21180 1352
rect 21232 1340 21238 1352
rect 21637 1343 21695 1349
rect 21637 1340 21649 1343
rect 21232 1312 21649 1340
rect 21232 1300 21238 1312
rect 21637 1309 21649 1312
rect 21683 1309 21695 1343
rect 21637 1303 21695 1309
rect 21818 1300 21824 1352
rect 21876 1340 21882 1352
rect 22005 1343 22063 1349
rect 21876 1336 21956 1340
rect 22005 1336 22017 1343
rect 21876 1312 22017 1336
rect 21876 1300 21882 1312
rect 21928 1309 22017 1312
rect 22051 1309 22063 1343
rect 21928 1308 22063 1309
rect 22005 1303 22063 1308
rect 22097 1343 22155 1349
rect 22097 1309 22109 1343
rect 22143 1309 22155 1343
rect 22204 1340 22232 1380
rect 22738 1368 22744 1420
rect 22796 1408 22802 1420
rect 22796 1380 23612 1408
rect 22796 1368 22802 1380
rect 22373 1343 22431 1349
rect 22373 1340 22385 1343
rect 22204 1312 22385 1340
rect 22097 1303 22155 1309
rect 22373 1309 22385 1312
rect 22419 1309 22431 1343
rect 22373 1303 22431 1309
rect 19337 1275 19395 1281
rect 19337 1241 19349 1275
rect 19383 1241 19395 1275
rect 19337 1235 19395 1241
rect 18923 1176 19288 1204
rect 19352 1204 19380 1235
rect 19702 1232 19708 1284
rect 19760 1272 19766 1284
rect 20441 1275 20499 1281
rect 20441 1272 20453 1275
rect 19760 1244 20453 1272
rect 19760 1232 19766 1244
rect 20441 1241 20453 1244
rect 20487 1241 20499 1275
rect 20441 1235 20499 1241
rect 20622 1232 20628 1284
rect 20680 1272 20686 1284
rect 22112 1272 22140 1303
rect 22646 1300 22652 1352
rect 22704 1300 22710 1352
rect 22925 1343 22983 1349
rect 22925 1309 22937 1343
rect 22971 1309 22983 1343
rect 22925 1303 22983 1309
rect 23385 1343 23443 1349
rect 23385 1309 23397 1343
rect 23431 1309 23443 1343
rect 23385 1303 23443 1309
rect 22940 1272 22968 1303
rect 20680 1244 22140 1272
rect 22204 1244 22968 1272
rect 23400 1272 23428 1303
rect 23474 1300 23480 1352
rect 23532 1300 23538 1352
rect 23584 1340 23612 1380
rect 24670 1368 24676 1420
rect 24728 1408 24734 1420
rect 25590 1408 25596 1420
rect 24728 1380 25596 1408
rect 24728 1368 24734 1380
rect 25590 1368 25596 1380
rect 25648 1368 25654 1420
rect 23753 1343 23811 1349
rect 23753 1340 23765 1343
rect 23584 1312 23765 1340
rect 23753 1309 23765 1312
rect 23799 1309 23811 1343
rect 23753 1303 23811 1309
rect 24026 1300 24032 1352
rect 24084 1300 24090 1352
rect 23566 1272 23572 1284
rect 23400 1244 23572 1272
rect 20680 1232 20686 1244
rect 19426 1204 19432 1216
rect 19352 1176 19432 1204
rect 18923 1173 18935 1176
rect 18877 1167 18935 1173
rect 19426 1164 19432 1176
rect 19484 1164 19490 1216
rect 20070 1164 20076 1216
rect 20128 1204 20134 1216
rect 21821 1207 21879 1213
rect 21821 1204 21833 1207
rect 20128 1176 21833 1204
rect 20128 1164 20134 1176
rect 21821 1173 21833 1176
rect 21867 1173 21879 1207
rect 21821 1167 21879 1173
rect 22002 1164 22008 1216
rect 22060 1204 22066 1216
rect 22204 1204 22232 1244
rect 23566 1232 23572 1244
rect 23624 1232 23630 1284
rect 22060 1176 22232 1204
rect 22060 1164 22066 1176
rect 22278 1164 22284 1216
rect 22336 1164 22342 1216
rect 22554 1164 22560 1216
rect 22612 1164 22618 1216
rect 22738 1164 22744 1216
rect 22796 1204 22802 1216
rect 22833 1207 22891 1213
rect 22833 1204 22845 1207
rect 22796 1176 22845 1204
rect 22796 1164 22802 1176
rect 22833 1173 22845 1176
rect 22879 1173 22891 1207
rect 22833 1167 22891 1173
rect 23106 1164 23112 1216
rect 23164 1164 23170 1216
rect 23290 1164 23296 1216
rect 23348 1204 23354 1216
rect 23661 1207 23719 1213
rect 23661 1204 23673 1207
rect 23348 1176 23673 1204
rect 23348 1164 23354 1176
rect 23661 1173 23673 1176
rect 23707 1173 23719 1207
rect 23661 1167 23719 1173
rect 23934 1164 23940 1216
rect 23992 1164 23998 1216
rect 24210 1164 24216 1216
rect 24268 1164 24274 1216
rect 1104 1114 25000 1136
rect 1104 1062 6884 1114
rect 6936 1062 6948 1114
rect 7000 1062 7012 1114
rect 7064 1062 7076 1114
rect 7128 1062 7140 1114
rect 7192 1062 12818 1114
rect 12870 1062 12882 1114
rect 12934 1062 12946 1114
rect 12998 1062 13010 1114
rect 13062 1062 13074 1114
rect 13126 1062 18752 1114
rect 18804 1062 18816 1114
rect 18868 1062 18880 1114
rect 18932 1062 18944 1114
rect 18996 1062 19008 1114
rect 19060 1062 24686 1114
rect 24738 1062 24750 1114
rect 24802 1062 24814 1114
rect 24866 1062 24878 1114
rect 24930 1062 24942 1114
rect 24994 1062 25000 1114
rect 1104 1040 25000 1062
rect 2038 960 2044 1012
rect 2096 960 2102 1012
rect 2314 960 2320 1012
rect 2372 1000 2378 1012
rect 2372 972 2774 1000
rect 2372 960 2378 972
rect 2056 796 2084 960
rect 2746 932 2774 972
rect 3326 960 3332 1012
rect 3384 1000 3390 1012
rect 5258 1000 5264 1012
rect 3384 972 5264 1000
rect 3384 960 3390 972
rect 5258 960 5264 972
rect 5316 960 5322 1012
rect 9214 960 9220 1012
rect 9272 1000 9278 1012
rect 13630 1000 13636 1012
rect 9272 972 13636 1000
rect 9272 960 9278 972
rect 13630 960 13636 972
rect 13688 960 13694 1012
rect 16666 960 16672 1012
rect 16724 1000 16730 1012
rect 17402 1000 17408 1012
rect 16724 972 17408 1000
rect 16724 960 16730 972
rect 17402 960 17408 972
rect 17460 960 17466 1012
rect 22278 1000 22284 1012
rect 22066 972 22284 1000
rect 5718 932 5724 944
rect 2746 904 5724 932
rect 5718 892 5724 904
rect 5776 892 5782 944
rect 5994 892 6000 944
rect 6052 932 6058 944
rect 10778 932 10784 944
rect 6052 904 10784 932
rect 6052 892 6058 904
rect 10778 892 10784 904
rect 10836 892 10842 944
rect 11238 892 11244 944
rect 11296 932 11302 944
rect 14918 932 14924 944
rect 11296 904 14924 932
rect 11296 892 11302 904
rect 14918 892 14924 904
rect 14976 892 14982 944
rect 15010 892 15016 944
rect 15068 932 15074 944
rect 22066 932 22094 972
rect 22278 960 22284 972
rect 22336 960 22342 1012
rect 22554 960 22560 1012
rect 22612 960 22618 1012
rect 23290 960 23296 1012
rect 23348 960 23354 1012
rect 15068 904 22094 932
rect 15068 892 15074 904
rect 7834 864 7840 876
rect 6012 836 7840 864
rect 2056 768 3924 796
rect 2774 688 2780 740
rect 2832 728 2838 740
rect 3510 728 3516 740
rect 2832 700 3516 728
rect 2832 688 2838 700
rect 3510 688 3516 700
rect 3568 688 3574 740
rect 3896 184 3924 768
rect 4522 756 4528 808
rect 4580 796 4586 808
rect 6012 796 6040 836
rect 7834 824 7840 836
rect 7892 824 7898 876
rect 8294 824 8300 876
rect 8352 824 8358 876
rect 9674 824 9680 876
rect 9732 864 9738 876
rect 9732 836 12434 864
rect 9732 824 9738 836
rect 4580 768 6040 796
rect 4580 756 4586 768
rect 6362 756 6368 808
rect 6420 756 6426 808
rect 7466 756 7472 808
rect 7524 756 7530 808
rect 4798 688 4804 740
rect 4856 728 4862 740
rect 5534 728 5540 740
rect 4856 700 5540 728
rect 4856 688 4862 700
rect 5534 688 5540 700
rect 5592 688 5598 740
rect 5166 620 5172 672
rect 5224 620 5230 672
rect 5184 456 5212 620
rect 6380 524 6408 756
rect 7484 592 7512 756
rect 8312 660 8340 824
rect 9122 756 9128 808
rect 9180 796 9186 808
rect 9766 796 9772 808
rect 9180 768 9772 796
rect 9180 756 9186 768
rect 9766 756 9772 768
rect 9824 756 9830 808
rect 12406 796 12434 836
rect 13630 824 13636 876
rect 13688 864 13694 876
rect 22572 864 22600 960
rect 23308 932 23336 960
rect 13688 836 22600 864
rect 22664 904 23336 932
rect 13688 824 13694 836
rect 14642 796 14648 808
rect 12406 768 14648 796
rect 14642 756 14648 768
rect 14700 756 14706 808
rect 22664 796 22692 904
rect 22738 824 22744 876
rect 22796 824 22802 876
rect 17052 768 22692 796
rect 8846 688 8852 740
rect 8904 728 8910 740
rect 9674 728 9680 740
rect 8904 700 9680 728
rect 8904 688 8910 700
rect 9674 688 9680 700
rect 9732 688 9738 740
rect 16942 660 16948 672
rect 8312 632 16948 660
rect 16942 620 16948 632
rect 17000 620 17006 672
rect 9950 592 9956 604
rect 7484 564 9956 592
rect 9950 552 9956 564
rect 10008 552 10014 604
rect 13906 552 13912 604
rect 13964 592 13970 604
rect 17052 592 17080 768
rect 21266 688 21272 740
rect 21324 728 21330 740
rect 22646 728 22652 740
rect 21324 700 22652 728
rect 21324 688 21330 700
rect 22646 688 22652 700
rect 22704 688 22710 740
rect 21450 620 21456 672
rect 21508 660 21514 672
rect 22002 660 22008 672
rect 21508 632 22008 660
rect 21508 620 21514 632
rect 22002 620 22008 632
rect 22060 620 22066 672
rect 22756 592 22784 824
rect 23474 688 23480 740
rect 23532 688 23538 740
rect 23492 592 23520 688
rect 13964 564 17080 592
rect 17328 564 22784 592
rect 22940 564 23520 592
rect 13964 552 13970 564
rect 11606 524 11612 536
rect 6380 496 11612 524
rect 11606 484 11612 496
rect 11664 484 11670 536
rect 13354 484 13360 536
rect 13412 524 13418 536
rect 17328 524 17356 564
rect 13412 496 17356 524
rect 13412 484 13418 496
rect 22002 484 22008 536
rect 22060 524 22066 536
rect 22940 524 22968 564
rect 24210 552 24216 604
rect 24268 552 24274 604
rect 24228 524 24256 552
rect 22060 496 22968 524
rect 23032 496 24256 524
rect 22060 484 22066 496
rect 10134 456 10140 468
rect 5184 428 10140 456
rect 10134 416 10140 428
rect 10192 416 10198 468
rect 16114 456 16120 468
rect 12406 428 16120 456
rect 4706 348 4712 400
rect 4764 388 4770 400
rect 7834 388 7840 400
rect 4764 360 7840 388
rect 4764 348 4770 360
rect 7834 348 7840 360
rect 7892 348 7898 400
rect 8018 348 8024 400
rect 8076 388 8082 400
rect 12406 388 12434 428
rect 16114 416 16120 428
rect 16172 416 16178 468
rect 16390 416 16396 468
rect 16448 456 16454 468
rect 23032 456 23060 496
rect 16448 428 23060 456
rect 16448 416 16454 428
rect 23106 416 23112 468
rect 23164 416 23170 468
rect 8076 360 12434 388
rect 8076 348 8082 360
rect 12526 348 12532 400
rect 12584 388 12590 400
rect 23124 388 23152 416
rect 12584 360 23152 388
rect 12584 348 12590 360
rect 11330 280 11336 332
rect 11388 280 11394 332
rect 22738 280 22744 332
rect 22796 320 22802 332
rect 24026 320 24032 332
rect 22796 292 24032 320
rect 22796 280 22802 292
rect 24026 280 24032 292
rect 24084 280 24090 332
rect 3970 212 3976 264
rect 4028 252 4034 264
rect 11348 252 11376 280
rect 4028 224 11376 252
rect 4028 212 4034 224
rect 10226 184 10232 196
rect 3896 156 10232 184
rect 10226 144 10232 156
rect 10284 144 10290 196
<< via1 >>
rect 6884 6502 6936 6554
rect 6948 6502 7000 6554
rect 7012 6502 7064 6554
rect 7076 6502 7128 6554
rect 7140 6502 7192 6554
rect 12818 6502 12870 6554
rect 12882 6502 12934 6554
rect 12946 6502 12998 6554
rect 13010 6502 13062 6554
rect 13074 6502 13126 6554
rect 18752 6502 18804 6554
rect 18816 6502 18868 6554
rect 18880 6502 18932 6554
rect 18944 6502 18996 6554
rect 19008 6502 19060 6554
rect 24686 6502 24738 6554
rect 24750 6502 24802 6554
rect 24814 6502 24866 6554
rect 24878 6502 24930 6554
rect 24942 6502 24994 6554
rect 2136 6400 2188 6452
rect 3792 6400 3844 6452
rect 4620 6443 4672 6452
rect 4620 6409 4629 6443
rect 4629 6409 4663 6443
rect 4663 6409 4672 6443
rect 4620 6400 4672 6409
rect 1400 6375 1452 6384
rect 1400 6341 1409 6375
rect 1409 6341 1443 6375
rect 1443 6341 1452 6375
rect 1400 6332 1452 6341
rect 2228 6307 2280 6316
rect 2228 6273 2237 6307
rect 2237 6273 2271 6307
rect 2271 6273 2280 6307
rect 2228 6264 2280 6273
rect 5632 6332 5684 6384
rect 7288 6400 7340 6452
rect 6092 6375 6144 6384
rect 6092 6341 6101 6375
rect 6101 6341 6135 6375
rect 6135 6341 6144 6375
rect 6092 6332 6144 6341
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 10600 6443 10652 6452
rect 10600 6409 10609 6443
rect 10609 6409 10643 6443
rect 10643 6409 10652 6443
rect 10600 6400 10652 6409
rect 11980 6443 12032 6452
rect 11980 6409 11989 6443
rect 11989 6409 12023 6443
rect 12023 6409 12032 6443
rect 11980 6400 12032 6409
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 9680 6264 9732 6316
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 12348 6307 12400 6316
rect 12348 6273 12357 6307
rect 12357 6273 12391 6307
rect 12391 6273 12400 6307
rect 12348 6264 12400 6273
rect 13176 6443 13228 6452
rect 13176 6409 13185 6443
rect 13185 6409 13219 6443
rect 13219 6409 13228 6443
rect 13176 6400 13228 6409
rect 12624 6307 12676 6316
rect 12624 6273 12633 6307
rect 12633 6273 12667 6307
rect 12667 6273 12676 6307
rect 12624 6264 12676 6273
rect 14280 6443 14332 6452
rect 14280 6409 14289 6443
rect 14289 6409 14323 6443
rect 14323 6409 14332 6443
rect 14280 6400 14332 6409
rect 15384 6443 15436 6452
rect 15384 6409 15393 6443
rect 15393 6409 15427 6443
rect 15427 6409 15436 6443
rect 15384 6400 15436 6409
rect 16856 6443 16908 6452
rect 16856 6409 16865 6443
rect 16865 6409 16899 6443
rect 16899 6409 16908 6443
rect 16856 6400 16908 6409
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 19432 6443 19484 6452
rect 19432 6409 19441 6443
rect 19441 6409 19475 6443
rect 19475 6409 19484 6443
rect 19432 6400 19484 6409
rect 20352 6443 20404 6452
rect 20352 6409 20361 6443
rect 20361 6409 20395 6443
rect 20395 6409 20404 6443
rect 20352 6400 20404 6409
rect 21548 6443 21600 6452
rect 21548 6409 21557 6443
rect 21557 6409 21591 6443
rect 21591 6409 21600 6443
rect 21548 6400 21600 6409
rect 13544 6307 13596 6316
rect 13544 6273 13553 6307
rect 13553 6273 13587 6307
rect 13587 6273 13596 6307
rect 13544 6264 13596 6273
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 15108 6307 15160 6316
rect 15108 6273 15117 6307
rect 15117 6273 15151 6307
rect 15151 6273 15160 6307
rect 15108 6264 15160 6273
rect 15660 6264 15712 6316
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 18328 6307 18380 6316
rect 18328 6273 18337 6307
rect 18337 6273 18371 6307
rect 18371 6273 18380 6307
rect 18328 6264 18380 6273
rect 19984 6307 20036 6316
rect 19984 6273 19993 6307
rect 19993 6273 20027 6307
rect 20027 6273 20036 6307
rect 19984 6264 20036 6273
rect 20536 6307 20588 6316
rect 20536 6273 20545 6307
rect 20545 6273 20579 6307
rect 20579 6273 20588 6307
rect 20536 6264 20588 6273
rect 23664 6400 23716 6452
rect 5632 6128 5684 6180
rect 21640 6196 21692 6248
rect 23112 6307 23164 6316
rect 23112 6273 23121 6307
rect 23121 6273 23155 6307
rect 23155 6273 23164 6307
rect 23112 6264 23164 6273
rect 23664 6307 23716 6316
rect 23664 6273 23673 6307
rect 23673 6273 23707 6307
rect 23707 6273 23716 6307
rect 23664 6264 23716 6273
rect 24216 6128 24268 6180
rect 22560 6103 22612 6112
rect 22560 6069 22569 6103
rect 22569 6069 22603 6103
rect 22603 6069 22612 6103
rect 22560 6060 22612 6069
rect 3917 5958 3969 6010
rect 3981 5958 4033 6010
rect 4045 5958 4097 6010
rect 4109 5958 4161 6010
rect 4173 5958 4225 6010
rect 9851 5958 9903 6010
rect 9915 5958 9967 6010
rect 9979 5958 10031 6010
rect 10043 5958 10095 6010
rect 10107 5958 10159 6010
rect 15785 5958 15837 6010
rect 15849 5958 15901 6010
rect 15913 5958 15965 6010
rect 15977 5958 16029 6010
rect 16041 5958 16093 6010
rect 21719 5958 21771 6010
rect 21783 5958 21835 6010
rect 21847 5958 21899 6010
rect 21911 5958 21963 6010
rect 21975 5958 22027 6010
rect 6552 5856 6604 5908
rect 7564 5856 7616 5908
rect 8760 5856 8812 5908
rect 9680 5899 9732 5908
rect 9680 5865 9689 5899
rect 9689 5865 9723 5899
rect 9723 5865 9732 5899
rect 9680 5856 9732 5865
rect 11152 5856 11204 5908
rect 12348 5856 12400 5908
rect 12624 5856 12676 5908
rect 13544 5856 13596 5908
rect 14648 5856 14700 5908
rect 15108 5856 15160 5908
rect 15660 5856 15712 5908
rect 17408 5856 17460 5908
rect 18328 5856 18380 5908
rect 20536 5856 20588 5908
rect 24492 5856 24544 5908
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 9864 5695 9916 5704
rect 9864 5661 9873 5695
rect 9873 5661 9907 5695
rect 9907 5661 9916 5695
rect 9864 5652 9916 5661
rect 11060 5695 11112 5704
rect 11060 5661 11069 5695
rect 11069 5661 11103 5695
rect 11103 5661 11112 5695
rect 11060 5652 11112 5661
rect 11980 5695 12032 5704
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 12440 5695 12492 5704
rect 12440 5661 12449 5695
rect 12449 5661 12483 5695
rect 12483 5661 12492 5695
rect 12440 5652 12492 5661
rect 13452 5695 13504 5704
rect 13452 5661 13461 5695
rect 13461 5661 13495 5695
rect 13495 5661 13504 5695
rect 13452 5652 13504 5661
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 14832 5695 14884 5704
rect 14832 5661 14841 5695
rect 14841 5661 14875 5695
rect 14875 5661 14884 5695
rect 14832 5652 14884 5661
rect 19984 5788 20036 5840
rect 24032 5788 24084 5840
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 17132 5695 17184 5704
rect 17132 5661 17141 5695
rect 17141 5661 17175 5695
rect 17175 5661 17184 5695
rect 17132 5652 17184 5661
rect 18420 5695 18472 5704
rect 18420 5661 18429 5695
rect 18429 5661 18463 5695
rect 18463 5661 18472 5695
rect 18420 5652 18472 5661
rect 19984 5695 20036 5704
rect 19984 5661 19993 5695
rect 19993 5661 20027 5695
rect 20027 5661 20036 5695
rect 19984 5652 20036 5661
rect 23848 5627 23900 5636
rect 23848 5593 23857 5627
rect 23857 5593 23891 5627
rect 23891 5593 23900 5627
rect 23848 5584 23900 5593
rect 6884 5414 6936 5466
rect 6948 5414 7000 5466
rect 7012 5414 7064 5466
rect 7076 5414 7128 5466
rect 7140 5414 7192 5466
rect 12818 5414 12870 5466
rect 12882 5414 12934 5466
rect 12946 5414 12998 5466
rect 13010 5414 13062 5466
rect 13074 5414 13126 5466
rect 18752 5414 18804 5466
rect 18816 5414 18868 5466
rect 18880 5414 18932 5466
rect 18944 5414 18996 5466
rect 19008 5414 19060 5466
rect 24686 5414 24738 5466
rect 24750 5414 24802 5466
rect 24814 5414 24866 5466
rect 24878 5414 24930 5466
rect 24942 5414 24994 5466
rect 6276 5312 6328 5364
rect 7564 5355 7616 5364
rect 7564 5321 7573 5355
rect 7573 5321 7607 5355
rect 7607 5321 7616 5355
rect 7564 5312 7616 5321
rect 8760 5355 8812 5364
rect 8760 5321 8769 5355
rect 8769 5321 8803 5355
rect 8803 5321 8812 5355
rect 8760 5312 8812 5321
rect 9864 5355 9916 5364
rect 9864 5321 9873 5355
rect 9873 5321 9907 5355
rect 9907 5321 9916 5355
rect 9864 5312 9916 5321
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 11980 5355 12032 5364
rect 11980 5321 11989 5355
rect 11989 5321 12023 5355
rect 12023 5321 12032 5355
rect 11980 5312 12032 5321
rect 12440 5355 12492 5364
rect 12440 5321 12449 5355
rect 12449 5321 12483 5355
rect 12483 5321 12492 5355
rect 12440 5312 12492 5321
rect 13452 5355 13504 5364
rect 13452 5321 13461 5355
rect 13461 5321 13495 5355
rect 13495 5321 13504 5355
rect 13452 5312 13504 5321
rect 14556 5355 14608 5364
rect 14556 5321 14565 5355
rect 14565 5321 14599 5355
rect 14599 5321 14608 5355
rect 14556 5312 14608 5321
rect 14832 5355 14884 5364
rect 14832 5321 14841 5355
rect 14841 5321 14875 5355
rect 14875 5321 14884 5355
rect 14832 5312 14884 5321
rect 15936 5355 15988 5364
rect 15936 5321 15945 5355
rect 15945 5321 15979 5355
rect 15979 5321 15988 5355
rect 15936 5312 15988 5321
rect 17132 5355 17184 5364
rect 17132 5321 17141 5355
rect 17141 5321 17175 5355
rect 17175 5321 17184 5355
rect 17132 5312 17184 5321
rect 18420 5355 18472 5364
rect 18420 5321 18429 5355
rect 18429 5321 18463 5355
rect 18463 5321 18472 5355
rect 18420 5312 18472 5321
rect 19984 5355 20036 5364
rect 19984 5321 19993 5355
rect 19993 5321 20027 5355
rect 20027 5321 20036 5355
rect 19984 5312 20036 5321
rect 23848 5312 23900 5364
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 13912 5244 13964 5296
rect 11244 5219 11296 5228
rect 11244 5185 11253 5219
rect 11253 5185 11287 5219
rect 11287 5185 11296 5219
rect 11244 5176 11296 5185
rect 9588 5108 9640 5160
rect 13728 5176 13780 5228
rect 14740 5219 14792 5228
rect 14740 5185 14749 5219
rect 14749 5185 14783 5219
rect 14783 5185 14792 5219
rect 14740 5176 14792 5185
rect 15016 5219 15068 5228
rect 15016 5185 15025 5219
rect 15025 5185 15059 5219
rect 15059 5185 15068 5219
rect 15016 5176 15068 5185
rect 13636 5040 13688 5092
rect 12624 4972 12676 5024
rect 17868 5176 17920 5228
rect 21456 5176 21508 5228
rect 24308 5219 24360 5228
rect 24308 5185 24317 5219
rect 24317 5185 24351 5219
rect 24351 5185 24360 5219
rect 24308 5176 24360 5185
rect 21364 5108 21416 5160
rect 21272 5040 21324 5092
rect 16396 4972 16448 5024
rect 3917 4870 3969 4922
rect 3981 4870 4033 4922
rect 4045 4870 4097 4922
rect 4109 4870 4161 4922
rect 4173 4870 4225 4922
rect 9851 4870 9903 4922
rect 9915 4870 9967 4922
rect 9979 4870 10031 4922
rect 10043 4870 10095 4922
rect 10107 4870 10159 4922
rect 15785 4870 15837 4922
rect 15849 4870 15901 4922
rect 15913 4870 15965 4922
rect 15977 4870 16029 4922
rect 16041 4870 16093 4922
rect 21719 4870 21771 4922
rect 21783 4870 21835 4922
rect 21847 4870 21899 4922
rect 21911 4870 21963 4922
rect 21975 4870 22027 4922
rect 6552 4768 6604 4820
rect 24308 4768 24360 4820
rect 13360 4632 13412 4684
rect 23940 4607 23992 4616
rect 23940 4573 23949 4607
rect 23949 4573 23983 4607
rect 23983 4573 23992 4607
rect 23940 4564 23992 4573
rect 6884 4326 6936 4378
rect 6948 4326 7000 4378
rect 7012 4326 7064 4378
rect 7076 4326 7128 4378
rect 7140 4326 7192 4378
rect 12818 4326 12870 4378
rect 12882 4326 12934 4378
rect 12946 4326 12998 4378
rect 13010 4326 13062 4378
rect 13074 4326 13126 4378
rect 18752 4326 18804 4378
rect 18816 4326 18868 4378
rect 18880 4326 18932 4378
rect 18944 4326 18996 4378
rect 19008 4326 19060 4378
rect 24686 4326 24738 4378
rect 24750 4326 24802 4378
rect 24814 4326 24866 4378
rect 24878 4326 24930 4378
rect 24942 4326 24994 4378
rect 3917 3782 3969 3834
rect 3981 3782 4033 3834
rect 4045 3782 4097 3834
rect 4109 3782 4161 3834
rect 4173 3782 4225 3834
rect 9851 3782 9903 3834
rect 9915 3782 9967 3834
rect 9979 3782 10031 3834
rect 10043 3782 10095 3834
rect 10107 3782 10159 3834
rect 15785 3782 15837 3834
rect 15849 3782 15901 3834
rect 15913 3782 15965 3834
rect 15977 3782 16029 3834
rect 16041 3782 16093 3834
rect 21719 3782 21771 3834
rect 21783 3782 21835 3834
rect 21847 3782 21899 3834
rect 21911 3782 21963 3834
rect 21975 3782 22027 3834
rect 23664 3680 23716 3732
rect 24124 3519 24176 3528
rect 24124 3485 24133 3519
rect 24133 3485 24167 3519
rect 24167 3485 24176 3519
rect 24124 3476 24176 3485
rect 23204 3340 23256 3392
rect 24308 3340 24360 3392
rect 6884 3238 6936 3290
rect 6948 3238 7000 3290
rect 7012 3238 7064 3290
rect 7076 3238 7128 3290
rect 7140 3238 7192 3290
rect 12818 3238 12870 3290
rect 12882 3238 12934 3290
rect 12946 3238 12998 3290
rect 13010 3238 13062 3290
rect 13074 3238 13126 3290
rect 18752 3238 18804 3290
rect 18816 3238 18868 3290
rect 18880 3238 18932 3290
rect 18944 3238 18996 3290
rect 19008 3238 19060 3290
rect 24686 3238 24738 3290
rect 24750 3238 24802 3290
rect 24814 3238 24866 3290
rect 24878 3238 24930 3290
rect 24942 3238 24994 3290
rect 24124 3179 24176 3188
rect 24124 3145 24133 3179
rect 24133 3145 24167 3179
rect 24167 3145 24176 3179
rect 24124 3136 24176 3145
rect 25044 3068 25096 3120
rect 1584 2932 1636 2984
rect 14372 2932 14424 2984
rect 17868 2864 17920 2916
rect 22652 2864 22704 2916
rect 24308 3043 24360 3052
rect 24308 3009 24317 3043
rect 24317 3009 24351 3043
rect 24351 3009 24360 3043
rect 24308 3000 24360 3009
rect 24492 2932 24544 2984
rect 24584 2864 24636 2916
rect 9496 2796 9548 2848
rect 12532 2796 12584 2848
rect 13176 2796 13228 2848
rect 15568 2796 15620 2848
rect 19616 2796 19668 2848
rect 20996 2796 21048 2848
rect 23020 2796 23072 2848
rect 23572 2839 23624 2848
rect 23572 2805 23581 2839
rect 23581 2805 23615 2839
rect 23615 2805 23624 2839
rect 23572 2796 23624 2805
rect 24032 2796 24084 2848
rect 3917 2694 3969 2746
rect 3981 2694 4033 2746
rect 4045 2694 4097 2746
rect 4109 2694 4161 2746
rect 4173 2694 4225 2746
rect 9851 2694 9903 2746
rect 9915 2694 9967 2746
rect 9979 2694 10031 2746
rect 10043 2694 10095 2746
rect 10107 2694 10159 2746
rect 15785 2694 15837 2746
rect 15849 2694 15901 2746
rect 15913 2694 15965 2746
rect 15977 2694 16029 2746
rect 16041 2694 16093 2746
rect 21719 2694 21771 2746
rect 21783 2694 21835 2746
rect 21847 2694 21899 2746
rect 21911 2694 21963 2746
rect 21975 2694 22027 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 2596 2592 2648 2644
rect 9128 2592 9180 2644
rect 5724 2524 5776 2576
rect 6276 2567 6328 2576
rect 6276 2533 6285 2567
rect 6285 2533 6319 2567
rect 6319 2533 6328 2567
rect 6276 2524 6328 2533
rect 7196 2567 7248 2576
rect 7196 2533 7205 2567
rect 7205 2533 7239 2567
rect 7239 2533 7248 2567
rect 7196 2524 7248 2533
rect 7564 2524 7616 2576
rect 480 2456 532 2508
rect 1308 2388 1360 2440
rect 4068 2456 4120 2508
rect 9036 2456 9088 2508
rect 204 2320 256 2372
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 6092 2431 6144 2440
rect 6092 2397 6101 2431
rect 6101 2397 6135 2431
rect 6135 2397 6144 2431
rect 6092 2388 6144 2397
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 1860 2252 1912 2304
rect 3332 2320 3384 2372
rect 6736 2320 6788 2372
rect 2412 2295 2464 2304
rect 2412 2261 2421 2295
rect 2421 2261 2455 2295
rect 2455 2261 2464 2295
rect 2412 2252 2464 2261
rect 3424 2252 3476 2304
rect 4436 2252 4488 2304
rect 5080 2252 5132 2304
rect 9496 2456 9548 2508
rect 13268 2524 13320 2576
rect 15016 2592 15068 2644
rect 22652 2592 22704 2644
rect 23204 2635 23256 2644
rect 23204 2601 23213 2635
rect 23213 2601 23247 2635
rect 23247 2601 23256 2635
rect 23204 2592 23256 2601
rect 9312 2388 9364 2440
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 9220 2320 9272 2372
rect 10692 2388 10744 2440
rect 11796 2388 11848 2440
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12164 2456 12216 2508
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 14188 2456 14240 2508
rect 11612 2320 11664 2372
rect 9404 2295 9456 2304
rect 9404 2261 9413 2295
rect 9413 2261 9447 2295
rect 9447 2261 9456 2295
rect 9404 2252 9456 2261
rect 9496 2252 9548 2304
rect 11244 2252 11296 2304
rect 11796 2295 11848 2304
rect 11796 2261 11805 2295
rect 11805 2261 11839 2295
rect 11839 2261 11848 2295
rect 11796 2252 11848 2261
rect 12440 2320 12492 2372
rect 15384 2388 15436 2440
rect 15568 2431 15620 2440
rect 15568 2397 15577 2431
rect 15577 2397 15611 2431
rect 15611 2397 15620 2431
rect 15568 2388 15620 2397
rect 19432 2524 19484 2576
rect 16028 2388 16080 2440
rect 16488 2431 16540 2440
rect 16488 2397 16497 2431
rect 16497 2397 16531 2431
rect 16531 2397 16540 2431
rect 16488 2388 16540 2397
rect 14556 2320 14608 2372
rect 16948 2388 17000 2440
rect 17592 2431 17644 2440
rect 17592 2397 17601 2431
rect 17601 2397 17635 2431
rect 17635 2397 17644 2431
rect 17592 2388 17644 2397
rect 17868 2431 17920 2440
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 17960 2388 18012 2440
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 19340 2456 19392 2508
rect 21364 2524 21416 2576
rect 18972 2431 19024 2440
rect 18972 2397 18981 2431
rect 18981 2397 19015 2431
rect 19015 2397 19024 2431
rect 18972 2388 19024 2397
rect 19708 2431 19760 2440
rect 19708 2397 19717 2431
rect 19717 2397 19751 2431
rect 19751 2397 19760 2431
rect 19708 2388 19760 2397
rect 20076 2388 20128 2440
rect 20260 2431 20312 2440
rect 20260 2397 20269 2431
rect 20269 2397 20303 2431
rect 20303 2397 20312 2431
rect 20260 2388 20312 2397
rect 12348 2295 12400 2304
rect 12348 2261 12357 2295
rect 12357 2261 12391 2295
rect 12391 2261 12400 2295
rect 12348 2252 12400 2261
rect 12716 2252 12768 2304
rect 14004 2252 14056 2304
rect 15292 2252 15344 2304
rect 15476 2252 15528 2304
rect 15568 2252 15620 2304
rect 16672 2252 16724 2304
rect 16856 2295 16908 2304
rect 16856 2261 16865 2295
rect 16865 2261 16899 2295
rect 16899 2261 16908 2295
rect 16856 2252 16908 2261
rect 17776 2252 17828 2304
rect 18052 2252 18104 2304
rect 18144 2252 18196 2304
rect 18236 2295 18288 2304
rect 18236 2261 18245 2295
rect 18245 2261 18279 2295
rect 18279 2261 18288 2295
rect 18236 2252 18288 2261
rect 19156 2252 19208 2304
rect 19248 2295 19300 2304
rect 19248 2261 19257 2295
rect 19257 2261 19291 2295
rect 19291 2261 19300 2295
rect 19248 2252 19300 2261
rect 19708 2252 19760 2304
rect 19984 2252 20036 2304
rect 20168 2320 20220 2372
rect 22376 2431 22428 2440
rect 22376 2397 22385 2431
rect 22385 2397 22419 2431
rect 22419 2397 22428 2431
rect 22376 2388 22428 2397
rect 22836 2431 22888 2440
rect 22836 2397 22845 2431
rect 22845 2397 22879 2431
rect 22879 2397 22888 2431
rect 22836 2388 22888 2397
rect 23296 2388 23348 2440
rect 25320 2456 25372 2508
rect 23756 2388 23808 2440
rect 24032 2388 24084 2440
rect 20352 2295 20404 2304
rect 20352 2261 20361 2295
rect 20361 2261 20395 2295
rect 20395 2261 20404 2295
rect 20352 2252 20404 2261
rect 20628 2295 20680 2304
rect 20628 2261 20637 2295
rect 20637 2261 20671 2295
rect 20671 2261 20680 2295
rect 20628 2252 20680 2261
rect 22652 2295 22704 2304
rect 22652 2261 22661 2295
rect 22661 2261 22695 2295
rect 22695 2261 22704 2295
rect 22652 2252 22704 2261
rect 23848 2320 23900 2372
rect 23940 2252 23992 2304
rect 24032 2295 24084 2304
rect 24032 2261 24041 2295
rect 24041 2261 24075 2295
rect 24075 2261 24084 2295
rect 24032 2252 24084 2261
rect 6884 2150 6936 2202
rect 6948 2150 7000 2202
rect 7012 2150 7064 2202
rect 7076 2150 7128 2202
rect 7140 2150 7192 2202
rect 12818 2150 12870 2202
rect 12882 2150 12934 2202
rect 12946 2150 12998 2202
rect 13010 2150 13062 2202
rect 13074 2150 13126 2202
rect 18752 2150 18804 2202
rect 18816 2150 18868 2202
rect 18880 2150 18932 2202
rect 18944 2150 18996 2202
rect 19008 2150 19060 2202
rect 24686 2150 24738 2202
rect 24750 2150 24802 2202
rect 24814 2150 24866 2202
rect 24878 2150 24930 2202
rect 24942 2150 24994 2202
rect 2320 2091 2372 2100
rect 2320 2057 2329 2091
rect 2329 2057 2363 2091
rect 2363 2057 2372 2091
rect 2320 2048 2372 2057
rect 756 1980 808 2032
rect 1768 1955 1820 1964
rect 1768 1921 1777 1955
rect 1777 1921 1811 1955
rect 1811 1921 1820 1955
rect 1768 1912 1820 1921
rect 2136 1955 2188 1964
rect 2136 1921 2145 1955
rect 2145 1921 2179 1955
rect 2179 1921 2188 1955
rect 2136 1912 2188 1921
rect 1032 1776 1084 1828
rect 1492 1751 1544 1760
rect 1492 1717 1501 1751
rect 1501 1717 1535 1751
rect 1535 1717 1544 1751
rect 1492 1708 1544 1717
rect 1952 1751 2004 1760
rect 1952 1717 1961 1751
rect 1961 1717 1995 1751
rect 1995 1717 2004 1751
rect 1952 1708 2004 1717
rect 3148 1955 3200 1964
rect 3148 1921 3157 1955
rect 3157 1921 3191 1955
rect 3191 1921 3200 1955
rect 3148 1912 3200 1921
rect 3608 1912 3660 1964
rect 3700 1955 3752 1964
rect 3700 1921 3709 1955
rect 3709 1921 3743 1955
rect 3743 1921 3752 1955
rect 3700 1912 3752 1921
rect 4160 1912 4212 1964
rect 3240 1844 3292 1896
rect 4712 1912 4764 1964
rect 4988 1912 5040 1964
rect 5448 1980 5500 2032
rect 5724 2048 5776 2100
rect 6828 2048 6880 2100
rect 7472 2048 7524 2100
rect 7564 2091 7616 2100
rect 7564 2057 7573 2091
rect 7573 2057 7607 2091
rect 7607 2057 7616 2091
rect 7564 2048 7616 2057
rect 7840 2091 7892 2100
rect 7840 2057 7849 2091
rect 7849 2057 7883 2091
rect 7883 2057 7892 2091
rect 7840 2048 7892 2057
rect 3056 1776 3108 1828
rect 4068 1819 4120 1828
rect 4068 1785 4077 1819
rect 4077 1785 4111 1819
rect 4111 1785 4120 1819
rect 4068 1776 4120 1785
rect 3424 1708 3476 1760
rect 3516 1751 3568 1760
rect 3516 1717 3525 1751
rect 3525 1717 3559 1751
rect 3559 1717 3568 1751
rect 3516 1708 3568 1717
rect 4252 1708 4304 1760
rect 6552 1912 6604 1964
rect 6644 1955 6696 1964
rect 6644 1921 6653 1955
rect 6653 1921 6687 1955
rect 6687 1921 6696 1955
rect 6644 1912 6696 1921
rect 6736 1912 6788 1964
rect 7380 1912 7432 1964
rect 7472 1955 7524 1964
rect 7472 1921 7481 1955
rect 7481 1921 7515 1955
rect 7515 1921 7524 1955
rect 7472 1912 7524 1921
rect 7748 1955 7800 1964
rect 7748 1921 7757 1955
rect 7757 1921 7791 1955
rect 7791 1921 7800 1955
rect 7748 1912 7800 1921
rect 8024 1955 8076 1964
rect 8024 1921 8033 1955
rect 8033 1921 8067 1955
rect 8067 1921 8076 1955
rect 8024 1912 8076 1921
rect 8484 1912 8536 1964
rect 8852 1955 8904 1964
rect 8852 1921 8861 1955
rect 8861 1921 8895 1955
rect 8895 1921 8904 1955
rect 8852 1912 8904 1921
rect 6276 1844 6328 1896
rect 9220 2091 9272 2100
rect 9220 2057 9229 2091
rect 9229 2057 9263 2091
rect 9263 2057 9272 2091
rect 9220 2048 9272 2057
rect 10876 2048 10928 2100
rect 9128 1955 9180 1964
rect 9128 1921 9137 1955
rect 9137 1921 9171 1955
rect 9171 1921 9180 1955
rect 9128 1912 9180 1921
rect 9220 1912 9272 1964
rect 9404 1955 9456 1964
rect 9404 1921 9413 1955
rect 9413 1921 9447 1955
rect 9447 1921 9456 1955
rect 9404 1912 9456 1921
rect 9772 1912 9824 1964
rect 10232 1955 10284 1964
rect 10232 1921 10241 1955
rect 10241 1921 10275 1955
rect 10275 1921 10284 1955
rect 10232 1912 10284 1921
rect 10324 1912 10376 1964
rect 11428 1980 11480 2032
rect 12716 1980 12768 2032
rect 11336 1912 11388 1964
rect 11612 1912 11664 1964
rect 12348 1912 12400 1964
rect 12808 1955 12860 1964
rect 12808 1921 12817 1955
rect 12817 1921 12851 1955
rect 12851 1921 12860 1955
rect 12808 1912 12860 1921
rect 14004 2048 14056 2100
rect 14188 2091 14240 2100
rect 14188 2057 14197 2091
rect 14197 2057 14231 2091
rect 14231 2057 14240 2091
rect 14188 2048 14240 2057
rect 14096 1955 14148 1964
rect 14096 1921 14105 1955
rect 14105 1921 14139 1955
rect 14139 1921 14148 1955
rect 14096 1912 14148 1921
rect 14372 1955 14424 1964
rect 14372 1921 14381 1955
rect 14381 1921 14415 1955
rect 14415 1921 14424 1955
rect 14372 1912 14424 1921
rect 15476 1980 15528 2032
rect 15384 1955 15436 1964
rect 15384 1921 15393 1955
rect 15393 1921 15427 1955
rect 15427 1921 15436 1955
rect 15384 1912 15436 1921
rect 17592 2048 17644 2100
rect 17868 2048 17920 2100
rect 17960 2048 18012 2100
rect 16028 1980 16080 2032
rect 16120 1912 16172 1964
rect 17776 1980 17828 2032
rect 18236 2048 18288 2100
rect 19156 2048 19208 2100
rect 19248 2048 19300 2100
rect 20352 2048 20404 2100
rect 20628 2048 20680 2100
rect 19340 1912 19392 1964
rect 20904 2091 20956 2100
rect 20904 2057 20913 2091
rect 20913 2057 20947 2091
rect 20947 2057 20956 2091
rect 20904 2048 20956 2057
rect 20996 2048 21048 2100
rect 21456 2091 21508 2100
rect 21456 2057 21465 2091
rect 21465 2057 21499 2091
rect 21499 2057 21508 2091
rect 21456 2048 21508 2057
rect 21640 2048 21692 2100
rect 22284 2091 22336 2100
rect 22284 2057 22293 2091
rect 22293 2057 22327 2091
rect 22327 2057 22336 2091
rect 22284 2048 22336 2057
rect 22652 2048 22704 2100
rect 23112 2048 23164 2100
rect 23204 2091 23256 2100
rect 23204 2057 23213 2091
rect 23213 2057 23247 2091
rect 23247 2057 23256 2091
rect 23204 2048 23256 2057
rect 23940 2048 23992 2100
rect 24032 2048 24084 2100
rect 5908 1819 5960 1828
rect 5908 1785 5917 1819
rect 5917 1785 5951 1819
rect 5951 1785 5960 1819
rect 5908 1776 5960 1785
rect 6368 1776 6420 1828
rect 5080 1708 5132 1760
rect 5172 1751 5224 1760
rect 5172 1717 5181 1751
rect 5181 1717 5215 1751
rect 5215 1717 5224 1751
rect 5172 1708 5224 1717
rect 5540 1708 5592 1760
rect 6000 1751 6052 1760
rect 6000 1717 6009 1751
rect 6009 1717 6043 1751
rect 6043 1717 6052 1751
rect 6000 1708 6052 1717
rect 6460 1751 6512 1760
rect 6460 1717 6469 1751
rect 6469 1717 6503 1751
rect 6503 1717 6512 1751
rect 6460 1708 6512 1717
rect 7840 1776 7892 1828
rect 7472 1708 7524 1760
rect 8024 1708 8076 1760
rect 8208 1708 8260 1760
rect 8668 1751 8720 1760
rect 8668 1717 8677 1751
rect 8677 1717 8711 1751
rect 8711 1717 8720 1751
rect 8668 1708 8720 1717
rect 8944 1776 8996 1828
rect 9496 1776 9548 1828
rect 10140 1776 10192 1828
rect 13176 1776 13228 1828
rect 14372 1776 14424 1828
rect 10508 1751 10560 1760
rect 10508 1717 10517 1751
rect 10517 1717 10551 1751
rect 10551 1717 10560 1751
rect 10508 1708 10560 1717
rect 11060 1751 11112 1760
rect 11060 1717 11069 1751
rect 11069 1717 11103 1751
rect 11103 1717 11112 1751
rect 11060 1708 11112 1717
rect 11704 1751 11756 1760
rect 11704 1717 11713 1751
rect 11713 1717 11747 1751
rect 11747 1717 11756 1751
rect 11704 1708 11756 1717
rect 11796 1708 11848 1760
rect 12440 1751 12492 1760
rect 12440 1717 12449 1751
rect 12449 1717 12483 1751
rect 12483 1717 12492 1751
rect 12440 1708 12492 1717
rect 12624 1708 12676 1760
rect 13544 1751 13596 1760
rect 13544 1717 13553 1751
rect 13553 1717 13587 1751
rect 13587 1717 13596 1751
rect 13544 1708 13596 1717
rect 14648 1751 14700 1760
rect 14648 1717 14657 1751
rect 14657 1717 14691 1751
rect 14691 1717 14700 1751
rect 14648 1708 14700 1717
rect 14740 1708 14792 1760
rect 15108 1708 15160 1760
rect 17776 1776 17828 1828
rect 19524 1776 19576 1828
rect 20444 1844 20496 1896
rect 21732 1912 21784 1964
rect 22100 1955 22152 1964
rect 22100 1921 22109 1955
rect 22109 1921 22143 1955
rect 22143 1921 22152 1955
rect 22100 1912 22152 1921
rect 23020 1955 23072 1964
rect 23020 1921 23029 1955
rect 23029 1921 23063 1955
rect 23063 1921 23072 1955
rect 23020 1912 23072 1921
rect 23388 1980 23440 2032
rect 15476 1751 15528 1760
rect 15476 1717 15485 1751
rect 15485 1717 15519 1751
rect 15519 1717 15528 1751
rect 15476 1708 15528 1717
rect 15660 1708 15712 1760
rect 16580 1708 16632 1760
rect 16764 1708 16816 1760
rect 17960 1708 18012 1760
rect 18236 1708 18288 1760
rect 19340 1708 19392 1760
rect 21456 1776 21508 1828
rect 24216 1776 24268 1828
rect 22376 1708 22428 1760
rect 23020 1708 23072 1760
rect 24124 1708 24176 1760
rect 3917 1606 3969 1658
rect 3981 1606 4033 1658
rect 4045 1606 4097 1658
rect 4109 1606 4161 1658
rect 4173 1606 4225 1658
rect 9851 1606 9903 1658
rect 9915 1606 9967 1658
rect 9979 1606 10031 1658
rect 10043 1606 10095 1658
rect 10107 1606 10159 1658
rect 15785 1606 15837 1658
rect 15849 1606 15901 1658
rect 15913 1606 15965 1658
rect 15977 1606 16029 1658
rect 16041 1606 16093 1658
rect 21719 1606 21771 1658
rect 21783 1606 21835 1658
rect 21847 1606 21899 1658
rect 21911 1606 21963 1658
rect 21975 1606 22027 1658
rect 2596 1547 2648 1556
rect 2596 1513 2605 1547
rect 2605 1513 2639 1547
rect 2639 1513 2648 1547
rect 2596 1504 2648 1513
rect 3240 1504 3292 1556
rect 2964 1436 3016 1488
rect 1492 1300 1544 1352
rect 3240 1368 3292 1420
rect 2780 1343 2832 1352
rect 2780 1309 2789 1343
rect 2789 1309 2823 1343
rect 2823 1309 2832 1343
rect 2780 1300 2832 1309
rect 3056 1343 3108 1352
rect 3056 1309 3065 1343
rect 3065 1309 3099 1343
rect 3099 1309 3108 1343
rect 3056 1300 3108 1309
rect 4436 1504 4488 1556
rect 6000 1504 6052 1556
rect 3516 1368 3568 1420
rect 3884 1300 3936 1352
rect 6368 1436 6420 1488
rect 7472 1504 7524 1556
rect 9220 1436 9272 1488
rect 9956 1504 10008 1556
rect 11428 1504 11480 1556
rect 12164 1504 12216 1556
rect 12440 1504 12492 1556
rect 13176 1504 13228 1556
rect 13820 1504 13872 1556
rect 15108 1504 15160 1556
rect 15384 1547 15436 1556
rect 15384 1513 15393 1547
rect 15393 1513 15427 1547
rect 15427 1513 15436 1547
rect 15384 1504 15436 1513
rect 15292 1436 15344 1488
rect 16120 1504 16172 1556
rect 16212 1504 16264 1556
rect 16488 1504 16540 1556
rect 1952 1207 2004 1216
rect 1952 1173 1961 1207
rect 1961 1173 1995 1207
rect 1995 1173 2004 1207
rect 1952 1164 2004 1173
rect 2044 1207 2096 1216
rect 2044 1173 2053 1207
rect 2053 1173 2087 1207
rect 2087 1173 2096 1207
rect 2044 1164 2096 1173
rect 2688 1232 2740 1284
rect 4804 1300 4856 1352
rect 5172 1300 5224 1352
rect 5540 1300 5592 1352
rect 6460 1300 6512 1352
rect 6828 1343 6880 1352
rect 6828 1309 6837 1343
rect 6837 1309 6871 1343
rect 6871 1309 6880 1343
rect 6828 1300 6880 1309
rect 2228 1164 2280 1216
rect 2320 1207 2372 1216
rect 2320 1173 2329 1207
rect 2329 1173 2363 1207
rect 2363 1173 2372 1207
rect 2320 1164 2372 1173
rect 3976 1164 4028 1216
rect 5264 1232 5316 1284
rect 7840 1300 7892 1352
rect 8576 1368 8628 1420
rect 8208 1343 8260 1352
rect 8208 1309 8217 1343
rect 8217 1309 8251 1343
rect 8251 1309 8260 1343
rect 8208 1300 8260 1309
rect 8668 1300 8720 1352
rect 8760 1343 8812 1352
rect 8760 1309 8769 1343
rect 8769 1309 8803 1343
rect 8803 1309 8812 1343
rect 8760 1300 8812 1309
rect 8944 1300 8996 1352
rect 4528 1164 4580 1216
rect 4712 1164 4764 1216
rect 5080 1207 5132 1216
rect 5080 1173 5089 1207
rect 5089 1173 5123 1207
rect 5123 1173 5132 1207
rect 5080 1164 5132 1173
rect 5172 1207 5224 1216
rect 5172 1173 5181 1207
rect 5181 1173 5215 1207
rect 5215 1173 5224 1207
rect 5172 1164 5224 1173
rect 5816 1164 5868 1216
rect 5908 1207 5960 1216
rect 5908 1173 5917 1207
rect 5917 1173 5951 1207
rect 5951 1173 5960 1207
rect 5908 1164 5960 1173
rect 6184 1207 6236 1216
rect 6184 1173 6193 1207
rect 6193 1173 6227 1207
rect 6227 1173 6236 1207
rect 6184 1164 6236 1173
rect 6368 1207 6420 1216
rect 6368 1173 6377 1207
rect 6377 1173 6411 1207
rect 6411 1173 6420 1207
rect 6368 1164 6420 1173
rect 7472 1207 7524 1216
rect 7472 1173 7481 1207
rect 7481 1173 7515 1207
rect 7515 1173 7524 1207
rect 7472 1164 7524 1173
rect 9956 1343 10008 1352
rect 9956 1309 9965 1343
rect 9965 1309 9999 1343
rect 9999 1309 10008 1343
rect 9956 1300 10008 1309
rect 10140 1300 10192 1352
rect 10508 1368 10560 1420
rect 10692 1368 10744 1420
rect 10876 1368 10928 1420
rect 11060 1411 11112 1420
rect 11060 1377 11069 1411
rect 11069 1377 11103 1411
rect 11103 1377 11112 1411
rect 11060 1368 11112 1377
rect 10600 1300 10652 1352
rect 8300 1207 8352 1216
rect 8300 1173 8309 1207
rect 8309 1173 8343 1207
rect 8343 1173 8352 1207
rect 8300 1164 8352 1173
rect 9128 1164 9180 1216
rect 9220 1207 9272 1216
rect 9220 1173 9229 1207
rect 9229 1173 9263 1207
rect 9263 1173 9272 1207
rect 9220 1164 9272 1173
rect 9680 1164 9732 1216
rect 10048 1164 10100 1216
rect 10692 1232 10744 1284
rect 10784 1275 10836 1284
rect 10784 1241 10793 1275
rect 10793 1241 10827 1275
rect 10827 1241 10836 1275
rect 10784 1232 10836 1241
rect 11612 1300 11664 1352
rect 11704 1343 11756 1352
rect 11704 1309 11713 1343
rect 11713 1309 11747 1343
rect 11747 1309 11756 1343
rect 11704 1300 11756 1309
rect 12256 1343 12308 1352
rect 12256 1309 12265 1343
rect 12265 1309 12299 1343
rect 12299 1309 12308 1343
rect 12256 1300 12308 1309
rect 13636 1368 13688 1420
rect 16304 1368 16356 1420
rect 17500 1504 17552 1556
rect 19800 1504 19852 1556
rect 21456 1547 21508 1556
rect 21456 1513 21465 1547
rect 21465 1513 21499 1547
rect 21499 1513 21508 1547
rect 21456 1504 21508 1513
rect 21640 1504 21692 1556
rect 23480 1504 23532 1556
rect 24676 1504 24728 1556
rect 17500 1368 17552 1420
rect 18696 1436 18748 1488
rect 18052 1368 18104 1420
rect 18604 1368 18656 1420
rect 21272 1436 21324 1488
rect 21088 1368 21140 1420
rect 11428 1164 11480 1216
rect 12348 1207 12400 1216
rect 12348 1173 12357 1207
rect 12357 1173 12391 1207
rect 12391 1173 12400 1207
rect 12348 1164 12400 1173
rect 13176 1300 13228 1352
rect 13268 1343 13320 1352
rect 13268 1309 13277 1343
rect 13277 1309 13311 1343
rect 13311 1309 13320 1343
rect 13268 1300 13320 1309
rect 14372 1300 14424 1352
rect 14648 1343 14700 1352
rect 14648 1309 14657 1343
rect 14657 1309 14691 1343
rect 14691 1309 14700 1343
rect 14648 1300 14700 1309
rect 14924 1300 14976 1352
rect 15384 1300 15436 1352
rect 15476 1300 15528 1352
rect 16120 1300 16172 1352
rect 16580 1300 16632 1352
rect 16856 1300 16908 1352
rect 12716 1164 12768 1216
rect 13084 1207 13136 1216
rect 13084 1173 13093 1207
rect 13093 1173 13127 1207
rect 13127 1173 13136 1207
rect 13084 1164 13136 1173
rect 13452 1207 13504 1216
rect 13452 1173 13461 1207
rect 13461 1173 13495 1207
rect 13495 1173 13504 1207
rect 13452 1164 13504 1173
rect 14004 1164 14056 1216
rect 14924 1164 14976 1216
rect 17408 1232 17460 1284
rect 16488 1164 16540 1216
rect 19984 1300 20036 1352
rect 21180 1300 21232 1352
rect 21824 1300 21876 1352
rect 22744 1368 22796 1420
rect 19708 1232 19760 1284
rect 20628 1232 20680 1284
rect 22652 1343 22704 1352
rect 22652 1309 22661 1343
rect 22661 1309 22695 1343
rect 22695 1309 22704 1343
rect 22652 1300 22704 1309
rect 23480 1343 23532 1352
rect 23480 1309 23489 1343
rect 23489 1309 23523 1343
rect 23523 1309 23532 1343
rect 23480 1300 23532 1309
rect 24676 1368 24728 1420
rect 25596 1368 25648 1420
rect 24032 1343 24084 1352
rect 24032 1309 24041 1343
rect 24041 1309 24075 1343
rect 24075 1309 24084 1343
rect 24032 1300 24084 1309
rect 19432 1164 19484 1216
rect 20076 1164 20128 1216
rect 22008 1164 22060 1216
rect 23572 1232 23624 1284
rect 22284 1207 22336 1216
rect 22284 1173 22293 1207
rect 22293 1173 22327 1207
rect 22327 1173 22336 1207
rect 22284 1164 22336 1173
rect 22560 1207 22612 1216
rect 22560 1173 22569 1207
rect 22569 1173 22603 1207
rect 22603 1173 22612 1207
rect 22560 1164 22612 1173
rect 22744 1164 22796 1216
rect 23112 1207 23164 1216
rect 23112 1173 23121 1207
rect 23121 1173 23155 1207
rect 23155 1173 23164 1207
rect 23112 1164 23164 1173
rect 23296 1164 23348 1216
rect 23940 1207 23992 1216
rect 23940 1173 23949 1207
rect 23949 1173 23983 1207
rect 23983 1173 23992 1207
rect 23940 1164 23992 1173
rect 24216 1207 24268 1216
rect 24216 1173 24225 1207
rect 24225 1173 24259 1207
rect 24259 1173 24268 1207
rect 24216 1164 24268 1173
rect 6884 1062 6936 1114
rect 6948 1062 7000 1114
rect 7012 1062 7064 1114
rect 7076 1062 7128 1114
rect 7140 1062 7192 1114
rect 12818 1062 12870 1114
rect 12882 1062 12934 1114
rect 12946 1062 12998 1114
rect 13010 1062 13062 1114
rect 13074 1062 13126 1114
rect 18752 1062 18804 1114
rect 18816 1062 18868 1114
rect 18880 1062 18932 1114
rect 18944 1062 18996 1114
rect 19008 1062 19060 1114
rect 24686 1062 24738 1114
rect 24750 1062 24802 1114
rect 24814 1062 24866 1114
rect 24878 1062 24930 1114
rect 24942 1062 24994 1114
rect 2044 960 2096 1012
rect 2320 960 2372 1012
rect 3332 960 3384 1012
rect 5264 960 5316 1012
rect 9220 960 9272 1012
rect 13636 960 13688 1012
rect 16672 960 16724 1012
rect 17408 960 17460 1012
rect 5724 892 5776 944
rect 6000 892 6052 944
rect 10784 892 10836 944
rect 11244 892 11296 944
rect 14924 892 14976 944
rect 15016 892 15068 944
rect 22284 960 22336 1012
rect 22560 960 22612 1012
rect 23296 960 23348 1012
rect 2780 688 2832 740
rect 3516 688 3568 740
rect 4528 756 4580 808
rect 7840 824 7892 876
rect 8300 824 8352 876
rect 9680 824 9732 876
rect 6368 756 6420 808
rect 7472 756 7524 808
rect 4804 688 4856 740
rect 5540 688 5592 740
rect 5172 620 5224 672
rect 9128 756 9180 808
rect 9772 756 9824 808
rect 13636 824 13688 876
rect 14648 756 14700 808
rect 22744 824 22796 876
rect 8852 688 8904 740
rect 9680 688 9732 740
rect 16948 620 17000 672
rect 9956 552 10008 604
rect 13912 552 13964 604
rect 21272 688 21324 740
rect 22652 688 22704 740
rect 21456 620 21508 672
rect 22008 620 22060 672
rect 23480 688 23532 740
rect 11612 484 11664 536
rect 13360 484 13412 536
rect 22008 484 22060 536
rect 24216 552 24268 604
rect 10140 416 10192 468
rect 4712 348 4764 400
rect 7840 348 7892 400
rect 8024 348 8076 400
rect 16120 416 16172 468
rect 16396 416 16448 468
rect 23112 416 23164 468
rect 12532 348 12584 400
rect 11336 280 11388 332
rect 22744 280 22796 332
rect 24032 280 24084 332
rect 3976 212 4028 264
rect 10232 144 10284 196
<< metal2 >>
rect 938 7970 994 8000
rect 938 7942 1440 7970
rect 938 7840 994 7942
rect 1412 6390 1440 7942
rect 2134 7840 2190 8000
rect 3330 7970 3386 8000
rect 4526 7970 4582 8000
rect 5722 7970 5778 8000
rect 6918 7970 6974 8000
rect 8114 7970 8170 8000
rect 9310 7970 9366 8000
rect 10506 7970 10562 8000
rect 11702 7970 11758 8000
rect 12898 7970 12954 8000
rect 14094 7970 14150 8000
rect 15290 7970 15346 8000
rect 16486 7970 16542 8000
rect 17682 7970 17738 8000
rect 18878 7970 18934 8000
rect 20074 7970 20130 8000
rect 21270 7970 21326 8000
rect 22466 7970 22522 8000
rect 3330 7942 3832 7970
rect 3330 7840 3386 7942
rect 2148 6458 2176 7840
rect 3804 6458 3832 7942
rect 4526 7942 4660 7970
rect 4526 7840 4582 7942
rect 4632 6458 4660 7942
rect 5722 7942 6132 7970
rect 5722 7840 5778 7942
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 6104 6390 6132 7942
rect 6918 7942 7328 7970
rect 6918 7840 6974 7942
rect 6884 6556 7192 6565
rect 6884 6554 6890 6556
rect 6946 6554 6970 6556
rect 7026 6554 7050 6556
rect 7106 6554 7130 6556
rect 7186 6554 7192 6556
rect 6946 6502 6948 6554
rect 7128 6502 7130 6554
rect 6884 6500 6890 6502
rect 6946 6500 6970 6502
rect 7026 6500 7050 6502
rect 7106 6500 7130 6502
rect 7186 6500 7192 6502
rect 6884 6491 7192 6500
rect 7300 6458 7328 7942
rect 8114 7942 8432 7970
rect 8114 7840 8170 7942
rect 8404 6458 8432 7942
rect 9310 7942 9444 7970
rect 9310 7840 9366 7942
rect 9416 6458 9444 7942
rect 10506 7942 10640 7970
rect 10506 7840 10562 7942
rect 10612 6458 10640 7942
rect 11702 7942 12020 7970
rect 11702 7840 11758 7942
rect 11992 6458 12020 7942
rect 12898 7942 13216 7970
rect 12898 7840 12954 7942
rect 12818 6556 13126 6565
rect 12818 6554 12824 6556
rect 12880 6554 12904 6556
rect 12960 6554 12984 6556
rect 13040 6554 13064 6556
rect 13120 6554 13126 6556
rect 12880 6502 12882 6554
rect 13062 6502 13064 6554
rect 12818 6500 12824 6502
rect 12880 6500 12904 6502
rect 12960 6500 12984 6502
rect 13040 6500 13064 6502
rect 13120 6500 13126 6502
rect 12818 6491 13126 6500
rect 13188 6458 13216 7942
rect 14094 7942 14320 7970
rect 14094 7840 14150 7942
rect 14292 6458 14320 7942
rect 15290 7942 15424 7970
rect 15290 7840 15346 7942
rect 15396 6458 15424 7942
rect 16486 7942 16896 7970
rect 16486 7840 16542 7942
rect 16868 6458 16896 7942
rect 17682 7942 17816 7970
rect 17682 7840 17738 7942
rect 17788 6458 17816 7942
rect 18878 7942 19472 7970
rect 18878 7840 18934 7942
rect 18752 6556 19060 6565
rect 18752 6554 18758 6556
rect 18814 6554 18838 6556
rect 18894 6554 18918 6556
rect 18974 6554 18998 6556
rect 19054 6554 19060 6556
rect 18814 6502 18816 6554
rect 18996 6502 18998 6554
rect 18752 6500 18758 6502
rect 18814 6500 18838 6502
rect 18894 6500 18918 6502
rect 18974 6500 18998 6502
rect 19054 6500 19060 6502
rect 18752 6491 19060 6500
rect 19444 6458 19472 7942
rect 20074 7942 20392 7970
rect 20074 7840 20130 7942
rect 20364 6458 20392 7942
rect 21270 7942 21588 7970
rect 21270 7840 21326 7942
rect 21560 6458 21588 7942
rect 22466 7942 22600 7970
rect 22466 7840 22522 7942
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 1400 6384 1452 6390
rect 5632 6384 5684 6390
rect 1400 6326 1452 6332
rect 2226 6352 2282 6361
rect 5632 6326 5684 6332
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 2226 6287 2228 6296
rect 2280 6287 2282 6296
rect 2228 6258 2280 6264
rect 5644 6186 5672 6326
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 3917 6012 4225 6021
rect 3917 6010 3923 6012
rect 3979 6010 4003 6012
rect 4059 6010 4083 6012
rect 4139 6010 4163 6012
rect 4219 6010 4225 6012
rect 3979 5958 3981 6010
rect 4161 5958 4163 6010
rect 3917 5956 3923 5958
rect 3979 5956 4003 5958
rect 4059 5956 4083 5958
rect 4139 5956 4163 5958
rect 4219 5956 4225 5958
rect 3917 5947 4225 5956
rect 6564 5914 6592 6258
rect 7576 5914 7604 6258
rect 8772 5914 8800 6258
rect 9692 5914 9720 6258
rect 9851 6012 10159 6021
rect 9851 6010 9857 6012
rect 9913 6010 9937 6012
rect 9993 6010 10017 6012
rect 10073 6010 10097 6012
rect 10153 6010 10159 6012
rect 9913 5958 9915 6010
rect 10095 5958 10097 6010
rect 9851 5956 9857 5958
rect 9913 5956 9937 5958
rect 9993 5956 10017 5958
rect 10073 5956 10097 5958
rect 10153 5956 10159 5958
rect 9851 5947 10159 5956
rect 11164 5914 11192 6258
rect 12360 5914 12388 6258
rect 12636 5914 12664 6258
rect 13556 5914 13584 6258
rect 14660 5914 14688 6258
rect 15120 5914 15148 6258
rect 15672 5914 15700 6258
rect 15785 6012 16093 6021
rect 15785 6010 15791 6012
rect 15847 6010 15871 6012
rect 15927 6010 15951 6012
rect 16007 6010 16031 6012
rect 16087 6010 16093 6012
rect 15847 5958 15849 6010
rect 16029 5958 16031 6010
rect 15785 5956 15791 5958
rect 15847 5956 15871 5958
rect 15927 5956 15951 5958
rect 16007 5956 16031 5958
rect 16087 5956 16093 5958
rect 15785 5947 16093 5956
rect 17420 5914 17448 6258
rect 18340 5914 18368 6258
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 19996 5846 20024 6258
rect 20548 5914 20576 6258
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 6288 5370 6316 5646
rect 6884 5468 7192 5477
rect 6884 5466 6890 5468
rect 6946 5466 6970 5468
rect 7026 5466 7050 5468
rect 7106 5466 7130 5468
rect 7186 5466 7192 5468
rect 6946 5414 6948 5466
rect 7128 5414 7130 5466
rect 6884 5412 6890 5414
rect 6946 5412 6970 5414
rect 7026 5412 7050 5414
rect 7106 5412 7130 5414
rect 7186 5412 7192 5414
rect 6884 5403 7192 5412
rect 7576 5370 7604 5646
rect 8772 5370 8800 5646
rect 9876 5370 9904 5646
rect 11072 5370 11100 5646
rect 11992 5370 12020 5646
rect 12452 5370 12480 5646
rect 12818 5468 13126 5477
rect 12818 5466 12824 5468
rect 12880 5466 12904 5468
rect 12960 5466 12984 5468
rect 13040 5466 13064 5468
rect 13120 5466 13126 5468
rect 12880 5414 12882 5466
rect 13062 5414 13064 5466
rect 12818 5412 12824 5414
rect 12880 5412 12904 5414
rect 12960 5412 12984 5414
rect 13040 5412 13064 5414
rect 13120 5412 13126 5414
rect 12818 5403 13126 5412
rect 13464 5370 13492 5646
rect 14568 5370 14596 5646
rect 14844 5370 14872 5646
rect 15948 5370 15976 5646
rect 17144 5370 17172 5646
rect 18432 5370 18460 5646
rect 18752 5468 19060 5477
rect 18752 5466 18758 5468
rect 18814 5466 18838 5468
rect 18894 5466 18918 5468
rect 18974 5466 18998 5468
rect 19054 5466 19060 5468
rect 18814 5414 18816 5466
rect 18996 5414 18998 5466
rect 18752 5412 18758 5414
rect 18814 5412 18838 5414
rect 18894 5412 18918 5414
rect 18974 5412 18998 5414
rect 19054 5412 19060 5414
rect 18752 5403 19060 5412
rect 19996 5370 20024 5646
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 13912 5296 13964 5302
rect 13912 5238 13964 5244
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 3917 4924 4225 4933
rect 3917 4922 3923 4924
rect 3979 4922 4003 4924
rect 4059 4922 4083 4924
rect 4139 4922 4163 4924
rect 4219 4922 4225 4924
rect 3979 4870 3981 4922
rect 4161 4870 4163 4922
rect 3917 4868 3923 4870
rect 3979 4868 4003 4870
rect 4059 4868 4083 4870
rect 4139 4868 4163 4870
rect 4219 4868 4225 4870
rect 3917 4859 4225 4868
rect 6564 4826 6592 5170
rect 9588 5160 9640 5166
rect 9586 5128 9588 5137
rect 9640 5128 9642 5137
rect 9586 5063 9642 5072
rect 9851 4924 10159 4933
rect 9851 4922 9857 4924
rect 9913 4922 9937 4924
rect 9993 4922 10017 4924
rect 10073 4922 10097 4924
rect 10153 4922 10159 4924
rect 9913 4870 9915 4922
rect 10095 4870 10097 4922
rect 9851 4868 9857 4870
rect 9913 4868 9937 4870
rect 9993 4868 10017 4870
rect 10073 4868 10097 4870
rect 10153 4868 10159 4870
rect 9851 4859 10159 4868
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6884 4380 7192 4389
rect 6884 4378 6890 4380
rect 6946 4378 6970 4380
rect 7026 4378 7050 4380
rect 7106 4378 7130 4380
rect 7186 4378 7192 4380
rect 6946 4326 6948 4378
rect 7128 4326 7130 4378
rect 6884 4324 6890 4326
rect 6946 4324 6970 4326
rect 7026 4324 7050 4326
rect 7106 4324 7130 4326
rect 7186 4324 7192 4326
rect 6884 4315 7192 4324
rect 11256 4185 11284 5170
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 11242 4176 11298 4185
rect 11242 4111 11298 4120
rect 3917 3836 4225 3845
rect 3917 3834 3923 3836
rect 3979 3834 4003 3836
rect 4059 3834 4083 3836
rect 4139 3834 4163 3836
rect 4219 3834 4225 3836
rect 3979 3782 3981 3834
rect 4161 3782 4163 3834
rect 3917 3780 3923 3782
rect 3979 3780 4003 3782
rect 4059 3780 4083 3782
rect 4139 3780 4163 3782
rect 4219 3780 4225 3782
rect 3917 3771 4225 3780
rect 9851 3836 10159 3845
rect 9851 3834 9857 3836
rect 9913 3834 9937 3836
rect 9993 3834 10017 3836
rect 10073 3834 10097 3836
rect 10153 3834 10159 3836
rect 9913 3782 9915 3834
rect 10095 3782 10097 3834
rect 9851 3780 9857 3782
rect 9913 3780 9937 3782
rect 9993 3780 10017 3782
rect 10073 3780 10097 3782
rect 10153 3780 10159 3782
rect 9851 3771 10159 3780
rect 6884 3292 7192 3301
rect 6884 3290 6890 3292
rect 6946 3290 6970 3292
rect 7026 3290 7050 3292
rect 7106 3290 7130 3292
rect 7186 3290 7192 3292
rect 6946 3238 6948 3290
rect 7128 3238 7130 3290
rect 6884 3236 6890 3238
rect 6946 3236 6970 3238
rect 7026 3236 7050 3238
rect 7106 3236 7130 3238
rect 7186 3236 7192 3238
rect 6884 3227 7192 3236
rect 7470 3088 7526 3097
rect 7470 3023 7526 3032
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1596 2650 1624 2926
rect 3917 2748 4225 2757
rect 3917 2746 3923 2748
rect 3979 2746 4003 2748
rect 4059 2746 4083 2748
rect 4139 2746 4163 2748
rect 4219 2746 4225 2748
rect 3979 2694 3981 2746
rect 4161 2694 4163 2746
rect 3917 2692 3923 2694
rect 3979 2692 4003 2694
rect 4059 2692 4083 2694
rect 4139 2692 4163 2694
rect 4219 2692 4225 2694
rect 3917 2683 4225 2692
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 480 2508 532 2514
rect 480 2450 532 2456
rect 204 2372 256 2378
rect 204 2314 256 2320
rect 216 160 244 2314
rect 492 160 520 2450
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 756 2032 808 2038
rect 756 1974 808 1980
rect 768 160 796 1974
rect 1032 1828 1084 1834
rect 1032 1770 1084 1776
rect 1044 160 1072 1770
rect 1320 160 1348 2382
rect 1860 2304 1912 2310
rect 1860 2246 1912 2252
rect 2412 2304 2464 2310
rect 2412 2246 2464 2252
rect 1768 1964 1820 1970
rect 1768 1906 1820 1912
rect 1492 1760 1544 1766
rect 1492 1702 1544 1708
rect 1504 1358 1532 1702
rect 1492 1352 1544 1358
rect 1492 1294 1544 1300
rect 202 0 258 160
rect 478 0 534 160
rect 754 0 810 160
rect 1030 0 1086 160
rect 1306 0 1362 160
rect 1582 82 1638 160
rect 1780 82 1808 1906
rect 1872 160 1900 2246
rect 2320 2100 2372 2106
rect 2320 2042 2372 2048
rect 2136 1964 2188 1970
rect 2136 1906 2188 1912
rect 1952 1760 2004 1766
rect 1950 1728 1952 1737
rect 2004 1728 2006 1737
rect 1950 1663 2006 1672
rect 1952 1216 2004 1222
rect 1952 1158 2004 1164
rect 2044 1216 2096 1222
rect 2044 1158 2096 1164
rect 1964 377 1992 1158
rect 2056 1018 2084 1158
rect 2044 1012 2096 1018
rect 2044 954 2096 960
rect 1950 368 2006 377
rect 1950 303 2006 312
rect 2148 160 2176 1906
rect 2332 1329 2360 2042
rect 2424 2009 2452 2246
rect 2410 2000 2466 2009
rect 2410 1935 2466 1944
rect 2608 1562 2636 2586
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 6276 2576 6328 2582
rect 7196 2576 7248 2582
rect 6276 2518 6328 2524
rect 7194 2544 7196 2553
rect 7248 2544 7250 2553
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 3148 1964 3200 1970
rect 3148 1906 3200 1912
rect 3056 1828 3108 1834
rect 3056 1770 3108 1776
rect 2596 1556 2648 1562
rect 2596 1498 2648 1504
rect 2964 1488 3016 1494
rect 2962 1456 2964 1465
rect 3016 1456 3018 1465
rect 2962 1391 3018 1400
rect 3068 1358 3096 1770
rect 2780 1352 2832 1358
rect 2318 1320 2374 1329
rect 2780 1294 2832 1300
rect 3056 1352 3108 1358
rect 3056 1294 3108 1300
rect 2318 1255 2374 1264
rect 2688 1284 2740 1290
rect 2688 1226 2740 1232
rect 2228 1216 2280 1222
rect 2228 1158 2280 1164
rect 2320 1216 2372 1222
rect 2320 1158 2372 1164
rect 1582 54 1808 82
rect 1582 0 1638 54
rect 1858 0 1914 160
rect 2134 0 2190 160
rect 2240 82 2268 1158
rect 2332 1018 2360 1158
rect 2320 1012 2372 1018
rect 2320 954 2372 960
rect 2700 160 2728 1226
rect 2792 746 2820 1294
rect 2780 740 2832 746
rect 2780 682 2832 688
rect 2410 82 2466 160
rect 2240 54 2466 82
rect 2410 0 2466 54
rect 2686 0 2742 160
rect 2962 82 3018 160
rect 3160 82 3188 1906
rect 3240 1896 3292 1902
rect 3240 1838 3292 1844
rect 3252 1562 3280 1838
rect 3240 1556 3292 1562
rect 3240 1498 3292 1504
rect 3240 1420 3292 1426
rect 3240 1362 3292 1368
rect 3252 160 3280 1362
rect 3344 1018 3372 2314
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 1766 3464 2246
rect 3608 1964 3660 1970
rect 3608 1906 3660 1912
rect 3700 1964 3752 1970
rect 3700 1906 3752 1912
rect 3424 1760 3476 1766
rect 3424 1702 3476 1708
rect 3516 1760 3568 1766
rect 3516 1702 3568 1708
rect 3528 1426 3556 1702
rect 3516 1420 3568 1426
rect 3516 1362 3568 1368
rect 3332 1012 3384 1018
rect 3332 954 3384 960
rect 3516 740 3568 746
rect 3516 682 3568 688
rect 3528 160 3556 682
rect 2962 54 3188 82
rect 2962 0 3018 54
rect 3238 0 3294 160
rect 3514 0 3570 160
rect 3620 82 3648 1906
rect 3712 218 3740 1906
rect 4080 1834 4108 2450
rect 4896 2440 4948 2446
rect 4632 2400 4896 2428
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4160 1964 4212 1970
rect 4212 1924 4384 1952
rect 4160 1906 4212 1912
rect 4068 1828 4120 1834
rect 4068 1770 4120 1776
rect 4252 1760 4304 1766
rect 4252 1702 4304 1708
rect 3917 1660 4225 1669
rect 3917 1658 3923 1660
rect 3979 1658 4003 1660
rect 4059 1658 4083 1660
rect 4139 1658 4163 1660
rect 4219 1658 4225 1660
rect 3979 1606 3981 1658
rect 4161 1606 4163 1658
rect 3917 1604 3923 1606
rect 3979 1604 4003 1606
rect 4059 1604 4083 1606
rect 4139 1604 4163 1606
rect 4219 1604 4225 1606
rect 3917 1595 4225 1604
rect 3884 1352 3936 1358
rect 4264 1306 4292 1702
rect 3936 1300 4292 1306
rect 3884 1294 4292 1300
rect 3896 1278 4292 1294
rect 3976 1216 4028 1222
rect 3976 1158 4028 1164
rect 3988 270 4016 1158
rect 3976 264 4028 270
rect 3712 190 3924 218
rect 3976 206 4028 212
rect 3790 82 3846 160
rect 3620 54 3846 82
rect 3896 82 3924 190
rect 4356 160 4384 1924
rect 4448 1562 4476 2246
rect 4436 1556 4488 1562
rect 4436 1498 4488 1504
rect 4528 1216 4580 1222
rect 4528 1158 4580 1164
rect 4540 814 4568 1158
rect 4528 808 4580 814
rect 4528 750 4580 756
rect 4632 160 4660 2400
rect 4896 2382 4948 2388
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 4712 1964 4764 1970
rect 4988 1964 5040 1970
rect 4764 1924 4936 1952
rect 4712 1906 4764 1912
rect 4804 1352 4856 1358
rect 4804 1294 4856 1300
rect 4712 1216 4764 1222
rect 4712 1158 4764 1164
rect 4724 406 4752 1158
rect 4816 746 4844 1294
rect 4804 740 4856 746
rect 4804 682 4856 688
rect 4712 400 4764 406
rect 4712 342 4764 348
rect 4908 160 4936 1924
rect 4988 1906 5040 1912
rect 4066 82 4122 160
rect 3896 54 4122 82
rect 3790 0 3846 54
rect 4066 0 4122 54
rect 4342 0 4398 160
rect 4618 0 4674 160
rect 4894 0 4950 160
rect 5000 82 5028 1906
rect 5092 1766 5120 2246
rect 5736 2106 5764 2518
rect 6092 2440 6144 2446
rect 6288 2417 6316 2518
rect 7194 2479 7250 2488
rect 7380 2440 7432 2446
rect 6092 2382 6144 2388
rect 6274 2408 6330 2417
rect 5724 2100 5776 2106
rect 5724 2042 5776 2048
rect 5448 2032 5500 2038
rect 5448 1974 5500 1980
rect 5080 1760 5132 1766
rect 5080 1702 5132 1708
rect 5172 1760 5224 1766
rect 5172 1702 5224 1708
rect 5184 1358 5212 1702
rect 5172 1352 5224 1358
rect 5078 1320 5134 1329
rect 5172 1294 5224 1300
rect 5078 1255 5134 1264
rect 5264 1284 5316 1290
rect 5092 1222 5120 1255
rect 5264 1226 5316 1232
rect 5080 1216 5132 1222
rect 5080 1158 5132 1164
rect 5172 1216 5224 1222
rect 5172 1158 5224 1164
rect 5184 678 5212 1158
rect 5276 1018 5304 1226
rect 5264 1012 5316 1018
rect 5264 954 5316 960
rect 5172 672 5224 678
rect 5172 614 5224 620
rect 5460 160 5488 1974
rect 5906 1864 5962 1873
rect 5906 1799 5908 1808
rect 5960 1799 5962 1808
rect 5908 1770 5960 1776
rect 5540 1760 5592 1766
rect 5540 1702 5592 1708
rect 6000 1760 6052 1766
rect 6000 1702 6052 1708
rect 5552 1358 5580 1702
rect 6012 1562 6040 1702
rect 6000 1556 6052 1562
rect 6000 1498 6052 1504
rect 5540 1352 5592 1358
rect 5540 1294 5592 1300
rect 5828 1278 6040 1306
rect 5828 1222 5856 1278
rect 5816 1216 5868 1222
rect 5816 1158 5868 1164
rect 5908 1216 5960 1222
rect 5908 1158 5960 1164
rect 5724 944 5776 950
rect 5776 892 5856 898
rect 5724 886 5856 892
rect 5736 870 5856 886
rect 5540 740 5592 746
rect 5540 682 5592 688
rect 5552 626 5580 682
rect 5552 598 5764 626
rect 5736 160 5764 598
rect 5828 354 5856 870
rect 5920 785 5948 1158
rect 6012 950 6040 1278
rect 6000 944 6052 950
rect 6000 886 6052 892
rect 5906 776 5962 785
rect 5906 711 5962 720
rect 6104 490 6132 2382
rect 7300 2400 7380 2428
rect 6274 2343 6330 2352
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 6748 1970 6776 2314
rect 6884 2204 7192 2213
rect 6884 2202 6890 2204
rect 6946 2202 6970 2204
rect 7026 2202 7050 2204
rect 7106 2202 7130 2204
rect 7186 2202 7192 2204
rect 6946 2150 6948 2202
rect 7128 2150 7130 2202
rect 6884 2148 6890 2150
rect 6946 2148 6970 2150
rect 7026 2148 7050 2150
rect 7106 2148 7130 2150
rect 7186 2148 7192 2150
rect 6884 2139 7192 2148
rect 6828 2100 6880 2106
rect 6828 2042 6880 2048
rect 6552 1964 6604 1970
rect 6552 1906 6604 1912
rect 6644 1964 6696 1970
rect 6644 1906 6696 1912
rect 6736 1964 6788 1970
rect 6736 1906 6788 1912
rect 6276 1896 6328 1902
rect 6276 1838 6328 1844
rect 6184 1216 6236 1222
rect 6184 1158 6236 1164
rect 6196 649 6224 1158
rect 6182 640 6238 649
rect 6182 575 6238 584
rect 6012 462 6132 490
rect 5906 368 5962 377
rect 5828 326 5906 354
rect 5906 303 5962 312
rect 6012 160 6040 462
rect 6288 160 6316 1838
rect 6368 1828 6420 1834
rect 6368 1770 6420 1776
rect 6380 1494 6408 1770
rect 6460 1760 6512 1766
rect 6460 1702 6512 1708
rect 6368 1488 6420 1494
rect 6368 1430 6420 1436
rect 6472 1358 6500 1702
rect 6460 1352 6512 1358
rect 6460 1294 6512 1300
rect 6368 1216 6420 1222
rect 6368 1158 6420 1164
rect 6380 814 6408 1158
rect 6368 808 6420 814
rect 6368 750 6420 756
rect 6564 160 6592 1906
rect 6656 1000 6684 1906
rect 6840 1358 6868 2042
rect 6828 1352 6880 1358
rect 6828 1294 6880 1300
rect 6884 1116 7192 1125
rect 6884 1114 6890 1116
rect 6946 1114 6970 1116
rect 7026 1114 7050 1116
rect 7106 1114 7130 1116
rect 7186 1114 7192 1116
rect 6946 1062 6948 1114
rect 7128 1062 7130 1114
rect 6884 1060 6890 1062
rect 6946 1060 6970 1062
rect 7026 1060 7050 1062
rect 7106 1060 7130 1062
rect 7186 1060 7192 1062
rect 6884 1051 7192 1060
rect 7300 1000 7328 2400
rect 7380 2382 7432 2388
rect 7484 2106 7512 3023
rect 9034 2952 9090 2961
rect 9034 2887 9090 2896
rect 12254 2952 12310 2961
rect 12254 2887 12310 2896
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7576 2106 7604 2518
rect 9048 2514 9076 2887
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 7838 2272 7894 2281
rect 7838 2207 7894 2216
rect 7852 2106 7880 2207
rect 8298 2136 8354 2145
rect 7472 2100 7524 2106
rect 7472 2042 7524 2048
rect 7564 2100 7616 2106
rect 7564 2042 7616 2048
rect 7840 2100 7892 2106
rect 8298 2071 8354 2080
rect 7840 2042 7892 2048
rect 7380 1964 7432 1970
rect 7380 1906 7432 1912
rect 7472 1964 7524 1970
rect 7748 1964 7800 1970
rect 7524 1924 7696 1952
rect 7472 1906 7524 1912
rect 6656 972 6868 1000
rect 6840 160 6868 972
rect 7116 972 7328 1000
rect 7116 160 7144 972
rect 7392 160 7420 1906
rect 7472 1760 7524 1766
rect 7472 1702 7524 1708
rect 7484 1562 7512 1702
rect 7472 1556 7524 1562
rect 7472 1498 7524 1504
rect 7472 1216 7524 1222
rect 7472 1158 7524 1164
rect 7484 814 7512 1158
rect 7472 808 7524 814
rect 7472 750 7524 756
rect 7668 160 7696 1924
rect 8024 1964 8076 1970
rect 7800 1924 7972 1952
rect 7748 1906 7800 1912
rect 7840 1828 7892 1834
rect 7840 1770 7892 1776
rect 7852 1358 7880 1770
rect 7840 1352 7892 1358
rect 7840 1294 7892 1300
rect 7838 1184 7894 1193
rect 7838 1119 7894 1128
rect 7852 882 7880 1119
rect 7840 876 7892 882
rect 7840 818 7892 824
rect 7838 504 7894 513
rect 7838 439 7894 448
rect 7852 406 7880 439
rect 7840 400 7892 406
rect 7840 342 7892 348
rect 7944 160 7972 1924
rect 8076 1924 8156 1952
rect 8024 1906 8076 1912
rect 8024 1760 8076 1766
rect 8024 1702 8076 1708
rect 8036 406 8064 1702
rect 8128 1000 8156 1924
rect 8208 1760 8260 1766
rect 8312 1737 8340 2071
rect 9140 1970 9168 2586
rect 9508 2514 9536 2790
rect 9851 2748 10159 2757
rect 9851 2746 9857 2748
rect 9913 2746 9937 2748
rect 9993 2746 10017 2748
rect 10073 2746 10097 2748
rect 10153 2746 10159 2748
rect 9913 2694 9915 2746
rect 10095 2694 10097 2746
rect 9851 2692 9857 2694
rect 9913 2692 9937 2694
rect 9993 2692 10017 2694
rect 10073 2692 10097 2694
rect 10153 2692 10159 2694
rect 9851 2683 10159 2692
rect 10230 2680 10286 2689
rect 10230 2615 10286 2624
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9312 2440 9364 2446
rect 9864 2440 9916 2446
rect 9312 2382 9364 2388
rect 9692 2400 9864 2428
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 9232 2106 9260 2314
rect 9220 2100 9272 2106
rect 9220 2042 9272 2048
rect 8484 1964 8536 1970
rect 8484 1906 8536 1912
rect 8852 1964 8904 1970
rect 9128 1964 9180 1970
rect 8904 1924 9076 1952
rect 8852 1906 8904 1912
rect 8208 1702 8260 1708
rect 8298 1728 8354 1737
rect 8220 1358 8248 1702
rect 8298 1663 8354 1672
rect 8208 1352 8260 1358
rect 8208 1294 8260 1300
rect 8300 1216 8352 1222
rect 8300 1158 8352 1164
rect 8128 972 8248 1000
rect 8024 400 8076 406
rect 8024 342 8076 348
rect 8220 160 8248 972
rect 8312 882 8340 1158
rect 8300 876 8352 882
rect 8300 818 8352 824
rect 8496 160 8524 1906
rect 8944 1828 8996 1834
rect 8944 1770 8996 1776
rect 8668 1760 8720 1766
rect 8668 1702 8720 1708
rect 8576 1420 8628 1426
rect 8576 1362 8628 1368
rect 8588 762 8616 1362
rect 8680 1358 8708 1702
rect 8956 1358 8984 1770
rect 8668 1352 8720 1358
rect 8668 1294 8720 1300
rect 8760 1352 8812 1358
rect 8760 1294 8812 1300
rect 8944 1352 8996 1358
rect 8944 1294 8996 1300
rect 8772 898 8800 1294
rect 8772 870 8892 898
rect 8588 734 8800 762
rect 8864 746 8892 870
rect 8772 160 8800 734
rect 8852 740 8904 746
rect 8852 682 8904 688
rect 9048 160 9076 1924
rect 9128 1906 9180 1912
rect 9220 1964 9272 1970
rect 9220 1906 9272 1912
rect 9232 1494 9260 1906
rect 9220 1488 9272 1494
rect 9220 1430 9272 1436
rect 9128 1216 9180 1222
rect 9128 1158 9180 1164
rect 9220 1216 9272 1222
rect 9220 1158 9272 1164
rect 9140 814 9168 1158
rect 9232 1018 9260 1158
rect 9220 1012 9272 1018
rect 9220 954 9272 960
rect 9128 808 9180 814
rect 9128 750 9180 756
rect 9324 160 9352 2382
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9416 1970 9444 2246
rect 9404 1964 9456 1970
rect 9404 1906 9456 1912
rect 9508 1834 9536 2246
rect 9496 1828 9548 1834
rect 9496 1770 9548 1776
rect 9692 1442 9720 2400
rect 9864 2382 9916 2388
rect 10244 2281 10272 2615
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 10230 2272 10286 2281
rect 10230 2207 10286 2216
rect 10152 2060 10640 2088
rect 9772 1964 9824 1970
rect 9772 1906 9824 1912
rect 9600 1414 9720 1442
rect 9600 160 9628 1414
rect 9680 1216 9732 1222
rect 9680 1158 9732 1164
rect 9692 882 9720 1158
rect 9680 876 9732 882
rect 9680 818 9732 824
rect 9784 814 9812 1906
rect 10152 1834 10180 2060
rect 10232 1964 10284 1970
rect 10232 1906 10284 1912
rect 10324 1964 10376 1970
rect 10324 1906 10376 1912
rect 10140 1828 10192 1834
rect 10140 1770 10192 1776
rect 9851 1660 10159 1669
rect 9851 1658 9857 1660
rect 9913 1658 9937 1660
rect 9993 1658 10017 1660
rect 10073 1658 10097 1660
rect 10153 1658 10159 1660
rect 9913 1606 9915 1658
rect 10095 1606 10097 1658
rect 9851 1604 9857 1606
rect 9913 1604 9937 1606
rect 9993 1604 10017 1606
rect 10073 1604 10097 1606
rect 10153 1604 10159 1606
rect 9851 1595 10159 1604
rect 9956 1556 10008 1562
rect 9956 1498 10008 1504
rect 9968 1442 9996 1498
rect 9876 1414 9996 1442
rect 9876 1193 9904 1414
rect 9956 1352 10008 1358
rect 9956 1294 10008 1300
rect 10140 1352 10192 1358
rect 10140 1294 10192 1300
rect 9862 1184 9918 1193
rect 9862 1119 9918 1128
rect 9772 808 9824 814
rect 9772 750 9824 756
rect 9680 740 9732 746
rect 9680 682 9732 688
rect 9692 626 9720 682
rect 9692 598 9904 626
rect 9968 610 9996 1294
rect 10048 1216 10100 1222
rect 10048 1158 10100 1164
rect 9876 160 9904 598
rect 9956 604 10008 610
rect 9956 546 10008 552
rect 5170 82 5226 160
rect 5000 54 5226 82
rect 5170 0 5226 54
rect 5446 0 5502 160
rect 5722 0 5778 160
rect 5998 0 6054 160
rect 6274 0 6330 160
rect 6550 0 6606 160
rect 6826 0 6882 160
rect 7102 0 7158 160
rect 7378 0 7434 160
rect 7654 0 7710 160
rect 7930 0 7986 160
rect 8206 0 8262 160
rect 8482 0 8538 160
rect 8758 0 8814 160
rect 9034 0 9090 160
rect 9310 0 9366 160
rect 9586 0 9642 160
rect 9862 0 9918 160
rect 10060 82 10088 1158
rect 10152 474 10180 1294
rect 10140 468 10192 474
rect 10140 410 10192 416
rect 10244 202 10272 1906
rect 10336 1465 10364 1906
rect 10508 1760 10560 1766
rect 10428 1720 10508 1748
rect 10322 1456 10378 1465
rect 10322 1391 10378 1400
rect 10232 196 10284 202
rect 10138 82 10194 160
rect 10428 160 10456 1720
rect 10508 1702 10560 1708
rect 10508 1420 10560 1426
rect 10508 1362 10560 1368
rect 10520 377 10548 1362
rect 10612 1358 10640 2060
rect 10704 1426 10732 2382
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 10888 1426 10916 2042
rect 11060 1760 11112 1766
rect 10980 1720 11060 1748
rect 10692 1420 10744 1426
rect 10692 1362 10744 1368
rect 10876 1420 10928 1426
rect 10876 1362 10928 1368
rect 10600 1352 10652 1358
rect 10600 1294 10652 1300
rect 10692 1284 10744 1290
rect 10692 1226 10744 1232
rect 10784 1284 10836 1290
rect 10784 1226 10836 1232
rect 10506 368 10562 377
rect 10506 303 10562 312
rect 10704 160 10732 1226
rect 10796 950 10824 1226
rect 10784 944 10836 950
rect 10784 886 10836 892
rect 10980 160 11008 1720
rect 11060 1702 11112 1708
rect 11060 1420 11112 1426
rect 11060 1362 11112 1368
rect 10232 138 10284 144
rect 10060 54 10194 82
rect 10138 0 10194 54
rect 10414 0 10470 160
rect 10690 0 10746 160
rect 10966 0 11022 160
rect 11072 82 11100 1362
rect 11256 950 11284 2246
rect 11428 2032 11480 2038
rect 11428 1974 11480 1980
rect 11336 1964 11388 1970
rect 11336 1906 11388 1912
rect 11244 944 11296 950
rect 11244 886 11296 892
rect 11348 338 11376 1906
rect 11440 1562 11468 1974
rect 11624 1970 11652 2314
rect 11808 2310 11836 2382
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 11992 1986 12020 2382
rect 11612 1964 11664 1970
rect 11992 1958 12112 1986
rect 11612 1906 11664 1912
rect 11716 1822 11928 1850
rect 11716 1766 11744 1822
rect 11704 1760 11756 1766
rect 11704 1702 11756 1708
rect 11796 1760 11848 1766
rect 11796 1702 11848 1708
rect 11428 1556 11480 1562
rect 11428 1498 11480 1504
rect 11612 1352 11664 1358
rect 11612 1294 11664 1300
rect 11704 1352 11756 1358
rect 11704 1294 11756 1300
rect 11428 1216 11480 1222
rect 11480 1176 11560 1204
rect 11428 1158 11480 1164
rect 11336 332 11388 338
rect 11336 274 11388 280
rect 11532 160 11560 1176
rect 11624 542 11652 1294
rect 11716 921 11744 1294
rect 11702 912 11758 921
rect 11702 847 11758 856
rect 11612 536 11664 542
rect 11612 478 11664 484
rect 11808 160 11836 1702
rect 11242 82 11298 160
rect 11072 54 11298 82
rect 11242 0 11298 54
rect 11518 0 11574 160
rect 11794 0 11850 160
rect 11900 82 11928 1822
rect 12084 388 12112 1958
rect 12176 1562 12204 2450
rect 12164 1556 12216 1562
rect 12164 1498 12216 1504
rect 12268 1358 12296 2887
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 12544 2446 12572 2790
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12360 1970 12388 2246
rect 12452 2009 12480 2314
rect 12636 2258 12664 4966
rect 13360 4684 13412 4690
rect 13360 4626 13412 4632
rect 12818 4380 13126 4389
rect 12818 4378 12824 4380
rect 12880 4378 12904 4380
rect 12960 4378 12984 4380
rect 13040 4378 13064 4380
rect 13120 4378 13126 4380
rect 12880 4326 12882 4378
rect 13062 4326 13064 4378
rect 12818 4324 12824 4326
rect 12880 4324 12904 4326
rect 12960 4324 12984 4326
rect 13040 4324 13064 4326
rect 13120 4324 13126 4326
rect 12818 4315 13126 4324
rect 12818 3292 13126 3301
rect 12818 3290 12824 3292
rect 12880 3290 12904 3292
rect 12960 3290 12984 3292
rect 13040 3290 13064 3292
rect 13120 3290 13126 3292
rect 12880 3238 12882 3290
rect 13062 3238 13064 3290
rect 12818 3236 12824 3238
rect 12880 3236 12904 3238
rect 12960 3236 12984 3238
rect 13040 3236 13064 3238
rect 13120 3236 13126 3238
rect 12818 3227 13126 3236
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 12544 2230 12664 2258
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 12438 2000 12494 2009
rect 12348 1964 12400 1970
rect 12438 1935 12494 1944
rect 12348 1906 12400 1912
rect 12440 1760 12492 1766
rect 12440 1702 12492 1708
rect 12452 1562 12480 1702
rect 12440 1556 12492 1562
rect 12440 1498 12492 1504
rect 12256 1352 12308 1358
rect 12256 1294 12308 1300
rect 12348 1216 12400 1222
rect 12348 1158 12400 1164
rect 11992 377 12112 388
rect 11978 368 12112 377
rect 12034 360 12112 368
rect 11978 303 12034 312
rect 12360 160 12388 1158
rect 12544 406 12572 2230
rect 12728 2038 12756 2246
rect 12818 2204 13126 2213
rect 12818 2202 12824 2204
rect 12880 2202 12904 2204
rect 12960 2202 12984 2204
rect 13040 2202 13064 2204
rect 13120 2202 13126 2204
rect 12880 2150 12882 2202
rect 13062 2150 13064 2202
rect 12818 2148 12824 2150
rect 12880 2148 12904 2150
rect 12960 2148 12984 2150
rect 13040 2148 13064 2150
rect 13120 2148 13126 2150
rect 12818 2139 13126 2148
rect 12716 2032 12768 2038
rect 12716 1974 12768 1980
rect 12808 1964 12860 1970
rect 12808 1906 12860 1912
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 12532 400 12584 406
rect 12532 342 12584 348
rect 12636 160 12664 1702
rect 12820 1329 12848 1906
rect 13188 1834 13216 2790
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 13176 1828 13228 1834
rect 13176 1770 13228 1776
rect 13176 1556 13228 1562
rect 13176 1498 13228 1504
rect 13188 1358 13216 1498
rect 13280 1358 13308 2518
rect 13176 1352 13228 1358
rect 12806 1320 12862 1329
rect 13176 1294 13228 1300
rect 13268 1352 13320 1358
rect 13268 1294 13320 1300
rect 12806 1255 12862 1264
rect 12716 1216 12768 1222
rect 12716 1158 12768 1164
rect 13084 1216 13136 1222
rect 13136 1176 13216 1204
rect 13084 1158 13136 1164
rect 12728 762 12756 1158
rect 12818 1116 13126 1125
rect 12818 1114 12824 1116
rect 12880 1114 12904 1116
rect 12960 1114 12984 1116
rect 13040 1114 13064 1116
rect 13120 1114 13126 1116
rect 12880 1062 12882 1114
rect 13062 1062 13064 1114
rect 12818 1060 12824 1062
rect 12880 1060 12904 1062
rect 12960 1060 12984 1062
rect 13040 1060 13064 1062
rect 13120 1060 13126 1062
rect 12818 1051 13126 1060
rect 12728 734 12940 762
rect 12912 160 12940 734
rect 13188 160 13216 1176
rect 13372 542 13400 4626
rect 13648 2496 13676 5034
rect 13740 4729 13768 5170
rect 13726 4720 13782 4729
rect 13726 4655 13782 4664
rect 13464 2468 13676 2496
rect 13464 1442 13492 2468
rect 13544 1760 13596 1766
rect 13542 1728 13544 1737
rect 13596 1728 13598 1737
rect 13542 1663 13598 1672
rect 13820 1556 13872 1562
rect 13740 1516 13820 1544
rect 13464 1414 13584 1442
rect 13452 1216 13504 1222
rect 13452 1158 13504 1164
rect 13360 536 13412 542
rect 13360 478 13412 484
rect 13464 160 13492 1158
rect 13556 898 13584 1414
rect 13636 1420 13688 1426
rect 13636 1362 13688 1368
rect 13648 1018 13676 1362
rect 13636 1012 13688 1018
rect 13636 954 13688 960
rect 13556 882 13676 898
rect 13556 876 13688 882
rect 13556 870 13636 876
rect 13636 818 13688 824
rect 13740 160 13768 1516
rect 13820 1498 13872 1504
rect 13924 610 13952 5238
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14004 2304 14056 2310
rect 14004 2246 14056 2252
rect 14016 2106 14044 2246
rect 14200 2106 14228 2450
rect 14004 2100 14056 2106
rect 14004 2042 14056 2048
rect 14188 2100 14240 2106
rect 14188 2042 14240 2048
rect 14094 2000 14150 2009
rect 14384 1970 14412 2926
rect 14752 2774 14780 5170
rect 14752 2746 14872 2774
rect 14554 2680 14610 2689
rect 14554 2615 14610 2624
rect 14568 2378 14596 2615
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 14094 1935 14096 1944
rect 14148 1935 14150 1944
rect 14372 1964 14424 1970
rect 14096 1906 14148 1912
rect 14372 1906 14424 1912
rect 14844 1850 14872 2746
rect 15028 2650 15056 5170
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 15785 4924 16093 4933
rect 15785 4922 15791 4924
rect 15847 4922 15871 4924
rect 15927 4922 15951 4924
rect 16007 4922 16031 4924
rect 16087 4922 16093 4924
rect 15847 4870 15849 4922
rect 16029 4870 16031 4922
rect 15785 4868 15791 4870
rect 15847 4868 15871 4870
rect 15927 4868 15951 4870
rect 16007 4868 16031 4870
rect 16087 4868 16093 4870
rect 15785 4859 16093 4868
rect 15785 3836 16093 3845
rect 15785 3834 15791 3836
rect 15847 3834 15871 3836
rect 15927 3834 15951 3836
rect 16007 3834 16031 3836
rect 16087 3834 16093 3836
rect 15847 3782 15849 3834
rect 16029 3782 16031 3834
rect 15785 3780 15791 3782
rect 15847 3780 15871 3782
rect 15927 3780 15951 3782
rect 16007 3780 16031 3782
rect 16087 3780 16093 3782
rect 15785 3771 16093 3780
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15016 2644 15068 2650
rect 15016 2586 15068 2592
rect 15580 2446 15608 2790
rect 15785 2748 16093 2757
rect 15785 2746 15791 2748
rect 15847 2746 15871 2748
rect 15927 2746 15951 2748
rect 16007 2746 16031 2748
rect 16087 2746 16093 2748
rect 15847 2694 15849 2746
rect 16029 2694 16031 2746
rect 15785 2692 15791 2694
rect 15847 2692 15871 2694
rect 15927 2692 15951 2694
rect 16007 2692 16031 2694
rect 16087 2692 16093 2694
rect 15785 2683 16093 2692
rect 15384 2440 15436 2446
rect 15304 2400 15384 2428
rect 15304 2310 15332 2400
rect 15384 2382 15436 2388
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 15488 2038 15516 2246
rect 15476 2032 15528 2038
rect 15476 1974 15528 1980
rect 15384 1964 15436 1970
rect 15384 1906 15436 1912
rect 14372 1828 14424 1834
rect 14844 1822 15056 1850
rect 14372 1770 14424 1776
rect 14384 1358 14412 1770
rect 14648 1760 14700 1766
rect 14648 1702 14700 1708
rect 14740 1760 14792 1766
rect 14740 1702 14792 1708
rect 14660 1442 14688 1702
rect 14476 1414 14688 1442
rect 14372 1352 14424 1358
rect 14372 1294 14424 1300
rect 14004 1216 14056 1222
rect 14004 1158 14056 1164
rect 13912 604 13964 610
rect 13912 546 13964 552
rect 14016 160 14044 1158
rect 12070 82 12126 160
rect 11900 54 12126 82
rect 12070 0 12126 54
rect 12346 0 12402 160
rect 12622 0 12678 160
rect 12898 0 12954 160
rect 13174 0 13230 160
rect 13450 0 13506 160
rect 13726 0 13782 160
rect 14002 0 14058 160
rect 14278 82 14334 160
rect 14476 82 14504 1414
rect 14648 1352 14700 1358
rect 14648 1294 14700 1300
rect 14660 814 14688 1294
rect 14648 808 14700 814
rect 14648 750 14700 756
rect 14278 54 14504 82
rect 14554 82 14610 160
rect 14752 82 14780 1702
rect 14924 1352 14976 1358
rect 14844 1300 14924 1306
rect 14844 1294 14976 1300
rect 14844 1278 14964 1294
rect 14844 160 14872 1278
rect 14924 1216 14976 1222
rect 14924 1158 14976 1164
rect 14936 950 14964 1158
rect 15028 950 15056 1822
rect 15108 1760 15160 1766
rect 15108 1702 15160 1708
rect 15198 1728 15254 1737
rect 15120 1562 15148 1702
rect 15396 1714 15424 1906
rect 15254 1686 15424 1714
rect 15476 1760 15528 1766
rect 15476 1702 15528 1708
rect 15198 1663 15254 1672
rect 15108 1556 15160 1562
rect 15108 1498 15160 1504
rect 15384 1556 15436 1562
rect 15384 1498 15436 1504
rect 15292 1488 15344 1494
rect 15120 1436 15292 1442
rect 15120 1430 15344 1436
rect 15120 1414 15332 1430
rect 14924 944 14976 950
rect 14924 886 14976 892
rect 15016 944 15068 950
rect 15016 886 15068 892
rect 15120 160 15148 1414
rect 15396 1358 15424 1498
rect 15488 1358 15516 1702
rect 15384 1352 15436 1358
rect 15384 1294 15436 1300
rect 15476 1352 15528 1358
rect 15476 1294 15528 1300
rect 15580 1170 15608 2246
rect 16040 2038 16068 2382
rect 16028 2032 16080 2038
rect 16028 1974 16080 1980
rect 16120 1964 16172 1970
rect 16120 1906 16172 1912
rect 15660 1760 15712 1766
rect 15660 1702 15712 1708
rect 15396 1142 15608 1170
rect 15396 160 15424 1142
rect 15672 160 15700 1702
rect 15785 1660 16093 1669
rect 15785 1658 15791 1660
rect 15847 1658 15871 1660
rect 15927 1658 15951 1660
rect 16007 1658 16031 1660
rect 16087 1658 16093 1660
rect 15847 1606 15849 1658
rect 16029 1606 16031 1658
rect 15785 1604 15791 1606
rect 15847 1604 15871 1606
rect 15927 1604 15951 1606
rect 16007 1604 16031 1606
rect 16087 1604 16093 1606
rect 15785 1595 16093 1604
rect 16132 1562 16160 1906
rect 16120 1556 16172 1562
rect 16120 1498 16172 1504
rect 16212 1556 16264 1562
rect 16212 1498 16264 1504
rect 16224 1442 16252 1498
rect 15948 1414 16252 1442
rect 16304 1420 16356 1426
rect 15948 160 15976 1414
rect 16304 1362 16356 1368
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 16132 474 16160 1294
rect 16120 468 16172 474
rect 16120 410 16172 416
rect 14554 54 14780 82
rect 14278 0 14334 54
rect 14554 0 14610 54
rect 14830 0 14886 160
rect 15106 0 15162 160
rect 15382 0 15438 160
rect 15658 0 15714 160
rect 15934 0 15990 160
rect 16210 82 16266 160
rect 16316 82 16344 1362
rect 16408 474 16436 4966
rect 17880 2922 17908 5170
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21272 5092 21324 5098
rect 21272 5034 21324 5040
rect 18752 4380 19060 4389
rect 18752 4378 18758 4380
rect 18814 4378 18838 4380
rect 18894 4378 18918 4380
rect 18974 4378 18998 4380
rect 19054 4378 19060 4380
rect 18814 4326 18816 4378
rect 18996 4326 18998 4378
rect 18752 4324 18758 4326
rect 18814 4324 18838 4326
rect 18894 4324 18918 4326
rect 18974 4324 18998 4326
rect 19054 4324 19060 4326
rect 18752 4315 19060 4324
rect 18752 3292 19060 3301
rect 18752 3290 18758 3292
rect 18814 3290 18838 3292
rect 18894 3290 18918 3292
rect 18974 3290 18998 3292
rect 19054 3290 19060 3292
rect 18814 3238 18816 3290
rect 18996 3238 18998 3290
rect 18752 3236 18758 3238
rect 18814 3236 18838 3238
rect 18894 3236 18918 3238
rect 18974 3236 18998 3238
rect 19054 3236 19060 3238
rect 18752 3227 19060 3236
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 19616 2848 19668 2854
rect 19616 2790 19668 2796
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 21178 2816 21234 2825
rect 19432 2576 19484 2582
rect 18142 2544 18198 2553
rect 19432 2518 19484 2524
rect 18142 2479 18198 2488
rect 19340 2508 19392 2514
rect 18156 2446 18184 2479
rect 19340 2450 19392 2456
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 18144 2440 18196 2446
rect 18972 2440 19024 2446
rect 18144 2382 18196 2388
rect 18340 2400 18972 2428
rect 16500 1562 16528 2382
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16580 1760 16632 1766
rect 16580 1702 16632 1708
rect 16488 1556 16540 1562
rect 16488 1498 16540 1504
rect 16592 1358 16620 1702
rect 16580 1352 16632 1358
rect 16580 1294 16632 1300
rect 16488 1216 16540 1222
rect 16488 1158 16540 1164
rect 16396 468 16448 474
rect 16396 410 16448 416
rect 16500 160 16528 1158
rect 16684 1018 16712 2246
rect 16764 1760 16816 1766
rect 16764 1702 16816 1708
rect 16672 1012 16724 1018
rect 16672 954 16724 960
rect 16776 160 16804 1702
rect 16868 1358 16896 2246
rect 16856 1352 16908 1358
rect 16856 1294 16908 1300
rect 16960 678 16988 2382
rect 17604 2106 17632 2382
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17592 2100 17644 2106
rect 17592 2042 17644 2048
rect 17788 2038 17816 2246
rect 17880 2106 17908 2382
rect 17972 2106 18000 2382
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18144 2304 18196 2310
rect 18144 2246 18196 2252
rect 18236 2304 18288 2310
rect 18236 2246 18288 2252
rect 17868 2100 17920 2106
rect 17868 2042 17920 2048
rect 17960 2100 18012 2106
rect 17960 2042 18012 2048
rect 17776 2032 17828 2038
rect 17776 1974 17828 1980
rect 17776 1828 17828 1834
rect 17604 1788 17776 1816
rect 17500 1556 17552 1562
rect 17052 1516 17500 1544
rect 16948 672 17000 678
rect 16948 614 17000 620
rect 17052 160 17080 1516
rect 17500 1498 17552 1504
rect 17500 1420 17552 1426
rect 17328 1380 17500 1408
rect 17328 160 17356 1380
rect 17500 1362 17552 1368
rect 17408 1284 17460 1290
rect 17408 1226 17460 1232
rect 17420 1018 17448 1226
rect 17408 1012 17460 1018
rect 17408 954 17460 960
rect 17604 160 17632 1788
rect 17776 1770 17828 1776
rect 17880 1822 18000 1850
rect 17880 160 17908 1822
rect 17972 1766 18000 1822
rect 17960 1760 18012 1766
rect 17960 1702 18012 1708
rect 18064 1426 18092 2246
rect 18052 1420 18104 1426
rect 18052 1362 18104 1368
rect 18156 1000 18184 2246
rect 18248 2106 18276 2246
rect 18236 2100 18288 2106
rect 18236 2042 18288 2048
rect 18236 1760 18288 1766
rect 18236 1702 18288 1708
rect 18064 972 18184 1000
rect 18064 649 18092 972
rect 18248 898 18276 1702
rect 18156 870 18276 898
rect 18050 640 18106 649
rect 18050 575 18106 584
rect 18156 160 18184 870
rect 18340 785 18368 2400
rect 18972 2382 19024 2388
rect 19156 2304 19208 2310
rect 19156 2246 19208 2252
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 18752 2204 19060 2213
rect 18752 2202 18758 2204
rect 18814 2202 18838 2204
rect 18894 2202 18918 2204
rect 18974 2202 18998 2204
rect 19054 2202 19060 2204
rect 18814 2150 18816 2202
rect 18996 2150 18998 2202
rect 18752 2148 18758 2150
rect 18814 2148 18838 2150
rect 18894 2148 18918 2150
rect 18974 2148 18998 2150
rect 19054 2148 19060 2150
rect 18752 2139 19060 2148
rect 19168 2106 19196 2246
rect 19260 2106 19288 2246
rect 19156 2100 19208 2106
rect 19156 2042 19208 2048
rect 19248 2100 19300 2106
rect 19248 2042 19300 2048
rect 19352 1970 19380 2450
rect 19340 1964 19392 1970
rect 19340 1906 19392 1912
rect 19340 1760 19392 1766
rect 19340 1702 19392 1708
rect 18432 1550 18736 1578
rect 18326 776 18382 785
rect 18326 711 18382 720
rect 18432 160 18460 1550
rect 18708 1494 18736 1550
rect 18696 1488 18748 1494
rect 18696 1430 18748 1436
rect 18604 1420 18656 1426
rect 19352 1408 19380 1702
rect 18604 1362 18656 1368
rect 19168 1380 19380 1408
rect 18616 626 18644 1362
rect 18752 1116 19060 1125
rect 18752 1114 18758 1116
rect 18814 1114 18838 1116
rect 18894 1114 18918 1116
rect 18974 1114 18998 1116
rect 19054 1114 19060 1116
rect 18814 1062 18816 1114
rect 18996 1062 18998 1114
rect 18752 1060 18758 1062
rect 18814 1060 18838 1062
rect 18894 1060 18918 1062
rect 18974 1060 18998 1062
rect 19054 1060 19060 1062
rect 18752 1051 19060 1060
rect 19168 898 19196 1380
rect 19444 1222 19472 2518
rect 19524 1828 19576 1834
rect 19524 1770 19576 1776
rect 19432 1216 19484 1222
rect 19432 1158 19484 1164
rect 19536 1034 19564 1770
rect 18984 870 19196 898
rect 19260 1006 19564 1034
rect 18616 598 18736 626
rect 18708 160 18736 598
rect 18984 160 19012 870
rect 19260 160 19288 1006
rect 16210 54 16344 82
rect 16210 0 16266 54
rect 16486 0 16542 160
rect 16762 0 16818 160
rect 17038 0 17094 160
rect 17314 0 17370 160
rect 17590 0 17646 160
rect 17866 0 17922 160
rect 18142 0 18198 160
rect 18418 0 18474 160
rect 18694 0 18750 160
rect 18970 0 19026 160
rect 19246 0 19302 160
rect 19522 82 19578 160
rect 19628 82 19656 2790
rect 19708 2440 19760 2446
rect 19706 2408 19708 2417
rect 20076 2440 20128 2446
rect 19760 2408 19762 2417
rect 20076 2382 20128 2388
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 19706 2343 19762 2352
rect 19708 2304 19760 2310
rect 19708 2246 19760 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19720 1290 19748 2246
rect 19800 1556 19852 1562
rect 19800 1498 19852 1504
rect 19708 1284 19760 1290
rect 19708 1226 19760 1232
rect 19812 160 19840 1498
rect 19996 1358 20024 2246
rect 19984 1352 20036 1358
rect 19984 1294 20036 1300
rect 20088 1222 20116 2382
rect 20168 2372 20220 2378
rect 20168 2314 20220 2320
rect 20076 1216 20128 1222
rect 20076 1158 20128 1164
rect 19522 54 19656 82
rect 19522 0 19578 54
rect 19798 0 19854 160
rect 20074 82 20130 160
rect 20180 82 20208 2314
rect 20272 1873 20300 2382
rect 20352 2304 20404 2310
rect 20352 2246 20404 2252
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 20902 2272 20958 2281
rect 20364 2106 20392 2246
rect 20640 2106 20668 2246
rect 20902 2207 20958 2216
rect 20916 2106 20944 2207
rect 21008 2106 21036 2790
rect 21178 2751 21234 2760
rect 20352 2100 20404 2106
rect 20352 2042 20404 2048
rect 20628 2100 20680 2106
rect 20628 2042 20680 2048
rect 20904 2100 20956 2106
rect 20904 2042 20956 2048
rect 20996 2100 21048 2106
rect 20996 2042 21048 2048
rect 20444 1896 20496 1902
rect 20258 1864 20314 1873
rect 20258 1799 20314 1808
rect 20364 1856 20444 1884
rect 20364 160 20392 1856
rect 20444 1838 20496 1844
rect 21088 1420 21140 1426
rect 21088 1362 21140 1368
rect 20628 1284 20680 1290
rect 20628 1226 20680 1232
rect 20640 160 20668 1226
rect 20074 54 20208 82
rect 20074 0 20130 54
rect 20350 0 20406 160
rect 20626 0 20682 160
rect 20902 82 20958 160
rect 21100 82 21128 1362
rect 21192 1358 21220 2751
rect 21284 1494 21312 5034
rect 21376 2582 21404 5102
rect 21364 2576 21416 2582
rect 21364 2518 21416 2524
rect 21468 2106 21496 5170
rect 21652 2106 21680 6190
rect 22572 6118 22600 7942
rect 23662 7840 23718 8000
rect 24858 7970 24914 8000
rect 24504 7942 24914 7970
rect 23676 6458 23704 7840
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 21719 6012 22027 6021
rect 21719 6010 21725 6012
rect 21781 6010 21805 6012
rect 21861 6010 21885 6012
rect 21941 6010 21965 6012
rect 22021 6010 22027 6012
rect 21781 5958 21783 6010
rect 21963 5958 21965 6010
rect 21719 5956 21725 5958
rect 21781 5956 21805 5958
rect 21861 5956 21885 5958
rect 21941 5956 21965 5958
rect 22021 5956 22027 5958
rect 21719 5947 22027 5956
rect 21719 4924 22027 4933
rect 21719 4922 21725 4924
rect 21781 4922 21805 4924
rect 21861 4922 21885 4924
rect 21941 4922 21965 4924
rect 22021 4922 22027 4924
rect 21781 4870 21783 4922
rect 21963 4870 21965 4922
rect 21719 4868 21725 4870
rect 21781 4868 21805 4870
rect 21861 4868 21885 4870
rect 21941 4868 21965 4870
rect 22021 4868 22027 4870
rect 21719 4859 22027 4868
rect 21719 3836 22027 3845
rect 21719 3834 21725 3836
rect 21781 3834 21805 3836
rect 21861 3834 21885 3836
rect 21941 3834 21965 3836
rect 22021 3834 22027 3836
rect 21781 3782 21783 3834
rect 21963 3782 21965 3834
rect 21719 3780 21725 3782
rect 21781 3780 21805 3782
rect 21861 3780 21885 3782
rect 21941 3780 21965 3782
rect 22021 3780 22027 3782
rect 21719 3771 22027 3780
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 21719 2748 22027 2757
rect 21719 2746 21725 2748
rect 21781 2746 21805 2748
rect 21861 2746 21885 2748
rect 21941 2746 21965 2748
rect 22021 2746 22027 2748
rect 21781 2694 21783 2746
rect 21963 2694 21965 2746
rect 21719 2692 21725 2694
rect 21781 2692 21805 2694
rect 21861 2692 21885 2694
rect 21941 2692 21965 2694
rect 22021 2692 22027 2694
rect 21719 2683 22027 2692
rect 22664 2650 22692 2858
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 23032 2666 23060 2790
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 22848 2638 23060 2666
rect 22848 2446 22876 2638
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 22836 2440 22888 2446
rect 22836 2382 22888 2388
rect 22282 2272 22338 2281
rect 22282 2207 22338 2216
rect 22296 2106 22324 2207
rect 21456 2100 21508 2106
rect 21456 2042 21508 2048
rect 21640 2100 21692 2106
rect 21640 2042 21692 2048
rect 22284 2100 22336 2106
rect 22284 2042 22336 2048
rect 21732 1964 21784 1970
rect 21652 1924 21732 1952
rect 21456 1828 21508 1834
rect 21456 1770 21508 1776
rect 21468 1562 21496 1770
rect 21652 1562 21680 1924
rect 21732 1906 21784 1912
rect 22100 1964 22152 1970
rect 22100 1906 22152 1912
rect 21719 1660 22027 1669
rect 21719 1658 21725 1660
rect 21781 1658 21805 1660
rect 21861 1658 21885 1660
rect 21941 1658 21965 1660
rect 22021 1658 22027 1660
rect 21781 1606 21783 1658
rect 21963 1606 21965 1658
rect 21719 1604 21725 1606
rect 21781 1604 21805 1606
rect 21861 1604 21885 1606
rect 21941 1604 21965 1606
rect 22021 1604 22027 1606
rect 21719 1595 22027 1604
rect 21456 1556 21508 1562
rect 21456 1498 21508 1504
rect 21640 1556 21692 1562
rect 21640 1498 21692 1504
rect 21272 1488 21324 1494
rect 21272 1430 21324 1436
rect 22112 1408 22140 1906
rect 22388 1766 22416 2382
rect 22652 2304 22704 2310
rect 22652 2246 22704 2252
rect 22664 2106 22692 2246
rect 23124 2106 23152 6258
rect 23676 3738 23704 6258
rect 24216 6180 24268 6186
rect 24216 6122 24268 6128
rect 24032 5840 24084 5846
rect 24032 5782 24084 5788
rect 23848 5636 23900 5642
rect 23848 5578 23900 5584
rect 23860 5370 23888 5578
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 23216 2650 23244 3334
rect 23572 2848 23624 2854
rect 23572 2790 23624 2796
rect 23204 2644 23256 2650
rect 23204 2586 23256 2592
rect 23296 2440 23348 2446
rect 23202 2408 23258 2417
rect 23348 2388 23520 2394
rect 23296 2382 23520 2388
rect 23308 2366 23520 2382
rect 23202 2343 23258 2352
rect 23216 2106 23244 2343
rect 22652 2100 22704 2106
rect 22652 2042 22704 2048
rect 23112 2100 23164 2106
rect 23112 2042 23164 2048
rect 23204 2100 23256 2106
rect 23204 2042 23256 2048
rect 23388 2032 23440 2038
rect 23388 1974 23440 1980
rect 23020 1964 23072 1970
rect 22848 1924 23020 1952
rect 22376 1760 22428 1766
rect 22376 1702 22428 1708
rect 21928 1380 22140 1408
rect 22480 1426 22784 1442
rect 22480 1420 22796 1426
rect 22480 1414 22744 1420
rect 21180 1352 21232 1358
rect 21180 1294 21232 1300
rect 21824 1352 21876 1358
rect 21824 1294 21876 1300
rect 21272 740 21324 746
rect 21272 682 21324 688
rect 21284 354 21312 682
rect 21456 672 21508 678
rect 21456 614 21508 620
rect 21192 326 21312 354
rect 21192 160 21220 326
rect 21468 160 21496 614
rect 21836 513 21864 1294
rect 21822 504 21878 513
rect 21822 439 21878 448
rect 20902 54 21128 82
rect 20902 0 20958 54
rect 21178 0 21234 160
rect 21454 0 21510 160
rect 21730 82 21786 160
rect 21928 82 21956 1380
rect 22008 1216 22060 1222
rect 22008 1158 22060 1164
rect 22284 1216 22336 1222
rect 22284 1158 22336 1164
rect 22020 678 22048 1158
rect 22296 1018 22324 1158
rect 22284 1012 22336 1018
rect 22284 954 22336 960
rect 22008 672 22060 678
rect 22008 614 22060 620
rect 22008 536 22060 542
rect 22008 478 22060 484
rect 22020 160 22048 478
rect 21730 54 21956 82
rect 21730 0 21786 54
rect 22006 0 22062 160
rect 22282 82 22338 160
rect 22480 82 22508 1414
rect 22744 1362 22796 1368
rect 22652 1352 22704 1358
rect 22652 1294 22704 1300
rect 22560 1216 22612 1222
rect 22560 1158 22612 1164
rect 22572 1018 22600 1158
rect 22560 1012 22612 1018
rect 22560 954 22612 960
rect 22664 746 22692 1294
rect 22744 1216 22796 1222
rect 22744 1158 22796 1164
rect 22756 882 22784 1158
rect 22744 876 22796 882
rect 22744 818 22796 824
rect 22652 740 22704 746
rect 22652 682 22704 688
rect 22744 332 22796 338
rect 22744 274 22796 280
rect 22282 54 22508 82
rect 22558 82 22614 160
rect 22756 82 22784 274
rect 22848 160 22876 1924
rect 23020 1906 23072 1912
rect 23020 1760 23072 1766
rect 23020 1702 23072 1708
rect 23032 354 23060 1702
rect 23112 1216 23164 1222
rect 23112 1158 23164 1164
rect 23296 1216 23348 1222
rect 23296 1158 23348 1164
rect 23124 474 23152 1158
rect 23308 1018 23336 1158
rect 23296 1012 23348 1018
rect 23296 954 23348 960
rect 23112 468 23164 474
rect 23112 410 23164 416
rect 23032 326 23152 354
rect 23124 160 23152 326
rect 23400 160 23428 1974
rect 23492 1562 23520 2366
rect 23480 1556 23532 1562
rect 23480 1498 23532 1504
rect 23480 1352 23532 1358
rect 23480 1294 23532 1300
rect 23492 746 23520 1294
rect 23584 1290 23612 2790
rect 23676 2502 23796 2530
rect 23572 1284 23624 1290
rect 23572 1226 23624 1232
rect 23480 740 23532 746
rect 23480 682 23532 688
rect 23676 160 23704 2502
rect 23768 2446 23796 2502
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23848 2372 23900 2378
rect 23848 2314 23900 2320
rect 23860 762 23888 2314
rect 23952 2310 23980 4558
rect 24044 2938 24072 5782
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 24136 3194 24164 3470
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 24044 2910 24164 2938
rect 24032 2848 24084 2854
rect 24032 2790 24084 2796
rect 24044 2446 24072 2790
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 23940 2304 23992 2310
rect 23940 2246 23992 2252
rect 24032 2304 24084 2310
rect 24032 2246 24084 2252
rect 24044 2106 24072 2246
rect 23940 2100 23992 2106
rect 23940 2042 23992 2048
rect 24032 2100 24084 2106
rect 24032 2042 24084 2048
rect 23952 1442 23980 2042
rect 24136 1766 24164 2910
rect 24228 1834 24256 6122
rect 24504 5914 24532 7942
rect 24858 7840 24914 7942
rect 24686 6556 24994 6565
rect 24686 6554 24692 6556
rect 24748 6554 24772 6556
rect 24828 6554 24852 6556
rect 24908 6554 24932 6556
rect 24988 6554 24994 6556
rect 24748 6502 24750 6554
rect 24930 6502 24932 6554
rect 24686 6500 24692 6502
rect 24748 6500 24772 6502
rect 24828 6500 24852 6502
rect 24908 6500 24932 6502
rect 24988 6500 24994 6502
rect 24686 6491 24994 6500
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24686 5468 24994 5477
rect 24686 5466 24692 5468
rect 24748 5466 24772 5468
rect 24828 5466 24852 5468
rect 24908 5466 24932 5468
rect 24988 5466 24994 5468
rect 24748 5414 24750 5466
rect 24930 5414 24932 5466
rect 24686 5412 24692 5414
rect 24748 5412 24772 5414
rect 24828 5412 24852 5414
rect 24908 5412 24932 5414
rect 24988 5412 24994 5414
rect 24686 5403 24994 5412
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24320 4826 24348 5170
rect 24308 4820 24360 4826
rect 24308 4762 24360 4768
rect 24686 4380 24994 4389
rect 24686 4378 24692 4380
rect 24748 4378 24772 4380
rect 24828 4378 24852 4380
rect 24908 4378 24932 4380
rect 24988 4378 24994 4380
rect 24748 4326 24750 4378
rect 24930 4326 24932 4378
rect 24686 4324 24692 4326
rect 24748 4324 24772 4326
rect 24828 4324 24852 4326
rect 24908 4324 24932 4326
rect 24988 4324 24994 4326
rect 24686 4315 24994 4324
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 24320 3058 24348 3334
rect 24686 3292 24994 3301
rect 24686 3290 24692 3292
rect 24748 3290 24772 3292
rect 24828 3290 24852 3292
rect 24908 3290 24932 3292
rect 24988 3290 24994 3292
rect 24748 3238 24750 3290
rect 24930 3238 24932 3290
rect 24686 3236 24692 3238
rect 24748 3236 24772 3238
rect 24828 3236 24852 3238
rect 24908 3236 24932 3238
rect 24988 3236 24994 3238
rect 24686 3227 24994 3236
rect 25044 3120 25096 3126
rect 25044 3062 25096 3068
rect 24308 3052 24360 3058
rect 24308 2994 24360 3000
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 24216 1828 24268 1834
rect 24216 1770 24268 1776
rect 24124 1760 24176 1766
rect 24124 1702 24176 1708
rect 23952 1414 24164 1442
rect 24032 1352 24084 1358
rect 24032 1294 24084 1300
rect 23940 1216 23992 1222
rect 23940 1158 23992 1164
rect 23952 921 23980 1158
rect 23938 912 23994 921
rect 23938 847 23994 856
rect 23860 734 23980 762
rect 23952 160 23980 734
rect 24044 338 24072 1294
rect 24136 490 24164 1414
rect 24216 1216 24268 1222
rect 24216 1158 24268 1164
rect 24228 610 24256 1158
rect 24216 604 24268 610
rect 24216 546 24268 552
rect 24136 462 24256 490
rect 24032 332 24084 338
rect 24032 274 24084 280
rect 24228 160 24256 462
rect 24504 160 24532 2926
rect 24584 2916 24636 2922
rect 24584 2858 24636 2864
rect 22558 54 22784 82
rect 22282 0 22338 54
rect 22558 0 22614 54
rect 22834 0 22890 160
rect 23110 0 23166 160
rect 23386 0 23442 160
rect 23662 0 23718 160
rect 23938 0 23994 160
rect 24214 0 24270 160
rect 24490 0 24546 160
rect 24596 82 24624 2858
rect 24686 2204 24994 2213
rect 24686 2202 24692 2204
rect 24748 2202 24772 2204
rect 24828 2202 24852 2204
rect 24908 2202 24932 2204
rect 24988 2202 24994 2204
rect 24748 2150 24750 2202
rect 24930 2150 24932 2202
rect 24686 2148 24692 2150
rect 24748 2148 24772 2150
rect 24828 2148 24852 2150
rect 24908 2148 24932 2150
rect 24988 2148 24994 2150
rect 24686 2139 24994 2148
rect 24676 1556 24728 1562
rect 24676 1498 24728 1504
rect 24688 1426 24716 1498
rect 24676 1420 24728 1426
rect 24676 1362 24728 1368
rect 24686 1116 24994 1125
rect 24686 1114 24692 1116
rect 24748 1114 24772 1116
rect 24828 1114 24852 1116
rect 24908 1114 24932 1116
rect 24988 1114 24994 1116
rect 24748 1062 24750 1114
rect 24930 1062 24932 1114
rect 24686 1060 24692 1062
rect 24748 1060 24772 1062
rect 24828 1060 24852 1062
rect 24908 1060 24932 1062
rect 24988 1060 24994 1062
rect 24686 1051 24994 1060
rect 25056 160 25084 3062
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 25332 160 25360 2450
rect 25596 1420 25648 1426
rect 25596 1362 25648 1368
rect 25608 160 25636 1362
rect 24766 82 24822 160
rect 24596 54 24822 82
rect 24766 0 24822 54
rect 25042 0 25098 160
rect 25318 0 25374 160
rect 25594 0 25650 160
<< via2 >>
rect 6890 6554 6946 6556
rect 6970 6554 7026 6556
rect 7050 6554 7106 6556
rect 7130 6554 7186 6556
rect 6890 6502 6936 6554
rect 6936 6502 6946 6554
rect 6970 6502 7000 6554
rect 7000 6502 7012 6554
rect 7012 6502 7026 6554
rect 7050 6502 7064 6554
rect 7064 6502 7076 6554
rect 7076 6502 7106 6554
rect 7130 6502 7140 6554
rect 7140 6502 7186 6554
rect 6890 6500 6946 6502
rect 6970 6500 7026 6502
rect 7050 6500 7106 6502
rect 7130 6500 7186 6502
rect 12824 6554 12880 6556
rect 12904 6554 12960 6556
rect 12984 6554 13040 6556
rect 13064 6554 13120 6556
rect 12824 6502 12870 6554
rect 12870 6502 12880 6554
rect 12904 6502 12934 6554
rect 12934 6502 12946 6554
rect 12946 6502 12960 6554
rect 12984 6502 12998 6554
rect 12998 6502 13010 6554
rect 13010 6502 13040 6554
rect 13064 6502 13074 6554
rect 13074 6502 13120 6554
rect 12824 6500 12880 6502
rect 12904 6500 12960 6502
rect 12984 6500 13040 6502
rect 13064 6500 13120 6502
rect 18758 6554 18814 6556
rect 18838 6554 18894 6556
rect 18918 6554 18974 6556
rect 18998 6554 19054 6556
rect 18758 6502 18804 6554
rect 18804 6502 18814 6554
rect 18838 6502 18868 6554
rect 18868 6502 18880 6554
rect 18880 6502 18894 6554
rect 18918 6502 18932 6554
rect 18932 6502 18944 6554
rect 18944 6502 18974 6554
rect 18998 6502 19008 6554
rect 19008 6502 19054 6554
rect 18758 6500 18814 6502
rect 18838 6500 18894 6502
rect 18918 6500 18974 6502
rect 18998 6500 19054 6502
rect 2226 6316 2282 6352
rect 2226 6296 2228 6316
rect 2228 6296 2280 6316
rect 2280 6296 2282 6316
rect 3923 6010 3979 6012
rect 4003 6010 4059 6012
rect 4083 6010 4139 6012
rect 4163 6010 4219 6012
rect 3923 5958 3969 6010
rect 3969 5958 3979 6010
rect 4003 5958 4033 6010
rect 4033 5958 4045 6010
rect 4045 5958 4059 6010
rect 4083 5958 4097 6010
rect 4097 5958 4109 6010
rect 4109 5958 4139 6010
rect 4163 5958 4173 6010
rect 4173 5958 4219 6010
rect 3923 5956 3979 5958
rect 4003 5956 4059 5958
rect 4083 5956 4139 5958
rect 4163 5956 4219 5958
rect 9857 6010 9913 6012
rect 9937 6010 9993 6012
rect 10017 6010 10073 6012
rect 10097 6010 10153 6012
rect 9857 5958 9903 6010
rect 9903 5958 9913 6010
rect 9937 5958 9967 6010
rect 9967 5958 9979 6010
rect 9979 5958 9993 6010
rect 10017 5958 10031 6010
rect 10031 5958 10043 6010
rect 10043 5958 10073 6010
rect 10097 5958 10107 6010
rect 10107 5958 10153 6010
rect 9857 5956 9913 5958
rect 9937 5956 9993 5958
rect 10017 5956 10073 5958
rect 10097 5956 10153 5958
rect 15791 6010 15847 6012
rect 15871 6010 15927 6012
rect 15951 6010 16007 6012
rect 16031 6010 16087 6012
rect 15791 5958 15837 6010
rect 15837 5958 15847 6010
rect 15871 5958 15901 6010
rect 15901 5958 15913 6010
rect 15913 5958 15927 6010
rect 15951 5958 15965 6010
rect 15965 5958 15977 6010
rect 15977 5958 16007 6010
rect 16031 5958 16041 6010
rect 16041 5958 16087 6010
rect 15791 5956 15847 5958
rect 15871 5956 15927 5958
rect 15951 5956 16007 5958
rect 16031 5956 16087 5958
rect 6890 5466 6946 5468
rect 6970 5466 7026 5468
rect 7050 5466 7106 5468
rect 7130 5466 7186 5468
rect 6890 5414 6936 5466
rect 6936 5414 6946 5466
rect 6970 5414 7000 5466
rect 7000 5414 7012 5466
rect 7012 5414 7026 5466
rect 7050 5414 7064 5466
rect 7064 5414 7076 5466
rect 7076 5414 7106 5466
rect 7130 5414 7140 5466
rect 7140 5414 7186 5466
rect 6890 5412 6946 5414
rect 6970 5412 7026 5414
rect 7050 5412 7106 5414
rect 7130 5412 7186 5414
rect 12824 5466 12880 5468
rect 12904 5466 12960 5468
rect 12984 5466 13040 5468
rect 13064 5466 13120 5468
rect 12824 5414 12870 5466
rect 12870 5414 12880 5466
rect 12904 5414 12934 5466
rect 12934 5414 12946 5466
rect 12946 5414 12960 5466
rect 12984 5414 12998 5466
rect 12998 5414 13010 5466
rect 13010 5414 13040 5466
rect 13064 5414 13074 5466
rect 13074 5414 13120 5466
rect 12824 5412 12880 5414
rect 12904 5412 12960 5414
rect 12984 5412 13040 5414
rect 13064 5412 13120 5414
rect 18758 5466 18814 5468
rect 18838 5466 18894 5468
rect 18918 5466 18974 5468
rect 18998 5466 19054 5468
rect 18758 5414 18804 5466
rect 18804 5414 18814 5466
rect 18838 5414 18868 5466
rect 18868 5414 18880 5466
rect 18880 5414 18894 5466
rect 18918 5414 18932 5466
rect 18932 5414 18944 5466
rect 18944 5414 18974 5466
rect 18998 5414 19008 5466
rect 19008 5414 19054 5466
rect 18758 5412 18814 5414
rect 18838 5412 18894 5414
rect 18918 5412 18974 5414
rect 18998 5412 19054 5414
rect 3923 4922 3979 4924
rect 4003 4922 4059 4924
rect 4083 4922 4139 4924
rect 4163 4922 4219 4924
rect 3923 4870 3969 4922
rect 3969 4870 3979 4922
rect 4003 4870 4033 4922
rect 4033 4870 4045 4922
rect 4045 4870 4059 4922
rect 4083 4870 4097 4922
rect 4097 4870 4109 4922
rect 4109 4870 4139 4922
rect 4163 4870 4173 4922
rect 4173 4870 4219 4922
rect 3923 4868 3979 4870
rect 4003 4868 4059 4870
rect 4083 4868 4139 4870
rect 4163 4868 4219 4870
rect 9586 5108 9588 5128
rect 9588 5108 9640 5128
rect 9640 5108 9642 5128
rect 9586 5072 9642 5108
rect 9857 4922 9913 4924
rect 9937 4922 9993 4924
rect 10017 4922 10073 4924
rect 10097 4922 10153 4924
rect 9857 4870 9903 4922
rect 9903 4870 9913 4922
rect 9937 4870 9967 4922
rect 9967 4870 9979 4922
rect 9979 4870 9993 4922
rect 10017 4870 10031 4922
rect 10031 4870 10043 4922
rect 10043 4870 10073 4922
rect 10097 4870 10107 4922
rect 10107 4870 10153 4922
rect 9857 4868 9913 4870
rect 9937 4868 9993 4870
rect 10017 4868 10073 4870
rect 10097 4868 10153 4870
rect 6890 4378 6946 4380
rect 6970 4378 7026 4380
rect 7050 4378 7106 4380
rect 7130 4378 7186 4380
rect 6890 4326 6936 4378
rect 6936 4326 6946 4378
rect 6970 4326 7000 4378
rect 7000 4326 7012 4378
rect 7012 4326 7026 4378
rect 7050 4326 7064 4378
rect 7064 4326 7076 4378
rect 7076 4326 7106 4378
rect 7130 4326 7140 4378
rect 7140 4326 7186 4378
rect 6890 4324 6946 4326
rect 6970 4324 7026 4326
rect 7050 4324 7106 4326
rect 7130 4324 7186 4326
rect 11242 4120 11298 4176
rect 3923 3834 3979 3836
rect 4003 3834 4059 3836
rect 4083 3834 4139 3836
rect 4163 3834 4219 3836
rect 3923 3782 3969 3834
rect 3969 3782 3979 3834
rect 4003 3782 4033 3834
rect 4033 3782 4045 3834
rect 4045 3782 4059 3834
rect 4083 3782 4097 3834
rect 4097 3782 4109 3834
rect 4109 3782 4139 3834
rect 4163 3782 4173 3834
rect 4173 3782 4219 3834
rect 3923 3780 3979 3782
rect 4003 3780 4059 3782
rect 4083 3780 4139 3782
rect 4163 3780 4219 3782
rect 9857 3834 9913 3836
rect 9937 3834 9993 3836
rect 10017 3834 10073 3836
rect 10097 3834 10153 3836
rect 9857 3782 9903 3834
rect 9903 3782 9913 3834
rect 9937 3782 9967 3834
rect 9967 3782 9979 3834
rect 9979 3782 9993 3834
rect 10017 3782 10031 3834
rect 10031 3782 10043 3834
rect 10043 3782 10073 3834
rect 10097 3782 10107 3834
rect 10107 3782 10153 3834
rect 9857 3780 9913 3782
rect 9937 3780 9993 3782
rect 10017 3780 10073 3782
rect 10097 3780 10153 3782
rect 6890 3290 6946 3292
rect 6970 3290 7026 3292
rect 7050 3290 7106 3292
rect 7130 3290 7186 3292
rect 6890 3238 6936 3290
rect 6936 3238 6946 3290
rect 6970 3238 7000 3290
rect 7000 3238 7012 3290
rect 7012 3238 7026 3290
rect 7050 3238 7064 3290
rect 7064 3238 7076 3290
rect 7076 3238 7106 3290
rect 7130 3238 7140 3290
rect 7140 3238 7186 3290
rect 6890 3236 6946 3238
rect 6970 3236 7026 3238
rect 7050 3236 7106 3238
rect 7130 3236 7186 3238
rect 7470 3032 7526 3088
rect 3923 2746 3979 2748
rect 4003 2746 4059 2748
rect 4083 2746 4139 2748
rect 4163 2746 4219 2748
rect 3923 2694 3969 2746
rect 3969 2694 3979 2746
rect 4003 2694 4033 2746
rect 4033 2694 4045 2746
rect 4045 2694 4059 2746
rect 4083 2694 4097 2746
rect 4097 2694 4109 2746
rect 4109 2694 4139 2746
rect 4163 2694 4173 2746
rect 4173 2694 4219 2746
rect 3923 2692 3979 2694
rect 4003 2692 4059 2694
rect 4083 2692 4139 2694
rect 4163 2692 4219 2694
rect 1950 1708 1952 1728
rect 1952 1708 2004 1728
rect 2004 1708 2006 1728
rect 1950 1672 2006 1708
rect 1950 312 2006 368
rect 2410 1944 2466 2000
rect 7194 2524 7196 2544
rect 7196 2524 7248 2544
rect 7248 2524 7250 2544
rect 2962 1436 2964 1456
rect 2964 1436 3016 1456
rect 3016 1436 3018 1456
rect 2962 1400 3018 1436
rect 2318 1264 2374 1320
rect 3923 1658 3979 1660
rect 4003 1658 4059 1660
rect 4083 1658 4139 1660
rect 4163 1658 4219 1660
rect 3923 1606 3969 1658
rect 3969 1606 3979 1658
rect 4003 1606 4033 1658
rect 4033 1606 4045 1658
rect 4045 1606 4059 1658
rect 4083 1606 4097 1658
rect 4097 1606 4109 1658
rect 4109 1606 4139 1658
rect 4163 1606 4173 1658
rect 4173 1606 4219 1658
rect 3923 1604 3979 1606
rect 4003 1604 4059 1606
rect 4083 1604 4139 1606
rect 4163 1604 4219 1606
rect 7194 2488 7250 2524
rect 5078 1264 5134 1320
rect 5906 1828 5962 1864
rect 5906 1808 5908 1828
rect 5908 1808 5960 1828
rect 5960 1808 5962 1828
rect 5906 720 5962 776
rect 6274 2352 6330 2408
rect 6890 2202 6946 2204
rect 6970 2202 7026 2204
rect 7050 2202 7106 2204
rect 7130 2202 7186 2204
rect 6890 2150 6936 2202
rect 6936 2150 6946 2202
rect 6970 2150 7000 2202
rect 7000 2150 7012 2202
rect 7012 2150 7026 2202
rect 7050 2150 7064 2202
rect 7064 2150 7076 2202
rect 7076 2150 7106 2202
rect 7130 2150 7140 2202
rect 7140 2150 7186 2202
rect 6890 2148 6946 2150
rect 6970 2148 7026 2150
rect 7050 2148 7106 2150
rect 7130 2148 7186 2150
rect 6182 584 6238 640
rect 5906 312 5962 368
rect 6890 1114 6946 1116
rect 6970 1114 7026 1116
rect 7050 1114 7106 1116
rect 7130 1114 7186 1116
rect 6890 1062 6936 1114
rect 6936 1062 6946 1114
rect 6970 1062 7000 1114
rect 7000 1062 7012 1114
rect 7012 1062 7026 1114
rect 7050 1062 7064 1114
rect 7064 1062 7076 1114
rect 7076 1062 7106 1114
rect 7130 1062 7140 1114
rect 7140 1062 7186 1114
rect 6890 1060 6946 1062
rect 6970 1060 7026 1062
rect 7050 1060 7106 1062
rect 7130 1060 7186 1062
rect 9034 2896 9090 2952
rect 12254 2896 12310 2952
rect 7838 2216 7894 2272
rect 8298 2080 8354 2136
rect 7838 1128 7894 1184
rect 7838 448 7894 504
rect 9857 2746 9913 2748
rect 9937 2746 9993 2748
rect 10017 2746 10073 2748
rect 10097 2746 10153 2748
rect 9857 2694 9903 2746
rect 9903 2694 9913 2746
rect 9937 2694 9967 2746
rect 9967 2694 9979 2746
rect 9979 2694 9993 2746
rect 10017 2694 10031 2746
rect 10031 2694 10043 2746
rect 10043 2694 10073 2746
rect 10097 2694 10107 2746
rect 10107 2694 10153 2746
rect 9857 2692 9913 2694
rect 9937 2692 9993 2694
rect 10017 2692 10073 2694
rect 10097 2692 10153 2694
rect 10230 2624 10286 2680
rect 8298 1672 8354 1728
rect 10230 2216 10286 2272
rect 9857 1658 9913 1660
rect 9937 1658 9993 1660
rect 10017 1658 10073 1660
rect 10097 1658 10153 1660
rect 9857 1606 9903 1658
rect 9903 1606 9913 1658
rect 9937 1606 9967 1658
rect 9967 1606 9979 1658
rect 9979 1606 9993 1658
rect 10017 1606 10031 1658
rect 10031 1606 10043 1658
rect 10043 1606 10073 1658
rect 10097 1606 10107 1658
rect 10107 1606 10153 1658
rect 9857 1604 9913 1606
rect 9937 1604 9993 1606
rect 10017 1604 10073 1606
rect 10097 1604 10153 1606
rect 9862 1128 9918 1184
rect 10322 1400 10378 1456
rect 10506 312 10562 368
rect 11702 856 11758 912
rect 12824 4378 12880 4380
rect 12904 4378 12960 4380
rect 12984 4378 13040 4380
rect 13064 4378 13120 4380
rect 12824 4326 12870 4378
rect 12870 4326 12880 4378
rect 12904 4326 12934 4378
rect 12934 4326 12946 4378
rect 12946 4326 12960 4378
rect 12984 4326 12998 4378
rect 12998 4326 13010 4378
rect 13010 4326 13040 4378
rect 13064 4326 13074 4378
rect 13074 4326 13120 4378
rect 12824 4324 12880 4326
rect 12904 4324 12960 4326
rect 12984 4324 13040 4326
rect 13064 4324 13120 4326
rect 12824 3290 12880 3292
rect 12904 3290 12960 3292
rect 12984 3290 13040 3292
rect 13064 3290 13120 3292
rect 12824 3238 12870 3290
rect 12870 3238 12880 3290
rect 12904 3238 12934 3290
rect 12934 3238 12946 3290
rect 12946 3238 12960 3290
rect 12984 3238 12998 3290
rect 12998 3238 13010 3290
rect 13010 3238 13040 3290
rect 13064 3238 13074 3290
rect 13074 3238 13120 3290
rect 12824 3236 12880 3238
rect 12904 3236 12960 3238
rect 12984 3236 13040 3238
rect 13064 3236 13120 3238
rect 12438 1944 12494 2000
rect 11978 312 12034 368
rect 12824 2202 12880 2204
rect 12904 2202 12960 2204
rect 12984 2202 13040 2204
rect 13064 2202 13120 2204
rect 12824 2150 12870 2202
rect 12870 2150 12880 2202
rect 12904 2150 12934 2202
rect 12934 2150 12946 2202
rect 12946 2150 12960 2202
rect 12984 2150 12998 2202
rect 12998 2150 13010 2202
rect 13010 2150 13040 2202
rect 13064 2150 13074 2202
rect 13074 2150 13120 2202
rect 12824 2148 12880 2150
rect 12904 2148 12960 2150
rect 12984 2148 13040 2150
rect 13064 2148 13120 2150
rect 12806 1264 12862 1320
rect 12824 1114 12880 1116
rect 12904 1114 12960 1116
rect 12984 1114 13040 1116
rect 13064 1114 13120 1116
rect 12824 1062 12870 1114
rect 12870 1062 12880 1114
rect 12904 1062 12934 1114
rect 12934 1062 12946 1114
rect 12946 1062 12960 1114
rect 12984 1062 12998 1114
rect 12998 1062 13010 1114
rect 13010 1062 13040 1114
rect 13064 1062 13074 1114
rect 13074 1062 13120 1114
rect 12824 1060 12880 1062
rect 12904 1060 12960 1062
rect 12984 1060 13040 1062
rect 13064 1060 13120 1062
rect 13726 4664 13782 4720
rect 13542 1708 13544 1728
rect 13544 1708 13596 1728
rect 13596 1708 13598 1728
rect 13542 1672 13598 1708
rect 14094 1964 14150 2000
rect 14554 2624 14610 2680
rect 14094 1944 14096 1964
rect 14096 1944 14148 1964
rect 14148 1944 14150 1964
rect 15791 4922 15847 4924
rect 15871 4922 15927 4924
rect 15951 4922 16007 4924
rect 16031 4922 16087 4924
rect 15791 4870 15837 4922
rect 15837 4870 15847 4922
rect 15871 4870 15901 4922
rect 15901 4870 15913 4922
rect 15913 4870 15927 4922
rect 15951 4870 15965 4922
rect 15965 4870 15977 4922
rect 15977 4870 16007 4922
rect 16031 4870 16041 4922
rect 16041 4870 16087 4922
rect 15791 4868 15847 4870
rect 15871 4868 15927 4870
rect 15951 4868 16007 4870
rect 16031 4868 16087 4870
rect 15791 3834 15847 3836
rect 15871 3834 15927 3836
rect 15951 3834 16007 3836
rect 16031 3834 16087 3836
rect 15791 3782 15837 3834
rect 15837 3782 15847 3834
rect 15871 3782 15901 3834
rect 15901 3782 15913 3834
rect 15913 3782 15927 3834
rect 15951 3782 15965 3834
rect 15965 3782 15977 3834
rect 15977 3782 16007 3834
rect 16031 3782 16041 3834
rect 16041 3782 16087 3834
rect 15791 3780 15847 3782
rect 15871 3780 15927 3782
rect 15951 3780 16007 3782
rect 16031 3780 16087 3782
rect 15791 2746 15847 2748
rect 15871 2746 15927 2748
rect 15951 2746 16007 2748
rect 16031 2746 16087 2748
rect 15791 2694 15837 2746
rect 15837 2694 15847 2746
rect 15871 2694 15901 2746
rect 15901 2694 15913 2746
rect 15913 2694 15927 2746
rect 15951 2694 15965 2746
rect 15965 2694 15977 2746
rect 15977 2694 16007 2746
rect 16031 2694 16041 2746
rect 16041 2694 16087 2746
rect 15791 2692 15847 2694
rect 15871 2692 15927 2694
rect 15951 2692 16007 2694
rect 16031 2692 16087 2694
rect 15198 1672 15254 1728
rect 15791 1658 15847 1660
rect 15871 1658 15927 1660
rect 15951 1658 16007 1660
rect 16031 1658 16087 1660
rect 15791 1606 15837 1658
rect 15837 1606 15847 1658
rect 15871 1606 15901 1658
rect 15901 1606 15913 1658
rect 15913 1606 15927 1658
rect 15951 1606 15965 1658
rect 15965 1606 15977 1658
rect 15977 1606 16007 1658
rect 16031 1606 16041 1658
rect 16041 1606 16087 1658
rect 15791 1604 15847 1606
rect 15871 1604 15927 1606
rect 15951 1604 16007 1606
rect 16031 1604 16087 1606
rect 18758 4378 18814 4380
rect 18838 4378 18894 4380
rect 18918 4378 18974 4380
rect 18998 4378 19054 4380
rect 18758 4326 18804 4378
rect 18804 4326 18814 4378
rect 18838 4326 18868 4378
rect 18868 4326 18880 4378
rect 18880 4326 18894 4378
rect 18918 4326 18932 4378
rect 18932 4326 18944 4378
rect 18944 4326 18974 4378
rect 18998 4326 19008 4378
rect 19008 4326 19054 4378
rect 18758 4324 18814 4326
rect 18838 4324 18894 4326
rect 18918 4324 18974 4326
rect 18998 4324 19054 4326
rect 18758 3290 18814 3292
rect 18838 3290 18894 3292
rect 18918 3290 18974 3292
rect 18998 3290 19054 3292
rect 18758 3238 18804 3290
rect 18804 3238 18814 3290
rect 18838 3238 18868 3290
rect 18868 3238 18880 3290
rect 18880 3238 18894 3290
rect 18918 3238 18932 3290
rect 18932 3238 18944 3290
rect 18944 3238 18974 3290
rect 18998 3238 19008 3290
rect 19008 3238 19054 3290
rect 18758 3236 18814 3238
rect 18838 3236 18894 3238
rect 18918 3236 18974 3238
rect 18998 3236 19054 3238
rect 18142 2488 18198 2544
rect 18050 584 18106 640
rect 18758 2202 18814 2204
rect 18838 2202 18894 2204
rect 18918 2202 18974 2204
rect 18998 2202 19054 2204
rect 18758 2150 18804 2202
rect 18804 2150 18814 2202
rect 18838 2150 18868 2202
rect 18868 2150 18880 2202
rect 18880 2150 18894 2202
rect 18918 2150 18932 2202
rect 18932 2150 18944 2202
rect 18944 2150 18974 2202
rect 18998 2150 19008 2202
rect 19008 2150 19054 2202
rect 18758 2148 18814 2150
rect 18838 2148 18894 2150
rect 18918 2148 18974 2150
rect 18998 2148 19054 2150
rect 18326 720 18382 776
rect 18758 1114 18814 1116
rect 18838 1114 18894 1116
rect 18918 1114 18974 1116
rect 18998 1114 19054 1116
rect 18758 1062 18804 1114
rect 18804 1062 18814 1114
rect 18838 1062 18868 1114
rect 18868 1062 18880 1114
rect 18880 1062 18894 1114
rect 18918 1062 18932 1114
rect 18932 1062 18944 1114
rect 18944 1062 18974 1114
rect 18998 1062 19008 1114
rect 19008 1062 19054 1114
rect 18758 1060 18814 1062
rect 18838 1060 18894 1062
rect 18918 1060 18974 1062
rect 18998 1060 19054 1062
rect 19706 2388 19708 2408
rect 19708 2388 19760 2408
rect 19760 2388 19762 2408
rect 19706 2352 19762 2388
rect 20902 2216 20958 2272
rect 21178 2760 21234 2816
rect 20258 1808 20314 1864
rect 21725 6010 21781 6012
rect 21805 6010 21861 6012
rect 21885 6010 21941 6012
rect 21965 6010 22021 6012
rect 21725 5958 21771 6010
rect 21771 5958 21781 6010
rect 21805 5958 21835 6010
rect 21835 5958 21847 6010
rect 21847 5958 21861 6010
rect 21885 5958 21899 6010
rect 21899 5958 21911 6010
rect 21911 5958 21941 6010
rect 21965 5958 21975 6010
rect 21975 5958 22021 6010
rect 21725 5956 21781 5958
rect 21805 5956 21861 5958
rect 21885 5956 21941 5958
rect 21965 5956 22021 5958
rect 21725 4922 21781 4924
rect 21805 4922 21861 4924
rect 21885 4922 21941 4924
rect 21965 4922 22021 4924
rect 21725 4870 21771 4922
rect 21771 4870 21781 4922
rect 21805 4870 21835 4922
rect 21835 4870 21847 4922
rect 21847 4870 21861 4922
rect 21885 4870 21899 4922
rect 21899 4870 21911 4922
rect 21911 4870 21941 4922
rect 21965 4870 21975 4922
rect 21975 4870 22021 4922
rect 21725 4868 21781 4870
rect 21805 4868 21861 4870
rect 21885 4868 21941 4870
rect 21965 4868 22021 4870
rect 21725 3834 21781 3836
rect 21805 3834 21861 3836
rect 21885 3834 21941 3836
rect 21965 3834 22021 3836
rect 21725 3782 21771 3834
rect 21771 3782 21781 3834
rect 21805 3782 21835 3834
rect 21835 3782 21847 3834
rect 21847 3782 21861 3834
rect 21885 3782 21899 3834
rect 21899 3782 21911 3834
rect 21911 3782 21941 3834
rect 21965 3782 21975 3834
rect 21975 3782 22021 3834
rect 21725 3780 21781 3782
rect 21805 3780 21861 3782
rect 21885 3780 21941 3782
rect 21965 3780 22021 3782
rect 21725 2746 21781 2748
rect 21805 2746 21861 2748
rect 21885 2746 21941 2748
rect 21965 2746 22021 2748
rect 21725 2694 21771 2746
rect 21771 2694 21781 2746
rect 21805 2694 21835 2746
rect 21835 2694 21847 2746
rect 21847 2694 21861 2746
rect 21885 2694 21899 2746
rect 21899 2694 21911 2746
rect 21911 2694 21941 2746
rect 21965 2694 21975 2746
rect 21975 2694 22021 2746
rect 21725 2692 21781 2694
rect 21805 2692 21861 2694
rect 21885 2692 21941 2694
rect 21965 2692 22021 2694
rect 22282 2216 22338 2272
rect 21725 1658 21781 1660
rect 21805 1658 21861 1660
rect 21885 1658 21941 1660
rect 21965 1658 22021 1660
rect 21725 1606 21771 1658
rect 21771 1606 21781 1658
rect 21805 1606 21835 1658
rect 21835 1606 21847 1658
rect 21847 1606 21861 1658
rect 21885 1606 21899 1658
rect 21899 1606 21911 1658
rect 21911 1606 21941 1658
rect 21965 1606 21975 1658
rect 21975 1606 22021 1658
rect 21725 1604 21781 1606
rect 21805 1604 21861 1606
rect 21885 1604 21941 1606
rect 21965 1604 22021 1606
rect 23202 2352 23258 2408
rect 21822 448 21878 504
rect 24692 6554 24748 6556
rect 24772 6554 24828 6556
rect 24852 6554 24908 6556
rect 24932 6554 24988 6556
rect 24692 6502 24738 6554
rect 24738 6502 24748 6554
rect 24772 6502 24802 6554
rect 24802 6502 24814 6554
rect 24814 6502 24828 6554
rect 24852 6502 24866 6554
rect 24866 6502 24878 6554
rect 24878 6502 24908 6554
rect 24932 6502 24942 6554
rect 24942 6502 24988 6554
rect 24692 6500 24748 6502
rect 24772 6500 24828 6502
rect 24852 6500 24908 6502
rect 24932 6500 24988 6502
rect 24692 5466 24748 5468
rect 24772 5466 24828 5468
rect 24852 5466 24908 5468
rect 24932 5466 24988 5468
rect 24692 5414 24738 5466
rect 24738 5414 24748 5466
rect 24772 5414 24802 5466
rect 24802 5414 24814 5466
rect 24814 5414 24828 5466
rect 24852 5414 24866 5466
rect 24866 5414 24878 5466
rect 24878 5414 24908 5466
rect 24932 5414 24942 5466
rect 24942 5414 24988 5466
rect 24692 5412 24748 5414
rect 24772 5412 24828 5414
rect 24852 5412 24908 5414
rect 24932 5412 24988 5414
rect 24692 4378 24748 4380
rect 24772 4378 24828 4380
rect 24852 4378 24908 4380
rect 24932 4378 24988 4380
rect 24692 4326 24738 4378
rect 24738 4326 24748 4378
rect 24772 4326 24802 4378
rect 24802 4326 24814 4378
rect 24814 4326 24828 4378
rect 24852 4326 24866 4378
rect 24866 4326 24878 4378
rect 24878 4326 24908 4378
rect 24932 4326 24942 4378
rect 24942 4326 24988 4378
rect 24692 4324 24748 4326
rect 24772 4324 24828 4326
rect 24852 4324 24908 4326
rect 24932 4324 24988 4326
rect 24692 3290 24748 3292
rect 24772 3290 24828 3292
rect 24852 3290 24908 3292
rect 24932 3290 24988 3292
rect 24692 3238 24738 3290
rect 24738 3238 24748 3290
rect 24772 3238 24802 3290
rect 24802 3238 24814 3290
rect 24814 3238 24828 3290
rect 24852 3238 24866 3290
rect 24866 3238 24878 3290
rect 24878 3238 24908 3290
rect 24932 3238 24942 3290
rect 24942 3238 24988 3290
rect 24692 3236 24748 3238
rect 24772 3236 24828 3238
rect 24852 3236 24908 3238
rect 24932 3236 24988 3238
rect 23938 856 23994 912
rect 24692 2202 24748 2204
rect 24772 2202 24828 2204
rect 24852 2202 24908 2204
rect 24932 2202 24988 2204
rect 24692 2150 24738 2202
rect 24738 2150 24748 2202
rect 24772 2150 24802 2202
rect 24802 2150 24814 2202
rect 24814 2150 24828 2202
rect 24852 2150 24866 2202
rect 24866 2150 24878 2202
rect 24878 2150 24908 2202
rect 24932 2150 24942 2202
rect 24942 2150 24988 2202
rect 24692 2148 24748 2150
rect 24772 2148 24828 2150
rect 24852 2148 24908 2150
rect 24932 2148 24988 2150
rect 24692 1114 24748 1116
rect 24772 1114 24828 1116
rect 24852 1114 24908 1116
rect 24932 1114 24988 1116
rect 24692 1062 24738 1114
rect 24738 1062 24748 1114
rect 24772 1062 24802 1114
rect 24802 1062 24814 1114
rect 24814 1062 24828 1114
rect 24852 1062 24866 1114
rect 24866 1062 24878 1114
rect 24878 1062 24908 1114
rect 24932 1062 24942 1114
rect 24942 1062 24988 1114
rect 24692 1060 24748 1062
rect 24772 1060 24828 1062
rect 24852 1060 24908 1062
rect 24932 1060 24988 1062
<< metal3 >>
rect 6880 6560 7196 6561
rect 6880 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7196 6560
rect 6880 6495 7196 6496
rect 12814 6560 13130 6561
rect 12814 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13130 6560
rect 12814 6495 13130 6496
rect 18748 6560 19064 6561
rect 18748 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19064 6560
rect 18748 6495 19064 6496
rect 24682 6560 24998 6561
rect 24682 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 24998 6560
rect 24682 6495 24998 6496
rect 2221 6354 2287 6357
rect 20662 6354 20668 6356
rect 2221 6352 20668 6354
rect 2221 6296 2226 6352
rect 2282 6296 20668 6352
rect 2221 6294 20668 6296
rect 2221 6291 2287 6294
rect 20662 6292 20668 6294
rect 20732 6292 20738 6356
rect 3913 6016 4229 6017
rect 3913 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4229 6016
rect 3913 5951 4229 5952
rect 9847 6016 10163 6017
rect 9847 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10163 6016
rect 9847 5951 10163 5952
rect 15781 6016 16097 6017
rect 15781 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16097 6016
rect 15781 5951 16097 5952
rect 21715 6016 22031 6017
rect 21715 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22031 6016
rect 21715 5951 22031 5952
rect 6880 5472 7196 5473
rect 6880 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7196 5472
rect 6880 5407 7196 5408
rect 12814 5472 13130 5473
rect 12814 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13130 5472
rect 12814 5407 13130 5408
rect 18748 5472 19064 5473
rect 18748 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19064 5472
rect 18748 5407 19064 5408
rect 24682 5472 24998 5473
rect 24682 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 24998 5472
rect 24682 5407 24998 5408
rect 9581 5130 9647 5133
rect 22134 5130 22140 5132
rect 9581 5128 22140 5130
rect 9581 5072 9586 5128
rect 9642 5072 22140 5128
rect 9581 5070 22140 5072
rect 9581 5067 9647 5070
rect 22134 5068 22140 5070
rect 22204 5068 22210 5132
rect 3913 4928 4229 4929
rect 3913 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4229 4928
rect 3913 4863 4229 4864
rect 9847 4928 10163 4929
rect 9847 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10163 4928
rect 9847 4863 10163 4864
rect 15781 4928 16097 4929
rect 15781 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16097 4928
rect 15781 4863 16097 4864
rect 21715 4928 22031 4929
rect 21715 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22031 4928
rect 21715 4863 22031 4864
rect 13721 4722 13787 4725
rect 22318 4722 22324 4724
rect 13721 4720 22324 4722
rect 13721 4664 13726 4720
rect 13782 4664 22324 4720
rect 13721 4662 22324 4664
rect 13721 4659 13787 4662
rect 22318 4660 22324 4662
rect 22388 4660 22394 4724
rect 6880 4384 7196 4385
rect 6880 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7196 4384
rect 6880 4319 7196 4320
rect 12814 4384 13130 4385
rect 12814 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13130 4384
rect 12814 4319 13130 4320
rect 18748 4384 19064 4385
rect 18748 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19064 4384
rect 18748 4319 19064 4320
rect 24682 4384 24998 4385
rect 24682 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 24998 4384
rect 24682 4319 24998 4320
rect 11237 4178 11303 4181
rect 15142 4178 15148 4180
rect 11237 4176 15148 4178
rect 11237 4120 11242 4176
rect 11298 4120 15148 4176
rect 11237 4118 15148 4120
rect 11237 4115 11303 4118
rect 15142 4116 15148 4118
rect 15212 4116 15218 4180
rect 3913 3840 4229 3841
rect 3913 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4229 3840
rect 3913 3775 4229 3776
rect 9847 3840 10163 3841
rect 9847 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10163 3840
rect 9847 3775 10163 3776
rect 15781 3840 16097 3841
rect 15781 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16097 3840
rect 15781 3775 16097 3776
rect 21715 3840 22031 3841
rect 21715 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22031 3840
rect 21715 3775 22031 3776
rect 6880 3296 7196 3297
rect 6880 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7196 3296
rect 6880 3231 7196 3232
rect 12814 3296 13130 3297
rect 12814 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13130 3296
rect 12814 3231 13130 3232
rect 18748 3296 19064 3297
rect 18748 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19064 3296
rect 18748 3231 19064 3232
rect 24682 3296 24998 3297
rect 24682 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 24998 3296
rect 24682 3231 24998 3232
rect 7465 3090 7531 3093
rect 7465 3088 16866 3090
rect 7465 3032 7470 3088
rect 7526 3032 16866 3088
rect 7465 3030 16866 3032
rect 7465 3027 7531 3030
rect 9029 2954 9095 2957
rect 12249 2954 12315 2957
rect 9029 2952 12315 2954
rect 9029 2896 9034 2952
rect 9090 2896 12254 2952
rect 12310 2896 12315 2952
rect 9029 2894 12315 2896
rect 9029 2891 9095 2894
rect 12249 2891 12315 2894
rect 16806 2818 16866 3030
rect 21173 2818 21239 2821
rect 16806 2816 21239 2818
rect 16806 2760 21178 2816
rect 21234 2760 21239 2816
rect 16806 2758 21239 2760
rect 21173 2755 21239 2758
rect 3913 2752 4229 2753
rect 3913 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4229 2752
rect 3913 2687 4229 2688
rect 9847 2752 10163 2753
rect 9847 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10163 2752
rect 9847 2687 10163 2688
rect 15781 2752 16097 2753
rect 15781 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16097 2752
rect 15781 2687 16097 2688
rect 21715 2752 22031 2753
rect 21715 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22031 2752
rect 21715 2687 22031 2688
rect 10225 2682 10291 2685
rect 14549 2682 14615 2685
rect 10225 2680 14615 2682
rect 10225 2624 10230 2680
rect 10286 2624 14554 2680
rect 14610 2624 14615 2680
rect 10225 2622 14615 2624
rect 10225 2619 10291 2622
rect 14549 2619 14615 2622
rect 7189 2546 7255 2549
rect 18137 2546 18203 2549
rect 7189 2544 18203 2546
rect 7189 2488 7194 2544
rect 7250 2488 18142 2544
rect 18198 2488 18203 2544
rect 7189 2486 18203 2488
rect 7189 2483 7255 2486
rect 18137 2483 18203 2486
rect 6269 2410 6335 2413
rect 19701 2410 19767 2413
rect 6269 2408 19767 2410
rect 6269 2352 6274 2408
rect 6330 2352 19706 2408
rect 19762 2352 19767 2408
rect 6269 2350 19767 2352
rect 6269 2347 6335 2350
rect 19701 2347 19767 2350
rect 22318 2348 22324 2412
rect 22388 2410 22394 2412
rect 23197 2410 23263 2413
rect 22388 2408 23263 2410
rect 22388 2352 23202 2408
rect 23258 2352 23263 2408
rect 22388 2350 23263 2352
rect 22388 2348 22394 2350
rect 23197 2347 23263 2350
rect 7833 2274 7899 2277
rect 10225 2274 10291 2277
rect 7833 2272 10291 2274
rect 7833 2216 7838 2272
rect 7894 2216 10230 2272
rect 10286 2216 10291 2272
rect 7833 2214 10291 2216
rect 7833 2211 7899 2214
rect 10225 2211 10291 2214
rect 20662 2212 20668 2276
rect 20732 2274 20738 2276
rect 20897 2274 20963 2277
rect 20732 2272 20963 2274
rect 20732 2216 20902 2272
rect 20958 2216 20963 2272
rect 20732 2214 20963 2216
rect 20732 2212 20738 2214
rect 20897 2211 20963 2214
rect 22134 2212 22140 2276
rect 22204 2274 22210 2276
rect 22277 2274 22343 2277
rect 22204 2272 22343 2274
rect 22204 2216 22282 2272
rect 22338 2216 22343 2272
rect 22204 2214 22343 2216
rect 22204 2212 22210 2214
rect 22277 2211 22343 2214
rect 6880 2208 7196 2209
rect 6880 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7196 2208
rect 6880 2143 7196 2144
rect 12814 2208 13130 2209
rect 12814 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13130 2208
rect 12814 2143 13130 2144
rect 18748 2208 19064 2209
rect 18748 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19064 2208
rect 18748 2143 19064 2144
rect 24682 2208 24998 2209
rect 24682 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 24998 2208
rect 24682 2143 24998 2144
rect 8293 2138 8359 2141
rect 8293 2136 12634 2138
rect 8293 2080 8298 2136
rect 8354 2080 12634 2136
rect 8293 2078 12634 2080
rect 8293 2075 8359 2078
rect 2405 2002 2471 2005
rect 12433 2002 12499 2005
rect 2405 2000 12499 2002
rect 2405 1944 2410 2000
rect 2466 1944 12438 2000
rect 12494 1944 12499 2000
rect 2405 1942 12499 1944
rect 12574 2002 12634 2078
rect 14089 2002 14155 2005
rect 12574 2000 14155 2002
rect 12574 1944 14094 2000
rect 14150 1944 14155 2000
rect 12574 1942 14155 1944
rect 2405 1939 2471 1942
rect 12433 1939 12499 1942
rect 14089 1939 14155 1942
rect 5901 1866 5967 1869
rect 20253 1866 20319 1869
rect 2730 1806 5090 1866
rect 1945 1730 2011 1733
rect 2730 1730 2790 1806
rect 1945 1728 2790 1730
rect 1945 1672 1950 1728
rect 2006 1672 2790 1728
rect 1945 1670 2790 1672
rect 5030 1730 5090 1806
rect 5901 1864 20319 1866
rect 5901 1808 5906 1864
rect 5962 1808 20258 1864
rect 20314 1808 20319 1864
rect 5901 1806 20319 1808
rect 5901 1803 5967 1806
rect 20253 1803 20319 1806
rect 8293 1730 8359 1733
rect 5030 1728 8359 1730
rect 5030 1672 8298 1728
rect 8354 1672 8359 1728
rect 5030 1670 8359 1672
rect 1945 1667 2011 1670
rect 8293 1667 8359 1670
rect 13537 1730 13603 1733
rect 15193 1730 15259 1733
rect 13537 1728 15259 1730
rect 13537 1672 13542 1728
rect 13598 1672 15198 1728
rect 15254 1672 15259 1728
rect 13537 1670 15259 1672
rect 13537 1667 13603 1670
rect 15193 1667 15259 1670
rect 3913 1664 4229 1665
rect 3913 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4229 1664
rect 3913 1599 4229 1600
rect 9847 1664 10163 1665
rect 9847 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10163 1664
rect 9847 1599 10163 1600
rect 15781 1664 16097 1665
rect 15781 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16097 1664
rect 15781 1599 16097 1600
rect 21715 1664 22031 1665
rect 21715 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22031 1664
rect 21715 1599 22031 1600
rect 2957 1458 3023 1461
rect 10317 1458 10383 1461
rect 2957 1456 10383 1458
rect 2957 1400 2962 1456
rect 3018 1400 10322 1456
rect 10378 1400 10383 1456
rect 2957 1398 10383 1400
rect 2957 1395 3023 1398
rect 10317 1395 10383 1398
rect 2313 1322 2379 1325
rect 5073 1322 5139 1325
rect 12801 1322 12867 1325
rect 2313 1320 2790 1322
rect 2313 1264 2318 1320
rect 2374 1264 2790 1320
rect 2313 1262 2790 1264
rect 2313 1259 2379 1262
rect 2730 914 2790 1262
rect 5073 1320 12867 1322
rect 5073 1264 5078 1320
rect 5134 1264 12806 1320
rect 12862 1264 12867 1320
rect 5073 1262 12867 1264
rect 5073 1259 5139 1262
rect 12801 1259 12867 1262
rect 7833 1186 7899 1189
rect 9857 1186 9923 1189
rect 7833 1184 9923 1186
rect 7833 1128 7838 1184
rect 7894 1128 9862 1184
rect 9918 1128 9923 1184
rect 7833 1126 9923 1128
rect 7833 1123 7899 1126
rect 9857 1123 9923 1126
rect 6880 1120 7196 1121
rect 6880 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7196 1120
rect 6880 1055 7196 1056
rect 12814 1120 13130 1121
rect 12814 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13130 1120
rect 12814 1055 13130 1056
rect 18748 1120 19064 1121
rect 18748 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19064 1120
rect 18748 1055 19064 1056
rect 24682 1120 24998 1121
rect 24682 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 24998 1120
rect 24682 1055 24998 1056
rect 11697 914 11763 917
rect 2730 912 11763 914
rect 2730 856 11702 912
rect 11758 856 11763 912
rect 2730 854 11763 856
rect 11697 851 11763 854
rect 15142 852 15148 916
rect 15212 914 15218 916
rect 23933 914 23999 917
rect 15212 912 23999 914
rect 15212 856 23938 912
rect 23994 856 23999 912
rect 15212 854 23999 856
rect 15212 852 15218 854
rect 23933 851 23999 854
rect 5901 778 5967 781
rect 18321 778 18387 781
rect 5901 776 18387 778
rect 5901 720 5906 776
rect 5962 720 18326 776
rect 18382 720 18387 776
rect 5901 718 18387 720
rect 5901 715 5967 718
rect 18321 715 18387 718
rect 6177 642 6243 645
rect 18045 642 18111 645
rect 6177 640 18111 642
rect 6177 584 6182 640
rect 6238 584 18050 640
rect 18106 584 18111 640
rect 6177 582 18111 584
rect 6177 579 6243 582
rect 18045 579 18111 582
rect 7833 506 7899 509
rect 21817 506 21883 509
rect 7833 504 21883 506
rect 7833 448 7838 504
rect 7894 448 21822 504
rect 21878 448 21883 504
rect 7833 446 21883 448
rect 7833 443 7899 446
rect 21817 443 21883 446
rect 1945 370 2011 373
rect 5901 370 5967 373
rect 10501 370 10567 373
rect 11973 370 12039 373
rect 1945 368 2790 370
rect 1945 312 1950 368
rect 2006 312 2790 368
rect 1945 310 2790 312
rect 1945 307 2011 310
rect 2730 234 2790 310
rect 5901 368 10567 370
rect 5901 312 5906 368
rect 5962 312 10506 368
rect 10562 312 10567 368
rect 5901 310 10567 312
rect 5901 307 5967 310
rect 10501 307 10567 310
rect 10734 368 12039 370
rect 10734 312 11978 368
rect 12034 312 12039 368
rect 10734 310 12039 312
rect 10734 234 10794 310
rect 11973 307 12039 310
rect 2730 174 10794 234
<< via3 >>
rect 6886 6556 6950 6560
rect 6886 6500 6890 6556
rect 6890 6500 6946 6556
rect 6946 6500 6950 6556
rect 6886 6496 6950 6500
rect 6966 6556 7030 6560
rect 6966 6500 6970 6556
rect 6970 6500 7026 6556
rect 7026 6500 7030 6556
rect 6966 6496 7030 6500
rect 7046 6556 7110 6560
rect 7046 6500 7050 6556
rect 7050 6500 7106 6556
rect 7106 6500 7110 6556
rect 7046 6496 7110 6500
rect 7126 6556 7190 6560
rect 7126 6500 7130 6556
rect 7130 6500 7186 6556
rect 7186 6500 7190 6556
rect 7126 6496 7190 6500
rect 12820 6556 12884 6560
rect 12820 6500 12824 6556
rect 12824 6500 12880 6556
rect 12880 6500 12884 6556
rect 12820 6496 12884 6500
rect 12900 6556 12964 6560
rect 12900 6500 12904 6556
rect 12904 6500 12960 6556
rect 12960 6500 12964 6556
rect 12900 6496 12964 6500
rect 12980 6556 13044 6560
rect 12980 6500 12984 6556
rect 12984 6500 13040 6556
rect 13040 6500 13044 6556
rect 12980 6496 13044 6500
rect 13060 6556 13124 6560
rect 13060 6500 13064 6556
rect 13064 6500 13120 6556
rect 13120 6500 13124 6556
rect 13060 6496 13124 6500
rect 18754 6556 18818 6560
rect 18754 6500 18758 6556
rect 18758 6500 18814 6556
rect 18814 6500 18818 6556
rect 18754 6496 18818 6500
rect 18834 6556 18898 6560
rect 18834 6500 18838 6556
rect 18838 6500 18894 6556
rect 18894 6500 18898 6556
rect 18834 6496 18898 6500
rect 18914 6556 18978 6560
rect 18914 6500 18918 6556
rect 18918 6500 18974 6556
rect 18974 6500 18978 6556
rect 18914 6496 18978 6500
rect 18994 6556 19058 6560
rect 18994 6500 18998 6556
rect 18998 6500 19054 6556
rect 19054 6500 19058 6556
rect 18994 6496 19058 6500
rect 24688 6556 24752 6560
rect 24688 6500 24692 6556
rect 24692 6500 24748 6556
rect 24748 6500 24752 6556
rect 24688 6496 24752 6500
rect 24768 6556 24832 6560
rect 24768 6500 24772 6556
rect 24772 6500 24828 6556
rect 24828 6500 24832 6556
rect 24768 6496 24832 6500
rect 24848 6556 24912 6560
rect 24848 6500 24852 6556
rect 24852 6500 24908 6556
rect 24908 6500 24912 6556
rect 24848 6496 24912 6500
rect 24928 6556 24992 6560
rect 24928 6500 24932 6556
rect 24932 6500 24988 6556
rect 24988 6500 24992 6556
rect 24928 6496 24992 6500
rect 20668 6292 20732 6356
rect 3919 6012 3983 6016
rect 3919 5956 3923 6012
rect 3923 5956 3979 6012
rect 3979 5956 3983 6012
rect 3919 5952 3983 5956
rect 3999 6012 4063 6016
rect 3999 5956 4003 6012
rect 4003 5956 4059 6012
rect 4059 5956 4063 6012
rect 3999 5952 4063 5956
rect 4079 6012 4143 6016
rect 4079 5956 4083 6012
rect 4083 5956 4139 6012
rect 4139 5956 4143 6012
rect 4079 5952 4143 5956
rect 4159 6012 4223 6016
rect 4159 5956 4163 6012
rect 4163 5956 4219 6012
rect 4219 5956 4223 6012
rect 4159 5952 4223 5956
rect 9853 6012 9917 6016
rect 9853 5956 9857 6012
rect 9857 5956 9913 6012
rect 9913 5956 9917 6012
rect 9853 5952 9917 5956
rect 9933 6012 9997 6016
rect 9933 5956 9937 6012
rect 9937 5956 9993 6012
rect 9993 5956 9997 6012
rect 9933 5952 9997 5956
rect 10013 6012 10077 6016
rect 10013 5956 10017 6012
rect 10017 5956 10073 6012
rect 10073 5956 10077 6012
rect 10013 5952 10077 5956
rect 10093 6012 10157 6016
rect 10093 5956 10097 6012
rect 10097 5956 10153 6012
rect 10153 5956 10157 6012
rect 10093 5952 10157 5956
rect 15787 6012 15851 6016
rect 15787 5956 15791 6012
rect 15791 5956 15847 6012
rect 15847 5956 15851 6012
rect 15787 5952 15851 5956
rect 15867 6012 15931 6016
rect 15867 5956 15871 6012
rect 15871 5956 15927 6012
rect 15927 5956 15931 6012
rect 15867 5952 15931 5956
rect 15947 6012 16011 6016
rect 15947 5956 15951 6012
rect 15951 5956 16007 6012
rect 16007 5956 16011 6012
rect 15947 5952 16011 5956
rect 16027 6012 16091 6016
rect 16027 5956 16031 6012
rect 16031 5956 16087 6012
rect 16087 5956 16091 6012
rect 16027 5952 16091 5956
rect 21721 6012 21785 6016
rect 21721 5956 21725 6012
rect 21725 5956 21781 6012
rect 21781 5956 21785 6012
rect 21721 5952 21785 5956
rect 21801 6012 21865 6016
rect 21801 5956 21805 6012
rect 21805 5956 21861 6012
rect 21861 5956 21865 6012
rect 21801 5952 21865 5956
rect 21881 6012 21945 6016
rect 21881 5956 21885 6012
rect 21885 5956 21941 6012
rect 21941 5956 21945 6012
rect 21881 5952 21945 5956
rect 21961 6012 22025 6016
rect 21961 5956 21965 6012
rect 21965 5956 22021 6012
rect 22021 5956 22025 6012
rect 21961 5952 22025 5956
rect 6886 5468 6950 5472
rect 6886 5412 6890 5468
rect 6890 5412 6946 5468
rect 6946 5412 6950 5468
rect 6886 5408 6950 5412
rect 6966 5468 7030 5472
rect 6966 5412 6970 5468
rect 6970 5412 7026 5468
rect 7026 5412 7030 5468
rect 6966 5408 7030 5412
rect 7046 5468 7110 5472
rect 7046 5412 7050 5468
rect 7050 5412 7106 5468
rect 7106 5412 7110 5468
rect 7046 5408 7110 5412
rect 7126 5468 7190 5472
rect 7126 5412 7130 5468
rect 7130 5412 7186 5468
rect 7186 5412 7190 5468
rect 7126 5408 7190 5412
rect 12820 5468 12884 5472
rect 12820 5412 12824 5468
rect 12824 5412 12880 5468
rect 12880 5412 12884 5468
rect 12820 5408 12884 5412
rect 12900 5468 12964 5472
rect 12900 5412 12904 5468
rect 12904 5412 12960 5468
rect 12960 5412 12964 5468
rect 12900 5408 12964 5412
rect 12980 5468 13044 5472
rect 12980 5412 12984 5468
rect 12984 5412 13040 5468
rect 13040 5412 13044 5468
rect 12980 5408 13044 5412
rect 13060 5468 13124 5472
rect 13060 5412 13064 5468
rect 13064 5412 13120 5468
rect 13120 5412 13124 5468
rect 13060 5408 13124 5412
rect 18754 5468 18818 5472
rect 18754 5412 18758 5468
rect 18758 5412 18814 5468
rect 18814 5412 18818 5468
rect 18754 5408 18818 5412
rect 18834 5468 18898 5472
rect 18834 5412 18838 5468
rect 18838 5412 18894 5468
rect 18894 5412 18898 5468
rect 18834 5408 18898 5412
rect 18914 5468 18978 5472
rect 18914 5412 18918 5468
rect 18918 5412 18974 5468
rect 18974 5412 18978 5468
rect 18914 5408 18978 5412
rect 18994 5468 19058 5472
rect 18994 5412 18998 5468
rect 18998 5412 19054 5468
rect 19054 5412 19058 5468
rect 18994 5408 19058 5412
rect 24688 5468 24752 5472
rect 24688 5412 24692 5468
rect 24692 5412 24748 5468
rect 24748 5412 24752 5468
rect 24688 5408 24752 5412
rect 24768 5468 24832 5472
rect 24768 5412 24772 5468
rect 24772 5412 24828 5468
rect 24828 5412 24832 5468
rect 24768 5408 24832 5412
rect 24848 5468 24912 5472
rect 24848 5412 24852 5468
rect 24852 5412 24908 5468
rect 24908 5412 24912 5468
rect 24848 5408 24912 5412
rect 24928 5468 24992 5472
rect 24928 5412 24932 5468
rect 24932 5412 24988 5468
rect 24988 5412 24992 5468
rect 24928 5408 24992 5412
rect 22140 5068 22204 5132
rect 3919 4924 3983 4928
rect 3919 4868 3923 4924
rect 3923 4868 3979 4924
rect 3979 4868 3983 4924
rect 3919 4864 3983 4868
rect 3999 4924 4063 4928
rect 3999 4868 4003 4924
rect 4003 4868 4059 4924
rect 4059 4868 4063 4924
rect 3999 4864 4063 4868
rect 4079 4924 4143 4928
rect 4079 4868 4083 4924
rect 4083 4868 4139 4924
rect 4139 4868 4143 4924
rect 4079 4864 4143 4868
rect 4159 4924 4223 4928
rect 4159 4868 4163 4924
rect 4163 4868 4219 4924
rect 4219 4868 4223 4924
rect 4159 4864 4223 4868
rect 9853 4924 9917 4928
rect 9853 4868 9857 4924
rect 9857 4868 9913 4924
rect 9913 4868 9917 4924
rect 9853 4864 9917 4868
rect 9933 4924 9997 4928
rect 9933 4868 9937 4924
rect 9937 4868 9993 4924
rect 9993 4868 9997 4924
rect 9933 4864 9997 4868
rect 10013 4924 10077 4928
rect 10013 4868 10017 4924
rect 10017 4868 10073 4924
rect 10073 4868 10077 4924
rect 10013 4864 10077 4868
rect 10093 4924 10157 4928
rect 10093 4868 10097 4924
rect 10097 4868 10153 4924
rect 10153 4868 10157 4924
rect 10093 4864 10157 4868
rect 15787 4924 15851 4928
rect 15787 4868 15791 4924
rect 15791 4868 15847 4924
rect 15847 4868 15851 4924
rect 15787 4864 15851 4868
rect 15867 4924 15931 4928
rect 15867 4868 15871 4924
rect 15871 4868 15927 4924
rect 15927 4868 15931 4924
rect 15867 4864 15931 4868
rect 15947 4924 16011 4928
rect 15947 4868 15951 4924
rect 15951 4868 16007 4924
rect 16007 4868 16011 4924
rect 15947 4864 16011 4868
rect 16027 4924 16091 4928
rect 16027 4868 16031 4924
rect 16031 4868 16087 4924
rect 16087 4868 16091 4924
rect 16027 4864 16091 4868
rect 21721 4924 21785 4928
rect 21721 4868 21725 4924
rect 21725 4868 21781 4924
rect 21781 4868 21785 4924
rect 21721 4864 21785 4868
rect 21801 4924 21865 4928
rect 21801 4868 21805 4924
rect 21805 4868 21861 4924
rect 21861 4868 21865 4924
rect 21801 4864 21865 4868
rect 21881 4924 21945 4928
rect 21881 4868 21885 4924
rect 21885 4868 21941 4924
rect 21941 4868 21945 4924
rect 21881 4864 21945 4868
rect 21961 4924 22025 4928
rect 21961 4868 21965 4924
rect 21965 4868 22021 4924
rect 22021 4868 22025 4924
rect 21961 4864 22025 4868
rect 22324 4660 22388 4724
rect 6886 4380 6950 4384
rect 6886 4324 6890 4380
rect 6890 4324 6946 4380
rect 6946 4324 6950 4380
rect 6886 4320 6950 4324
rect 6966 4380 7030 4384
rect 6966 4324 6970 4380
rect 6970 4324 7026 4380
rect 7026 4324 7030 4380
rect 6966 4320 7030 4324
rect 7046 4380 7110 4384
rect 7046 4324 7050 4380
rect 7050 4324 7106 4380
rect 7106 4324 7110 4380
rect 7046 4320 7110 4324
rect 7126 4380 7190 4384
rect 7126 4324 7130 4380
rect 7130 4324 7186 4380
rect 7186 4324 7190 4380
rect 7126 4320 7190 4324
rect 12820 4380 12884 4384
rect 12820 4324 12824 4380
rect 12824 4324 12880 4380
rect 12880 4324 12884 4380
rect 12820 4320 12884 4324
rect 12900 4380 12964 4384
rect 12900 4324 12904 4380
rect 12904 4324 12960 4380
rect 12960 4324 12964 4380
rect 12900 4320 12964 4324
rect 12980 4380 13044 4384
rect 12980 4324 12984 4380
rect 12984 4324 13040 4380
rect 13040 4324 13044 4380
rect 12980 4320 13044 4324
rect 13060 4380 13124 4384
rect 13060 4324 13064 4380
rect 13064 4324 13120 4380
rect 13120 4324 13124 4380
rect 13060 4320 13124 4324
rect 18754 4380 18818 4384
rect 18754 4324 18758 4380
rect 18758 4324 18814 4380
rect 18814 4324 18818 4380
rect 18754 4320 18818 4324
rect 18834 4380 18898 4384
rect 18834 4324 18838 4380
rect 18838 4324 18894 4380
rect 18894 4324 18898 4380
rect 18834 4320 18898 4324
rect 18914 4380 18978 4384
rect 18914 4324 18918 4380
rect 18918 4324 18974 4380
rect 18974 4324 18978 4380
rect 18914 4320 18978 4324
rect 18994 4380 19058 4384
rect 18994 4324 18998 4380
rect 18998 4324 19054 4380
rect 19054 4324 19058 4380
rect 18994 4320 19058 4324
rect 24688 4380 24752 4384
rect 24688 4324 24692 4380
rect 24692 4324 24748 4380
rect 24748 4324 24752 4380
rect 24688 4320 24752 4324
rect 24768 4380 24832 4384
rect 24768 4324 24772 4380
rect 24772 4324 24828 4380
rect 24828 4324 24832 4380
rect 24768 4320 24832 4324
rect 24848 4380 24912 4384
rect 24848 4324 24852 4380
rect 24852 4324 24908 4380
rect 24908 4324 24912 4380
rect 24848 4320 24912 4324
rect 24928 4380 24992 4384
rect 24928 4324 24932 4380
rect 24932 4324 24988 4380
rect 24988 4324 24992 4380
rect 24928 4320 24992 4324
rect 15148 4116 15212 4180
rect 3919 3836 3983 3840
rect 3919 3780 3923 3836
rect 3923 3780 3979 3836
rect 3979 3780 3983 3836
rect 3919 3776 3983 3780
rect 3999 3836 4063 3840
rect 3999 3780 4003 3836
rect 4003 3780 4059 3836
rect 4059 3780 4063 3836
rect 3999 3776 4063 3780
rect 4079 3836 4143 3840
rect 4079 3780 4083 3836
rect 4083 3780 4139 3836
rect 4139 3780 4143 3836
rect 4079 3776 4143 3780
rect 4159 3836 4223 3840
rect 4159 3780 4163 3836
rect 4163 3780 4219 3836
rect 4219 3780 4223 3836
rect 4159 3776 4223 3780
rect 9853 3836 9917 3840
rect 9853 3780 9857 3836
rect 9857 3780 9913 3836
rect 9913 3780 9917 3836
rect 9853 3776 9917 3780
rect 9933 3836 9997 3840
rect 9933 3780 9937 3836
rect 9937 3780 9993 3836
rect 9993 3780 9997 3836
rect 9933 3776 9997 3780
rect 10013 3836 10077 3840
rect 10013 3780 10017 3836
rect 10017 3780 10073 3836
rect 10073 3780 10077 3836
rect 10013 3776 10077 3780
rect 10093 3836 10157 3840
rect 10093 3780 10097 3836
rect 10097 3780 10153 3836
rect 10153 3780 10157 3836
rect 10093 3776 10157 3780
rect 15787 3836 15851 3840
rect 15787 3780 15791 3836
rect 15791 3780 15847 3836
rect 15847 3780 15851 3836
rect 15787 3776 15851 3780
rect 15867 3836 15931 3840
rect 15867 3780 15871 3836
rect 15871 3780 15927 3836
rect 15927 3780 15931 3836
rect 15867 3776 15931 3780
rect 15947 3836 16011 3840
rect 15947 3780 15951 3836
rect 15951 3780 16007 3836
rect 16007 3780 16011 3836
rect 15947 3776 16011 3780
rect 16027 3836 16091 3840
rect 16027 3780 16031 3836
rect 16031 3780 16087 3836
rect 16087 3780 16091 3836
rect 16027 3776 16091 3780
rect 21721 3836 21785 3840
rect 21721 3780 21725 3836
rect 21725 3780 21781 3836
rect 21781 3780 21785 3836
rect 21721 3776 21785 3780
rect 21801 3836 21865 3840
rect 21801 3780 21805 3836
rect 21805 3780 21861 3836
rect 21861 3780 21865 3836
rect 21801 3776 21865 3780
rect 21881 3836 21945 3840
rect 21881 3780 21885 3836
rect 21885 3780 21941 3836
rect 21941 3780 21945 3836
rect 21881 3776 21945 3780
rect 21961 3836 22025 3840
rect 21961 3780 21965 3836
rect 21965 3780 22021 3836
rect 22021 3780 22025 3836
rect 21961 3776 22025 3780
rect 6886 3292 6950 3296
rect 6886 3236 6890 3292
rect 6890 3236 6946 3292
rect 6946 3236 6950 3292
rect 6886 3232 6950 3236
rect 6966 3292 7030 3296
rect 6966 3236 6970 3292
rect 6970 3236 7026 3292
rect 7026 3236 7030 3292
rect 6966 3232 7030 3236
rect 7046 3292 7110 3296
rect 7046 3236 7050 3292
rect 7050 3236 7106 3292
rect 7106 3236 7110 3292
rect 7046 3232 7110 3236
rect 7126 3292 7190 3296
rect 7126 3236 7130 3292
rect 7130 3236 7186 3292
rect 7186 3236 7190 3292
rect 7126 3232 7190 3236
rect 12820 3292 12884 3296
rect 12820 3236 12824 3292
rect 12824 3236 12880 3292
rect 12880 3236 12884 3292
rect 12820 3232 12884 3236
rect 12900 3292 12964 3296
rect 12900 3236 12904 3292
rect 12904 3236 12960 3292
rect 12960 3236 12964 3292
rect 12900 3232 12964 3236
rect 12980 3292 13044 3296
rect 12980 3236 12984 3292
rect 12984 3236 13040 3292
rect 13040 3236 13044 3292
rect 12980 3232 13044 3236
rect 13060 3292 13124 3296
rect 13060 3236 13064 3292
rect 13064 3236 13120 3292
rect 13120 3236 13124 3292
rect 13060 3232 13124 3236
rect 18754 3292 18818 3296
rect 18754 3236 18758 3292
rect 18758 3236 18814 3292
rect 18814 3236 18818 3292
rect 18754 3232 18818 3236
rect 18834 3292 18898 3296
rect 18834 3236 18838 3292
rect 18838 3236 18894 3292
rect 18894 3236 18898 3292
rect 18834 3232 18898 3236
rect 18914 3292 18978 3296
rect 18914 3236 18918 3292
rect 18918 3236 18974 3292
rect 18974 3236 18978 3292
rect 18914 3232 18978 3236
rect 18994 3292 19058 3296
rect 18994 3236 18998 3292
rect 18998 3236 19054 3292
rect 19054 3236 19058 3292
rect 18994 3232 19058 3236
rect 24688 3292 24752 3296
rect 24688 3236 24692 3292
rect 24692 3236 24748 3292
rect 24748 3236 24752 3292
rect 24688 3232 24752 3236
rect 24768 3292 24832 3296
rect 24768 3236 24772 3292
rect 24772 3236 24828 3292
rect 24828 3236 24832 3292
rect 24768 3232 24832 3236
rect 24848 3292 24912 3296
rect 24848 3236 24852 3292
rect 24852 3236 24908 3292
rect 24908 3236 24912 3292
rect 24848 3232 24912 3236
rect 24928 3292 24992 3296
rect 24928 3236 24932 3292
rect 24932 3236 24988 3292
rect 24988 3236 24992 3292
rect 24928 3232 24992 3236
rect 3919 2748 3983 2752
rect 3919 2692 3923 2748
rect 3923 2692 3979 2748
rect 3979 2692 3983 2748
rect 3919 2688 3983 2692
rect 3999 2748 4063 2752
rect 3999 2692 4003 2748
rect 4003 2692 4059 2748
rect 4059 2692 4063 2748
rect 3999 2688 4063 2692
rect 4079 2748 4143 2752
rect 4079 2692 4083 2748
rect 4083 2692 4139 2748
rect 4139 2692 4143 2748
rect 4079 2688 4143 2692
rect 4159 2748 4223 2752
rect 4159 2692 4163 2748
rect 4163 2692 4219 2748
rect 4219 2692 4223 2748
rect 4159 2688 4223 2692
rect 9853 2748 9917 2752
rect 9853 2692 9857 2748
rect 9857 2692 9913 2748
rect 9913 2692 9917 2748
rect 9853 2688 9917 2692
rect 9933 2748 9997 2752
rect 9933 2692 9937 2748
rect 9937 2692 9993 2748
rect 9993 2692 9997 2748
rect 9933 2688 9997 2692
rect 10013 2748 10077 2752
rect 10013 2692 10017 2748
rect 10017 2692 10073 2748
rect 10073 2692 10077 2748
rect 10013 2688 10077 2692
rect 10093 2748 10157 2752
rect 10093 2692 10097 2748
rect 10097 2692 10153 2748
rect 10153 2692 10157 2748
rect 10093 2688 10157 2692
rect 15787 2748 15851 2752
rect 15787 2692 15791 2748
rect 15791 2692 15847 2748
rect 15847 2692 15851 2748
rect 15787 2688 15851 2692
rect 15867 2748 15931 2752
rect 15867 2692 15871 2748
rect 15871 2692 15927 2748
rect 15927 2692 15931 2748
rect 15867 2688 15931 2692
rect 15947 2748 16011 2752
rect 15947 2692 15951 2748
rect 15951 2692 16007 2748
rect 16007 2692 16011 2748
rect 15947 2688 16011 2692
rect 16027 2748 16091 2752
rect 16027 2692 16031 2748
rect 16031 2692 16087 2748
rect 16087 2692 16091 2748
rect 16027 2688 16091 2692
rect 21721 2748 21785 2752
rect 21721 2692 21725 2748
rect 21725 2692 21781 2748
rect 21781 2692 21785 2748
rect 21721 2688 21785 2692
rect 21801 2748 21865 2752
rect 21801 2692 21805 2748
rect 21805 2692 21861 2748
rect 21861 2692 21865 2748
rect 21801 2688 21865 2692
rect 21881 2748 21945 2752
rect 21881 2692 21885 2748
rect 21885 2692 21941 2748
rect 21941 2692 21945 2748
rect 21881 2688 21945 2692
rect 21961 2748 22025 2752
rect 21961 2692 21965 2748
rect 21965 2692 22021 2748
rect 22021 2692 22025 2748
rect 21961 2688 22025 2692
rect 22324 2348 22388 2412
rect 20668 2212 20732 2276
rect 22140 2212 22204 2276
rect 6886 2204 6950 2208
rect 6886 2148 6890 2204
rect 6890 2148 6946 2204
rect 6946 2148 6950 2204
rect 6886 2144 6950 2148
rect 6966 2204 7030 2208
rect 6966 2148 6970 2204
rect 6970 2148 7026 2204
rect 7026 2148 7030 2204
rect 6966 2144 7030 2148
rect 7046 2204 7110 2208
rect 7046 2148 7050 2204
rect 7050 2148 7106 2204
rect 7106 2148 7110 2204
rect 7046 2144 7110 2148
rect 7126 2204 7190 2208
rect 7126 2148 7130 2204
rect 7130 2148 7186 2204
rect 7186 2148 7190 2204
rect 7126 2144 7190 2148
rect 12820 2204 12884 2208
rect 12820 2148 12824 2204
rect 12824 2148 12880 2204
rect 12880 2148 12884 2204
rect 12820 2144 12884 2148
rect 12900 2204 12964 2208
rect 12900 2148 12904 2204
rect 12904 2148 12960 2204
rect 12960 2148 12964 2204
rect 12900 2144 12964 2148
rect 12980 2204 13044 2208
rect 12980 2148 12984 2204
rect 12984 2148 13040 2204
rect 13040 2148 13044 2204
rect 12980 2144 13044 2148
rect 13060 2204 13124 2208
rect 13060 2148 13064 2204
rect 13064 2148 13120 2204
rect 13120 2148 13124 2204
rect 13060 2144 13124 2148
rect 18754 2204 18818 2208
rect 18754 2148 18758 2204
rect 18758 2148 18814 2204
rect 18814 2148 18818 2204
rect 18754 2144 18818 2148
rect 18834 2204 18898 2208
rect 18834 2148 18838 2204
rect 18838 2148 18894 2204
rect 18894 2148 18898 2204
rect 18834 2144 18898 2148
rect 18914 2204 18978 2208
rect 18914 2148 18918 2204
rect 18918 2148 18974 2204
rect 18974 2148 18978 2204
rect 18914 2144 18978 2148
rect 18994 2204 19058 2208
rect 18994 2148 18998 2204
rect 18998 2148 19054 2204
rect 19054 2148 19058 2204
rect 18994 2144 19058 2148
rect 24688 2204 24752 2208
rect 24688 2148 24692 2204
rect 24692 2148 24748 2204
rect 24748 2148 24752 2204
rect 24688 2144 24752 2148
rect 24768 2204 24832 2208
rect 24768 2148 24772 2204
rect 24772 2148 24828 2204
rect 24828 2148 24832 2204
rect 24768 2144 24832 2148
rect 24848 2204 24912 2208
rect 24848 2148 24852 2204
rect 24852 2148 24908 2204
rect 24908 2148 24912 2204
rect 24848 2144 24912 2148
rect 24928 2204 24992 2208
rect 24928 2148 24932 2204
rect 24932 2148 24988 2204
rect 24988 2148 24992 2204
rect 24928 2144 24992 2148
rect 3919 1660 3983 1664
rect 3919 1604 3923 1660
rect 3923 1604 3979 1660
rect 3979 1604 3983 1660
rect 3919 1600 3983 1604
rect 3999 1660 4063 1664
rect 3999 1604 4003 1660
rect 4003 1604 4059 1660
rect 4059 1604 4063 1660
rect 3999 1600 4063 1604
rect 4079 1660 4143 1664
rect 4079 1604 4083 1660
rect 4083 1604 4139 1660
rect 4139 1604 4143 1660
rect 4079 1600 4143 1604
rect 4159 1660 4223 1664
rect 4159 1604 4163 1660
rect 4163 1604 4219 1660
rect 4219 1604 4223 1660
rect 4159 1600 4223 1604
rect 9853 1660 9917 1664
rect 9853 1604 9857 1660
rect 9857 1604 9913 1660
rect 9913 1604 9917 1660
rect 9853 1600 9917 1604
rect 9933 1660 9997 1664
rect 9933 1604 9937 1660
rect 9937 1604 9993 1660
rect 9993 1604 9997 1660
rect 9933 1600 9997 1604
rect 10013 1660 10077 1664
rect 10013 1604 10017 1660
rect 10017 1604 10073 1660
rect 10073 1604 10077 1660
rect 10013 1600 10077 1604
rect 10093 1660 10157 1664
rect 10093 1604 10097 1660
rect 10097 1604 10153 1660
rect 10153 1604 10157 1660
rect 10093 1600 10157 1604
rect 15787 1660 15851 1664
rect 15787 1604 15791 1660
rect 15791 1604 15847 1660
rect 15847 1604 15851 1660
rect 15787 1600 15851 1604
rect 15867 1660 15931 1664
rect 15867 1604 15871 1660
rect 15871 1604 15927 1660
rect 15927 1604 15931 1660
rect 15867 1600 15931 1604
rect 15947 1660 16011 1664
rect 15947 1604 15951 1660
rect 15951 1604 16007 1660
rect 16007 1604 16011 1660
rect 15947 1600 16011 1604
rect 16027 1660 16091 1664
rect 16027 1604 16031 1660
rect 16031 1604 16087 1660
rect 16087 1604 16091 1660
rect 16027 1600 16091 1604
rect 21721 1660 21785 1664
rect 21721 1604 21725 1660
rect 21725 1604 21781 1660
rect 21781 1604 21785 1660
rect 21721 1600 21785 1604
rect 21801 1660 21865 1664
rect 21801 1604 21805 1660
rect 21805 1604 21861 1660
rect 21861 1604 21865 1660
rect 21801 1600 21865 1604
rect 21881 1660 21945 1664
rect 21881 1604 21885 1660
rect 21885 1604 21941 1660
rect 21941 1604 21945 1660
rect 21881 1600 21945 1604
rect 21961 1660 22025 1664
rect 21961 1604 21965 1660
rect 21965 1604 22021 1660
rect 22021 1604 22025 1660
rect 21961 1600 22025 1604
rect 6886 1116 6950 1120
rect 6886 1060 6890 1116
rect 6890 1060 6946 1116
rect 6946 1060 6950 1116
rect 6886 1056 6950 1060
rect 6966 1116 7030 1120
rect 6966 1060 6970 1116
rect 6970 1060 7026 1116
rect 7026 1060 7030 1116
rect 6966 1056 7030 1060
rect 7046 1116 7110 1120
rect 7046 1060 7050 1116
rect 7050 1060 7106 1116
rect 7106 1060 7110 1116
rect 7046 1056 7110 1060
rect 7126 1116 7190 1120
rect 7126 1060 7130 1116
rect 7130 1060 7186 1116
rect 7186 1060 7190 1116
rect 7126 1056 7190 1060
rect 12820 1116 12884 1120
rect 12820 1060 12824 1116
rect 12824 1060 12880 1116
rect 12880 1060 12884 1116
rect 12820 1056 12884 1060
rect 12900 1116 12964 1120
rect 12900 1060 12904 1116
rect 12904 1060 12960 1116
rect 12960 1060 12964 1116
rect 12900 1056 12964 1060
rect 12980 1116 13044 1120
rect 12980 1060 12984 1116
rect 12984 1060 13040 1116
rect 13040 1060 13044 1116
rect 12980 1056 13044 1060
rect 13060 1116 13124 1120
rect 13060 1060 13064 1116
rect 13064 1060 13120 1116
rect 13120 1060 13124 1116
rect 13060 1056 13124 1060
rect 18754 1116 18818 1120
rect 18754 1060 18758 1116
rect 18758 1060 18814 1116
rect 18814 1060 18818 1116
rect 18754 1056 18818 1060
rect 18834 1116 18898 1120
rect 18834 1060 18838 1116
rect 18838 1060 18894 1116
rect 18894 1060 18898 1116
rect 18834 1056 18898 1060
rect 18914 1116 18978 1120
rect 18914 1060 18918 1116
rect 18918 1060 18974 1116
rect 18974 1060 18978 1116
rect 18914 1056 18978 1060
rect 18994 1116 19058 1120
rect 18994 1060 18998 1116
rect 18998 1060 19054 1116
rect 19054 1060 19058 1116
rect 18994 1056 19058 1060
rect 24688 1116 24752 1120
rect 24688 1060 24692 1116
rect 24692 1060 24748 1116
rect 24748 1060 24752 1116
rect 24688 1056 24752 1060
rect 24768 1116 24832 1120
rect 24768 1060 24772 1116
rect 24772 1060 24828 1116
rect 24828 1060 24832 1116
rect 24768 1056 24832 1060
rect 24848 1116 24912 1120
rect 24848 1060 24852 1116
rect 24852 1060 24908 1116
rect 24908 1060 24912 1116
rect 24848 1056 24912 1060
rect 24928 1116 24992 1120
rect 24928 1060 24932 1116
rect 24932 1060 24988 1116
rect 24988 1060 24992 1116
rect 24928 1056 24992 1060
rect 15148 852 15212 916
<< metal4 >>
rect 3911 6016 4231 6576
rect 3911 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4231 6016
rect 3911 4928 4231 5952
rect 3911 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4231 4928
rect 3911 3840 4231 4864
rect 3911 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4231 3840
rect 3911 2752 4231 3776
rect 3911 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4231 2752
rect 3911 1664 4231 2688
rect 3911 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4231 1664
rect 3911 1040 4231 1600
rect 6878 6560 7198 6576
rect 6878 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7198 6560
rect 6878 5472 7198 6496
rect 6878 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7198 5472
rect 6878 4384 7198 5408
rect 6878 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7198 4384
rect 6878 3296 7198 4320
rect 6878 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7198 3296
rect 6878 2208 7198 3232
rect 6878 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7198 2208
rect 6878 1120 7198 2144
rect 6878 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7198 1120
rect 6878 1040 7198 1056
rect 9845 6016 10165 6576
rect 9845 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10165 6016
rect 9845 4928 10165 5952
rect 9845 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10165 4928
rect 9845 3840 10165 4864
rect 9845 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10165 3840
rect 9845 2752 10165 3776
rect 9845 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10165 2752
rect 9845 1664 10165 2688
rect 9845 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10165 1664
rect 9845 1040 10165 1600
rect 12812 6560 13132 6576
rect 12812 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13132 6560
rect 12812 5472 13132 6496
rect 12812 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13132 5472
rect 12812 4384 13132 5408
rect 12812 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13132 4384
rect 12812 3296 13132 4320
rect 15779 6016 16099 6576
rect 15779 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16099 6016
rect 15779 4928 16099 5952
rect 15779 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16099 4928
rect 15147 4180 15213 4181
rect 15147 4116 15148 4180
rect 15212 4116 15213 4180
rect 15147 4115 15213 4116
rect 12812 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13132 3296
rect 12812 2208 13132 3232
rect 12812 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13132 2208
rect 12812 1120 13132 2144
rect 12812 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13132 1120
rect 12812 1040 13132 1056
rect 15150 917 15210 4115
rect 15779 3840 16099 4864
rect 15779 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16099 3840
rect 15779 2752 16099 3776
rect 15779 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16099 2752
rect 15779 1664 16099 2688
rect 15779 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16099 1664
rect 15779 1040 16099 1600
rect 18746 6560 19066 6576
rect 18746 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19066 6560
rect 18746 5472 19066 6496
rect 20667 6356 20733 6357
rect 20667 6292 20668 6356
rect 20732 6292 20733 6356
rect 20667 6291 20733 6292
rect 18746 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19066 5472
rect 18746 4384 19066 5408
rect 18746 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19066 4384
rect 18746 3296 19066 4320
rect 18746 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19066 3296
rect 18746 2208 19066 3232
rect 20670 2277 20730 6291
rect 21713 6016 22033 6576
rect 21713 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22033 6016
rect 21713 4928 22033 5952
rect 24680 6560 25000 6576
rect 24680 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 25000 6560
rect 24680 5472 25000 6496
rect 24680 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 25000 5472
rect 22139 5132 22205 5133
rect 22139 5068 22140 5132
rect 22204 5068 22205 5132
rect 22139 5067 22205 5068
rect 21713 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22033 4928
rect 21713 3840 22033 4864
rect 21713 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22033 3840
rect 21713 2752 22033 3776
rect 21713 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22033 2752
rect 20667 2276 20733 2277
rect 20667 2212 20668 2276
rect 20732 2212 20733 2276
rect 20667 2211 20733 2212
rect 18746 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19066 2208
rect 18746 1120 19066 2144
rect 18746 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19066 1120
rect 18746 1040 19066 1056
rect 21713 1664 22033 2688
rect 22142 2277 22202 5067
rect 22323 4724 22389 4725
rect 22323 4660 22324 4724
rect 22388 4660 22389 4724
rect 22323 4659 22389 4660
rect 22326 2413 22386 4659
rect 24680 4384 25000 5408
rect 24680 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 25000 4384
rect 24680 3296 25000 4320
rect 24680 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 25000 3296
rect 22323 2412 22389 2413
rect 22323 2348 22324 2412
rect 22388 2348 22389 2412
rect 22323 2347 22389 2348
rect 22139 2276 22205 2277
rect 22139 2212 22140 2276
rect 22204 2212 22205 2276
rect 22139 2211 22205 2212
rect 21713 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22033 1664
rect 21713 1040 22033 1600
rect 24680 2208 25000 3232
rect 24680 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 25000 2208
rect 24680 1120 25000 2144
rect 24680 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 25000 1120
rect 24680 1040 25000 1056
rect 15147 916 15213 917
rect 15147 852 15148 916
rect 15212 852 15213 916
rect 15147 851 15213 852
use sky130_fd_sc_hd__clkbuf_1  _00_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _01_
timestamp 1688980957
transform 1 0 1472 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _02_
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _03_
timestamp 1688980957
transform 1 0 7176 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _04_
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _05_
timestamp 1688980957
transform 1 0 12420 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp 1688980957
transform 1 0 9292 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1688980957
transform 1 0 13064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1688980957
transform 1 0 13248 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1688980957
transform 1 0 15456 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _11_
timestamp 1688980957
transform 1 0 15088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1688980957
transform 1 0 5428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1688980957
transform 1 0 4324 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1688980957
transform 1 0 4048 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _17_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1688980957
transform 1 0 9476 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1688980957
transform 1 0 15364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1688980957
transform 1 0 16284 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1688980957
transform 1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1688980957
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1688980957
transform 1 0 17112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1688980957
transform 1 0 17664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1688980957
transform 1 0 18216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1688980957
transform 1 0 18768 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1688980957
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _36_
timestamp 1688980957
transform 1 0 20516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _37_
timestamp 1688980957
transform 1 0 14628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1688980957
transform 1 0 12420 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1688980957
transform 1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1688980957
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1688980957
transform 1 0 12144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1688980957
transform 1 0 13340 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1688980957
transform 1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1688980957
transform 1 0 17204 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1688980957
transform 1 0 18124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1688980957
transform 1 0 19780 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1688980957
transform 1 0 20792 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1688980957
transform 1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1688980957
transform 1 0 24104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8372 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 13064 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform -1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_126
timestamp 1688980957
transform 1 0 12696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_136 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13616 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_151
timestamp 1688980957
transform 1 0 14996 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_10
timestamp 1688980957
transform 1 0 2024 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_138
timestamp 1688980957
transform 1 0 13800 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_231
timestamp 1688980957
transform 1 0 22356 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_241
timestamp 1688980957
transform 1 0 23276 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_254
timestamp 1688980957
transform 1 0 24472 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_42
timestamp 1688980957
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_89
timestamp 1688980957
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_96
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_102
timestamp 1688980957
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_106
timestamp 1688980957
transform 1 0 10856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_110
timestamp 1688980957
transform 1 0 11224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_128
timestamp 1688980957
transform 1 0 12880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_149
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_158
timestamp 1688980957
transform 1 0 15640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_215
timestamp 1688980957
transform 1 0 20884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_227
timestamp 1688980957
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_253
timestamp 1688980957
transform 1 0 24380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_60
timestamp 1688980957
transform 1 0 6624 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_68
timestamp 1688980957
transform 1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_73
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_86
timestamp 1688980957
transform 1 0 9016 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_94
timestamp 1688980957
transform 1 0 9752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_98
timestamp 1688980957
transform 1 0 10120 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_106
timestamp 1688980957
transform 1 0 10856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_117
timestamp 1688980957
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_121
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_126
timestamp 1688980957
transform 1 0 12696 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_132
timestamp 1688980957
transform 1 0 13248 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_145
timestamp 1688980957
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_152
timestamp 1688980957
transform 1 0 15088 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_160
timestamp 1688980957
transform 1 0 15824 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_164
timestamp 1688980957
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_173
timestamp 1688980957
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_177
timestamp 1688980957
transform 1 0 17388 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_185
timestamp 1688980957
transform 1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_191
timestamp 1688980957
transform 1 0 18676 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_203
timestamp 1688980957
transform 1 0 19780 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_208
timestamp 1688980957
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_220
timestamp 1688980957
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_253
timestamp 1688980957
transform 1 0 24380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_57
timestamp 1688980957
transform 1 0 6348 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_71
timestamp 1688980957
transform 1 0 7636 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_79
timestamp 1688980957
transform 1 0 8372 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_96
timestamp 1688980957
transform 1 0 9936 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_104
timestamp 1688980957
transform 1 0 10672 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_115
timestamp 1688980957
transform 1 0 11684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_119
timestamp 1688980957
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_124
timestamp 1688980957
transform 1 0 12512 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_135
timestamp 1688980957
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_150
timestamp 1688980957
transform 1 0 14904 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_158
timestamp 1688980957
transform 1 0 15640 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_162
timestamp 1688980957
transform 1 0 16008 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_170
timestamp 1688980957
transform 1 0 16744 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_175
timestamp 1688980957
transform 1 0 17204 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_183
timestamp 1688980957
transform 1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_206
timestamp 1688980957
transform 1 0 20056 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_218
timestamp 1688980957
transform 1 0 21160 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_230
timestamp 1688980957
transform 1 0 22264 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_242
timestamp 1688980957
transform 1 0 23368 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_17
timestamp 1688980957
transform 1 0 2668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_25
timestamp 1688980957
transform 1 0 3404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_35
timestamp 1688980957
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_42
timestamp 1688980957
transform 1 0 4968 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_48
timestamp 1688980957
transform 1 0 5520 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_60
timestamp 1688980957
transform 1 0 6624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_71
timestamp 1688980957
transform 1 0 7636 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_85
timestamp 1688980957
transform 1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_97
timestamp 1688980957
transform 1 0 10028 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_126
timestamp 1688980957
transform 1 0 12696 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_136
timestamp 1688980957
transform 1 0 13616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_162
timestamp 1688980957
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_178
timestamp 1688980957
transform 1 0 17480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_188
timestamp 1688980957
transform 1 0 18400 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_206
timestamp 1688980957
transform 1 0 20056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_228
timestamp 1688980957
transform 1 0 22080 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_240
timestamp 1688980957
transform 1 0 23184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_253
timestamp 1688980957
transform 1 0 24380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 21436 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 24196 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 23736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 22448 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 23276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 23184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 22080 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 22356 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 22632 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 22908 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 22080 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 23460 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 23736 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 24012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 23000 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 2392 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 2668 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 2576 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 3220 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 3496 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 3772 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 4324 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 4600 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 4876 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 1748 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 2116 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 1748 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 2024 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 2944 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 2300 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 4600 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 8096 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 8648 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 6072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 5704 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 5980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 6440 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 6992 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 7268 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 7544 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 7820 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20700 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._00_
timestamp 1688980957
transform 1 0 8372 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._01_
timestamp 1688980957
transform 1 0 1472 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._02_
timestamp 1688980957
transform 1 0 6900 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._03_
timestamp 1688980957
transform 1 0 6624 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._04_
timestamp 1688980957
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._05_
timestamp 1688980957
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._06_
timestamp 1688980957
transform 1 0 10028 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._07_
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._08_
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._09_
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._10_
timestamp 1688980957
transform 1 0 13892 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._11_
timestamp 1688980957
transform 1 0 14168 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._12_
timestamp 1688980957
transform 1 0 5428 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._13_
timestamp 1688980957
transform 1 0 5152 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._14_
timestamp 1688980957
transform 1 0 3404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._15_
timestamp 1688980957
transform 1 0 3128 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._16_
timestamp 1688980957
transform 1 0 2852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._17_
timestamp 1688980957
transform 1 0 4048 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._18_
timestamp 1688980957
transform 1 0 6716 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._19_
timestamp 1688980957
transform 1 0 8924 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._20_
timestamp 1688980957
transform 1 0 9752 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_RAM_IO_switch_matrix._21_
timestamp 1688980957
transform 1 0 9016 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._22_
timestamp 1688980957
transform 1 0 17940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_RAM_IO_switch_matrix._23_
timestamp 1688980957
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_RAM_IO_switch_matrix._24_
timestamp 1688980957
transform 1 0 5704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._25_
timestamp 1688980957
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._26_
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._27_
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._28_
timestamp 1688980957
transform 1 0 9200 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._29_
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._30_
timestamp 1688980957
transform 1 0 13524 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._31_
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._32_
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._33_
timestamp 1688980957
transform 1 0 17388 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._34_
timestamp 1688980957
transform 1 0 17664 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._35_
timestamp 1688980957
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output58 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output59 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output60
timestamp 1688980957
transform 1 0 15180 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output62
timestamp 1688980957
transform 1 0 17572 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output63
timestamp 1688980957
transform 1 0 19228 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1688980957
transform 1 0 20148 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1688980957
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output66
timestamp 1688980957
transform 1 0 22356 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output67
timestamp 1688980957
transform 1 0 23736 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output68
timestamp 1688980957
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output69
timestamp 1688980957
transform 1 0 3772 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output70
timestamp 1688980957
transform 1 0 4416 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output71
timestamp 1688980957
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1688980957
transform 1 0 6808 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 1688980957
transform 1 0 8004 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output74
timestamp 1688980957
transform 1 0 9200 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 10396 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1688980957
transform 1 0 11776 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1688980957
transform 1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1688980957
transform 1 0 9568 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 10304 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1688980957
transform 1 0 9936 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 10856 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1688980957
transform 1 0 13248 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1688980957
transform 1 0 14628 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1688980957
transform 1 0 14444 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1688980957
transform 1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 10672 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1688980957
transform 1 0 10304 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 11868 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 12144 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 12696 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform 1 0 11776 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 15732 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 19780 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 20332 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output101
timestamp 1688980957
transform 1 0 19596 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 20148 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1688980957
transform 1 0 21068 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 20884 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 16836 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 19044 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 17940 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 18492 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform -1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 24840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 24840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 24840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 24840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 24840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0._0_
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1._0_
timestamp 1688980957
transform 1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2._0_
timestamp 1688980957
transform 1 0 11960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3._0_
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4._0_
timestamp 1688980957
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5._0_
timestamp 1688980957
transform 1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6._0_
timestamp 1688980957
transform 1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7._0_
timestamp 1688980957
transform 1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8._0_
timestamp 1688980957
transform 1 0 12420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9._0_
timestamp 1688980957
transform 1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10._0_
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11._0_
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12._0_
timestamp 1688980957
transform 1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13._0_
timestamp 1688980957
transform 1 0 18400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14._0_
timestamp 1688980957
transform 1 0 23368 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15._0_
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16._0_
timestamp 1688980957
transform 1 0 23184 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17._0_
timestamp 1688980957
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18._0_
timestamp 1688980957
transform 1 0 24104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19._0_
timestamp 1688980957
transform 1 0 23736 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0._0_
timestamp 1688980957
transform 1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1._0_
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_2._0_
timestamp 1688980957
transform 1 0 11776 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3._0_
timestamp 1688980957
transform 1 0 6072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4._0_
timestamp 1688980957
transform 1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5._0_
timestamp 1688980957
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6._0_
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7._0_
timestamp 1688980957
transform 1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8._0_
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9._0_
timestamp 1688980957
transform 1 0 13248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10._0_
timestamp 1688980957
transform 1 0 14628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11._0_
timestamp 1688980957
transform 1 0 15732 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12._0_
timestamp 1688980957
transform 1 0 16928 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13._0_
timestamp 1688980957
transform 1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14._0_
timestamp 1688980957
transform 1 0 23644 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15._0_
timestamp 1688980957
transform 1 0 23920 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16._0_
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17._0_
timestamp 1688980957
transform 1 0 22724 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18._0_
timestamp 1688980957
transform 1 0 23920 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19._0_
timestamp 1688980957
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 3680 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 8832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 13984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 19136 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 24288 0 -1 6528
box -38 -48 130 592
<< labels >>
flabel metal2 s 20350 0 20406 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 23110 0 23166 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 23386 0 23442 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 23662 0 23718 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 23938 0 23994 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 24214 0 24270 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 24490 0 24546 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 24766 0 24822 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 25042 0 25098 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 25318 0 25374 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 25594 0 25650 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 20626 0 20682 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 20902 0 20958 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 21178 0 21234 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 21454 0 21510 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 21730 0 21786 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 22006 0 22062 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 22282 0 22338 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 22558 0 22614 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 22834 0 22890 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 2134 7840 2190 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 14094 7840 14150 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 15290 7840 15346 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 16486 7840 16542 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 17682 7840 17738 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 18878 7840 18934 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 20074 7840 20130 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 21270 7840 21326 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 22466 7840 22522 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 23662 7840 23718 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 24858 7840 24914 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 3330 7840 3386 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 4526 7840 4582 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 5722 7840 5778 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 6918 7840 6974 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 8114 7840 8170 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 9310 7840 9366 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 10506 7840 10562 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 11702 7840 11758 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 12898 7840 12954 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 202 0 258 160 0 FreeSans 224 90 0 0 N1END[0]
port 40 nsew signal input
flabel metal2 s 478 0 534 160 0 FreeSans 224 90 0 0 N1END[1]
port 41 nsew signal input
flabel metal2 s 754 0 810 160 0 FreeSans 224 90 0 0 N1END[2]
port 42 nsew signal input
flabel metal2 s 1030 0 1086 160 0 FreeSans 224 90 0 0 N1END[3]
port 43 nsew signal input
flabel metal2 s 3514 0 3570 160 0 FreeSans 224 90 0 0 N2END[0]
port 44 nsew signal input
flabel metal2 s 3790 0 3846 160 0 FreeSans 224 90 0 0 N2END[1]
port 45 nsew signal input
flabel metal2 s 4066 0 4122 160 0 FreeSans 224 90 0 0 N2END[2]
port 46 nsew signal input
flabel metal2 s 4342 0 4398 160 0 FreeSans 224 90 0 0 N2END[3]
port 47 nsew signal input
flabel metal2 s 4618 0 4674 160 0 FreeSans 224 90 0 0 N2END[4]
port 48 nsew signal input
flabel metal2 s 4894 0 4950 160 0 FreeSans 224 90 0 0 N2END[5]
port 49 nsew signal input
flabel metal2 s 5170 0 5226 160 0 FreeSans 224 90 0 0 N2END[6]
port 50 nsew signal input
flabel metal2 s 5446 0 5502 160 0 FreeSans 224 90 0 0 N2END[7]
port 51 nsew signal input
flabel metal2 s 1306 0 1362 160 0 FreeSans 224 90 0 0 N2MID[0]
port 52 nsew signal input
flabel metal2 s 1582 0 1638 160 0 FreeSans 224 90 0 0 N2MID[1]
port 53 nsew signal input
flabel metal2 s 1858 0 1914 160 0 FreeSans 224 90 0 0 N2MID[2]
port 54 nsew signal input
flabel metal2 s 2134 0 2190 160 0 FreeSans 224 90 0 0 N2MID[3]
port 55 nsew signal input
flabel metal2 s 2410 0 2466 160 0 FreeSans 224 90 0 0 N2MID[4]
port 56 nsew signal input
flabel metal2 s 2686 0 2742 160 0 FreeSans 224 90 0 0 N2MID[5]
port 57 nsew signal input
flabel metal2 s 2962 0 3018 160 0 FreeSans 224 90 0 0 N2MID[6]
port 58 nsew signal input
flabel metal2 s 3238 0 3294 160 0 FreeSans 224 90 0 0 N2MID[7]
port 59 nsew signal input
flabel metal2 s 5722 0 5778 160 0 FreeSans 224 90 0 0 N4END[0]
port 60 nsew signal input
flabel metal2 s 8482 0 8538 160 0 FreeSans 224 90 0 0 N4END[10]
port 61 nsew signal input
flabel metal2 s 8758 0 8814 160 0 FreeSans 224 90 0 0 N4END[11]
port 62 nsew signal input
flabel metal2 s 9034 0 9090 160 0 FreeSans 224 90 0 0 N4END[12]
port 63 nsew signal input
flabel metal2 s 9310 0 9366 160 0 FreeSans 224 90 0 0 N4END[13]
port 64 nsew signal input
flabel metal2 s 9586 0 9642 160 0 FreeSans 224 90 0 0 N4END[14]
port 65 nsew signal input
flabel metal2 s 9862 0 9918 160 0 FreeSans 224 90 0 0 N4END[15]
port 66 nsew signal input
flabel metal2 s 5998 0 6054 160 0 FreeSans 224 90 0 0 N4END[1]
port 67 nsew signal input
flabel metal2 s 6274 0 6330 160 0 FreeSans 224 90 0 0 N4END[2]
port 68 nsew signal input
flabel metal2 s 6550 0 6606 160 0 FreeSans 224 90 0 0 N4END[3]
port 69 nsew signal input
flabel metal2 s 6826 0 6882 160 0 FreeSans 224 90 0 0 N4END[4]
port 70 nsew signal input
flabel metal2 s 7102 0 7158 160 0 FreeSans 224 90 0 0 N4END[5]
port 71 nsew signal input
flabel metal2 s 7378 0 7434 160 0 FreeSans 224 90 0 0 N4END[6]
port 72 nsew signal input
flabel metal2 s 7654 0 7710 160 0 FreeSans 224 90 0 0 N4END[7]
port 73 nsew signal input
flabel metal2 s 7930 0 7986 160 0 FreeSans 224 90 0 0 N4END[8]
port 74 nsew signal input
flabel metal2 s 8206 0 8262 160 0 FreeSans 224 90 0 0 N4END[9]
port 75 nsew signal input
flabel metal2 s 10138 0 10194 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 76 nsew signal tristate
flabel metal2 s 10414 0 10470 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 77 nsew signal tristate
flabel metal2 s 10690 0 10746 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 78 nsew signal tristate
flabel metal2 s 10966 0 11022 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 79 nsew signal tristate
flabel metal2 s 13450 0 13506 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 80 nsew signal tristate
flabel metal2 s 13726 0 13782 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 81 nsew signal tristate
flabel metal2 s 14002 0 14058 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 82 nsew signal tristate
flabel metal2 s 14278 0 14334 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 83 nsew signal tristate
flabel metal2 s 14554 0 14610 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 84 nsew signal tristate
flabel metal2 s 14830 0 14886 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 85 nsew signal tristate
flabel metal2 s 15106 0 15162 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 86 nsew signal tristate
flabel metal2 s 15382 0 15438 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 87 nsew signal tristate
flabel metal2 s 11242 0 11298 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 88 nsew signal tristate
flabel metal2 s 11518 0 11574 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 89 nsew signal tristate
flabel metal2 s 11794 0 11850 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 90 nsew signal tristate
flabel metal2 s 12070 0 12126 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 91 nsew signal tristate
flabel metal2 s 12346 0 12402 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 92 nsew signal tristate
flabel metal2 s 12622 0 12678 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 93 nsew signal tristate
flabel metal2 s 12898 0 12954 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 94 nsew signal tristate
flabel metal2 s 13174 0 13230 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 95 nsew signal tristate
flabel metal2 s 15658 0 15714 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 96 nsew signal tristate
flabel metal2 s 18418 0 18474 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 97 nsew signal tristate
flabel metal2 s 18694 0 18750 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 98 nsew signal tristate
flabel metal2 s 18970 0 19026 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 99 nsew signal tristate
flabel metal2 s 19246 0 19302 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 100 nsew signal tristate
flabel metal2 s 19522 0 19578 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 101 nsew signal tristate
flabel metal2 s 19798 0 19854 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 102 nsew signal tristate
flabel metal2 s 15934 0 15990 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 103 nsew signal tristate
flabel metal2 s 16210 0 16266 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 104 nsew signal tristate
flabel metal2 s 16486 0 16542 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 105 nsew signal tristate
flabel metal2 s 16762 0 16818 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 106 nsew signal tristate
flabel metal2 s 17038 0 17094 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 107 nsew signal tristate
flabel metal2 s 17314 0 17370 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 108 nsew signal tristate
flabel metal2 s 17590 0 17646 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 109 nsew signal tristate
flabel metal2 s 17866 0 17922 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 110 nsew signal tristate
flabel metal2 s 18142 0 18198 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 111 nsew signal tristate
flabel metal2 s 20074 0 20130 160 0 FreeSans 224 90 0 0 UserCLK
port 112 nsew signal input
flabel metal2 s 938 7840 994 8000 0 FreeSans 224 90 0 0 UserCLKo
port 113 nsew signal tristate
flabel metal4 s 6878 1040 7198 6576 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 12812 1040 13132 6576 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 18746 1040 19066 6576 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 24680 1040 25000 6576 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 3911 1040 4231 6576 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 9845 1040 10165 6576 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 15779 1040 16099 6576 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 21713 1040 22033 6576 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
rlabel via1 13052 6528 13052 6528 0 VGND
rlabel metal1 12972 5984 12972 5984 0 VPWR
rlabel metal2 20378 976 20378 976 0 FrameStrobe[0]
rlabel metal2 23138 211 23138 211 0 FrameStrobe[10]
rlabel metal2 23414 1044 23414 1044 0 FrameStrobe[11]
rlabel metal2 23690 1299 23690 1299 0 FrameStrobe[12]
rlabel metal2 23966 415 23966 415 0 FrameStrobe[13]
rlabel metal2 24242 279 24242 279 0 FrameStrobe[14]
rlabel metal1 24288 2958 24288 2958 0 FrameStrobe[15]
rlabel metal1 24196 2890 24196 2890 0 FrameStrobe[16]
rlabel metal1 24288 3094 24288 3094 0 FrameStrobe[17]
rlabel metal2 25346 1282 25346 1282 0 FrameStrobe[18]
rlabel metal2 25622 738 25622 738 0 FrameStrobe[19]
rlabel metal2 20654 670 20654 670 0 FrameStrobe[1]
rlabel metal2 21029 68 21029 68 0 FrameStrobe[2]
rlabel metal2 21206 211 21206 211 0 FrameStrobe[3]
rlabel metal2 21482 364 21482 364 0 FrameStrobe[4]
rlabel metal2 21857 68 21857 68 0 FrameStrobe[5]
rlabel metal2 22034 296 22034 296 0 FrameStrobe[6]
rlabel metal2 22409 68 22409 68 0 FrameStrobe[7]
rlabel metal2 22685 68 22685 68 0 FrameStrobe[8]
rlabel metal2 22862 1010 22862 1010 0 FrameStrobe[9]
rlabel metal1 2346 6426 2346 6426 0 FrameStrobe_O[0]
rlabel metal2 14221 7956 14221 7956 0 FrameStrobe_O[10]
rlabel metal2 15371 7956 15371 7956 0 FrameStrobe_O[11]
rlabel metal2 16705 7956 16705 7956 0 FrameStrobe_O[12]
rlabel metal2 17763 7956 17763 7956 0 FrameStrobe_O[13]
rlabel metal2 19189 7956 19189 7956 0 FrameStrobe_O[14]
rlabel metal2 20378 7191 20378 7191 0 FrameStrobe_O[15]
rlabel metal2 21574 7191 21574 7191 0 FrameStrobe_O[16]
rlabel metal2 22547 7956 22547 7956 0 FrameStrobe_O[17]
rlabel metal2 23690 7184 23690 7184 0 FrameStrobe_O[18]
rlabel metal1 24334 5882 24334 5882 0 FrameStrobe_O[19]
rlabel metal2 3595 7956 3595 7956 0 FrameStrobe_O[1]
rlabel metal2 4607 7956 4607 7956 0 FrameStrobe_O[2]
rlabel metal2 5941 7956 5941 7956 0 FrameStrobe_O[3]
rlabel metal2 7137 7956 7137 7956 0 FrameStrobe_O[4]
rlabel metal2 8287 7956 8287 7956 0 FrameStrobe_O[5]
rlabel metal2 9391 7956 9391 7956 0 FrameStrobe_O[6]
rlabel metal2 10587 7956 10587 7956 0 FrameStrobe_O[7]
rlabel metal2 12006 7191 12006 7191 0 FrameStrobe_O[8]
rlabel metal2 13202 7191 13202 7191 0 FrameStrobe_O[9]
rlabel metal2 8234 1530 8234 1530 0 Inst_N_term_RAM_IO_switch_matrix.S1BEG0
rlabel metal1 1610 1326 1610 1326 0 Inst_N_term_RAM_IO_switch_matrix.S1BEG1
rlabel metal1 7682 1292 7682 1292 0 Inst_N_term_RAM_IO_switch_matrix.S1BEG2
rlabel metal1 7314 1326 7314 1326 0 Inst_N_term_RAM_IO_switch_matrix.S1BEG3
rlabel metal1 11730 2448 11730 2448 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG0
rlabel metal2 12374 2108 12374 2108 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG1
rlabel viali 9522 1324 9522 1324 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG2
rlabel metal1 12190 2414 12190 2414 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG3
rlabel metal1 13294 2448 13294 2448 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG4
rlabel metal1 13478 1972 13478 1972 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG5
rlabel metal1 15824 1938 15824 1938 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG6
rlabel metal2 14214 2278 14214 2278 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG7
rlabel metal1 5612 1326 5612 1326 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb0
rlabel metal1 5290 1326 5290 1326 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb1
rlabel metal1 4462 1326 4462 1326 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb2
rlabel metal1 4002 1292 4002 1292 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb3
rlabel metal1 3082 1530 3082 1530 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb4
rlabel metal1 4922 1292 4922 1292 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb5
rlabel metal1 6578 1360 6578 1360 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb6
rlabel metal1 9614 1938 9614 1938 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb7
rlabel metal1 10120 1734 10120 1734 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG0
rlabel metal2 13662 1190 13662 1190 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG1
rlabel metal1 18584 1326 18584 1326 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG10
rlabel metal2 18078 799 18078 799 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG11
rlabel metal2 18354 1581 18354 1581 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG12
rlabel metal1 19458 2380 19458 2380 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG13
rlabel metal1 20562 2448 20562 2448 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG14
rlabel metal1 20976 1190 20976 1190 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG15
rlabel metal2 9246 2210 9246 2210 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG2
rlabel metal2 16974 1530 16974 1530 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG3
rlabel metal2 15410 1819 15410 1819 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG4
rlabel metal1 16422 1530 16422 1530 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG5
rlabel metal1 17342 2448 17342 2448 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG6
rlabel metal1 17526 2074 17526 2074 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG7
rlabel metal1 17802 2074 17802 2074 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG8
rlabel metal2 21482 1666 21482 1666 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG9
rlabel metal2 230 1214 230 1214 0 N1END[0]
rlabel metal2 506 1282 506 1282 0 N1END[1]
rlabel metal2 782 1044 782 1044 0 N1END[2]
rlabel metal2 1058 942 1058 942 0 N1END[3]
rlabel metal2 3542 398 3542 398 0 N2END[0]
rlabel metal2 3719 68 3719 68 0 N2END[1]
rlabel metal2 3995 68 3995 68 0 N2END[2]
rlabel metal2 4370 1010 4370 1010 0 N2END[3]
rlabel metal2 4646 1248 4646 1248 0 N2END[4]
rlabel metal2 4922 1010 4922 1010 0 N2END[5]
rlabel metal2 5099 68 5099 68 0 N2END[6]
rlabel metal2 5474 1044 5474 1044 0 N2END[7]
rlabel metal2 1334 1248 1334 1248 0 N2MID[0]
rlabel metal2 1709 68 1709 68 0 N2MID[1]
rlabel metal2 1886 1180 1886 1180 0 N2MID[2]
rlabel metal2 2162 1010 2162 1010 0 N2MID[3]
rlabel metal2 2339 68 2339 68 0 N2MID[4]
rlabel metal2 2714 670 2714 670 0 N2MID[5]
rlabel metal2 3089 68 3089 68 0 N2MID[6]
rlabel metal1 2714 1360 2714 1360 0 N2MID[7]
rlabel metal2 5750 347 5750 347 0 N4END[0]
rlabel metal2 8510 1010 8510 1010 0 N4END[10]
rlabel metal2 8786 415 8786 415 0 N4END[11]
rlabel metal2 9062 1010 9062 1010 0 N4END[12]
rlabel metal2 9338 1248 9338 1248 0 N4END[13]
rlabel metal2 9614 755 9614 755 0 N4END[14]
rlabel metal2 9890 347 9890 347 0 N4END[15]
rlabel metal2 6026 279 6026 279 0 N4END[1]
rlabel metal2 6302 976 6302 976 0 N4END[2]
rlabel metal2 6578 1010 6578 1010 0 N4END[3]
rlabel metal2 6854 534 6854 534 0 N4END[4]
rlabel metal2 7130 534 7130 534 0 N4END[5]
rlabel metal2 7406 1010 7406 1010 0 N4END[6]
rlabel metal2 7682 1010 7682 1010 0 N4END[7]
rlabel metal2 7958 1010 7958 1010 0 N4END[8]
rlabel metal2 8234 534 8234 534 0 N4END[9]
rlabel metal2 10113 68 10113 68 0 S1BEG[0]
rlabel metal2 10442 908 10442 908 0 S1BEG[1]
rlabel metal2 10718 670 10718 670 0 S1BEG[2]
rlabel metal2 10994 908 10994 908 0 S1BEG[3]
rlabel metal2 13478 636 13478 636 0 S2BEG[0]
rlabel metal2 13754 806 13754 806 0 S2BEG[1]
rlabel metal2 14030 636 14030 636 0 S2BEG[2]
rlabel metal2 14405 68 14405 68 0 S2BEG[3]
rlabel metal2 14681 68 14681 68 0 S2BEG[4]
rlabel metal2 14858 687 14858 687 0 S2BEG[5]
rlabel metal2 15134 755 15134 755 0 S2BEG[6]
rlabel metal2 15410 619 15410 619 0 S2BEG[7]
rlabel metal2 11171 68 11171 68 0 S2BEGb[0]
rlabel metal2 11546 636 11546 636 0 S2BEGb[1]
rlabel metal2 11822 908 11822 908 0 S2BEGb[2]
rlabel metal2 11999 68 11999 68 0 S2BEGb[3]
rlabel metal2 12374 636 12374 636 0 S2BEGb[4]
rlabel metal2 12650 908 12650 908 0 S2BEGb[5]
rlabel metal2 12926 415 12926 415 0 S2BEGb[6]
rlabel metal2 13202 636 13202 636 0 S2BEGb[7]
rlabel metal2 15686 908 15686 908 0 S4BEG[0]
rlabel metal2 18446 823 18446 823 0 S4BEG[10]
rlabel metal2 18722 347 18722 347 0 S4BEG[11]
rlabel metal2 18998 483 18998 483 0 S4BEG[12]
rlabel metal2 19274 551 19274 551 0 S4BEG[13]
rlabel metal1 21160 2074 21160 2074 0 S4BEG[14]
rlabel metal2 19826 806 19826 806 0 S4BEG[15]
rlabel metal2 15962 755 15962 755 0 S4BEG[1]
rlabel metal2 16291 68 16291 68 0 S4BEG[2]
rlabel metal2 16514 636 16514 636 0 S4BEG[3]
rlabel metal2 16790 908 16790 908 0 S4BEG[4]
rlabel metal2 17066 806 17066 806 0 S4BEG[5]
rlabel metal2 17342 738 17342 738 0 S4BEG[6]
rlabel metal2 17618 942 17618 942 0 S4BEG[7]
rlabel metal2 17894 959 17894 959 0 S4BEG[8]
rlabel metal2 18170 483 18170 483 0 S4BEG[9]
rlabel metal2 20155 68 20155 68 0 UserCLK
rlabel metal2 1203 7956 1203 7956 0 UserCLKo
rlabel metal1 20838 5202 20838 5202 0 net1
rlabel metal2 23230 2992 23230 2992 0 net10
rlabel metal1 20102 1258 20102 1258 0 net100
rlabel metal1 19458 2006 19458 2006 0 net101
rlabel metal1 20286 2040 20286 2040 0 net102
rlabel metal1 20746 1938 20746 1938 0 net103
rlabel metal1 20516 1326 20516 1326 0 net104
rlabel metal1 16698 1326 16698 1326 0 net105
rlabel metal2 14950 1054 14950 1054 0 net106
rlabel metal1 17388 1326 17388 1326 0 net107
rlabel metal1 16974 1904 16974 1904 0 net108
rlabel metal1 17940 1258 17940 1258 0 net109
rlabel metal1 22954 2312 22954 2312 0 net11
rlabel metal1 19366 1224 19366 1224 0 net110
rlabel metal1 18676 1938 18676 1938 0 net111
rlabel metal1 17940 2006 17940 2006 0 net112
rlabel metal1 18630 2040 18630 2040 0 net113
rlabel via2 2254 6307 2254 6307 0 net114
rlabel metal2 14950 1836 14950 1836 0 net12
rlabel metal2 13570 2482 13570 2482 0 net13
rlabel metal1 15364 510 15364 510 0 net14
rlabel metal2 12604 2244 12604 2244 0 net15
rlabel metal2 22310 2159 22310 2159 0 net16
rlabel metal1 15502 578 15502 578 0 net17
rlabel metal4 15180 2516 15180 2516 0 net18
rlabel metal1 16192 4998 16192 4998 0 net19
rlabel metal2 15042 3910 15042 3910 0 net2
rlabel metal1 13708 5202 13708 5202 0 net20
rlabel metal2 5750 2312 5750 2312 0 net21
rlabel metal1 2346 2312 2346 2312 0 net22
rlabel metal1 1702 1904 1702 1904 0 net23
rlabel metal1 2714 2040 2714 2040 0 net24
rlabel metal2 2622 2074 2622 2074 0 net25
rlabel metal1 6854 1938 6854 1938 0 net26
rlabel metal1 4186 1326 4186 1326 0 net27
rlabel metal2 3082 1564 3082 1564 0 net28
rlabel metal1 3358 1428 3358 1428 0 net29
rlabel metal1 18722 5066 18722 5066 0 net3
rlabel metal1 3772 1326 3772 1326 0 net30
rlabel metal1 5382 1904 5382 1904 0 net31
rlabel metal1 5658 1870 5658 1870 0 net32
rlabel metal2 1610 2788 1610 2788 0 net33
rlabel via2 1978 1717 1978 1717 0 net34
rlabel metal2 2438 2125 2438 2125 0 net35
rlabel metal2 2346 1683 2346 1683 0 net36
rlabel metal2 1978 765 1978 765 0 net37
rlabel metal1 2070 884 2070 884 0 net38
rlabel metal2 12558 2618 12558 2618 0 net39
rlabel metal2 17894 4046 17894 4046 0 net4
rlabel metal2 2346 1088 2346 1088 0 net40
rlabel metal2 21850 901 21850 901 0 net41
rlabel metal2 16146 884 16146 884 0 net42
rlabel metal1 13754 2006 13754 2006 0 net43
rlabel metal1 8602 1326 8602 1326 0 net44
rlabel metal2 9430 2108 9430 2108 0 net45
rlabel metal2 9522 2040 9522 2040 0 net46
rlabel metal1 8878 1190 8878 1190 0 net47
rlabel via2 19734 2397 19734 2397 0 net48
rlabel metal2 20286 2125 20286 2125 0 net49
rlabel metal1 18630 5168 18630 5168 0 net5
rlabel metal1 5750 1360 5750 1360 0 net50
rlabel metal1 6256 1326 6256 1326 0 net51
rlabel metal2 18170 2465 18170 2465 0 net52
rlabel metal1 21436 1326 21436 1326 0 net53
rlabel metal1 15134 1496 15134 1496 0 net54
rlabel metal1 14950 2584 14950 2584 0 net55
rlabel metal2 14582 2499 14582 2499 0 net56
rlabel metal1 20838 2040 20838 2040 0 net57
rlabel metal2 5658 6256 5658 6256 0 net58
rlabel metal1 14582 6358 14582 6358 0 net59
rlabel metal1 23460 1938 23460 1938 0 net6
rlabel metal1 15548 6358 15548 6358 0 net60
rlabel metal1 17020 6358 17020 6358 0 net61
rlabel metal1 17940 6358 17940 6358 0 net62
rlabel metal1 19596 6358 19596 6358 0 net63
rlabel metal1 20194 6324 20194 6324 0 net64
rlabel metal1 21620 6290 21620 6290 0 net65
rlabel metal1 22494 6392 22494 6392 0 net66
rlabel metal1 23690 6358 23690 6358 0 net67
rlabel metal1 24012 5338 24012 5338 0 net68
rlabel metal1 3910 6188 3910 6188 0 net69
rlabel metal1 23966 2822 23966 2822 0 net7
rlabel metal1 12466 6324 12466 6324 0 net70
rlabel metal1 5750 6392 5750 6392 0 net71
rlabel metal1 7176 6358 7176 6358 0 net72
rlabel metal1 8372 6358 8372 6358 0 net73
rlabel metal1 9568 6358 9568 6358 0 net74
rlabel metal1 10764 6358 10764 6358 0 net75
rlabel metal1 12006 6290 12006 6290 0 net76
rlabel metal1 13202 6290 13202 6290 0 net77
rlabel metal1 9614 1292 9614 1292 0 net78
rlabel via2 2990 1445 2990 1445 0 net79
rlabel metal1 23506 1258 23506 1258 0 net8
rlabel metal1 7498 680 7498 680 0 net80
rlabel metal1 8234 1462 8234 1462 0 net81
rlabel metal2 13294 1938 13294 1938 0 net82
rlabel metal1 13708 1258 13708 1258 0 net83
rlabel metal2 14674 1054 14674 1054 0 net84
rlabel metal1 14490 1904 14490 1904 0 net85
rlabel metal1 14858 1972 14858 1972 0 net86
rlabel metal1 14858 1258 14858 1258 0 net87
rlabel metal1 15686 1326 15686 1326 0 net88
rlabel metal1 15962 2448 15962 2448 0 net89
rlabel metal1 23184 2822 23184 2822 0 net9
rlabel metal2 10810 1088 10810 1088 0 net90
rlabel metal1 10258 1326 10258 1326 0 net91
rlabel metal1 4462 1190 4462 1190 0 net92
rlabel metal1 3910 1190 3910 1190 0 net93
rlabel metal2 4094 2142 4094 2142 0 net94
rlabel metal2 12834 1615 12834 1615 0 net95
rlabel metal1 11822 1360 11822 1360 0 net96
rlabel metal1 12558 1360 12558 1360 0 net97
rlabel metal1 15686 2006 15686 2006 0 net98
rlabel metal1 19596 1326 19596 1326 0 net99
rlabel metal2 20010 5508 20010 5508 0 strobe_inbuf_0.X
rlabel metal2 14582 5508 14582 5508 0 strobe_inbuf_1.X
rlabel metal2 14858 5508 14858 5508 0 strobe_inbuf_10.X
rlabel metal2 15962 5508 15962 5508 0 strobe_inbuf_11.X
rlabel metal2 17158 5508 17158 5508 0 strobe_inbuf_12.X
rlabel metal2 18446 5508 18446 5508 0 strobe_inbuf_13.X
rlabel metal1 23874 1904 23874 1904 0 strobe_inbuf_14.X
rlabel metal1 24104 1938 24104 1938 0 strobe_inbuf_15.X
rlabel metal2 21666 1734 21666 1734 0 strobe_inbuf_16.X
rlabel metal1 22954 1972 22954 1972 0 strobe_inbuf_17.X
rlabel metal2 24150 3332 24150 3332 0 strobe_inbuf_18.X
rlabel metal1 24242 4624 24242 4624 0 strobe_inbuf_19.X
rlabel metal2 12006 5508 12006 5508 0 strobe_inbuf_2.X
rlabel metal1 6348 5338 6348 5338 0 strobe_inbuf_3.X
rlabel metal2 7590 5508 7590 5508 0 strobe_inbuf_4.X
rlabel metal2 8786 5508 8786 5508 0 strobe_inbuf_5.X
rlabel metal2 9890 5508 9890 5508 0 strobe_inbuf_6.X
rlabel metal2 11086 5508 11086 5508 0 strobe_inbuf_7.X
rlabel metal2 12466 5508 12466 5508 0 strobe_inbuf_8.X
rlabel metal2 13478 5508 13478 5508 0 strobe_inbuf_9.X
rlabel metal1 20194 5882 20194 5882 0 strobe_outbuf_0.X
rlabel metal1 14536 5882 14536 5882 0 strobe_outbuf_1.X
rlabel metal1 14904 5542 14904 5542 0 strobe_outbuf_10.X
rlabel metal1 15732 5882 15732 5882 0 strobe_outbuf_11.X
rlabel metal1 17204 5882 17204 5882 0 strobe_outbuf_12.X
rlabel metal1 18308 5882 18308 5882 0 strobe_outbuf_13.X
rlabel metal2 24104 2924 24104 2924 0 strobe_outbuf_14.X
rlabel metal1 21022 6222 21022 6222 0 strobe_outbuf_15.X
rlabel metal1 21758 2074 21758 2074 0 strobe_outbuf_16.X
rlabel metal1 22954 2074 22954 2074 0 strobe_outbuf_17.X
rlabel metal1 23828 3706 23828 3706 0 strobe_outbuf_18.X
rlabel metal1 24196 4794 24196 4794 0 strobe_outbuf_19.X
rlabel metal1 12650 5848 12650 5848 0 strobe_outbuf_2.X
rlabel metal1 6348 5882 6348 5882 0 strobe_outbuf_3.X
rlabel metal1 7498 5882 7498 5882 0 strobe_outbuf_4.X
rlabel metal1 8694 5882 8694 5882 0 strobe_outbuf_5.X
rlabel metal2 9706 6086 9706 6086 0 strobe_outbuf_6.X
rlabel metal1 11040 5882 11040 5882 0 strobe_outbuf_7.X
rlabel metal1 12328 5882 12328 5882 0 strobe_outbuf_8.X
rlabel metal1 13432 5882 13432 5882 0 strobe_outbuf_9.X
<< properties >>
string FIXED_BBOX 0 0 26000 8000
<< end >>
