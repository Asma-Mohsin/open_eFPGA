magic
tech sky130A
magscale 1 2
timestamp 1733326700
<< obsli1 >>
rect 460 1071 44528 43537
<< obsm1 >>
rect 14 76 44974 44804
<< metal2 >>
rect 5170 44840 5226 45000
rect 5446 44840 5502 45000
rect 5722 44840 5778 45000
rect 5998 44840 6054 45000
rect 6274 44840 6330 45000
rect 6550 44840 6606 45000
rect 6826 44840 6882 45000
rect 7102 44840 7158 45000
rect 7378 44840 7434 45000
rect 7654 44840 7710 45000
rect 7930 44840 7986 45000
rect 8206 44840 8262 45000
rect 8482 44840 8538 45000
rect 8758 44840 8814 45000
rect 9034 44840 9090 45000
rect 9310 44840 9366 45000
rect 9586 44840 9642 45000
rect 9862 44840 9918 45000
rect 10138 44840 10194 45000
rect 10414 44840 10470 45000
rect 10690 44840 10746 45000
rect 10966 44840 11022 45000
rect 11242 44840 11298 45000
rect 11518 44840 11574 45000
rect 11794 44840 11850 45000
rect 12070 44840 12126 45000
rect 12346 44840 12402 45000
rect 12622 44840 12678 45000
rect 12898 44840 12954 45000
rect 13174 44840 13230 45000
rect 13450 44840 13506 45000
rect 13726 44840 13782 45000
rect 14002 44840 14058 45000
rect 14278 44840 14334 45000
rect 14554 44840 14610 45000
rect 14830 44840 14886 45000
rect 15106 44840 15162 45000
rect 15382 44840 15438 45000
rect 15658 44840 15714 45000
rect 15934 44840 15990 45000
rect 16210 44840 16266 45000
rect 16486 44840 16542 45000
rect 16762 44840 16818 45000
rect 17038 44840 17094 45000
rect 17314 44840 17370 45000
rect 17590 44840 17646 45000
rect 17866 44840 17922 45000
rect 18142 44840 18198 45000
rect 18418 44840 18474 45000
rect 18694 44840 18750 45000
rect 18970 44840 19026 45000
rect 19246 44840 19302 45000
rect 19522 44840 19578 45000
rect 19798 44840 19854 45000
rect 20074 44840 20130 45000
rect 20350 44840 20406 45000
rect 20626 44840 20682 45000
rect 20902 44840 20958 45000
rect 21178 44840 21234 45000
rect 21454 44840 21510 45000
rect 21730 44840 21786 45000
rect 22006 44840 22062 45000
rect 22282 44840 22338 45000
rect 22558 44840 22614 45000
rect 22834 44840 22890 45000
rect 23110 44840 23166 45000
rect 23386 44840 23442 45000
rect 23662 44840 23718 45000
rect 23938 44840 23994 45000
rect 24214 44840 24270 45000
rect 24490 44840 24546 45000
rect 24766 44840 24822 45000
rect 25042 44840 25098 45000
rect 25318 44840 25374 45000
rect 25594 44840 25650 45000
rect 25870 44840 25926 45000
rect 26146 44840 26202 45000
rect 26422 44840 26478 45000
rect 26698 44840 26754 45000
rect 26974 44840 27030 45000
rect 27250 44840 27306 45000
rect 27526 44840 27582 45000
rect 27802 44840 27858 45000
rect 28078 44840 28134 45000
rect 28354 44840 28410 45000
rect 28630 44840 28686 45000
rect 28906 44840 28962 45000
rect 29182 44840 29238 45000
rect 29458 44840 29514 45000
rect 29734 44840 29790 45000
rect 30010 44840 30066 45000
rect 30286 44840 30342 45000
rect 30562 44840 30618 45000
rect 30838 44840 30894 45000
rect 31114 44840 31170 45000
rect 31390 44840 31446 45000
rect 31666 44840 31722 45000
rect 31942 44840 31998 45000
rect 32218 44840 32274 45000
rect 32494 44840 32550 45000
rect 32770 44840 32826 45000
rect 33046 44840 33102 45000
rect 33322 44840 33378 45000
rect 33598 44840 33654 45000
rect 33874 44840 33930 45000
rect 34150 44840 34206 45000
rect 34426 44840 34482 45000
rect 34702 44840 34758 45000
rect 34978 44840 35034 45000
rect 35254 44840 35310 45000
rect 35530 44840 35586 45000
rect 35806 44840 35862 45000
rect 36082 44840 36138 45000
rect 36358 44840 36414 45000
rect 36634 44840 36690 45000
rect 36910 44840 36966 45000
rect 37186 44840 37242 45000
rect 37462 44840 37518 45000
rect 37738 44840 37794 45000
rect 38014 44840 38070 45000
rect 38290 44840 38346 45000
rect 38566 44840 38622 45000
rect 38842 44840 38898 45000
rect 39118 44840 39174 45000
rect 39394 44840 39450 45000
rect 39670 44840 39726 45000
rect 5170 0 5226 160
rect 5446 0 5502 160
rect 5722 0 5778 160
rect 5998 0 6054 160
rect 6274 0 6330 160
rect 6550 0 6606 160
rect 6826 0 6882 160
rect 7102 0 7158 160
rect 7378 0 7434 160
rect 7654 0 7710 160
rect 7930 0 7986 160
rect 8206 0 8262 160
rect 8482 0 8538 160
rect 8758 0 8814 160
rect 9034 0 9090 160
rect 9310 0 9366 160
rect 9586 0 9642 160
rect 9862 0 9918 160
rect 10138 0 10194 160
rect 10414 0 10470 160
rect 10690 0 10746 160
rect 10966 0 11022 160
rect 11242 0 11298 160
rect 11518 0 11574 160
rect 11794 0 11850 160
rect 12070 0 12126 160
rect 12346 0 12402 160
rect 12622 0 12678 160
rect 12898 0 12954 160
rect 13174 0 13230 160
rect 13450 0 13506 160
rect 13726 0 13782 160
rect 14002 0 14058 160
rect 14278 0 14334 160
rect 14554 0 14610 160
rect 14830 0 14886 160
rect 15106 0 15162 160
rect 15382 0 15438 160
rect 15658 0 15714 160
rect 15934 0 15990 160
rect 16210 0 16266 160
rect 16486 0 16542 160
rect 16762 0 16818 160
rect 17038 0 17094 160
rect 17314 0 17370 160
rect 17590 0 17646 160
rect 17866 0 17922 160
rect 18142 0 18198 160
rect 18418 0 18474 160
rect 18694 0 18750 160
rect 18970 0 19026 160
rect 19246 0 19302 160
rect 19522 0 19578 160
rect 19798 0 19854 160
rect 20074 0 20130 160
rect 20350 0 20406 160
rect 20626 0 20682 160
rect 20902 0 20958 160
rect 21178 0 21234 160
rect 21454 0 21510 160
rect 21730 0 21786 160
rect 22006 0 22062 160
rect 22282 0 22338 160
rect 22558 0 22614 160
rect 22834 0 22890 160
rect 23110 0 23166 160
rect 23386 0 23442 160
rect 23662 0 23718 160
rect 23938 0 23994 160
rect 24214 0 24270 160
rect 24490 0 24546 160
rect 24766 0 24822 160
rect 25042 0 25098 160
rect 25318 0 25374 160
rect 25594 0 25650 160
rect 25870 0 25926 160
rect 26146 0 26202 160
rect 26422 0 26478 160
rect 26698 0 26754 160
rect 26974 0 27030 160
rect 27250 0 27306 160
rect 27526 0 27582 160
rect 27802 0 27858 160
rect 28078 0 28134 160
rect 28354 0 28410 160
rect 28630 0 28686 160
rect 28906 0 28962 160
rect 29182 0 29238 160
rect 29458 0 29514 160
rect 29734 0 29790 160
rect 30010 0 30066 160
rect 30286 0 30342 160
rect 30562 0 30618 160
rect 30838 0 30894 160
rect 31114 0 31170 160
rect 31390 0 31446 160
rect 31666 0 31722 160
rect 31942 0 31998 160
rect 32218 0 32274 160
rect 32494 0 32550 160
rect 32770 0 32826 160
rect 33046 0 33102 160
rect 33322 0 33378 160
rect 33598 0 33654 160
rect 33874 0 33930 160
rect 34150 0 34206 160
rect 34426 0 34482 160
rect 34702 0 34758 160
rect 34978 0 35034 160
rect 35254 0 35310 160
rect 35530 0 35586 160
rect 35806 0 35862 160
rect 36082 0 36138 160
rect 36358 0 36414 160
rect 36634 0 36690 160
rect 36910 0 36966 160
rect 37186 0 37242 160
rect 37462 0 37518 160
rect 37738 0 37794 160
rect 38014 0 38070 160
rect 38290 0 38346 160
rect 38566 0 38622 160
rect 38842 0 38898 160
rect 39118 0 39174 160
rect 39394 0 39450 160
rect 39670 0 39726 160
<< obsm2 >>
rect 20 44784 5114 44962
rect 5282 44784 5390 44962
rect 5558 44784 5666 44962
rect 5834 44784 5942 44962
rect 6110 44784 6218 44962
rect 6386 44784 6494 44962
rect 6662 44784 6770 44962
rect 6938 44784 7046 44962
rect 7214 44784 7322 44962
rect 7490 44784 7598 44962
rect 7766 44784 7874 44962
rect 8042 44784 8150 44962
rect 8318 44784 8426 44962
rect 8594 44784 8702 44962
rect 8870 44784 8978 44962
rect 9146 44784 9254 44962
rect 9422 44784 9530 44962
rect 9698 44784 9806 44962
rect 9974 44784 10082 44962
rect 10250 44784 10358 44962
rect 10526 44784 10634 44962
rect 10802 44784 10910 44962
rect 11078 44784 11186 44962
rect 11354 44784 11462 44962
rect 11630 44784 11738 44962
rect 11906 44784 12014 44962
rect 12182 44784 12290 44962
rect 12458 44784 12566 44962
rect 12734 44784 12842 44962
rect 13010 44784 13118 44962
rect 13286 44784 13394 44962
rect 13562 44784 13670 44962
rect 13838 44784 13946 44962
rect 14114 44784 14222 44962
rect 14390 44784 14498 44962
rect 14666 44784 14774 44962
rect 14942 44784 15050 44962
rect 15218 44784 15326 44962
rect 15494 44784 15602 44962
rect 15770 44784 15878 44962
rect 16046 44784 16154 44962
rect 16322 44784 16430 44962
rect 16598 44784 16706 44962
rect 16874 44784 16982 44962
rect 17150 44784 17258 44962
rect 17426 44784 17534 44962
rect 17702 44784 17810 44962
rect 17978 44784 18086 44962
rect 18254 44784 18362 44962
rect 18530 44784 18638 44962
rect 18806 44784 18914 44962
rect 19082 44784 19190 44962
rect 19358 44784 19466 44962
rect 19634 44784 19742 44962
rect 19910 44784 20018 44962
rect 20186 44784 20294 44962
rect 20462 44784 20570 44962
rect 20738 44784 20846 44962
rect 21014 44784 21122 44962
rect 21290 44784 21398 44962
rect 21566 44784 21674 44962
rect 21842 44784 21950 44962
rect 22118 44784 22226 44962
rect 22394 44784 22502 44962
rect 22670 44784 22778 44962
rect 22946 44784 23054 44962
rect 23222 44784 23330 44962
rect 23498 44784 23606 44962
rect 23774 44784 23882 44962
rect 24050 44784 24158 44962
rect 24326 44784 24434 44962
rect 24602 44784 24710 44962
rect 24878 44784 24986 44962
rect 25154 44784 25262 44962
rect 25430 44784 25538 44962
rect 25706 44784 25814 44962
rect 25982 44784 26090 44962
rect 26258 44784 26366 44962
rect 26534 44784 26642 44962
rect 26810 44784 26918 44962
rect 27086 44784 27194 44962
rect 27362 44784 27470 44962
rect 27638 44784 27746 44962
rect 27914 44784 28022 44962
rect 28190 44784 28298 44962
rect 28466 44784 28574 44962
rect 28742 44784 28850 44962
rect 29018 44784 29126 44962
rect 29294 44784 29402 44962
rect 29570 44784 29678 44962
rect 29846 44784 29954 44962
rect 30122 44784 30230 44962
rect 30398 44784 30506 44962
rect 30674 44784 30782 44962
rect 30950 44784 31058 44962
rect 31226 44784 31334 44962
rect 31502 44784 31610 44962
rect 31778 44784 31886 44962
rect 32054 44784 32162 44962
rect 32330 44784 32438 44962
rect 32606 44784 32714 44962
rect 32882 44784 32990 44962
rect 33158 44784 33266 44962
rect 33434 44784 33542 44962
rect 33710 44784 33818 44962
rect 33986 44784 34094 44962
rect 34262 44784 34370 44962
rect 34538 44784 34646 44962
rect 34814 44784 34922 44962
rect 35090 44784 35198 44962
rect 35366 44784 35474 44962
rect 35642 44784 35750 44962
rect 35918 44784 36026 44962
rect 36194 44784 36302 44962
rect 36470 44784 36578 44962
rect 36746 44784 36854 44962
rect 37022 44784 37130 44962
rect 37298 44784 37406 44962
rect 37574 44784 37682 44962
rect 37850 44784 37958 44962
rect 38126 44784 38234 44962
rect 38402 44784 38510 44962
rect 38678 44784 38786 44962
rect 38954 44784 39062 44962
rect 39230 44784 39338 44962
rect 39506 44784 39614 44962
rect 39782 44784 44968 44962
rect 20 216 44968 44784
rect 20 31 5114 216
rect 5282 31 5390 216
rect 5558 31 5666 216
rect 5834 31 5942 216
rect 6110 31 6218 216
rect 6386 31 6494 216
rect 6662 31 6770 216
rect 6938 31 7046 216
rect 7214 31 7322 216
rect 7490 31 7598 216
rect 7766 31 7874 216
rect 8042 31 8150 216
rect 8318 31 8426 216
rect 8594 31 8702 216
rect 8870 31 8978 216
rect 9146 31 9254 216
rect 9422 31 9530 216
rect 9698 31 9806 216
rect 9974 31 10082 216
rect 10250 31 10358 216
rect 10526 31 10634 216
rect 10802 31 10910 216
rect 11078 31 11186 216
rect 11354 31 11462 216
rect 11630 31 11738 216
rect 11906 31 12014 216
rect 12182 31 12290 216
rect 12458 31 12566 216
rect 12734 31 12842 216
rect 13010 31 13118 216
rect 13286 31 13394 216
rect 13562 31 13670 216
rect 13838 31 13946 216
rect 14114 31 14222 216
rect 14390 31 14498 216
rect 14666 31 14774 216
rect 14942 31 15050 216
rect 15218 31 15326 216
rect 15494 31 15602 216
rect 15770 31 15878 216
rect 16046 31 16154 216
rect 16322 31 16430 216
rect 16598 31 16706 216
rect 16874 31 16982 216
rect 17150 31 17258 216
rect 17426 31 17534 216
rect 17702 31 17810 216
rect 17978 31 18086 216
rect 18254 31 18362 216
rect 18530 31 18638 216
rect 18806 31 18914 216
rect 19082 31 19190 216
rect 19358 31 19466 216
rect 19634 31 19742 216
rect 19910 31 20018 216
rect 20186 31 20294 216
rect 20462 31 20570 216
rect 20738 31 20846 216
rect 21014 31 21122 216
rect 21290 31 21398 216
rect 21566 31 21674 216
rect 21842 31 21950 216
rect 22118 31 22226 216
rect 22394 31 22502 216
rect 22670 31 22778 216
rect 22946 31 23054 216
rect 23222 31 23330 216
rect 23498 31 23606 216
rect 23774 31 23882 216
rect 24050 31 24158 216
rect 24326 31 24434 216
rect 24602 31 24710 216
rect 24878 31 24986 216
rect 25154 31 25262 216
rect 25430 31 25538 216
rect 25706 31 25814 216
rect 25982 31 26090 216
rect 26258 31 26366 216
rect 26534 31 26642 216
rect 26810 31 26918 216
rect 27086 31 27194 216
rect 27362 31 27470 216
rect 27638 31 27746 216
rect 27914 31 28022 216
rect 28190 31 28298 216
rect 28466 31 28574 216
rect 28742 31 28850 216
rect 29018 31 29126 216
rect 29294 31 29402 216
rect 29570 31 29678 216
rect 29846 31 29954 216
rect 30122 31 30230 216
rect 30398 31 30506 216
rect 30674 31 30782 216
rect 30950 31 31058 216
rect 31226 31 31334 216
rect 31502 31 31610 216
rect 31778 31 31886 216
rect 32054 31 32162 216
rect 32330 31 32438 216
rect 32606 31 32714 216
rect 32882 31 32990 216
rect 33158 31 33266 216
rect 33434 31 33542 216
rect 33710 31 33818 216
rect 33986 31 34094 216
rect 34262 31 34370 216
rect 34538 31 34646 216
rect 34814 31 34922 216
rect 35090 31 35198 216
rect 35366 31 35474 216
rect 35642 31 35750 216
rect 35918 31 36026 216
rect 36194 31 36302 216
rect 36470 31 36578 216
rect 36746 31 36854 216
rect 37022 31 37130 216
rect 37298 31 37406 216
rect 37574 31 37682 216
rect 37850 31 37958 216
rect 38126 31 38234 216
rect 38402 31 38510 216
rect 38678 31 38786 216
rect 38954 31 39062 216
rect 39230 31 39338 216
rect 39506 31 39614 216
rect 39782 31 44968 216
<< metal3 >>
rect 0 39720 160 39840
rect 0 39448 160 39568
rect 0 39176 160 39296
rect 0 38904 160 39024
rect 0 38632 160 38752
rect 0 38360 160 38480
rect 0 38088 160 38208
rect 0 37816 160 37936
rect 0 37544 160 37664
rect 0 37272 160 37392
rect 0 37000 160 37120
rect 0 36728 160 36848
rect 0 36456 160 36576
rect 0 36184 160 36304
rect 0 35912 160 36032
rect 0 35640 160 35760
rect 0 35368 160 35488
rect 0 35096 160 35216
rect 0 34824 160 34944
rect 0 34552 160 34672
rect 0 34280 160 34400
rect 0 34008 160 34128
rect 0 33736 160 33856
rect 0 33464 160 33584
rect 0 33192 160 33312
rect 0 32920 160 33040
rect 0 32648 160 32768
rect 0 32376 160 32496
rect 0 32104 160 32224
rect 0 31832 160 31952
rect 0 31560 160 31680
rect 0 31288 160 31408
rect 0 31016 160 31136
rect 0 30744 160 30864
rect 0 30472 160 30592
rect 0 30200 160 30320
rect 0 29928 160 30048
rect 0 29656 160 29776
rect 0 29384 160 29504
rect 0 29112 160 29232
rect 0 28840 160 28960
rect 0 28568 160 28688
rect 0 28296 160 28416
rect 0 28024 160 28144
rect 0 27752 160 27872
rect 0 27480 160 27600
rect 0 27208 160 27328
rect 0 26936 160 27056
rect 0 26664 160 26784
rect 0 26392 160 26512
rect 0 26120 160 26240
rect 0 25848 160 25968
rect 0 25576 160 25696
rect 0 25304 160 25424
rect 0 25032 160 25152
rect 0 24760 160 24880
rect 0 24488 160 24608
rect 0 24216 160 24336
rect 0 23944 160 24064
rect 0 23672 160 23792
rect 0 23400 160 23520
rect 0 23128 160 23248
rect 0 22856 160 22976
rect 0 22584 160 22704
rect 0 22312 160 22432
rect 0 22040 160 22160
rect 0 21768 160 21888
rect 0 21496 160 21616
rect 0 21224 160 21344
rect 0 20952 160 21072
rect 0 20680 160 20800
rect 0 20408 160 20528
rect 0 20136 160 20256
rect 0 19864 160 19984
rect 0 19592 160 19712
rect 0 19320 160 19440
rect 0 19048 160 19168
rect 0 18776 160 18896
rect 0 18504 160 18624
rect 0 18232 160 18352
rect 0 17960 160 18080
rect 0 17688 160 17808
rect 0 17416 160 17536
rect 0 17144 160 17264
rect 0 16872 160 16992
rect 0 16600 160 16720
rect 0 16328 160 16448
rect 0 16056 160 16176
rect 0 15784 160 15904
rect 0 15512 160 15632
rect 0 15240 160 15360
rect 0 14968 160 15088
rect 0 14696 160 14816
rect 0 14424 160 14544
rect 0 14152 160 14272
rect 0 13880 160 14000
rect 0 13608 160 13728
rect 0 13336 160 13456
rect 0 13064 160 13184
rect 0 12792 160 12912
rect 0 12520 160 12640
rect 0 12248 160 12368
rect 0 11976 160 12096
rect 0 11704 160 11824
rect 0 11432 160 11552
rect 0 11160 160 11280
rect 0 10888 160 11008
rect 0 10616 160 10736
rect 0 10344 160 10464
rect 0 10072 160 10192
rect 0 9800 160 9920
rect 0 9528 160 9648
rect 0 9256 160 9376
rect 0 8984 160 9104
rect 0 8712 160 8832
rect 0 8440 160 8560
rect 0 8168 160 8288
rect 0 7896 160 8016
rect 0 7624 160 7744
rect 0 7352 160 7472
rect 0 7080 160 7200
rect 0 6808 160 6928
rect 0 6536 160 6656
rect 0 6264 160 6384
rect 0 5992 160 6112
rect 0 5720 160 5840
rect 0 5448 160 5568
rect 0 5176 160 5296
rect 44840 39720 45000 39840
rect 44840 39448 45000 39568
rect 44840 39176 45000 39296
rect 44840 38904 45000 39024
rect 44840 38632 45000 38752
rect 44840 38360 45000 38480
rect 44840 38088 45000 38208
rect 44840 37816 45000 37936
rect 44840 37544 45000 37664
rect 44840 37272 45000 37392
rect 44840 37000 45000 37120
rect 44840 36728 45000 36848
rect 44840 36456 45000 36576
rect 44840 36184 45000 36304
rect 44840 35912 45000 36032
rect 44840 35640 45000 35760
rect 44840 35368 45000 35488
rect 44840 35096 45000 35216
rect 44840 34824 45000 34944
rect 44840 34552 45000 34672
rect 44840 34280 45000 34400
rect 44840 34008 45000 34128
rect 44840 33736 45000 33856
rect 44840 33464 45000 33584
rect 44840 33192 45000 33312
rect 44840 32920 45000 33040
rect 44840 32648 45000 32768
rect 44840 32376 45000 32496
rect 44840 32104 45000 32224
rect 44840 31832 45000 31952
rect 44840 31560 45000 31680
rect 44840 31288 45000 31408
rect 44840 31016 45000 31136
rect 44840 30744 45000 30864
rect 44840 30472 45000 30592
rect 44840 30200 45000 30320
rect 44840 29928 45000 30048
rect 44840 29656 45000 29776
rect 44840 29384 45000 29504
rect 44840 29112 45000 29232
rect 44840 28840 45000 28960
rect 44840 28568 45000 28688
rect 44840 28296 45000 28416
rect 44840 28024 45000 28144
rect 44840 27752 45000 27872
rect 44840 27480 45000 27600
rect 44840 27208 45000 27328
rect 44840 26936 45000 27056
rect 44840 26664 45000 26784
rect 44840 26392 45000 26512
rect 44840 26120 45000 26240
rect 44840 25848 45000 25968
rect 44840 25576 45000 25696
rect 44840 25304 45000 25424
rect 44840 25032 45000 25152
rect 44840 24760 45000 24880
rect 44840 24488 45000 24608
rect 44840 24216 45000 24336
rect 44840 23944 45000 24064
rect 44840 23672 45000 23792
rect 44840 23400 45000 23520
rect 44840 23128 45000 23248
rect 44840 22856 45000 22976
rect 44840 22584 45000 22704
rect 44840 22312 45000 22432
rect 44840 22040 45000 22160
rect 44840 21768 45000 21888
rect 44840 21496 45000 21616
rect 44840 21224 45000 21344
rect 44840 20952 45000 21072
rect 44840 20680 45000 20800
rect 44840 20408 45000 20528
rect 44840 20136 45000 20256
rect 44840 19864 45000 19984
rect 44840 19592 45000 19712
rect 44840 19320 45000 19440
rect 44840 19048 45000 19168
rect 44840 18776 45000 18896
rect 44840 18504 45000 18624
rect 44840 18232 45000 18352
rect 44840 17960 45000 18080
rect 44840 17688 45000 17808
rect 44840 17416 45000 17536
rect 44840 17144 45000 17264
rect 44840 16872 45000 16992
rect 44840 16600 45000 16720
rect 44840 16328 45000 16448
rect 44840 16056 45000 16176
rect 44840 15784 45000 15904
rect 44840 15512 45000 15632
rect 44840 15240 45000 15360
rect 44840 14968 45000 15088
rect 44840 14696 45000 14816
rect 44840 14424 45000 14544
rect 44840 14152 45000 14272
rect 44840 13880 45000 14000
rect 44840 13608 45000 13728
rect 44840 13336 45000 13456
rect 44840 13064 45000 13184
rect 44840 12792 45000 12912
rect 44840 12520 45000 12640
rect 44840 12248 45000 12368
rect 44840 11976 45000 12096
rect 44840 11704 45000 11824
rect 44840 11432 45000 11552
rect 44840 11160 45000 11280
rect 44840 10888 45000 11008
rect 44840 10616 45000 10736
rect 44840 10344 45000 10464
rect 44840 10072 45000 10192
rect 44840 9800 45000 9920
rect 44840 9528 45000 9648
rect 44840 9256 45000 9376
rect 44840 8984 45000 9104
rect 44840 8712 45000 8832
rect 44840 8440 45000 8560
rect 44840 8168 45000 8288
rect 44840 7896 45000 8016
rect 44840 7624 45000 7744
rect 44840 7352 45000 7472
rect 44840 7080 45000 7200
rect 44840 6808 45000 6928
rect 44840 6536 45000 6656
rect 44840 6264 45000 6384
rect 44840 5992 45000 6112
rect 44840 5720 45000 5840
rect 44840 5448 45000 5568
rect 44840 5176 45000 5296
<< obsm3 >>
rect 160 39920 44883 43892
rect 240 5096 44760 39920
rect 160 35 44883 5096
<< metal4 >>
rect 3564 1040 3884 43568
rect 11064 1040 11384 43568
rect 18564 1040 18884 43568
rect 26064 1040 26384 43568
rect 33564 1040 33884 43568
rect 41064 1040 41384 43568
<< obsm4 >>
rect 427 43648 44469 43893
rect 427 960 3484 43648
rect 3964 960 10984 43648
rect 11464 960 18484 43648
rect 18964 960 25984 43648
rect 26464 960 33484 43648
rect 33964 960 40984 43648
rect 41464 960 44469 43648
rect 427 35 44469 960
<< labels >>
rlabel metal2 s 34150 0 34206 160 6 Ci
port 1 nsew signal input
rlabel metal2 s 34150 44840 34206 45000 6 Co
port 2 nsew signal output
rlabel metal3 s 44840 18232 45000 18352 6 E1BEG[0]
port 3 nsew signal output
rlabel metal3 s 44840 18504 45000 18624 6 E1BEG[1]
port 4 nsew signal output
rlabel metal3 s 44840 18776 45000 18896 6 E1BEG[2]
port 5 nsew signal output
rlabel metal3 s 44840 19048 45000 19168 6 E1BEG[3]
port 6 nsew signal output
rlabel metal3 s 0 18232 160 18352 6 E1END[0]
port 7 nsew signal input
rlabel metal3 s 0 18504 160 18624 6 E1END[1]
port 8 nsew signal input
rlabel metal3 s 0 18776 160 18896 6 E1END[2]
port 9 nsew signal input
rlabel metal3 s 0 19048 160 19168 6 E1END[3]
port 10 nsew signal input
rlabel metal3 s 44840 19320 45000 19440 6 E2BEG[0]
port 11 nsew signal output
rlabel metal3 s 44840 19592 45000 19712 6 E2BEG[1]
port 12 nsew signal output
rlabel metal3 s 44840 19864 45000 19984 6 E2BEG[2]
port 13 nsew signal output
rlabel metal3 s 44840 20136 45000 20256 6 E2BEG[3]
port 14 nsew signal output
rlabel metal3 s 44840 20408 45000 20528 6 E2BEG[4]
port 15 nsew signal output
rlabel metal3 s 44840 20680 45000 20800 6 E2BEG[5]
port 16 nsew signal output
rlabel metal3 s 44840 20952 45000 21072 6 E2BEG[6]
port 17 nsew signal output
rlabel metal3 s 44840 21224 45000 21344 6 E2BEG[7]
port 18 nsew signal output
rlabel metal3 s 44840 21496 45000 21616 6 E2BEGb[0]
port 19 nsew signal output
rlabel metal3 s 44840 21768 45000 21888 6 E2BEGb[1]
port 20 nsew signal output
rlabel metal3 s 44840 22040 45000 22160 6 E2BEGb[2]
port 21 nsew signal output
rlabel metal3 s 44840 22312 45000 22432 6 E2BEGb[3]
port 22 nsew signal output
rlabel metal3 s 44840 22584 45000 22704 6 E2BEGb[4]
port 23 nsew signal output
rlabel metal3 s 44840 22856 45000 22976 6 E2BEGb[5]
port 24 nsew signal output
rlabel metal3 s 44840 23128 45000 23248 6 E2BEGb[6]
port 25 nsew signal output
rlabel metal3 s 44840 23400 45000 23520 6 E2BEGb[7]
port 26 nsew signal output
rlabel metal3 s 0 21496 160 21616 6 E2END[0]
port 27 nsew signal input
rlabel metal3 s 0 21768 160 21888 6 E2END[1]
port 28 nsew signal input
rlabel metal3 s 0 22040 160 22160 6 E2END[2]
port 29 nsew signal input
rlabel metal3 s 0 22312 160 22432 6 E2END[3]
port 30 nsew signal input
rlabel metal3 s 0 22584 160 22704 6 E2END[4]
port 31 nsew signal input
rlabel metal3 s 0 22856 160 22976 6 E2END[5]
port 32 nsew signal input
rlabel metal3 s 0 23128 160 23248 6 E2END[6]
port 33 nsew signal input
rlabel metal3 s 0 23400 160 23520 6 E2END[7]
port 34 nsew signal input
rlabel metal3 s 0 19320 160 19440 6 E2MID[0]
port 35 nsew signal input
rlabel metal3 s 0 19592 160 19712 6 E2MID[1]
port 36 nsew signal input
rlabel metal3 s 0 19864 160 19984 6 E2MID[2]
port 37 nsew signal input
rlabel metal3 s 0 20136 160 20256 6 E2MID[3]
port 38 nsew signal input
rlabel metal3 s 0 20408 160 20528 6 E2MID[4]
port 39 nsew signal input
rlabel metal3 s 0 20680 160 20800 6 E2MID[5]
port 40 nsew signal input
rlabel metal3 s 0 20952 160 21072 6 E2MID[6]
port 41 nsew signal input
rlabel metal3 s 0 21224 160 21344 6 E2MID[7]
port 42 nsew signal input
rlabel metal3 s 44840 28024 45000 28144 6 E6BEG[0]
port 43 nsew signal output
rlabel metal3 s 44840 30744 45000 30864 6 E6BEG[10]
port 44 nsew signal output
rlabel metal3 s 44840 31016 45000 31136 6 E6BEG[11]
port 45 nsew signal output
rlabel metal3 s 44840 28296 45000 28416 6 E6BEG[1]
port 46 nsew signal output
rlabel metal3 s 44840 28568 45000 28688 6 E6BEG[2]
port 47 nsew signal output
rlabel metal3 s 44840 28840 45000 28960 6 E6BEG[3]
port 48 nsew signal output
rlabel metal3 s 44840 29112 45000 29232 6 E6BEG[4]
port 49 nsew signal output
rlabel metal3 s 44840 29384 45000 29504 6 E6BEG[5]
port 50 nsew signal output
rlabel metal3 s 44840 29656 45000 29776 6 E6BEG[6]
port 51 nsew signal output
rlabel metal3 s 44840 29928 45000 30048 6 E6BEG[7]
port 52 nsew signal output
rlabel metal3 s 44840 30200 45000 30320 6 E6BEG[8]
port 53 nsew signal output
rlabel metal3 s 44840 30472 45000 30592 6 E6BEG[9]
port 54 nsew signal output
rlabel metal3 s 0 28024 160 28144 6 E6END[0]
port 55 nsew signal input
rlabel metal3 s 0 30744 160 30864 6 E6END[10]
port 56 nsew signal input
rlabel metal3 s 0 31016 160 31136 6 E6END[11]
port 57 nsew signal input
rlabel metal3 s 0 28296 160 28416 6 E6END[1]
port 58 nsew signal input
rlabel metal3 s 0 28568 160 28688 6 E6END[2]
port 59 nsew signal input
rlabel metal3 s 0 28840 160 28960 6 E6END[3]
port 60 nsew signal input
rlabel metal3 s 0 29112 160 29232 6 E6END[4]
port 61 nsew signal input
rlabel metal3 s 0 29384 160 29504 6 E6END[5]
port 62 nsew signal input
rlabel metal3 s 0 29656 160 29776 6 E6END[6]
port 63 nsew signal input
rlabel metal3 s 0 29928 160 30048 6 E6END[7]
port 64 nsew signal input
rlabel metal3 s 0 30200 160 30320 6 E6END[8]
port 65 nsew signal input
rlabel metal3 s 0 30472 160 30592 6 E6END[9]
port 66 nsew signal input
rlabel metal3 s 44840 23672 45000 23792 6 EE4BEG[0]
port 67 nsew signal output
rlabel metal3 s 44840 26392 45000 26512 6 EE4BEG[10]
port 68 nsew signal output
rlabel metal3 s 44840 26664 45000 26784 6 EE4BEG[11]
port 69 nsew signal output
rlabel metal3 s 44840 26936 45000 27056 6 EE4BEG[12]
port 70 nsew signal output
rlabel metal3 s 44840 27208 45000 27328 6 EE4BEG[13]
port 71 nsew signal output
rlabel metal3 s 44840 27480 45000 27600 6 EE4BEG[14]
port 72 nsew signal output
rlabel metal3 s 44840 27752 45000 27872 6 EE4BEG[15]
port 73 nsew signal output
rlabel metal3 s 44840 23944 45000 24064 6 EE4BEG[1]
port 74 nsew signal output
rlabel metal3 s 44840 24216 45000 24336 6 EE4BEG[2]
port 75 nsew signal output
rlabel metal3 s 44840 24488 45000 24608 6 EE4BEG[3]
port 76 nsew signal output
rlabel metal3 s 44840 24760 45000 24880 6 EE4BEG[4]
port 77 nsew signal output
rlabel metal3 s 44840 25032 45000 25152 6 EE4BEG[5]
port 78 nsew signal output
rlabel metal3 s 44840 25304 45000 25424 6 EE4BEG[6]
port 79 nsew signal output
rlabel metal3 s 44840 25576 45000 25696 6 EE4BEG[7]
port 80 nsew signal output
rlabel metal3 s 44840 25848 45000 25968 6 EE4BEG[8]
port 81 nsew signal output
rlabel metal3 s 44840 26120 45000 26240 6 EE4BEG[9]
port 82 nsew signal output
rlabel metal3 s 0 23672 160 23792 6 EE4END[0]
port 83 nsew signal input
rlabel metal3 s 0 26392 160 26512 6 EE4END[10]
port 84 nsew signal input
rlabel metal3 s 0 26664 160 26784 6 EE4END[11]
port 85 nsew signal input
rlabel metal3 s 0 26936 160 27056 6 EE4END[12]
port 86 nsew signal input
rlabel metal3 s 0 27208 160 27328 6 EE4END[13]
port 87 nsew signal input
rlabel metal3 s 0 27480 160 27600 6 EE4END[14]
port 88 nsew signal input
rlabel metal3 s 0 27752 160 27872 6 EE4END[15]
port 89 nsew signal input
rlabel metal3 s 0 23944 160 24064 6 EE4END[1]
port 90 nsew signal input
rlabel metal3 s 0 24216 160 24336 6 EE4END[2]
port 91 nsew signal input
rlabel metal3 s 0 24488 160 24608 6 EE4END[3]
port 92 nsew signal input
rlabel metal3 s 0 24760 160 24880 6 EE4END[4]
port 93 nsew signal input
rlabel metal3 s 0 25032 160 25152 6 EE4END[5]
port 94 nsew signal input
rlabel metal3 s 0 25304 160 25424 6 EE4END[6]
port 95 nsew signal input
rlabel metal3 s 0 25576 160 25696 6 EE4END[7]
port 96 nsew signal input
rlabel metal3 s 0 25848 160 25968 6 EE4END[8]
port 97 nsew signal input
rlabel metal3 s 0 26120 160 26240 6 EE4END[9]
port 98 nsew signal input
rlabel metal3 s 0 31288 160 31408 6 FrameData[0]
port 99 nsew signal input
rlabel metal3 s 0 34008 160 34128 6 FrameData[10]
port 100 nsew signal input
rlabel metal3 s 0 34280 160 34400 6 FrameData[11]
port 101 nsew signal input
rlabel metal3 s 0 34552 160 34672 6 FrameData[12]
port 102 nsew signal input
rlabel metal3 s 0 34824 160 34944 6 FrameData[13]
port 103 nsew signal input
rlabel metal3 s 0 35096 160 35216 6 FrameData[14]
port 104 nsew signal input
rlabel metal3 s 0 35368 160 35488 6 FrameData[15]
port 105 nsew signal input
rlabel metal3 s 0 35640 160 35760 6 FrameData[16]
port 106 nsew signal input
rlabel metal3 s 0 35912 160 36032 6 FrameData[17]
port 107 nsew signal input
rlabel metal3 s 0 36184 160 36304 6 FrameData[18]
port 108 nsew signal input
rlabel metal3 s 0 36456 160 36576 6 FrameData[19]
port 109 nsew signal input
rlabel metal3 s 0 31560 160 31680 6 FrameData[1]
port 110 nsew signal input
rlabel metal3 s 0 36728 160 36848 6 FrameData[20]
port 111 nsew signal input
rlabel metal3 s 0 37000 160 37120 6 FrameData[21]
port 112 nsew signal input
rlabel metal3 s 0 37272 160 37392 6 FrameData[22]
port 113 nsew signal input
rlabel metal3 s 0 37544 160 37664 6 FrameData[23]
port 114 nsew signal input
rlabel metal3 s 0 37816 160 37936 6 FrameData[24]
port 115 nsew signal input
rlabel metal3 s 0 38088 160 38208 6 FrameData[25]
port 116 nsew signal input
rlabel metal3 s 0 38360 160 38480 6 FrameData[26]
port 117 nsew signal input
rlabel metal3 s 0 38632 160 38752 6 FrameData[27]
port 118 nsew signal input
rlabel metal3 s 0 38904 160 39024 6 FrameData[28]
port 119 nsew signal input
rlabel metal3 s 0 39176 160 39296 6 FrameData[29]
port 120 nsew signal input
rlabel metal3 s 0 31832 160 31952 6 FrameData[2]
port 121 nsew signal input
rlabel metal3 s 0 39448 160 39568 6 FrameData[30]
port 122 nsew signal input
rlabel metal3 s 0 39720 160 39840 6 FrameData[31]
port 123 nsew signal input
rlabel metal3 s 0 32104 160 32224 6 FrameData[3]
port 124 nsew signal input
rlabel metal3 s 0 32376 160 32496 6 FrameData[4]
port 125 nsew signal input
rlabel metal3 s 0 32648 160 32768 6 FrameData[5]
port 126 nsew signal input
rlabel metal3 s 0 32920 160 33040 6 FrameData[6]
port 127 nsew signal input
rlabel metal3 s 0 33192 160 33312 6 FrameData[7]
port 128 nsew signal input
rlabel metal3 s 0 33464 160 33584 6 FrameData[8]
port 129 nsew signal input
rlabel metal3 s 0 33736 160 33856 6 FrameData[9]
port 130 nsew signal input
rlabel metal3 s 44840 31288 45000 31408 6 FrameData_O[0]
port 131 nsew signal output
rlabel metal3 s 44840 34008 45000 34128 6 FrameData_O[10]
port 132 nsew signal output
rlabel metal3 s 44840 34280 45000 34400 6 FrameData_O[11]
port 133 nsew signal output
rlabel metal3 s 44840 34552 45000 34672 6 FrameData_O[12]
port 134 nsew signal output
rlabel metal3 s 44840 34824 45000 34944 6 FrameData_O[13]
port 135 nsew signal output
rlabel metal3 s 44840 35096 45000 35216 6 FrameData_O[14]
port 136 nsew signal output
rlabel metal3 s 44840 35368 45000 35488 6 FrameData_O[15]
port 137 nsew signal output
rlabel metal3 s 44840 35640 45000 35760 6 FrameData_O[16]
port 138 nsew signal output
rlabel metal3 s 44840 35912 45000 36032 6 FrameData_O[17]
port 139 nsew signal output
rlabel metal3 s 44840 36184 45000 36304 6 FrameData_O[18]
port 140 nsew signal output
rlabel metal3 s 44840 36456 45000 36576 6 FrameData_O[19]
port 141 nsew signal output
rlabel metal3 s 44840 31560 45000 31680 6 FrameData_O[1]
port 142 nsew signal output
rlabel metal3 s 44840 36728 45000 36848 6 FrameData_O[20]
port 143 nsew signal output
rlabel metal3 s 44840 37000 45000 37120 6 FrameData_O[21]
port 144 nsew signal output
rlabel metal3 s 44840 37272 45000 37392 6 FrameData_O[22]
port 145 nsew signal output
rlabel metal3 s 44840 37544 45000 37664 6 FrameData_O[23]
port 146 nsew signal output
rlabel metal3 s 44840 37816 45000 37936 6 FrameData_O[24]
port 147 nsew signal output
rlabel metal3 s 44840 38088 45000 38208 6 FrameData_O[25]
port 148 nsew signal output
rlabel metal3 s 44840 38360 45000 38480 6 FrameData_O[26]
port 149 nsew signal output
rlabel metal3 s 44840 38632 45000 38752 6 FrameData_O[27]
port 150 nsew signal output
rlabel metal3 s 44840 38904 45000 39024 6 FrameData_O[28]
port 151 nsew signal output
rlabel metal3 s 44840 39176 45000 39296 6 FrameData_O[29]
port 152 nsew signal output
rlabel metal3 s 44840 31832 45000 31952 6 FrameData_O[2]
port 153 nsew signal output
rlabel metal3 s 44840 39448 45000 39568 6 FrameData_O[30]
port 154 nsew signal output
rlabel metal3 s 44840 39720 45000 39840 6 FrameData_O[31]
port 155 nsew signal output
rlabel metal3 s 44840 32104 45000 32224 6 FrameData_O[3]
port 156 nsew signal output
rlabel metal3 s 44840 32376 45000 32496 6 FrameData_O[4]
port 157 nsew signal output
rlabel metal3 s 44840 32648 45000 32768 6 FrameData_O[5]
port 158 nsew signal output
rlabel metal3 s 44840 32920 45000 33040 6 FrameData_O[6]
port 159 nsew signal output
rlabel metal3 s 44840 33192 45000 33312 6 FrameData_O[7]
port 160 nsew signal output
rlabel metal3 s 44840 33464 45000 33584 6 FrameData_O[8]
port 161 nsew signal output
rlabel metal3 s 44840 33736 45000 33856 6 FrameData_O[9]
port 162 nsew signal output
rlabel metal2 s 34426 0 34482 160 6 FrameStrobe[0]
port 163 nsew signal input
rlabel metal2 s 37186 0 37242 160 6 FrameStrobe[10]
port 164 nsew signal input
rlabel metal2 s 37462 0 37518 160 6 FrameStrobe[11]
port 165 nsew signal input
rlabel metal2 s 37738 0 37794 160 6 FrameStrobe[12]
port 166 nsew signal input
rlabel metal2 s 38014 0 38070 160 6 FrameStrobe[13]
port 167 nsew signal input
rlabel metal2 s 38290 0 38346 160 6 FrameStrobe[14]
port 168 nsew signal input
rlabel metal2 s 38566 0 38622 160 6 FrameStrobe[15]
port 169 nsew signal input
rlabel metal2 s 38842 0 38898 160 6 FrameStrobe[16]
port 170 nsew signal input
rlabel metal2 s 39118 0 39174 160 6 FrameStrobe[17]
port 171 nsew signal input
rlabel metal2 s 39394 0 39450 160 6 FrameStrobe[18]
port 172 nsew signal input
rlabel metal2 s 39670 0 39726 160 6 FrameStrobe[19]
port 173 nsew signal input
rlabel metal2 s 34702 0 34758 160 6 FrameStrobe[1]
port 174 nsew signal input
rlabel metal2 s 34978 0 35034 160 6 FrameStrobe[2]
port 175 nsew signal input
rlabel metal2 s 35254 0 35310 160 6 FrameStrobe[3]
port 176 nsew signal input
rlabel metal2 s 35530 0 35586 160 6 FrameStrobe[4]
port 177 nsew signal input
rlabel metal2 s 35806 0 35862 160 6 FrameStrobe[5]
port 178 nsew signal input
rlabel metal2 s 36082 0 36138 160 6 FrameStrobe[6]
port 179 nsew signal input
rlabel metal2 s 36358 0 36414 160 6 FrameStrobe[7]
port 180 nsew signal input
rlabel metal2 s 36634 0 36690 160 6 FrameStrobe[8]
port 181 nsew signal input
rlabel metal2 s 36910 0 36966 160 6 FrameStrobe[9]
port 182 nsew signal input
rlabel metal2 s 34426 44840 34482 45000 6 FrameStrobe_O[0]
port 183 nsew signal output
rlabel metal2 s 37186 44840 37242 45000 6 FrameStrobe_O[10]
port 184 nsew signal output
rlabel metal2 s 37462 44840 37518 45000 6 FrameStrobe_O[11]
port 185 nsew signal output
rlabel metal2 s 37738 44840 37794 45000 6 FrameStrobe_O[12]
port 186 nsew signal output
rlabel metal2 s 38014 44840 38070 45000 6 FrameStrobe_O[13]
port 187 nsew signal output
rlabel metal2 s 38290 44840 38346 45000 6 FrameStrobe_O[14]
port 188 nsew signal output
rlabel metal2 s 38566 44840 38622 45000 6 FrameStrobe_O[15]
port 189 nsew signal output
rlabel metal2 s 38842 44840 38898 45000 6 FrameStrobe_O[16]
port 190 nsew signal output
rlabel metal2 s 39118 44840 39174 45000 6 FrameStrobe_O[17]
port 191 nsew signal output
rlabel metal2 s 39394 44840 39450 45000 6 FrameStrobe_O[18]
port 192 nsew signal output
rlabel metal2 s 39670 44840 39726 45000 6 FrameStrobe_O[19]
port 193 nsew signal output
rlabel metal2 s 34702 44840 34758 45000 6 FrameStrobe_O[1]
port 194 nsew signal output
rlabel metal2 s 34978 44840 35034 45000 6 FrameStrobe_O[2]
port 195 nsew signal output
rlabel metal2 s 35254 44840 35310 45000 6 FrameStrobe_O[3]
port 196 nsew signal output
rlabel metal2 s 35530 44840 35586 45000 6 FrameStrobe_O[4]
port 197 nsew signal output
rlabel metal2 s 35806 44840 35862 45000 6 FrameStrobe_O[5]
port 198 nsew signal output
rlabel metal2 s 36082 44840 36138 45000 6 FrameStrobe_O[6]
port 199 nsew signal output
rlabel metal2 s 36358 44840 36414 45000 6 FrameStrobe_O[7]
port 200 nsew signal output
rlabel metal2 s 36634 44840 36690 45000 6 FrameStrobe_O[8]
port 201 nsew signal output
rlabel metal2 s 36910 44840 36966 45000 6 FrameStrobe_O[9]
port 202 nsew signal output
rlabel metal2 s 5170 44840 5226 45000 6 N1BEG[0]
port 203 nsew signal output
rlabel metal2 s 5446 44840 5502 45000 6 N1BEG[1]
port 204 nsew signal output
rlabel metal2 s 5722 44840 5778 45000 6 N1BEG[2]
port 205 nsew signal output
rlabel metal2 s 5998 44840 6054 45000 6 N1BEG[3]
port 206 nsew signal output
rlabel metal2 s 5170 0 5226 160 6 N1END[0]
port 207 nsew signal input
rlabel metal2 s 5446 0 5502 160 6 N1END[1]
port 208 nsew signal input
rlabel metal2 s 5722 0 5778 160 6 N1END[2]
port 209 nsew signal input
rlabel metal2 s 5998 0 6054 160 6 N1END[3]
port 210 nsew signal input
rlabel metal2 s 6274 44840 6330 45000 6 N2BEG[0]
port 211 nsew signal output
rlabel metal2 s 6550 44840 6606 45000 6 N2BEG[1]
port 212 nsew signal output
rlabel metal2 s 6826 44840 6882 45000 6 N2BEG[2]
port 213 nsew signal output
rlabel metal2 s 7102 44840 7158 45000 6 N2BEG[3]
port 214 nsew signal output
rlabel metal2 s 7378 44840 7434 45000 6 N2BEG[4]
port 215 nsew signal output
rlabel metal2 s 7654 44840 7710 45000 6 N2BEG[5]
port 216 nsew signal output
rlabel metal2 s 7930 44840 7986 45000 6 N2BEG[6]
port 217 nsew signal output
rlabel metal2 s 8206 44840 8262 45000 6 N2BEG[7]
port 218 nsew signal output
rlabel metal2 s 8482 44840 8538 45000 6 N2BEGb[0]
port 219 nsew signal output
rlabel metal2 s 8758 44840 8814 45000 6 N2BEGb[1]
port 220 nsew signal output
rlabel metal2 s 9034 44840 9090 45000 6 N2BEGb[2]
port 221 nsew signal output
rlabel metal2 s 9310 44840 9366 45000 6 N2BEGb[3]
port 222 nsew signal output
rlabel metal2 s 9586 44840 9642 45000 6 N2BEGb[4]
port 223 nsew signal output
rlabel metal2 s 9862 44840 9918 45000 6 N2BEGb[5]
port 224 nsew signal output
rlabel metal2 s 10138 44840 10194 45000 6 N2BEGb[6]
port 225 nsew signal output
rlabel metal2 s 10414 44840 10470 45000 6 N2BEGb[7]
port 226 nsew signal output
rlabel metal2 s 8482 0 8538 160 6 N2END[0]
port 227 nsew signal input
rlabel metal2 s 8758 0 8814 160 6 N2END[1]
port 228 nsew signal input
rlabel metal2 s 9034 0 9090 160 6 N2END[2]
port 229 nsew signal input
rlabel metal2 s 9310 0 9366 160 6 N2END[3]
port 230 nsew signal input
rlabel metal2 s 9586 0 9642 160 6 N2END[4]
port 231 nsew signal input
rlabel metal2 s 9862 0 9918 160 6 N2END[5]
port 232 nsew signal input
rlabel metal2 s 10138 0 10194 160 6 N2END[6]
port 233 nsew signal input
rlabel metal2 s 10414 0 10470 160 6 N2END[7]
port 234 nsew signal input
rlabel metal2 s 6274 0 6330 160 6 N2MID[0]
port 235 nsew signal input
rlabel metal2 s 6550 0 6606 160 6 N2MID[1]
port 236 nsew signal input
rlabel metal2 s 6826 0 6882 160 6 N2MID[2]
port 237 nsew signal input
rlabel metal2 s 7102 0 7158 160 6 N2MID[3]
port 238 nsew signal input
rlabel metal2 s 7378 0 7434 160 6 N2MID[4]
port 239 nsew signal input
rlabel metal2 s 7654 0 7710 160 6 N2MID[5]
port 240 nsew signal input
rlabel metal2 s 7930 0 7986 160 6 N2MID[6]
port 241 nsew signal input
rlabel metal2 s 8206 0 8262 160 6 N2MID[7]
port 242 nsew signal input
rlabel metal2 s 10690 44840 10746 45000 6 N4BEG[0]
port 243 nsew signal output
rlabel metal2 s 13450 44840 13506 45000 6 N4BEG[10]
port 244 nsew signal output
rlabel metal2 s 13726 44840 13782 45000 6 N4BEG[11]
port 245 nsew signal output
rlabel metal2 s 14002 44840 14058 45000 6 N4BEG[12]
port 246 nsew signal output
rlabel metal2 s 14278 44840 14334 45000 6 N4BEG[13]
port 247 nsew signal output
rlabel metal2 s 14554 44840 14610 45000 6 N4BEG[14]
port 248 nsew signal output
rlabel metal2 s 14830 44840 14886 45000 6 N4BEG[15]
port 249 nsew signal output
rlabel metal2 s 10966 44840 11022 45000 6 N4BEG[1]
port 250 nsew signal output
rlabel metal2 s 11242 44840 11298 45000 6 N4BEG[2]
port 251 nsew signal output
rlabel metal2 s 11518 44840 11574 45000 6 N4BEG[3]
port 252 nsew signal output
rlabel metal2 s 11794 44840 11850 45000 6 N4BEG[4]
port 253 nsew signal output
rlabel metal2 s 12070 44840 12126 45000 6 N4BEG[5]
port 254 nsew signal output
rlabel metal2 s 12346 44840 12402 45000 6 N4BEG[6]
port 255 nsew signal output
rlabel metal2 s 12622 44840 12678 45000 6 N4BEG[7]
port 256 nsew signal output
rlabel metal2 s 12898 44840 12954 45000 6 N4BEG[8]
port 257 nsew signal output
rlabel metal2 s 13174 44840 13230 45000 6 N4BEG[9]
port 258 nsew signal output
rlabel metal2 s 10690 0 10746 160 6 N4END[0]
port 259 nsew signal input
rlabel metal2 s 13450 0 13506 160 6 N4END[10]
port 260 nsew signal input
rlabel metal2 s 13726 0 13782 160 6 N4END[11]
port 261 nsew signal input
rlabel metal2 s 14002 0 14058 160 6 N4END[12]
port 262 nsew signal input
rlabel metal2 s 14278 0 14334 160 6 N4END[13]
port 263 nsew signal input
rlabel metal2 s 14554 0 14610 160 6 N4END[14]
port 264 nsew signal input
rlabel metal2 s 14830 0 14886 160 6 N4END[15]
port 265 nsew signal input
rlabel metal2 s 10966 0 11022 160 6 N4END[1]
port 266 nsew signal input
rlabel metal2 s 11242 0 11298 160 6 N4END[2]
port 267 nsew signal input
rlabel metal2 s 11518 0 11574 160 6 N4END[3]
port 268 nsew signal input
rlabel metal2 s 11794 0 11850 160 6 N4END[4]
port 269 nsew signal input
rlabel metal2 s 12070 0 12126 160 6 N4END[5]
port 270 nsew signal input
rlabel metal2 s 12346 0 12402 160 6 N4END[6]
port 271 nsew signal input
rlabel metal2 s 12622 0 12678 160 6 N4END[7]
port 272 nsew signal input
rlabel metal2 s 12898 0 12954 160 6 N4END[8]
port 273 nsew signal input
rlabel metal2 s 13174 0 13230 160 6 N4END[9]
port 274 nsew signal input
rlabel metal2 s 15106 44840 15162 45000 6 NN4BEG[0]
port 275 nsew signal output
rlabel metal2 s 17866 44840 17922 45000 6 NN4BEG[10]
port 276 nsew signal output
rlabel metal2 s 18142 44840 18198 45000 6 NN4BEG[11]
port 277 nsew signal output
rlabel metal2 s 18418 44840 18474 45000 6 NN4BEG[12]
port 278 nsew signal output
rlabel metal2 s 18694 44840 18750 45000 6 NN4BEG[13]
port 279 nsew signal output
rlabel metal2 s 18970 44840 19026 45000 6 NN4BEG[14]
port 280 nsew signal output
rlabel metal2 s 19246 44840 19302 45000 6 NN4BEG[15]
port 281 nsew signal output
rlabel metal2 s 15382 44840 15438 45000 6 NN4BEG[1]
port 282 nsew signal output
rlabel metal2 s 15658 44840 15714 45000 6 NN4BEG[2]
port 283 nsew signal output
rlabel metal2 s 15934 44840 15990 45000 6 NN4BEG[3]
port 284 nsew signal output
rlabel metal2 s 16210 44840 16266 45000 6 NN4BEG[4]
port 285 nsew signal output
rlabel metal2 s 16486 44840 16542 45000 6 NN4BEG[5]
port 286 nsew signal output
rlabel metal2 s 16762 44840 16818 45000 6 NN4BEG[6]
port 287 nsew signal output
rlabel metal2 s 17038 44840 17094 45000 6 NN4BEG[7]
port 288 nsew signal output
rlabel metal2 s 17314 44840 17370 45000 6 NN4BEG[8]
port 289 nsew signal output
rlabel metal2 s 17590 44840 17646 45000 6 NN4BEG[9]
port 290 nsew signal output
rlabel metal2 s 15106 0 15162 160 6 NN4END[0]
port 291 nsew signal input
rlabel metal2 s 17866 0 17922 160 6 NN4END[10]
port 292 nsew signal input
rlabel metal2 s 18142 0 18198 160 6 NN4END[11]
port 293 nsew signal input
rlabel metal2 s 18418 0 18474 160 6 NN4END[12]
port 294 nsew signal input
rlabel metal2 s 18694 0 18750 160 6 NN4END[13]
port 295 nsew signal input
rlabel metal2 s 18970 0 19026 160 6 NN4END[14]
port 296 nsew signal input
rlabel metal2 s 19246 0 19302 160 6 NN4END[15]
port 297 nsew signal input
rlabel metal2 s 15382 0 15438 160 6 NN4END[1]
port 298 nsew signal input
rlabel metal2 s 15658 0 15714 160 6 NN4END[2]
port 299 nsew signal input
rlabel metal2 s 15934 0 15990 160 6 NN4END[3]
port 300 nsew signal input
rlabel metal2 s 16210 0 16266 160 6 NN4END[4]
port 301 nsew signal input
rlabel metal2 s 16486 0 16542 160 6 NN4END[5]
port 302 nsew signal input
rlabel metal2 s 16762 0 16818 160 6 NN4END[6]
port 303 nsew signal input
rlabel metal2 s 17038 0 17094 160 6 NN4END[7]
port 304 nsew signal input
rlabel metal2 s 17314 0 17370 160 6 NN4END[8]
port 305 nsew signal input
rlabel metal2 s 17590 0 17646 160 6 NN4END[9]
port 306 nsew signal input
rlabel metal2 s 19522 0 19578 160 6 S1BEG[0]
port 307 nsew signal output
rlabel metal2 s 19798 0 19854 160 6 S1BEG[1]
port 308 nsew signal output
rlabel metal2 s 20074 0 20130 160 6 S1BEG[2]
port 309 nsew signal output
rlabel metal2 s 20350 0 20406 160 6 S1BEG[3]
port 310 nsew signal output
rlabel metal2 s 19522 44840 19578 45000 6 S1END[0]
port 311 nsew signal input
rlabel metal2 s 19798 44840 19854 45000 6 S1END[1]
port 312 nsew signal input
rlabel metal2 s 20074 44840 20130 45000 6 S1END[2]
port 313 nsew signal input
rlabel metal2 s 20350 44840 20406 45000 6 S1END[3]
port 314 nsew signal input
rlabel metal2 s 22834 0 22890 160 6 S2BEG[0]
port 315 nsew signal output
rlabel metal2 s 23110 0 23166 160 6 S2BEG[1]
port 316 nsew signal output
rlabel metal2 s 23386 0 23442 160 6 S2BEG[2]
port 317 nsew signal output
rlabel metal2 s 23662 0 23718 160 6 S2BEG[3]
port 318 nsew signal output
rlabel metal2 s 23938 0 23994 160 6 S2BEG[4]
port 319 nsew signal output
rlabel metal2 s 24214 0 24270 160 6 S2BEG[5]
port 320 nsew signal output
rlabel metal2 s 24490 0 24546 160 6 S2BEG[6]
port 321 nsew signal output
rlabel metal2 s 24766 0 24822 160 6 S2BEG[7]
port 322 nsew signal output
rlabel metal2 s 20626 0 20682 160 6 S2BEGb[0]
port 323 nsew signal output
rlabel metal2 s 20902 0 20958 160 6 S2BEGb[1]
port 324 nsew signal output
rlabel metal2 s 21178 0 21234 160 6 S2BEGb[2]
port 325 nsew signal output
rlabel metal2 s 21454 0 21510 160 6 S2BEGb[3]
port 326 nsew signal output
rlabel metal2 s 21730 0 21786 160 6 S2BEGb[4]
port 327 nsew signal output
rlabel metal2 s 22006 0 22062 160 6 S2BEGb[5]
port 328 nsew signal output
rlabel metal2 s 22282 0 22338 160 6 S2BEGb[6]
port 329 nsew signal output
rlabel metal2 s 22558 0 22614 160 6 S2BEGb[7]
port 330 nsew signal output
rlabel metal2 s 20626 44840 20682 45000 6 S2END[0]
port 331 nsew signal input
rlabel metal2 s 20902 44840 20958 45000 6 S2END[1]
port 332 nsew signal input
rlabel metal2 s 21178 44840 21234 45000 6 S2END[2]
port 333 nsew signal input
rlabel metal2 s 21454 44840 21510 45000 6 S2END[3]
port 334 nsew signal input
rlabel metal2 s 21730 44840 21786 45000 6 S2END[4]
port 335 nsew signal input
rlabel metal2 s 22006 44840 22062 45000 6 S2END[5]
port 336 nsew signal input
rlabel metal2 s 22282 44840 22338 45000 6 S2END[6]
port 337 nsew signal input
rlabel metal2 s 22558 44840 22614 45000 6 S2END[7]
port 338 nsew signal input
rlabel metal2 s 22834 44840 22890 45000 6 S2MID[0]
port 339 nsew signal input
rlabel metal2 s 23110 44840 23166 45000 6 S2MID[1]
port 340 nsew signal input
rlabel metal2 s 23386 44840 23442 45000 6 S2MID[2]
port 341 nsew signal input
rlabel metal2 s 23662 44840 23718 45000 6 S2MID[3]
port 342 nsew signal input
rlabel metal2 s 23938 44840 23994 45000 6 S2MID[4]
port 343 nsew signal input
rlabel metal2 s 24214 44840 24270 45000 6 S2MID[5]
port 344 nsew signal input
rlabel metal2 s 24490 44840 24546 45000 6 S2MID[6]
port 345 nsew signal input
rlabel metal2 s 24766 44840 24822 45000 6 S2MID[7]
port 346 nsew signal input
rlabel metal2 s 25042 0 25098 160 6 S4BEG[0]
port 347 nsew signal output
rlabel metal2 s 27802 0 27858 160 6 S4BEG[10]
port 348 nsew signal output
rlabel metal2 s 28078 0 28134 160 6 S4BEG[11]
port 349 nsew signal output
rlabel metal2 s 28354 0 28410 160 6 S4BEG[12]
port 350 nsew signal output
rlabel metal2 s 28630 0 28686 160 6 S4BEG[13]
port 351 nsew signal output
rlabel metal2 s 28906 0 28962 160 6 S4BEG[14]
port 352 nsew signal output
rlabel metal2 s 29182 0 29238 160 6 S4BEG[15]
port 353 nsew signal output
rlabel metal2 s 25318 0 25374 160 6 S4BEG[1]
port 354 nsew signal output
rlabel metal2 s 25594 0 25650 160 6 S4BEG[2]
port 355 nsew signal output
rlabel metal2 s 25870 0 25926 160 6 S4BEG[3]
port 356 nsew signal output
rlabel metal2 s 26146 0 26202 160 6 S4BEG[4]
port 357 nsew signal output
rlabel metal2 s 26422 0 26478 160 6 S4BEG[5]
port 358 nsew signal output
rlabel metal2 s 26698 0 26754 160 6 S4BEG[6]
port 359 nsew signal output
rlabel metal2 s 26974 0 27030 160 6 S4BEG[7]
port 360 nsew signal output
rlabel metal2 s 27250 0 27306 160 6 S4BEG[8]
port 361 nsew signal output
rlabel metal2 s 27526 0 27582 160 6 S4BEG[9]
port 362 nsew signal output
rlabel metal2 s 25042 44840 25098 45000 6 S4END[0]
port 363 nsew signal input
rlabel metal2 s 27802 44840 27858 45000 6 S4END[10]
port 364 nsew signal input
rlabel metal2 s 28078 44840 28134 45000 6 S4END[11]
port 365 nsew signal input
rlabel metal2 s 28354 44840 28410 45000 6 S4END[12]
port 366 nsew signal input
rlabel metal2 s 28630 44840 28686 45000 6 S4END[13]
port 367 nsew signal input
rlabel metal2 s 28906 44840 28962 45000 6 S4END[14]
port 368 nsew signal input
rlabel metal2 s 29182 44840 29238 45000 6 S4END[15]
port 369 nsew signal input
rlabel metal2 s 25318 44840 25374 45000 6 S4END[1]
port 370 nsew signal input
rlabel metal2 s 25594 44840 25650 45000 6 S4END[2]
port 371 nsew signal input
rlabel metal2 s 25870 44840 25926 45000 6 S4END[3]
port 372 nsew signal input
rlabel metal2 s 26146 44840 26202 45000 6 S4END[4]
port 373 nsew signal input
rlabel metal2 s 26422 44840 26478 45000 6 S4END[5]
port 374 nsew signal input
rlabel metal2 s 26698 44840 26754 45000 6 S4END[6]
port 375 nsew signal input
rlabel metal2 s 26974 44840 27030 45000 6 S4END[7]
port 376 nsew signal input
rlabel metal2 s 27250 44840 27306 45000 6 S4END[8]
port 377 nsew signal input
rlabel metal2 s 27526 44840 27582 45000 6 S4END[9]
port 378 nsew signal input
rlabel metal2 s 29458 0 29514 160 6 SS4BEG[0]
port 379 nsew signal output
rlabel metal2 s 32218 0 32274 160 6 SS4BEG[10]
port 380 nsew signal output
rlabel metal2 s 32494 0 32550 160 6 SS4BEG[11]
port 381 nsew signal output
rlabel metal2 s 32770 0 32826 160 6 SS4BEG[12]
port 382 nsew signal output
rlabel metal2 s 33046 0 33102 160 6 SS4BEG[13]
port 383 nsew signal output
rlabel metal2 s 33322 0 33378 160 6 SS4BEG[14]
port 384 nsew signal output
rlabel metal2 s 33598 0 33654 160 6 SS4BEG[15]
port 385 nsew signal output
rlabel metal2 s 29734 0 29790 160 6 SS4BEG[1]
port 386 nsew signal output
rlabel metal2 s 30010 0 30066 160 6 SS4BEG[2]
port 387 nsew signal output
rlabel metal2 s 30286 0 30342 160 6 SS4BEG[3]
port 388 nsew signal output
rlabel metal2 s 30562 0 30618 160 6 SS4BEG[4]
port 389 nsew signal output
rlabel metal2 s 30838 0 30894 160 6 SS4BEG[5]
port 390 nsew signal output
rlabel metal2 s 31114 0 31170 160 6 SS4BEG[6]
port 391 nsew signal output
rlabel metal2 s 31390 0 31446 160 6 SS4BEG[7]
port 392 nsew signal output
rlabel metal2 s 31666 0 31722 160 6 SS4BEG[8]
port 393 nsew signal output
rlabel metal2 s 31942 0 31998 160 6 SS4BEG[9]
port 394 nsew signal output
rlabel metal2 s 29458 44840 29514 45000 6 SS4END[0]
port 395 nsew signal input
rlabel metal2 s 32218 44840 32274 45000 6 SS4END[10]
port 396 nsew signal input
rlabel metal2 s 32494 44840 32550 45000 6 SS4END[11]
port 397 nsew signal input
rlabel metal2 s 32770 44840 32826 45000 6 SS4END[12]
port 398 nsew signal input
rlabel metal2 s 33046 44840 33102 45000 6 SS4END[13]
port 399 nsew signal input
rlabel metal2 s 33322 44840 33378 45000 6 SS4END[14]
port 400 nsew signal input
rlabel metal2 s 33598 44840 33654 45000 6 SS4END[15]
port 401 nsew signal input
rlabel metal2 s 29734 44840 29790 45000 6 SS4END[1]
port 402 nsew signal input
rlabel metal2 s 30010 44840 30066 45000 6 SS4END[2]
port 403 nsew signal input
rlabel metal2 s 30286 44840 30342 45000 6 SS4END[3]
port 404 nsew signal input
rlabel metal2 s 30562 44840 30618 45000 6 SS4END[4]
port 405 nsew signal input
rlabel metal2 s 30838 44840 30894 45000 6 SS4END[5]
port 406 nsew signal input
rlabel metal2 s 31114 44840 31170 45000 6 SS4END[6]
port 407 nsew signal input
rlabel metal2 s 31390 44840 31446 45000 6 SS4END[7]
port 408 nsew signal input
rlabel metal2 s 31666 44840 31722 45000 6 SS4END[8]
port 409 nsew signal input
rlabel metal2 s 31942 44840 31998 45000 6 SS4END[9]
port 410 nsew signal input
rlabel metal2 s 33874 0 33930 160 6 UserCLK
port 411 nsew signal input
rlabel metal2 s 33874 44840 33930 45000 6 UserCLKo
port 412 nsew signal output
rlabel metal3 s 0 5176 160 5296 6 W1BEG[0]
port 413 nsew signal output
rlabel metal3 s 0 5448 160 5568 6 W1BEG[1]
port 414 nsew signal output
rlabel metal3 s 0 5720 160 5840 6 W1BEG[2]
port 415 nsew signal output
rlabel metal3 s 0 5992 160 6112 6 W1BEG[3]
port 416 nsew signal output
rlabel metal3 s 44840 5176 45000 5296 6 W1END[0]
port 417 nsew signal input
rlabel metal3 s 44840 5448 45000 5568 6 W1END[1]
port 418 nsew signal input
rlabel metal3 s 44840 5720 45000 5840 6 W1END[2]
port 419 nsew signal input
rlabel metal3 s 44840 5992 45000 6112 6 W1END[3]
port 420 nsew signal input
rlabel metal3 s 0 6264 160 6384 6 W2BEG[0]
port 421 nsew signal output
rlabel metal3 s 0 6536 160 6656 6 W2BEG[1]
port 422 nsew signal output
rlabel metal3 s 0 6808 160 6928 6 W2BEG[2]
port 423 nsew signal output
rlabel metal3 s 0 7080 160 7200 6 W2BEG[3]
port 424 nsew signal output
rlabel metal3 s 0 7352 160 7472 6 W2BEG[4]
port 425 nsew signal output
rlabel metal3 s 0 7624 160 7744 6 W2BEG[5]
port 426 nsew signal output
rlabel metal3 s 0 7896 160 8016 6 W2BEG[6]
port 427 nsew signal output
rlabel metal3 s 0 8168 160 8288 6 W2BEG[7]
port 428 nsew signal output
rlabel metal3 s 0 8440 160 8560 6 W2BEGb[0]
port 429 nsew signal output
rlabel metal3 s 0 8712 160 8832 6 W2BEGb[1]
port 430 nsew signal output
rlabel metal3 s 0 8984 160 9104 6 W2BEGb[2]
port 431 nsew signal output
rlabel metal3 s 0 9256 160 9376 6 W2BEGb[3]
port 432 nsew signal output
rlabel metal3 s 0 9528 160 9648 6 W2BEGb[4]
port 433 nsew signal output
rlabel metal3 s 0 9800 160 9920 6 W2BEGb[5]
port 434 nsew signal output
rlabel metal3 s 0 10072 160 10192 6 W2BEGb[6]
port 435 nsew signal output
rlabel metal3 s 0 10344 160 10464 6 W2BEGb[7]
port 436 nsew signal output
rlabel metal3 s 44840 8440 45000 8560 6 W2END[0]
port 437 nsew signal input
rlabel metal3 s 44840 8712 45000 8832 6 W2END[1]
port 438 nsew signal input
rlabel metal3 s 44840 8984 45000 9104 6 W2END[2]
port 439 nsew signal input
rlabel metal3 s 44840 9256 45000 9376 6 W2END[3]
port 440 nsew signal input
rlabel metal3 s 44840 9528 45000 9648 6 W2END[4]
port 441 nsew signal input
rlabel metal3 s 44840 9800 45000 9920 6 W2END[5]
port 442 nsew signal input
rlabel metal3 s 44840 10072 45000 10192 6 W2END[6]
port 443 nsew signal input
rlabel metal3 s 44840 10344 45000 10464 6 W2END[7]
port 444 nsew signal input
rlabel metal3 s 44840 6264 45000 6384 6 W2MID[0]
port 445 nsew signal input
rlabel metal3 s 44840 6536 45000 6656 6 W2MID[1]
port 446 nsew signal input
rlabel metal3 s 44840 6808 45000 6928 6 W2MID[2]
port 447 nsew signal input
rlabel metal3 s 44840 7080 45000 7200 6 W2MID[3]
port 448 nsew signal input
rlabel metal3 s 44840 7352 45000 7472 6 W2MID[4]
port 449 nsew signal input
rlabel metal3 s 44840 7624 45000 7744 6 W2MID[5]
port 450 nsew signal input
rlabel metal3 s 44840 7896 45000 8016 6 W2MID[6]
port 451 nsew signal input
rlabel metal3 s 44840 8168 45000 8288 6 W2MID[7]
port 452 nsew signal input
rlabel metal3 s 0 14968 160 15088 6 W6BEG[0]
port 453 nsew signal output
rlabel metal3 s 0 17688 160 17808 6 W6BEG[10]
port 454 nsew signal output
rlabel metal3 s 0 17960 160 18080 6 W6BEG[11]
port 455 nsew signal output
rlabel metal3 s 0 15240 160 15360 6 W6BEG[1]
port 456 nsew signal output
rlabel metal3 s 0 15512 160 15632 6 W6BEG[2]
port 457 nsew signal output
rlabel metal3 s 0 15784 160 15904 6 W6BEG[3]
port 458 nsew signal output
rlabel metal3 s 0 16056 160 16176 6 W6BEG[4]
port 459 nsew signal output
rlabel metal3 s 0 16328 160 16448 6 W6BEG[5]
port 460 nsew signal output
rlabel metal3 s 0 16600 160 16720 6 W6BEG[6]
port 461 nsew signal output
rlabel metal3 s 0 16872 160 16992 6 W6BEG[7]
port 462 nsew signal output
rlabel metal3 s 0 17144 160 17264 6 W6BEG[8]
port 463 nsew signal output
rlabel metal3 s 0 17416 160 17536 6 W6BEG[9]
port 464 nsew signal output
rlabel metal3 s 44840 14968 45000 15088 6 W6END[0]
port 465 nsew signal input
rlabel metal3 s 44840 17688 45000 17808 6 W6END[10]
port 466 nsew signal input
rlabel metal3 s 44840 17960 45000 18080 6 W6END[11]
port 467 nsew signal input
rlabel metal3 s 44840 15240 45000 15360 6 W6END[1]
port 468 nsew signal input
rlabel metal3 s 44840 15512 45000 15632 6 W6END[2]
port 469 nsew signal input
rlabel metal3 s 44840 15784 45000 15904 6 W6END[3]
port 470 nsew signal input
rlabel metal3 s 44840 16056 45000 16176 6 W6END[4]
port 471 nsew signal input
rlabel metal3 s 44840 16328 45000 16448 6 W6END[5]
port 472 nsew signal input
rlabel metal3 s 44840 16600 45000 16720 6 W6END[6]
port 473 nsew signal input
rlabel metal3 s 44840 16872 45000 16992 6 W6END[7]
port 474 nsew signal input
rlabel metal3 s 44840 17144 45000 17264 6 W6END[8]
port 475 nsew signal input
rlabel metal3 s 44840 17416 45000 17536 6 W6END[9]
port 476 nsew signal input
rlabel metal3 s 0 10616 160 10736 6 WW4BEG[0]
port 477 nsew signal output
rlabel metal3 s 0 13336 160 13456 6 WW4BEG[10]
port 478 nsew signal output
rlabel metal3 s 0 13608 160 13728 6 WW4BEG[11]
port 479 nsew signal output
rlabel metal3 s 0 13880 160 14000 6 WW4BEG[12]
port 480 nsew signal output
rlabel metal3 s 0 14152 160 14272 6 WW4BEG[13]
port 481 nsew signal output
rlabel metal3 s 0 14424 160 14544 6 WW4BEG[14]
port 482 nsew signal output
rlabel metal3 s 0 14696 160 14816 6 WW4BEG[15]
port 483 nsew signal output
rlabel metal3 s 0 10888 160 11008 6 WW4BEG[1]
port 484 nsew signal output
rlabel metal3 s 0 11160 160 11280 6 WW4BEG[2]
port 485 nsew signal output
rlabel metal3 s 0 11432 160 11552 6 WW4BEG[3]
port 486 nsew signal output
rlabel metal3 s 0 11704 160 11824 6 WW4BEG[4]
port 487 nsew signal output
rlabel metal3 s 0 11976 160 12096 6 WW4BEG[5]
port 488 nsew signal output
rlabel metal3 s 0 12248 160 12368 6 WW4BEG[6]
port 489 nsew signal output
rlabel metal3 s 0 12520 160 12640 6 WW4BEG[7]
port 490 nsew signal output
rlabel metal3 s 0 12792 160 12912 6 WW4BEG[8]
port 491 nsew signal output
rlabel metal3 s 0 13064 160 13184 6 WW4BEG[9]
port 492 nsew signal output
rlabel metal3 s 44840 10616 45000 10736 6 WW4END[0]
port 493 nsew signal input
rlabel metal3 s 44840 13336 45000 13456 6 WW4END[10]
port 494 nsew signal input
rlabel metal3 s 44840 13608 45000 13728 6 WW4END[11]
port 495 nsew signal input
rlabel metal3 s 44840 13880 45000 14000 6 WW4END[12]
port 496 nsew signal input
rlabel metal3 s 44840 14152 45000 14272 6 WW4END[13]
port 497 nsew signal input
rlabel metal3 s 44840 14424 45000 14544 6 WW4END[14]
port 498 nsew signal input
rlabel metal3 s 44840 14696 45000 14816 6 WW4END[15]
port 499 nsew signal input
rlabel metal3 s 44840 10888 45000 11008 6 WW4END[1]
port 500 nsew signal input
rlabel metal3 s 44840 11160 45000 11280 6 WW4END[2]
port 501 nsew signal input
rlabel metal3 s 44840 11432 45000 11552 6 WW4END[3]
port 502 nsew signal input
rlabel metal3 s 44840 11704 45000 11824 6 WW4END[4]
port 503 nsew signal input
rlabel metal3 s 44840 11976 45000 12096 6 WW4END[5]
port 504 nsew signal input
rlabel metal3 s 44840 12248 45000 12368 6 WW4END[6]
port 505 nsew signal input
rlabel metal3 s 44840 12520 45000 12640 6 WW4END[7]
port 506 nsew signal input
rlabel metal3 s 44840 12792 45000 12912 6 WW4END[8]
port 507 nsew signal input
rlabel metal3 s 44840 13064 45000 13184 6 WW4END[9]
port 508 nsew signal input
rlabel metal4 s 3564 1040 3884 43568 6 vccd1
port 509 nsew power bidirectional
rlabel metal4 s 18564 1040 18884 43568 6 vccd1
port 509 nsew power bidirectional
rlabel metal4 s 33564 1040 33884 43568 6 vccd1
port 509 nsew power bidirectional
rlabel metal4 s 11064 1040 11384 43568 6 vssd1
port 510 nsew ground bidirectional
rlabel metal4 s 26064 1040 26384 43568 6 vssd1
port 510 nsew ground bidirectional
rlabel metal4 s 41064 1040 41384 43568 6 vssd1
port 510 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 45000 45000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9457560
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/LUT4AB/runs/24_12_04_15_33/results/signoff/LUT4AB.magic.gds
string GDS_START 221380
<< end >>

