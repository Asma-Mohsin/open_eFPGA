magic
tech sky130A
magscale 1 2
timestamp 1733308832
<< nwell >>
rect 1066 6789 43922 7355
rect 1066 5701 43922 6267
rect 1066 4613 43922 5179
rect 1066 3525 43922 4091
rect 1066 2437 43922 3003
<< obsli1 >>
rect 1104 2159 43884 7633
<< obsm1 >>
rect 1104 892 44040 7812
<< metal2 >>
rect 1306 9840 1362 10000
rect 3422 9840 3478 10000
rect 5538 9840 5594 10000
rect 7654 9840 7710 10000
rect 9770 9840 9826 10000
rect 11886 9840 11942 10000
rect 14002 9840 14058 10000
rect 16118 9840 16174 10000
rect 18234 9840 18290 10000
rect 20350 9840 20406 10000
rect 22466 9840 22522 10000
rect 24582 9840 24638 10000
rect 26698 9840 26754 10000
rect 28814 9840 28870 10000
rect 30930 9840 30986 10000
rect 33046 9840 33102 10000
rect 35162 9840 35218 10000
rect 37278 9840 37334 10000
rect 39394 9840 39450 10000
rect 41510 9840 41566 10000
rect 43626 9840 43682 10000
rect 5170 0 5226 160
rect 5446 0 5502 160
rect 5722 0 5778 160
rect 5998 0 6054 160
rect 6274 0 6330 160
rect 6550 0 6606 160
rect 6826 0 6882 160
rect 7102 0 7158 160
rect 7378 0 7434 160
rect 7654 0 7710 160
rect 7930 0 7986 160
rect 8206 0 8262 160
rect 8482 0 8538 160
rect 8758 0 8814 160
rect 9034 0 9090 160
rect 9310 0 9366 160
rect 9586 0 9642 160
rect 9862 0 9918 160
rect 10138 0 10194 160
rect 10414 0 10470 160
rect 10690 0 10746 160
rect 10966 0 11022 160
rect 11242 0 11298 160
rect 11518 0 11574 160
rect 11794 0 11850 160
rect 12070 0 12126 160
rect 12346 0 12402 160
rect 12622 0 12678 160
rect 12898 0 12954 160
rect 13174 0 13230 160
rect 13450 0 13506 160
rect 13726 0 13782 160
rect 14002 0 14058 160
rect 14278 0 14334 160
rect 14554 0 14610 160
rect 14830 0 14886 160
rect 15106 0 15162 160
rect 15382 0 15438 160
rect 15658 0 15714 160
rect 15934 0 15990 160
rect 16210 0 16266 160
rect 16486 0 16542 160
rect 16762 0 16818 160
rect 17038 0 17094 160
rect 17314 0 17370 160
rect 17590 0 17646 160
rect 17866 0 17922 160
rect 18142 0 18198 160
rect 18418 0 18474 160
rect 18694 0 18750 160
rect 18970 0 19026 160
rect 19246 0 19302 160
rect 19522 0 19578 160
rect 19798 0 19854 160
rect 20074 0 20130 160
rect 20350 0 20406 160
rect 20626 0 20682 160
rect 20902 0 20958 160
rect 21178 0 21234 160
rect 21454 0 21510 160
rect 21730 0 21786 160
rect 22006 0 22062 160
rect 22282 0 22338 160
rect 22558 0 22614 160
rect 22834 0 22890 160
rect 23110 0 23166 160
rect 23386 0 23442 160
rect 23662 0 23718 160
rect 23938 0 23994 160
rect 24214 0 24270 160
rect 24490 0 24546 160
rect 24766 0 24822 160
rect 25042 0 25098 160
rect 25318 0 25374 160
rect 25594 0 25650 160
rect 25870 0 25926 160
rect 26146 0 26202 160
rect 26422 0 26478 160
rect 26698 0 26754 160
rect 26974 0 27030 160
rect 27250 0 27306 160
rect 27526 0 27582 160
rect 27802 0 27858 160
rect 28078 0 28134 160
rect 28354 0 28410 160
rect 28630 0 28686 160
rect 28906 0 28962 160
rect 29182 0 29238 160
rect 29458 0 29514 160
rect 29734 0 29790 160
rect 30010 0 30066 160
rect 30286 0 30342 160
rect 30562 0 30618 160
rect 30838 0 30894 160
rect 31114 0 31170 160
rect 31390 0 31446 160
rect 31666 0 31722 160
rect 31942 0 31998 160
rect 32218 0 32274 160
rect 32494 0 32550 160
rect 32770 0 32826 160
rect 33046 0 33102 160
rect 33322 0 33378 160
rect 33598 0 33654 160
rect 33874 0 33930 160
rect 34150 0 34206 160
rect 34426 0 34482 160
rect 34702 0 34758 160
rect 34978 0 35034 160
rect 35254 0 35310 160
rect 35530 0 35586 160
rect 35806 0 35862 160
rect 36082 0 36138 160
rect 36358 0 36414 160
rect 36634 0 36690 160
rect 36910 0 36966 160
rect 37186 0 37242 160
rect 37462 0 37518 160
rect 37738 0 37794 160
rect 38014 0 38070 160
rect 38290 0 38346 160
rect 38566 0 38622 160
rect 38842 0 38898 160
rect 39118 0 39174 160
rect 39394 0 39450 160
rect 39670 0 39726 160
<< obsm2 >>
rect 1418 9784 3366 9874
rect 3534 9784 5482 9874
rect 5650 9784 7598 9874
rect 7766 9784 9714 9874
rect 9882 9784 11830 9874
rect 11998 9784 13946 9874
rect 14114 9784 16062 9874
rect 16230 9784 18178 9874
rect 18346 9784 20294 9874
rect 20462 9784 22410 9874
rect 22578 9784 24526 9874
rect 24694 9784 26642 9874
rect 26810 9784 28758 9874
rect 28926 9784 30874 9874
rect 31042 9784 32990 9874
rect 33158 9784 35106 9874
rect 35274 9784 37222 9874
rect 37390 9784 39338 9874
rect 39506 9784 41454 9874
rect 41622 9784 43570 9874
rect 43738 9784 44034 9874
rect 1308 216 44034 9784
rect 1308 54 5114 216
rect 5282 54 5390 216
rect 5558 54 5666 216
rect 5834 54 5942 216
rect 6110 54 6218 216
rect 6386 54 6494 216
rect 6662 54 6770 216
rect 6938 54 7046 216
rect 7214 54 7322 216
rect 7490 54 7598 216
rect 7766 54 7874 216
rect 8042 54 8150 216
rect 8318 54 8426 216
rect 8594 54 8702 216
rect 8870 54 8978 216
rect 9146 54 9254 216
rect 9422 54 9530 216
rect 9698 54 9806 216
rect 9974 54 10082 216
rect 10250 54 10358 216
rect 10526 54 10634 216
rect 10802 54 10910 216
rect 11078 54 11186 216
rect 11354 54 11462 216
rect 11630 54 11738 216
rect 11906 54 12014 216
rect 12182 54 12290 216
rect 12458 54 12566 216
rect 12734 54 12842 216
rect 13010 54 13118 216
rect 13286 54 13394 216
rect 13562 54 13670 216
rect 13838 54 13946 216
rect 14114 54 14222 216
rect 14390 54 14498 216
rect 14666 54 14774 216
rect 14942 54 15050 216
rect 15218 54 15326 216
rect 15494 54 15602 216
rect 15770 54 15878 216
rect 16046 54 16154 216
rect 16322 54 16430 216
rect 16598 54 16706 216
rect 16874 54 16982 216
rect 17150 54 17258 216
rect 17426 54 17534 216
rect 17702 54 17810 216
rect 17978 54 18086 216
rect 18254 54 18362 216
rect 18530 54 18638 216
rect 18806 54 18914 216
rect 19082 54 19190 216
rect 19358 54 19466 216
rect 19634 54 19742 216
rect 19910 54 20018 216
rect 20186 54 20294 216
rect 20462 54 20570 216
rect 20738 54 20846 216
rect 21014 54 21122 216
rect 21290 54 21398 216
rect 21566 54 21674 216
rect 21842 54 21950 216
rect 22118 54 22226 216
rect 22394 54 22502 216
rect 22670 54 22778 216
rect 22946 54 23054 216
rect 23222 54 23330 216
rect 23498 54 23606 216
rect 23774 54 23882 216
rect 24050 54 24158 216
rect 24326 54 24434 216
rect 24602 54 24710 216
rect 24878 54 24986 216
rect 25154 54 25262 216
rect 25430 54 25538 216
rect 25706 54 25814 216
rect 25982 54 26090 216
rect 26258 54 26366 216
rect 26534 54 26642 216
rect 26810 54 26918 216
rect 27086 54 27194 216
rect 27362 54 27470 216
rect 27638 54 27746 216
rect 27914 54 28022 216
rect 28190 54 28298 216
rect 28466 54 28574 216
rect 28742 54 28850 216
rect 29018 54 29126 216
rect 29294 54 29402 216
rect 29570 54 29678 216
rect 29846 54 29954 216
rect 30122 54 30230 216
rect 30398 54 30506 216
rect 30674 54 30782 216
rect 30950 54 31058 216
rect 31226 54 31334 216
rect 31502 54 31610 216
rect 31778 54 31886 216
rect 32054 54 32162 216
rect 32330 54 32438 216
rect 32606 54 32714 216
rect 32882 54 32990 216
rect 33158 54 33266 216
rect 33434 54 33542 216
rect 33710 54 33818 216
rect 33986 54 34094 216
rect 34262 54 34370 216
rect 34538 54 34646 216
rect 34814 54 34922 216
rect 35090 54 35198 216
rect 35366 54 35474 216
rect 35642 54 35750 216
rect 35918 54 36026 216
rect 36194 54 36302 216
rect 36470 54 36578 216
rect 36746 54 36854 216
rect 37022 54 37130 216
rect 37298 54 37406 216
rect 37574 54 37682 216
rect 37850 54 37958 216
rect 38126 54 38234 216
rect 38402 54 38510 216
rect 38678 54 38786 216
rect 38954 54 39062 216
rect 39230 54 39338 216
rect 39506 54 39614 216
rect 39782 54 44034 216
<< obsm3 >>
rect 6293 851 44038 7649
<< metal4 >>
rect 6291 2128 6611 7664
rect 11638 2128 11958 7664
rect 16985 2128 17305 7664
rect 22332 2128 22652 7664
rect 27679 2128 27999 7664
rect 33026 2128 33346 7664
rect 38373 2128 38693 7664
rect 43720 2128 44040 7664
<< obsm4 >>
rect 30235 2048 32946 5677
rect 33426 2048 36925 5677
rect 30235 851 36925 2048
<< labels >>
rlabel metal2 s 34150 0 34206 160 6 Ci
port 1 nsew signal input
rlabel metal2 s 34426 0 34482 160 6 FrameStrobe[0]
port 2 nsew signal input
rlabel metal2 s 37186 0 37242 160 6 FrameStrobe[10]
port 3 nsew signal input
rlabel metal2 s 37462 0 37518 160 6 FrameStrobe[11]
port 4 nsew signal input
rlabel metal2 s 37738 0 37794 160 6 FrameStrobe[12]
port 5 nsew signal input
rlabel metal2 s 38014 0 38070 160 6 FrameStrobe[13]
port 6 nsew signal input
rlabel metal2 s 38290 0 38346 160 6 FrameStrobe[14]
port 7 nsew signal input
rlabel metal2 s 38566 0 38622 160 6 FrameStrobe[15]
port 8 nsew signal input
rlabel metal2 s 38842 0 38898 160 6 FrameStrobe[16]
port 9 nsew signal input
rlabel metal2 s 39118 0 39174 160 6 FrameStrobe[17]
port 10 nsew signal input
rlabel metal2 s 39394 0 39450 160 6 FrameStrobe[18]
port 11 nsew signal input
rlabel metal2 s 39670 0 39726 160 6 FrameStrobe[19]
port 12 nsew signal input
rlabel metal2 s 34702 0 34758 160 6 FrameStrobe[1]
port 13 nsew signal input
rlabel metal2 s 34978 0 35034 160 6 FrameStrobe[2]
port 14 nsew signal input
rlabel metal2 s 35254 0 35310 160 6 FrameStrobe[3]
port 15 nsew signal input
rlabel metal2 s 35530 0 35586 160 6 FrameStrobe[4]
port 16 nsew signal input
rlabel metal2 s 35806 0 35862 160 6 FrameStrobe[5]
port 17 nsew signal input
rlabel metal2 s 36082 0 36138 160 6 FrameStrobe[6]
port 18 nsew signal input
rlabel metal2 s 36358 0 36414 160 6 FrameStrobe[7]
port 19 nsew signal input
rlabel metal2 s 36634 0 36690 160 6 FrameStrobe[8]
port 20 nsew signal input
rlabel metal2 s 36910 0 36966 160 6 FrameStrobe[9]
port 21 nsew signal input
rlabel metal2 s 3422 9840 3478 10000 6 FrameStrobe_O[0]
port 22 nsew signal output
rlabel metal2 s 24582 9840 24638 10000 6 FrameStrobe_O[10]
port 23 nsew signal output
rlabel metal2 s 26698 9840 26754 10000 6 FrameStrobe_O[11]
port 24 nsew signal output
rlabel metal2 s 28814 9840 28870 10000 6 FrameStrobe_O[12]
port 25 nsew signal output
rlabel metal2 s 30930 9840 30986 10000 6 FrameStrobe_O[13]
port 26 nsew signal output
rlabel metal2 s 33046 9840 33102 10000 6 FrameStrobe_O[14]
port 27 nsew signal output
rlabel metal2 s 35162 9840 35218 10000 6 FrameStrobe_O[15]
port 28 nsew signal output
rlabel metal2 s 37278 9840 37334 10000 6 FrameStrobe_O[16]
port 29 nsew signal output
rlabel metal2 s 39394 9840 39450 10000 6 FrameStrobe_O[17]
port 30 nsew signal output
rlabel metal2 s 41510 9840 41566 10000 6 FrameStrobe_O[18]
port 31 nsew signal output
rlabel metal2 s 43626 9840 43682 10000 6 FrameStrobe_O[19]
port 32 nsew signal output
rlabel metal2 s 5538 9840 5594 10000 6 FrameStrobe_O[1]
port 33 nsew signal output
rlabel metal2 s 7654 9840 7710 10000 6 FrameStrobe_O[2]
port 34 nsew signal output
rlabel metal2 s 9770 9840 9826 10000 6 FrameStrobe_O[3]
port 35 nsew signal output
rlabel metal2 s 11886 9840 11942 10000 6 FrameStrobe_O[4]
port 36 nsew signal output
rlabel metal2 s 14002 9840 14058 10000 6 FrameStrobe_O[5]
port 37 nsew signal output
rlabel metal2 s 16118 9840 16174 10000 6 FrameStrobe_O[6]
port 38 nsew signal output
rlabel metal2 s 18234 9840 18290 10000 6 FrameStrobe_O[7]
port 39 nsew signal output
rlabel metal2 s 20350 9840 20406 10000 6 FrameStrobe_O[8]
port 40 nsew signal output
rlabel metal2 s 22466 9840 22522 10000 6 FrameStrobe_O[9]
port 41 nsew signal output
rlabel metal2 s 5170 0 5226 160 6 N1END[0]
port 42 nsew signal input
rlabel metal2 s 5446 0 5502 160 6 N1END[1]
port 43 nsew signal input
rlabel metal2 s 5722 0 5778 160 6 N1END[2]
port 44 nsew signal input
rlabel metal2 s 5998 0 6054 160 6 N1END[3]
port 45 nsew signal input
rlabel metal2 s 8482 0 8538 160 6 N2END[0]
port 46 nsew signal input
rlabel metal2 s 8758 0 8814 160 6 N2END[1]
port 47 nsew signal input
rlabel metal2 s 9034 0 9090 160 6 N2END[2]
port 48 nsew signal input
rlabel metal2 s 9310 0 9366 160 6 N2END[3]
port 49 nsew signal input
rlabel metal2 s 9586 0 9642 160 6 N2END[4]
port 50 nsew signal input
rlabel metal2 s 9862 0 9918 160 6 N2END[5]
port 51 nsew signal input
rlabel metal2 s 10138 0 10194 160 6 N2END[6]
port 52 nsew signal input
rlabel metal2 s 10414 0 10470 160 6 N2END[7]
port 53 nsew signal input
rlabel metal2 s 6274 0 6330 160 6 N2MID[0]
port 54 nsew signal input
rlabel metal2 s 6550 0 6606 160 6 N2MID[1]
port 55 nsew signal input
rlabel metal2 s 6826 0 6882 160 6 N2MID[2]
port 56 nsew signal input
rlabel metal2 s 7102 0 7158 160 6 N2MID[3]
port 57 nsew signal input
rlabel metal2 s 7378 0 7434 160 6 N2MID[4]
port 58 nsew signal input
rlabel metal2 s 7654 0 7710 160 6 N2MID[5]
port 59 nsew signal input
rlabel metal2 s 7930 0 7986 160 6 N2MID[6]
port 60 nsew signal input
rlabel metal2 s 8206 0 8262 160 6 N2MID[7]
port 61 nsew signal input
rlabel metal2 s 10690 0 10746 160 6 N4END[0]
port 62 nsew signal input
rlabel metal2 s 13450 0 13506 160 6 N4END[10]
port 63 nsew signal input
rlabel metal2 s 13726 0 13782 160 6 N4END[11]
port 64 nsew signal input
rlabel metal2 s 14002 0 14058 160 6 N4END[12]
port 65 nsew signal input
rlabel metal2 s 14278 0 14334 160 6 N4END[13]
port 66 nsew signal input
rlabel metal2 s 14554 0 14610 160 6 N4END[14]
port 67 nsew signal input
rlabel metal2 s 14830 0 14886 160 6 N4END[15]
port 68 nsew signal input
rlabel metal2 s 10966 0 11022 160 6 N4END[1]
port 69 nsew signal input
rlabel metal2 s 11242 0 11298 160 6 N4END[2]
port 70 nsew signal input
rlabel metal2 s 11518 0 11574 160 6 N4END[3]
port 71 nsew signal input
rlabel metal2 s 11794 0 11850 160 6 N4END[4]
port 72 nsew signal input
rlabel metal2 s 12070 0 12126 160 6 N4END[5]
port 73 nsew signal input
rlabel metal2 s 12346 0 12402 160 6 N4END[6]
port 74 nsew signal input
rlabel metal2 s 12622 0 12678 160 6 N4END[7]
port 75 nsew signal input
rlabel metal2 s 12898 0 12954 160 6 N4END[8]
port 76 nsew signal input
rlabel metal2 s 13174 0 13230 160 6 N4END[9]
port 77 nsew signal input
rlabel metal2 s 15106 0 15162 160 6 NN4END[0]
port 78 nsew signal input
rlabel metal2 s 17866 0 17922 160 6 NN4END[10]
port 79 nsew signal input
rlabel metal2 s 18142 0 18198 160 6 NN4END[11]
port 80 nsew signal input
rlabel metal2 s 18418 0 18474 160 6 NN4END[12]
port 81 nsew signal input
rlabel metal2 s 18694 0 18750 160 6 NN4END[13]
port 82 nsew signal input
rlabel metal2 s 18970 0 19026 160 6 NN4END[14]
port 83 nsew signal input
rlabel metal2 s 19246 0 19302 160 6 NN4END[15]
port 84 nsew signal input
rlabel metal2 s 15382 0 15438 160 6 NN4END[1]
port 85 nsew signal input
rlabel metal2 s 15658 0 15714 160 6 NN4END[2]
port 86 nsew signal input
rlabel metal2 s 15934 0 15990 160 6 NN4END[3]
port 87 nsew signal input
rlabel metal2 s 16210 0 16266 160 6 NN4END[4]
port 88 nsew signal input
rlabel metal2 s 16486 0 16542 160 6 NN4END[5]
port 89 nsew signal input
rlabel metal2 s 16762 0 16818 160 6 NN4END[6]
port 90 nsew signal input
rlabel metal2 s 17038 0 17094 160 6 NN4END[7]
port 91 nsew signal input
rlabel metal2 s 17314 0 17370 160 6 NN4END[8]
port 92 nsew signal input
rlabel metal2 s 17590 0 17646 160 6 NN4END[9]
port 93 nsew signal input
rlabel metal2 s 19522 0 19578 160 6 S1BEG[0]
port 94 nsew signal output
rlabel metal2 s 19798 0 19854 160 6 S1BEG[1]
port 95 nsew signal output
rlabel metal2 s 20074 0 20130 160 6 S1BEG[2]
port 96 nsew signal output
rlabel metal2 s 20350 0 20406 160 6 S1BEG[3]
port 97 nsew signal output
rlabel metal2 s 22834 0 22890 160 6 S2BEG[0]
port 98 nsew signal output
rlabel metal2 s 23110 0 23166 160 6 S2BEG[1]
port 99 nsew signal output
rlabel metal2 s 23386 0 23442 160 6 S2BEG[2]
port 100 nsew signal output
rlabel metal2 s 23662 0 23718 160 6 S2BEG[3]
port 101 nsew signal output
rlabel metal2 s 23938 0 23994 160 6 S2BEG[4]
port 102 nsew signal output
rlabel metal2 s 24214 0 24270 160 6 S2BEG[5]
port 103 nsew signal output
rlabel metal2 s 24490 0 24546 160 6 S2BEG[6]
port 104 nsew signal output
rlabel metal2 s 24766 0 24822 160 6 S2BEG[7]
port 105 nsew signal output
rlabel metal2 s 20626 0 20682 160 6 S2BEGb[0]
port 106 nsew signal output
rlabel metal2 s 20902 0 20958 160 6 S2BEGb[1]
port 107 nsew signal output
rlabel metal2 s 21178 0 21234 160 6 S2BEGb[2]
port 108 nsew signal output
rlabel metal2 s 21454 0 21510 160 6 S2BEGb[3]
port 109 nsew signal output
rlabel metal2 s 21730 0 21786 160 6 S2BEGb[4]
port 110 nsew signal output
rlabel metal2 s 22006 0 22062 160 6 S2BEGb[5]
port 111 nsew signal output
rlabel metal2 s 22282 0 22338 160 6 S2BEGb[6]
port 112 nsew signal output
rlabel metal2 s 22558 0 22614 160 6 S2BEGb[7]
port 113 nsew signal output
rlabel metal2 s 25042 0 25098 160 6 S4BEG[0]
port 114 nsew signal output
rlabel metal2 s 27802 0 27858 160 6 S4BEG[10]
port 115 nsew signal output
rlabel metal2 s 28078 0 28134 160 6 S4BEG[11]
port 116 nsew signal output
rlabel metal2 s 28354 0 28410 160 6 S4BEG[12]
port 117 nsew signal output
rlabel metal2 s 28630 0 28686 160 6 S4BEG[13]
port 118 nsew signal output
rlabel metal2 s 28906 0 28962 160 6 S4BEG[14]
port 119 nsew signal output
rlabel metal2 s 29182 0 29238 160 6 S4BEG[15]
port 120 nsew signal output
rlabel metal2 s 25318 0 25374 160 6 S4BEG[1]
port 121 nsew signal output
rlabel metal2 s 25594 0 25650 160 6 S4BEG[2]
port 122 nsew signal output
rlabel metal2 s 25870 0 25926 160 6 S4BEG[3]
port 123 nsew signal output
rlabel metal2 s 26146 0 26202 160 6 S4BEG[4]
port 124 nsew signal output
rlabel metal2 s 26422 0 26478 160 6 S4BEG[5]
port 125 nsew signal output
rlabel metal2 s 26698 0 26754 160 6 S4BEG[6]
port 126 nsew signal output
rlabel metal2 s 26974 0 27030 160 6 S4BEG[7]
port 127 nsew signal output
rlabel metal2 s 27250 0 27306 160 6 S4BEG[8]
port 128 nsew signal output
rlabel metal2 s 27526 0 27582 160 6 S4BEG[9]
port 129 nsew signal output
rlabel metal2 s 29458 0 29514 160 6 SS4BEG[0]
port 130 nsew signal output
rlabel metal2 s 32218 0 32274 160 6 SS4BEG[10]
port 131 nsew signal output
rlabel metal2 s 32494 0 32550 160 6 SS4BEG[11]
port 132 nsew signal output
rlabel metal2 s 32770 0 32826 160 6 SS4BEG[12]
port 133 nsew signal output
rlabel metal2 s 33046 0 33102 160 6 SS4BEG[13]
port 134 nsew signal output
rlabel metal2 s 33322 0 33378 160 6 SS4BEG[14]
port 135 nsew signal output
rlabel metal2 s 33598 0 33654 160 6 SS4BEG[15]
port 136 nsew signal output
rlabel metal2 s 29734 0 29790 160 6 SS4BEG[1]
port 137 nsew signal output
rlabel metal2 s 30010 0 30066 160 6 SS4BEG[2]
port 138 nsew signal output
rlabel metal2 s 30286 0 30342 160 6 SS4BEG[3]
port 139 nsew signal output
rlabel metal2 s 30562 0 30618 160 6 SS4BEG[4]
port 140 nsew signal output
rlabel metal2 s 30838 0 30894 160 6 SS4BEG[5]
port 141 nsew signal output
rlabel metal2 s 31114 0 31170 160 6 SS4BEG[6]
port 142 nsew signal output
rlabel metal2 s 31390 0 31446 160 6 SS4BEG[7]
port 143 nsew signal output
rlabel metal2 s 31666 0 31722 160 6 SS4BEG[8]
port 144 nsew signal output
rlabel metal2 s 31942 0 31998 160 6 SS4BEG[9]
port 145 nsew signal output
rlabel metal2 s 33874 0 33930 160 6 UserCLK
port 146 nsew signal input
rlabel metal2 s 1306 9840 1362 10000 6 UserCLKo
port 147 nsew signal output
rlabel metal4 s 6291 2128 6611 7664 6 vccd1
port 148 nsew power bidirectional
rlabel metal4 s 16985 2128 17305 7664 6 vccd1
port 148 nsew power bidirectional
rlabel metal4 s 27679 2128 27999 7664 6 vccd1
port 148 nsew power bidirectional
rlabel metal4 s 38373 2128 38693 7664 6 vccd1
port 148 nsew power bidirectional
rlabel metal4 s 11638 2128 11958 7664 6 vssd1
port 149 nsew ground bidirectional
rlabel metal4 s 22332 2128 22652 7664 6 vssd1
port 149 nsew ground bidirectional
rlabel metal4 s 33026 2128 33346 7664 6 vssd1
port 149 nsew ground bidirectional
rlabel metal4 s 43720 2128 44040 7664 6 vssd1
port 149 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 45000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 507530
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/N_term_single/runs/24_12_04_10_39/results/signoff/N_term_single.magic.gds
string GDS_START 41474
<< end >>

