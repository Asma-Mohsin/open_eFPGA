magic
tech sky130A
magscale 1 2
timestamp 1733405999
<< viali >>
rect 1593 8585 1627 8619
rect 3985 8585 4019 8619
rect 5641 8585 5675 8619
rect 7941 8585 7975 8619
rect 10057 8585 10091 8619
rect 12173 8585 12207 8619
rect 14289 8585 14323 8619
rect 16405 8585 16439 8619
rect 18521 8585 18555 8619
rect 20637 8585 20671 8619
rect 22753 8585 22787 8619
rect 24685 8585 24719 8619
rect 27169 8585 27203 8619
rect 28917 8585 28951 8619
rect 31217 8585 31251 8619
rect 33149 8585 33183 8619
rect 35449 8585 35483 8619
rect 37473 8585 37507 8619
rect 40049 8585 40083 8619
rect 41797 8585 41831 8619
rect 43453 8585 43487 8619
rect 1501 8517 1535 8551
rect 3801 8449 3835 8483
rect 5181 8449 5215 8483
rect 5549 8449 5583 8483
rect 7757 8449 7791 8483
rect 9763 8449 9797 8483
rect 11989 8449 12023 8483
rect 14105 8449 14139 8483
rect 16221 8449 16255 8483
rect 18337 8449 18371 8483
rect 20453 8449 20487 8483
rect 22569 8449 22603 8483
rect 24593 8449 24627 8483
rect 26985 8449 27019 8483
rect 28825 8449 28859 8483
rect 31033 8449 31067 8483
rect 33057 8449 33091 8483
rect 35265 8449 35299 8483
rect 37381 8449 37415 8483
rect 39957 8449 39991 8483
rect 41705 8449 41739 8483
rect 43269 8449 43303 8483
rect 4445 8313 4479 8347
rect 9413 8313 9447 8347
rect 27537 3145 27571 3179
rect 19625 3009 19659 3043
rect 21925 3009 21959 3043
rect 27169 3009 27203 3043
rect 27445 3009 27479 3043
rect 27721 3009 27755 3043
rect 28273 3009 28307 3043
rect 28549 3009 28583 3043
rect 28825 3009 28859 3043
rect 29285 3009 29319 3043
rect 29561 3009 29595 3043
rect 22109 2873 22143 2907
rect 19441 2805 19475 2839
rect 26985 2805 27019 2839
rect 27261 2805 27295 2839
rect 28089 2805 28123 2839
rect 28365 2805 28399 2839
rect 28641 2805 28675 2839
rect 29101 2805 29135 2839
rect 29377 2805 29411 2839
rect 14105 2601 14139 2635
rect 16313 2601 16347 2635
rect 16497 2601 16531 2635
rect 18521 2601 18555 2635
rect 20545 2601 20579 2635
rect 20821 2601 20855 2635
rect 22937 2601 22971 2635
rect 24593 2601 24627 2635
rect 24961 2601 24995 2635
rect 25053 2601 25087 2635
rect 26617 2601 26651 2635
rect 27261 2601 27295 2635
rect 31401 2601 31435 2635
rect 33517 2601 33551 2635
rect 36369 2601 36403 2635
rect 37749 2601 37783 2635
rect 39497 2601 39531 2635
rect 40693 2601 40727 2635
rect 42257 2601 42291 2635
rect 17141 2533 17175 2567
rect 19441 2533 19475 2567
rect 20269 2533 20303 2567
rect 25329 2533 25363 2567
rect 25605 2533 25639 2567
rect 25881 2533 25915 2567
rect 14289 2397 14323 2431
rect 16129 2397 16163 2431
rect 16681 2397 16715 2431
rect 16957 2397 16991 2431
rect 18337 2397 18371 2431
rect 18797 2397 18831 2431
rect 18889 2397 18923 2431
rect 19625 2397 19659 2431
rect 19901 2397 19935 2431
rect 20177 2397 20211 2431
rect 20453 2397 20487 2431
rect 20729 2397 20763 2431
rect 21005 2397 21039 2431
rect 21281 2397 21315 2431
rect 21373 2397 21407 2431
rect 22109 2397 22143 2431
rect 22385 2397 22419 2431
rect 22661 2397 22695 2431
rect 23121 2397 23155 2431
rect 24409 2397 24443 2431
rect 24777 2397 24811 2431
rect 25237 2397 25271 2431
rect 25513 2397 25547 2431
rect 25789 2373 25823 2407
rect 26065 2397 26099 2431
rect 26341 2397 26375 2431
rect 26433 2397 26467 2431
rect 26893 2397 26927 2431
rect 27169 2397 27203 2431
rect 27445 2397 27479 2431
rect 27721 2397 27755 2431
rect 28181 2397 28215 2431
rect 28365 2397 28399 2431
rect 28733 2397 28767 2431
rect 29193 2397 29227 2431
rect 29745 2397 29779 2431
rect 30021 2397 30055 2431
rect 30297 2397 30331 2431
rect 30573 2397 30607 2431
rect 31577 2393 31611 2427
rect 31953 2397 31987 2431
rect 32873 2397 32907 2431
rect 33701 2397 33735 2431
rect 36553 2397 36587 2431
rect 37933 2397 37967 2431
rect 39681 2397 39715 2431
rect 40877 2397 40911 2431
rect 42441 2397 42475 2431
rect 18613 2261 18647 2295
rect 19073 2261 19107 2295
rect 19717 2261 19751 2295
rect 19993 2261 20027 2295
rect 21097 2261 21131 2295
rect 21557 2261 21591 2295
rect 21925 2261 21959 2295
rect 22201 2261 22235 2295
rect 22477 2261 22511 2295
rect 26157 2261 26191 2295
rect 26709 2261 26743 2295
rect 26985 2261 27019 2295
rect 27813 2261 27847 2295
rect 27997 2261 28031 2295
rect 28549 2261 28583 2295
rect 28917 2261 28951 2295
rect 29009 2261 29043 2295
rect 29561 2261 29595 2295
rect 29837 2261 29871 2295
rect 30113 2261 30147 2295
rect 30389 2261 30423 2295
rect 31769 2261 31803 2295
rect 33057 2261 33091 2295
rect 6745 2057 6779 2091
rect 14197 2057 14231 2091
rect 15393 2057 15427 2091
rect 15669 2057 15703 2091
rect 15945 2057 15979 2091
rect 16037 2057 16071 2091
rect 16497 2057 16531 2091
rect 16957 2057 16991 2091
rect 17233 2057 17267 2091
rect 17877 2057 17911 2091
rect 18153 2057 18187 2091
rect 18981 2057 19015 2091
rect 20637 2057 20671 2091
rect 23029 2057 23063 2091
rect 23857 2057 23891 2091
rect 24685 2057 24719 2091
rect 37289 2057 37323 2091
rect 37565 2057 37599 2091
rect 38117 2057 38151 2091
rect 38761 2057 38795 2091
rect 39957 2057 39991 2091
rect 20177 1989 20211 2023
rect 21281 1989 21315 2023
rect 25421 1989 25455 2023
rect 25973 1989 26007 2023
rect 27077 1989 27111 2023
rect 28181 1989 28215 2023
rect 28825 1989 28859 2023
rect 32229 1989 32263 2023
rect 32781 1989 32815 2023
rect 33333 1989 33367 2023
rect 34437 1989 34471 2023
rect 6561 1921 6595 1955
rect 13737 1921 13771 1955
rect 14381 1921 14415 1955
rect 15117 1921 15151 1955
rect 15209 1921 15243 1955
rect 15485 1921 15519 1955
rect 15761 1921 15795 1955
rect 16221 1921 16255 1955
rect 16313 1921 16347 1955
rect 16773 1921 16807 1955
rect 17049 1921 17083 1955
rect 17325 1921 17359 1955
rect 17601 1921 17635 1955
rect 18061 1921 18095 1955
rect 18337 1921 18371 1955
rect 18429 1921 18463 1955
rect 18705 1921 18739 1955
rect 19165 1921 19199 1955
rect 19441 1921 19475 1955
rect 19533 1921 19567 1955
rect 20821 1921 20855 1955
rect 21097 1921 21131 1955
rect 22109 1921 22143 1955
rect 22937 1921 22971 1955
rect 23213 1921 23247 1955
rect 23489 1921 23523 1955
rect 23765 1921 23799 1955
rect 24041 1921 24075 1955
rect 24317 1921 24351 1955
rect 24593 1921 24627 1955
rect 24869 1921 24903 1955
rect 25145 1921 25179 1955
rect 26801 1921 26835 1955
rect 27629 1921 27663 1955
rect 29285 1921 29319 1955
rect 29837 1921 29871 1955
rect 30297 1921 30331 1955
rect 30941 1921 30975 1955
rect 31493 1921 31527 1955
rect 33885 1921 33919 1955
rect 34897 1921 34931 1955
rect 36369 1921 36403 1955
rect 37473 1921 37507 1955
rect 37749 1921 37783 1955
rect 38301 1921 38335 1955
rect 38945 1921 38979 1955
rect 40141 1921 40175 1955
rect 41061 1921 41095 1955
rect 27353 1853 27387 1887
rect 17509 1785 17543 1819
rect 18613 1785 18647 1819
rect 22753 1785 22787 1819
rect 24961 1785 24995 1819
rect 28365 1785 28399 1819
rect 29009 1785 29043 1819
rect 36553 1785 36587 1819
rect 40877 1785 40911 1819
rect 13921 1717 13955 1751
rect 14933 1717 14967 1751
rect 17785 1717 17819 1751
rect 18889 1717 18923 1751
rect 19257 1717 19291 1751
rect 19717 1717 19751 1751
rect 20269 1717 20303 1751
rect 20913 1717 20947 1751
rect 21373 1717 21407 1751
rect 22201 1717 22235 1751
rect 23305 1717 23339 1751
rect 23581 1717 23615 1751
rect 24133 1717 24167 1751
rect 24409 1717 24443 1751
rect 25513 1717 25547 1751
rect 26249 1717 26283 1751
rect 26617 1717 26651 1751
rect 27721 1717 27755 1751
rect 29469 1717 29503 1751
rect 29929 1717 29963 1751
rect 30481 1717 30515 1751
rect 31033 1717 31067 1751
rect 31769 1717 31803 1751
rect 32321 1717 32355 1751
rect 32873 1717 32907 1751
rect 33425 1717 33459 1751
rect 33977 1717 34011 1751
rect 34529 1717 34563 1751
rect 35081 1717 35115 1751
rect 6837 1513 6871 1547
rect 7941 1513 7975 1547
rect 9413 1513 9447 1547
rect 10793 1513 10827 1547
rect 11989 1513 12023 1547
rect 12265 1513 12299 1547
rect 13921 1513 13955 1547
rect 14657 1513 14691 1547
rect 14933 1513 14967 1547
rect 15209 1513 15243 1547
rect 16037 1513 16071 1547
rect 16957 1513 16991 1547
rect 17233 1513 17267 1547
rect 17785 1513 17819 1547
rect 18613 1513 18647 1547
rect 23489 1513 23523 1547
rect 24961 1513 24995 1547
rect 25513 1513 25547 1547
rect 27169 1513 27203 1547
rect 28273 1513 28307 1547
rect 31401 1513 31435 1547
rect 32321 1513 32355 1547
rect 32873 1513 32907 1547
rect 33425 1513 33459 1547
rect 34897 1513 34931 1547
rect 39221 1513 39255 1547
rect 41245 1513 41279 1547
rect 41521 1513 41555 1547
rect 7389 1445 7423 1479
rect 9689 1445 9723 1479
rect 9965 1445 9999 1479
rect 10241 1445 10275 1479
rect 14381 1445 14415 1479
rect 15485 1445 15519 1479
rect 16313 1445 16347 1479
rect 17509 1445 17543 1479
rect 26709 1445 26743 1479
rect 30941 1445 30975 1479
rect 35909 1445 35943 1479
rect 37749 1445 37783 1479
rect 39865 1445 39899 1479
rect 40969 1445 41003 1479
rect 22201 1377 22235 1411
rect 30481 1377 30515 1411
rect 4905 1309 4939 1343
rect 5181 1309 5215 1343
rect 5457 1309 5491 1343
rect 5733 1309 5767 1343
rect 6009 1309 6043 1343
rect 6377 1309 6411 1343
rect 6653 1309 6687 1343
rect 6929 1309 6963 1343
rect 7205 1309 7239 1343
rect 7481 1309 7515 1343
rect 7757 1309 7791 1343
rect 8033 1309 8067 1343
rect 8309 1309 8343 1343
rect 8585 1309 8619 1343
rect 8953 1309 8987 1343
rect 9229 1309 9263 1343
rect 9505 1309 9539 1343
rect 9781 1309 9815 1343
rect 10057 1309 10091 1343
rect 10333 1309 10367 1343
rect 10609 1309 10643 1343
rect 10911 1309 10945 1343
rect 11161 1309 11195 1343
rect 11529 1309 11563 1343
rect 11805 1309 11839 1343
rect 12081 1309 12115 1343
rect 12357 1309 12391 1343
rect 12633 1309 12667 1343
rect 12909 1309 12943 1343
rect 13185 1309 13219 1343
rect 13461 1309 13495 1343
rect 13737 1309 13771 1343
rect 14105 1309 14139 1343
rect 14565 1309 14599 1343
rect 14841 1309 14875 1343
rect 15117 1309 15151 1343
rect 15393 1309 15427 1343
rect 15669 1309 15703 1343
rect 15945 1309 15979 1343
rect 16221 1309 16255 1343
rect 16497 1309 16531 1343
rect 16865 1309 16899 1343
rect 17141 1309 17175 1343
rect 17417 1309 17451 1343
rect 17693 1309 17727 1343
rect 17969 1309 18003 1343
rect 18245 1309 18279 1343
rect 18521 1309 18555 1343
rect 18797 1309 18831 1343
rect 19073 1309 19107 1343
rect 19257 1309 19291 1343
rect 19533 1309 19567 1343
rect 19901 1309 19935 1343
rect 20269 1309 20303 1343
rect 20729 1309 20763 1343
rect 21373 1309 21407 1343
rect 22569 1309 22603 1343
rect 22937 1309 22971 1343
rect 23397 1309 23431 1343
rect 23857 1309 23891 1343
rect 24409 1309 24443 1343
rect 25973 1309 26007 1343
rect 26525 1309 26559 1343
rect 27077 1309 27111 1343
rect 27611 1309 27645 1343
rect 28181 1309 28215 1343
rect 29377 1309 29411 1343
rect 30205 1309 30239 1343
rect 31953 1309 31987 1343
rect 33333 1309 33367 1343
rect 33885 1309 33919 1343
rect 34345 1309 34379 1343
rect 35725 1309 35759 1343
rect 36369 1309 36403 1343
rect 36461 1309 36495 1343
rect 36737 1309 36771 1343
rect 37473 1309 37507 1343
rect 37565 1309 37599 1343
rect 37841 1309 37875 1343
rect 38117 1309 38151 1343
rect 38393 1309 38427 1343
rect 38669 1309 38703 1343
rect 38945 1309 38979 1343
rect 39405 1309 39439 1343
rect 39497 1309 39531 1343
rect 40049 1309 40083 1343
rect 40325 1309 40359 1343
rect 40601 1309 40635 1343
rect 40877 1309 40911 1343
rect 41153 1309 41187 1343
rect 41429 1309 41463 1343
rect 41705 1309 41739 1343
rect 21925 1241 21959 1275
rect 24869 1241 24903 1275
rect 25421 1241 25455 1275
rect 29653 1241 29687 1275
rect 30757 1241 30791 1275
rect 31309 1241 31343 1275
rect 32229 1241 32263 1275
rect 32781 1241 32815 1275
rect 34805 1241 34839 1275
rect 5089 1173 5123 1207
rect 5365 1173 5399 1207
rect 5641 1173 5675 1207
rect 5917 1173 5951 1207
rect 6193 1173 6227 1207
rect 6561 1173 6595 1207
rect 7113 1173 7147 1207
rect 7665 1173 7699 1207
rect 8217 1173 8251 1207
rect 8493 1173 8527 1207
rect 8769 1173 8803 1207
rect 9137 1173 9171 1207
rect 10517 1173 10551 1207
rect 11069 1173 11103 1207
rect 11345 1173 11379 1207
rect 11713 1173 11747 1207
rect 12541 1173 12575 1207
rect 12817 1173 12851 1207
rect 13093 1173 13127 1207
rect 13369 1173 13403 1207
rect 13645 1173 13679 1207
rect 14289 1173 14323 1207
rect 15761 1173 15795 1207
rect 16681 1173 16715 1207
rect 18061 1173 18095 1207
rect 18337 1173 18371 1207
rect 18889 1173 18923 1207
rect 19441 1173 19475 1207
rect 19717 1173 19751 1207
rect 20085 1173 20119 1207
rect 20453 1173 20487 1207
rect 20821 1173 20855 1207
rect 21557 1173 21591 1207
rect 22753 1173 22787 1207
rect 23121 1173 23155 1207
rect 24041 1173 24075 1207
rect 24593 1173 24627 1207
rect 26065 1173 26099 1207
rect 27905 1173 27939 1207
rect 28825 1173 28859 1207
rect 29193 1173 29227 1207
rect 29745 1173 29779 1207
rect 31769 1173 31803 1207
rect 33977 1173 34011 1207
rect 34529 1173 34563 1207
rect 35449 1173 35483 1207
rect 36185 1173 36219 1207
rect 36645 1173 36679 1207
rect 36921 1173 36955 1207
rect 37289 1173 37323 1207
rect 38025 1173 38059 1207
rect 38301 1173 38335 1207
rect 38577 1173 38611 1207
rect 38853 1173 38887 1207
rect 39129 1173 39163 1207
rect 39681 1173 39715 1207
rect 40141 1173 40175 1207
rect 40417 1173 40451 1207
rect 40693 1173 40727 1207
<< metal1 >>
rect 13906 8780 13912 8832
rect 13964 8820 13970 8832
rect 23566 8820 23572 8832
rect 13964 8792 23572 8820
rect 13964 8780 13970 8792
rect 23566 8780 23572 8792
rect 23624 8780 23630 8832
rect 1104 8730 44040 8752
rect 1104 8678 11644 8730
rect 11696 8678 11708 8730
rect 11760 8678 11772 8730
rect 11824 8678 11836 8730
rect 11888 8678 11900 8730
rect 11952 8678 22338 8730
rect 22390 8678 22402 8730
rect 22454 8678 22466 8730
rect 22518 8678 22530 8730
rect 22582 8678 22594 8730
rect 22646 8678 33032 8730
rect 33084 8678 33096 8730
rect 33148 8678 33160 8730
rect 33212 8678 33224 8730
rect 33276 8678 33288 8730
rect 33340 8678 43726 8730
rect 43778 8678 43790 8730
rect 43842 8678 43854 8730
rect 43906 8678 43918 8730
rect 43970 8678 43982 8730
rect 44034 8678 44040 8730
rect 1104 8656 44040 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1452 8588 1593 8616
rect 1452 8576 1458 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 1581 8579 1639 8585
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3476 8588 3985 8616
rect 3476 8576 3482 8588
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 3973 8579 4031 8585
rect 5626 8576 5632 8628
rect 5684 8576 5690 8628
rect 7650 8576 7656 8628
rect 7708 8616 7714 8628
rect 7929 8619 7987 8625
rect 7929 8616 7941 8619
rect 7708 8588 7941 8616
rect 7708 8576 7714 8588
rect 7929 8585 7941 8588
rect 7975 8585 7987 8619
rect 7929 8579 7987 8585
rect 9600 8588 9904 8616
rect 1489 8551 1547 8557
rect 1489 8517 1501 8551
rect 1535 8548 1547 8551
rect 9600 8548 9628 8588
rect 1535 8520 9628 8548
rect 9876 8548 9904 8588
rect 10042 8576 10048 8628
rect 10100 8576 10106 8628
rect 11974 8576 11980 8628
rect 12032 8616 12038 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 12032 8588 12173 8616
rect 12032 8576 12038 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12161 8579 12219 8585
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14277 8619 14335 8625
rect 14277 8616 14289 8619
rect 14056 8588 14289 8616
rect 14056 8576 14062 8588
rect 14277 8585 14289 8588
rect 14323 8585 14335 8619
rect 14277 8579 14335 8585
rect 16114 8576 16120 8628
rect 16172 8616 16178 8628
rect 16393 8619 16451 8625
rect 16393 8616 16405 8619
rect 16172 8588 16405 8616
rect 16172 8576 16178 8588
rect 16393 8585 16405 8588
rect 16439 8585 16451 8619
rect 16393 8579 16451 8585
rect 18230 8576 18236 8628
rect 18288 8616 18294 8628
rect 18509 8619 18567 8625
rect 18509 8616 18521 8619
rect 18288 8588 18521 8616
rect 18288 8576 18294 8588
rect 18509 8585 18521 8588
rect 18555 8585 18567 8619
rect 18509 8579 18567 8585
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 20625 8619 20683 8625
rect 20625 8616 20637 8619
rect 20404 8588 20637 8616
rect 20404 8576 20410 8588
rect 20625 8585 20637 8588
rect 20671 8585 20683 8619
rect 20625 8579 20683 8585
rect 22738 8576 22744 8628
rect 22796 8576 22802 8628
rect 24670 8576 24676 8628
rect 24728 8576 24734 8628
rect 26694 8576 26700 8628
rect 26752 8616 26758 8628
rect 27157 8619 27215 8625
rect 27157 8616 27169 8619
rect 26752 8588 27169 8616
rect 26752 8576 26758 8588
rect 27157 8585 27169 8588
rect 27203 8585 27215 8619
rect 27157 8579 27215 8585
rect 28902 8576 28908 8628
rect 28960 8576 28966 8628
rect 30926 8576 30932 8628
rect 30984 8616 30990 8628
rect 31205 8619 31263 8625
rect 31205 8616 31217 8619
rect 30984 8588 31217 8616
rect 30984 8576 30990 8588
rect 31205 8585 31217 8588
rect 31251 8585 31263 8619
rect 31205 8579 31263 8585
rect 32950 8576 32956 8628
rect 33008 8616 33014 8628
rect 33137 8619 33195 8625
rect 33137 8616 33149 8619
rect 33008 8588 33149 8616
rect 33008 8576 33014 8588
rect 33137 8585 33149 8588
rect 33183 8585 33195 8619
rect 33137 8579 33195 8585
rect 35158 8576 35164 8628
rect 35216 8616 35222 8628
rect 35437 8619 35495 8625
rect 35437 8616 35449 8619
rect 35216 8588 35449 8616
rect 35216 8576 35222 8588
rect 35437 8585 35449 8588
rect 35483 8585 35495 8619
rect 35437 8579 35495 8585
rect 37458 8576 37464 8628
rect 37516 8576 37522 8628
rect 39390 8576 39396 8628
rect 39448 8616 39454 8628
rect 40037 8619 40095 8625
rect 40037 8616 40049 8619
rect 39448 8588 40049 8616
rect 39448 8576 39454 8588
rect 40037 8585 40049 8588
rect 40083 8585 40095 8619
rect 40037 8579 40095 8585
rect 41506 8576 41512 8628
rect 41564 8616 41570 8628
rect 41785 8619 41843 8625
rect 41785 8616 41797 8619
rect 41564 8588 41797 8616
rect 41564 8576 41570 8588
rect 41785 8585 41797 8588
rect 41831 8585 41843 8619
rect 41785 8579 41843 8585
rect 43441 8619 43499 8625
rect 43441 8585 43453 8619
rect 43487 8616 43499 8619
rect 43622 8616 43628 8628
rect 43487 8588 43628 8616
rect 43487 8585 43499 8588
rect 43441 8579 43499 8585
rect 43622 8576 43628 8588
rect 43680 8576 43686 8628
rect 22094 8548 22100 8560
rect 9876 8520 22100 8548
rect 1535 8517 1547 8520
rect 1489 8511 1547 8517
rect 22094 8508 22100 8520
rect 22152 8508 22158 8560
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8480 3847 8483
rect 5169 8483 5227 8489
rect 3835 8452 4476 8480
rect 3835 8449 3847 8452
rect 3789 8443 3847 8449
rect 4448 8356 4476 8452
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5534 8480 5540 8492
rect 5215 8452 5540 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 9766 8489 9772 8492
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 9751 8483 9772 8489
rect 9751 8449 9763 8483
rect 9751 8443 9772 8449
rect 7760 8412 7788 8443
rect 9766 8440 9772 8443
rect 9824 8440 9830 8492
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8480 12035 8483
rect 13906 8480 13912 8492
rect 12023 8452 13912 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 14090 8440 14096 8492
rect 14148 8440 14154 8492
rect 16206 8440 16212 8492
rect 16264 8440 16270 8492
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 18598 8480 18604 8492
rect 18371 8452 18604 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 20438 8440 20444 8492
rect 20496 8440 20502 8492
rect 22557 8483 22615 8489
rect 22557 8449 22569 8483
rect 22603 8480 22615 8483
rect 22922 8480 22928 8492
rect 22603 8452 22928 8480
rect 22603 8449 22615 8452
rect 22557 8443 22615 8449
rect 22922 8440 22928 8452
rect 22980 8440 22986 8492
rect 24581 8483 24639 8489
rect 24581 8449 24593 8483
rect 24627 8480 24639 8483
rect 25038 8480 25044 8492
rect 24627 8452 25044 8480
rect 24627 8449 24639 8452
rect 24581 8443 24639 8449
rect 25038 8440 25044 8452
rect 25096 8440 25102 8492
rect 26970 8440 26976 8492
rect 27028 8440 27034 8492
rect 28813 8483 28871 8489
rect 28813 8449 28825 8483
rect 28859 8480 28871 8483
rect 30098 8480 30104 8492
rect 28859 8452 30104 8480
rect 28859 8449 28871 8452
rect 28813 8443 28871 8449
rect 30098 8440 30104 8452
rect 30156 8440 30162 8492
rect 31018 8440 31024 8492
rect 31076 8440 31082 8492
rect 33045 8483 33103 8489
rect 33045 8449 33057 8483
rect 33091 8480 33103 8483
rect 33502 8480 33508 8492
rect 33091 8452 33508 8480
rect 33091 8449 33103 8452
rect 33045 8443 33103 8449
rect 33502 8440 33508 8452
rect 33560 8440 33566 8492
rect 35253 8483 35311 8489
rect 35253 8449 35265 8483
rect 35299 8480 35311 8483
rect 35299 8452 35894 8480
rect 35299 8449 35311 8452
rect 35253 8443 35311 8449
rect 26326 8412 26332 8424
rect 7760 8384 26332 8412
rect 26326 8372 26332 8384
rect 26384 8372 26390 8424
rect 4430 8304 4436 8356
rect 4488 8304 4494 8356
rect 9401 8347 9459 8353
rect 9401 8313 9413 8347
rect 9447 8344 9459 8347
rect 9766 8344 9772 8356
rect 9447 8316 9772 8344
rect 9447 8313 9459 8316
rect 9401 8307 9459 8313
rect 9766 8304 9772 8316
rect 9824 8344 9830 8356
rect 23290 8344 23296 8356
rect 9824 8316 23296 8344
rect 9824 8304 9830 8316
rect 23290 8304 23296 8316
rect 23348 8304 23354 8356
rect 35866 8344 35894 8452
rect 37366 8440 37372 8492
rect 37424 8440 37430 8492
rect 39942 8440 39948 8492
rect 40000 8440 40006 8492
rect 40678 8440 40684 8492
rect 40736 8480 40742 8492
rect 41693 8483 41751 8489
rect 41693 8480 41705 8483
rect 40736 8452 41705 8480
rect 40736 8440 40742 8452
rect 41693 8449 41705 8452
rect 41739 8449 41751 8483
rect 41693 8443 41751 8449
rect 43254 8440 43260 8492
rect 43312 8440 43318 8492
rect 36354 8344 36360 8356
rect 35866 8316 36360 8344
rect 36354 8304 36360 8316
rect 36412 8304 36418 8356
rect 1104 8186 43884 8208
rect 1104 8134 6297 8186
rect 6349 8134 6361 8186
rect 6413 8134 6425 8186
rect 6477 8134 6489 8186
rect 6541 8134 6553 8186
rect 6605 8134 16991 8186
rect 17043 8134 17055 8186
rect 17107 8134 17119 8186
rect 17171 8134 17183 8186
rect 17235 8134 17247 8186
rect 17299 8134 27685 8186
rect 27737 8134 27749 8186
rect 27801 8134 27813 8186
rect 27865 8134 27877 8186
rect 27929 8134 27941 8186
rect 27993 8134 38379 8186
rect 38431 8134 38443 8186
rect 38495 8134 38507 8186
rect 38559 8134 38571 8186
rect 38623 8134 38635 8186
rect 38687 8134 43884 8186
rect 1104 8112 43884 8134
rect 1104 7642 44040 7664
rect 1104 7590 11644 7642
rect 11696 7590 11708 7642
rect 11760 7590 11772 7642
rect 11824 7590 11836 7642
rect 11888 7590 11900 7642
rect 11952 7590 22338 7642
rect 22390 7590 22402 7642
rect 22454 7590 22466 7642
rect 22518 7590 22530 7642
rect 22582 7590 22594 7642
rect 22646 7590 33032 7642
rect 33084 7590 33096 7642
rect 33148 7590 33160 7642
rect 33212 7590 33224 7642
rect 33276 7590 33288 7642
rect 33340 7590 43726 7642
rect 43778 7590 43790 7642
rect 43842 7590 43854 7642
rect 43906 7590 43918 7642
rect 43970 7590 43982 7642
rect 44034 7590 44040 7642
rect 1104 7568 44040 7590
rect 1104 7098 43884 7120
rect 1104 7046 6297 7098
rect 6349 7046 6361 7098
rect 6413 7046 6425 7098
rect 6477 7046 6489 7098
rect 6541 7046 6553 7098
rect 6605 7046 16991 7098
rect 17043 7046 17055 7098
rect 17107 7046 17119 7098
rect 17171 7046 17183 7098
rect 17235 7046 17247 7098
rect 17299 7046 27685 7098
rect 27737 7046 27749 7098
rect 27801 7046 27813 7098
rect 27865 7046 27877 7098
rect 27929 7046 27941 7098
rect 27993 7046 38379 7098
rect 38431 7046 38443 7098
rect 38495 7046 38507 7098
rect 38559 7046 38571 7098
rect 38623 7046 38635 7098
rect 38687 7046 43884 7098
rect 1104 7024 43884 7046
rect 1104 6554 44040 6576
rect 1104 6502 11644 6554
rect 11696 6502 11708 6554
rect 11760 6502 11772 6554
rect 11824 6502 11836 6554
rect 11888 6502 11900 6554
rect 11952 6502 22338 6554
rect 22390 6502 22402 6554
rect 22454 6502 22466 6554
rect 22518 6502 22530 6554
rect 22582 6502 22594 6554
rect 22646 6502 33032 6554
rect 33084 6502 33096 6554
rect 33148 6502 33160 6554
rect 33212 6502 33224 6554
rect 33276 6502 33288 6554
rect 33340 6502 43726 6554
rect 43778 6502 43790 6554
rect 43842 6502 43854 6554
rect 43906 6502 43918 6554
rect 43970 6502 43982 6554
rect 44034 6502 44040 6554
rect 1104 6480 44040 6502
rect 1104 6010 43884 6032
rect 1104 5958 6297 6010
rect 6349 5958 6361 6010
rect 6413 5958 6425 6010
rect 6477 5958 6489 6010
rect 6541 5958 6553 6010
rect 6605 5958 16991 6010
rect 17043 5958 17055 6010
rect 17107 5958 17119 6010
rect 17171 5958 17183 6010
rect 17235 5958 17247 6010
rect 17299 5958 27685 6010
rect 27737 5958 27749 6010
rect 27801 5958 27813 6010
rect 27865 5958 27877 6010
rect 27929 5958 27941 6010
rect 27993 5958 38379 6010
rect 38431 5958 38443 6010
rect 38495 5958 38507 6010
rect 38559 5958 38571 6010
rect 38623 5958 38635 6010
rect 38687 5958 43884 6010
rect 1104 5936 43884 5958
rect 1104 5466 44040 5488
rect 1104 5414 11644 5466
rect 11696 5414 11708 5466
rect 11760 5414 11772 5466
rect 11824 5414 11836 5466
rect 11888 5414 11900 5466
rect 11952 5414 22338 5466
rect 22390 5414 22402 5466
rect 22454 5414 22466 5466
rect 22518 5414 22530 5466
rect 22582 5414 22594 5466
rect 22646 5414 33032 5466
rect 33084 5414 33096 5466
rect 33148 5414 33160 5466
rect 33212 5414 33224 5466
rect 33276 5414 33288 5466
rect 33340 5414 43726 5466
rect 43778 5414 43790 5466
rect 43842 5414 43854 5466
rect 43906 5414 43918 5466
rect 43970 5414 43982 5466
rect 44034 5414 44040 5466
rect 1104 5392 44040 5414
rect 1104 4922 43884 4944
rect 1104 4870 6297 4922
rect 6349 4870 6361 4922
rect 6413 4870 6425 4922
rect 6477 4870 6489 4922
rect 6541 4870 6553 4922
rect 6605 4870 16991 4922
rect 17043 4870 17055 4922
rect 17107 4870 17119 4922
rect 17171 4870 17183 4922
rect 17235 4870 17247 4922
rect 17299 4870 27685 4922
rect 27737 4870 27749 4922
rect 27801 4870 27813 4922
rect 27865 4870 27877 4922
rect 27929 4870 27941 4922
rect 27993 4870 38379 4922
rect 38431 4870 38443 4922
rect 38495 4870 38507 4922
rect 38559 4870 38571 4922
rect 38623 4870 38635 4922
rect 38687 4870 43884 4922
rect 1104 4848 43884 4870
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 23474 4672 23480 4684
rect 6880 4644 23480 4672
rect 6880 4632 6886 4644
rect 23474 4632 23480 4644
rect 23532 4632 23538 4684
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 23934 4604 23940 4616
rect 6788 4576 23940 4604
rect 6788 4564 6794 4576
rect 23934 4564 23940 4576
rect 23992 4564 23998 4616
rect 11974 4496 11980 4548
rect 12032 4536 12038 4548
rect 28074 4536 28080 4548
rect 12032 4508 28080 4536
rect 12032 4496 12038 4508
rect 28074 4496 28080 4508
rect 28132 4496 28138 4548
rect 11330 4428 11336 4480
rect 11388 4468 11394 4480
rect 28810 4468 28816 4480
rect 11388 4440 28816 4468
rect 11388 4428 11394 4440
rect 28810 4428 28816 4440
rect 28868 4428 28874 4480
rect 1104 4378 44040 4400
rect 1104 4326 11644 4378
rect 11696 4326 11708 4378
rect 11760 4326 11772 4378
rect 11824 4326 11836 4378
rect 11888 4326 11900 4378
rect 11952 4326 22338 4378
rect 22390 4326 22402 4378
rect 22454 4326 22466 4378
rect 22518 4326 22530 4378
rect 22582 4326 22594 4378
rect 22646 4326 33032 4378
rect 33084 4326 33096 4378
rect 33148 4326 33160 4378
rect 33212 4326 33224 4378
rect 33276 4326 33288 4378
rect 33340 4326 43726 4378
rect 43778 4326 43790 4378
rect 43842 4326 43854 4378
rect 43906 4326 43918 4378
rect 43970 4326 43982 4378
rect 44034 4326 44040 4378
rect 1104 4304 44040 4326
rect 16482 4224 16488 4276
rect 16540 4264 16546 4276
rect 33778 4264 33784 4276
rect 16540 4236 33784 4264
rect 16540 4224 16546 4236
rect 33778 4224 33784 4236
rect 33836 4224 33842 4276
rect 15654 4156 15660 4208
rect 15712 4196 15718 4208
rect 34882 4196 34888 4208
rect 15712 4168 34888 4196
rect 15712 4156 15718 4168
rect 34882 4156 34888 4168
rect 34940 4156 34946 4208
rect 1104 3834 43884 3856
rect 1104 3782 6297 3834
rect 6349 3782 6361 3834
rect 6413 3782 6425 3834
rect 6477 3782 6489 3834
rect 6541 3782 6553 3834
rect 6605 3782 16991 3834
rect 17043 3782 17055 3834
rect 17107 3782 17119 3834
rect 17171 3782 17183 3834
rect 17235 3782 17247 3834
rect 17299 3782 27685 3834
rect 27737 3782 27749 3834
rect 27801 3782 27813 3834
rect 27865 3782 27877 3834
rect 27929 3782 27941 3834
rect 27993 3782 38379 3834
rect 38431 3782 38443 3834
rect 38495 3782 38507 3834
rect 38559 3782 38571 3834
rect 38623 3782 38635 3834
rect 38687 3782 43884 3834
rect 1104 3760 43884 3782
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 30374 3448 30380 3460
rect 16356 3420 30380 3448
rect 16356 3408 16362 3420
rect 30374 3408 30380 3420
rect 30432 3408 30438 3460
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 21450 3380 21456 3392
rect 8076 3352 21456 3380
rect 8076 3340 8082 3352
rect 21450 3340 21456 3352
rect 21508 3340 21514 3392
rect 1104 3290 44040 3312
rect 1104 3238 11644 3290
rect 11696 3238 11708 3290
rect 11760 3238 11772 3290
rect 11824 3238 11836 3290
rect 11888 3238 11900 3290
rect 11952 3238 22338 3290
rect 22390 3238 22402 3290
rect 22454 3238 22466 3290
rect 22518 3238 22530 3290
rect 22582 3238 22594 3290
rect 22646 3238 33032 3290
rect 33084 3238 33096 3290
rect 33148 3238 33160 3290
rect 33212 3238 33224 3290
rect 33276 3238 33288 3290
rect 33340 3238 43726 3290
rect 43778 3238 43790 3290
rect 43842 3238 43854 3290
rect 43906 3238 43918 3290
rect 43970 3238 43982 3290
rect 44034 3238 44040 3290
rect 1104 3216 44040 3238
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 26142 3176 26148 3188
rect 18012 3148 26148 3176
rect 18012 3136 18018 3148
rect 26142 3136 26148 3148
rect 26200 3136 26206 3188
rect 27525 3179 27583 3185
rect 27525 3145 27537 3179
rect 27571 3176 27583 3179
rect 29914 3176 29920 3188
rect 27571 3148 29920 3176
rect 27571 3145 27583 3148
rect 27525 3139 27583 3145
rect 29914 3136 29920 3148
rect 29972 3136 29978 3188
rect 17678 3068 17684 3120
rect 17736 3108 17742 3120
rect 37274 3108 37280 3120
rect 17736 3080 26096 3108
rect 17736 3068 17742 3080
rect 26068 3052 26096 3080
rect 27172 3080 29224 3108
rect 5350 3000 5356 3052
rect 5408 3040 5414 3052
rect 19613 3043 19671 3049
rect 19613 3040 19625 3043
rect 5408 3012 19625 3040
rect 5408 3000 5414 3012
rect 19613 3009 19625 3012
rect 19659 3009 19671 3043
rect 19613 3003 19671 3009
rect 21913 3043 21971 3049
rect 21913 3009 21925 3043
rect 21959 3040 21971 3043
rect 25406 3040 25412 3052
rect 21959 3012 25412 3040
rect 21959 3009 21971 3012
rect 21913 3003 21971 3009
rect 25406 3000 25412 3012
rect 25464 3000 25470 3052
rect 26050 3000 26056 3052
rect 26108 3000 26114 3052
rect 27172 3049 27200 3080
rect 27157 3043 27215 3049
rect 27157 3009 27169 3043
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 27433 3043 27491 3049
rect 27433 3009 27445 3043
rect 27479 3009 27491 3043
rect 27433 3003 27491 3009
rect 27709 3043 27767 3049
rect 27709 3009 27721 3043
rect 27755 3040 27767 3043
rect 28074 3040 28080 3052
rect 27755 3012 28080 3040
rect 27755 3009 27767 3012
rect 27709 3003 27767 3009
rect 12250 2932 12256 2984
rect 12308 2972 12314 2984
rect 27448 2972 27476 3003
rect 28074 3000 28080 3012
rect 28132 3000 28138 3052
rect 28258 3000 28264 3052
rect 28316 3000 28322 3052
rect 28537 3043 28595 3049
rect 28537 3009 28549 3043
rect 28583 3009 28595 3043
rect 28537 3003 28595 3009
rect 12308 2944 27476 2972
rect 12308 2932 12314 2944
rect 27614 2932 27620 2984
rect 27672 2972 27678 2984
rect 28552 2972 28580 3003
rect 28810 3000 28816 3052
rect 28868 3000 28874 3052
rect 27672 2944 28580 2972
rect 27672 2932 27678 2944
rect 16574 2864 16580 2916
rect 16632 2904 16638 2916
rect 16632 2876 22048 2904
rect 16632 2864 16638 2876
rect 11514 2796 11520 2848
rect 11572 2836 11578 2848
rect 19334 2836 19340 2848
rect 11572 2808 19340 2836
rect 11572 2796 11578 2808
rect 19334 2796 19340 2808
rect 19392 2796 19398 2848
rect 19426 2796 19432 2848
rect 19484 2796 19490 2848
rect 22020 2836 22048 2876
rect 22094 2864 22100 2916
rect 22152 2864 22158 2916
rect 24670 2864 24676 2916
rect 24728 2864 24734 2916
rect 25222 2864 25228 2916
rect 25280 2904 25286 2916
rect 25866 2904 25872 2916
rect 25280 2876 25872 2904
rect 25280 2864 25286 2876
rect 25866 2864 25872 2876
rect 25924 2864 25930 2916
rect 27430 2864 27436 2916
rect 27488 2904 27494 2916
rect 29196 2904 29224 3080
rect 31726 3080 37280 3108
rect 29273 3043 29331 3049
rect 29273 3009 29285 3043
rect 29319 3009 29331 3043
rect 29273 3003 29331 3009
rect 29549 3043 29607 3049
rect 29549 3009 29561 3043
rect 29595 3040 29607 3043
rect 31726 3040 31754 3080
rect 37274 3068 37280 3080
rect 37332 3068 37338 3120
rect 39206 3040 39212 3052
rect 29595 3012 31754 3040
rect 35866 3012 39212 3040
rect 29595 3009 29607 3012
rect 29549 3003 29607 3009
rect 29288 2972 29316 3003
rect 35866 2972 35894 3012
rect 39206 3000 39212 3012
rect 39264 3000 39270 3052
rect 29288 2944 35894 2972
rect 31754 2904 31760 2916
rect 27488 2876 29132 2904
rect 29196 2876 31760 2904
rect 27488 2864 27494 2876
rect 24688 2836 24716 2864
rect 22020 2808 24716 2836
rect 25314 2796 25320 2848
rect 25372 2836 25378 2848
rect 26234 2836 26240 2848
rect 25372 2808 26240 2836
rect 25372 2796 25378 2808
rect 26234 2796 26240 2808
rect 26292 2796 26298 2848
rect 26418 2796 26424 2848
rect 26476 2836 26482 2848
rect 26973 2839 27031 2845
rect 26973 2836 26985 2839
rect 26476 2808 26985 2836
rect 26476 2796 26482 2808
rect 26973 2805 26985 2808
rect 27019 2805 27031 2839
rect 26973 2799 27031 2805
rect 27246 2796 27252 2848
rect 27304 2796 27310 2848
rect 28074 2796 28080 2848
rect 28132 2796 28138 2848
rect 28350 2796 28356 2848
rect 28408 2796 28414 2848
rect 28626 2796 28632 2848
rect 28684 2796 28690 2848
rect 29104 2845 29132 2876
rect 31754 2864 31760 2876
rect 31812 2864 31818 2916
rect 29089 2839 29147 2845
rect 29089 2805 29101 2839
rect 29135 2805 29147 2839
rect 29089 2799 29147 2805
rect 29362 2796 29368 2848
rect 29420 2796 29426 2848
rect 31110 2796 31116 2848
rect 31168 2836 31174 2848
rect 32950 2836 32956 2848
rect 31168 2808 32956 2836
rect 31168 2796 31174 2808
rect 32950 2796 32956 2808
rect 33008 2796 33014 2848
rect 1104 2746 43884 2768
rect 1104 2694 6297 2746
rect 6349 2694 6361 2746
rect 6413 2694 6425 2746
rect 6477 2694 6489 2746
rect 6541 2694 6553 2746
rect 6605 2694 16991 2746
rect 17043 2694 17055 2746
rect 17107 2694 17119 2746
rect 17171 2694 17183 2746
rect 17235 2694 17247 2746
rect 17299 2694 27685 2746
rect 27737 2694 27749 2746
rect 27801 2694 27813 2746
rect 27865 2694 27877 2746
rect 27929 2694 27941 2746
rect 27993 2694 38379 2746
rect 38431 2694 38443 2746
rect 38495 2694 38507 2746
rect 38559 2694 38571 2746
rect 38623 2694 38635 2746
rect 38687 2694 43884 2746
rect 1104 2672 43884 2694
rect 14090 2592 14096 2644
rect 14148 2592 14154 2644
rect 16298 2592 16304 2644
rect 16356 2592 16362 2644
rect 16390 2592 16396 2644
rect 16448 2632 16454 2644
rect 16485 2635 16543 2641
rect 16485 2632 16497 2635
rect 16448 2604 16497 2632
rect 16448 2592 16454 2604
rect 16485 2601 16497 2604
rect 16531 2601 16543 2635
rect 16485 2595 16543 2601
rect 18506 2592 18512 2644
rect 18564 2592 18570 2644
rect 18598 2592 18604 2644
rect 18656 2592 18662 2644
rect 18966 2592 18972 2644
rect 19024 2632 19030 2644
rect 19024 2604 20484 2632
rect 19024 2592 19030 2604
rect 17129 2567 17187 2573
rect 17129 2533 17141 2567
rect 17175 2564 17187 2567
rect 17770 2564 17776 2576
rect 17175 2536 17776 2564
rect 17175 2533 17187 2536
rect 17129 2527 17187 2533
rect 17770 2524 17776 2536
rect 17828 2524 17834 2576
rect 14274 2388 14280 2440
rect 14332 2388 14338 2440
rect 14642 2388 14648 2440
rect 14700 2428 14706 2440
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 14700 2400 16129 2428
rect 14700 2388 14706 2400
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16356 2400 16681 2428
rect 16356 2388 16362 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 16945 2431 17003 2437
rect 16945 2428 16957 2431
rect 16816 2400 16957 2428
rect 16816 2388 16822 2400
rect 16945 2397 16957 2400
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 18325 2431 18383 2437
rect 18325 2397 18337 2431
rect 18371 2428 18383 2431
rect 18414 2428 18420 2440
rect 18371 2400 18420 2428
rect 18371 2397 18383 2400
rect 18325 2391 18383 2397
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 18506 2388 18512 2440
rect 18564 2388 18570 2440
rect 10410 2320 10416 2372
rect 10468 2360 10474 2372
rect 18524 2360 18552 2388
rect 10468 2332 18552 2360
rect 10468 2320 10474 2332
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 18506 2292 18512 2304
rect 9732 2264 18512 2292
rect 9732 2252 9738 2264
rect 18506 2252 18512 2264
rect 18564 2252 18570 2304
rect 18616 2301 18644 2592
rect 19429 2567 19487 2573
rect 19429 2533 19441 2567
rect 19475 2564 19487 2567
rect 19794 2564 19800 2576
rect 19475 2536 19800 2564
rect 19475 2533 19487 2536
rect 19429 2527 19487 2533
rect 19794 2524 19800 2536
rect 19852 2524 19858 2576
rect 20257 2567 20315 2573
rect 20257 2533 20269 2567
rect 20303 2564 20315 2567
rect 20456 2564 20484 2604
rect 20530 2592 20536 2644
rect 20588 2592 20594 2644
rect 20806 2592 20812 2644
rect 20864 2592 20870 2644
rect 22922 2592 22928 2644
rect 22980 2592 22986 2644
rect 23566 2592 23572 2644
rect 23624 2632 23630 2644
rect 24581 2635 24639 2641
rect 24581 2632 24593 2635
rect 23624 2604 24593 2632
rect 23624 2592 23630 2604
rect 24581 2601 24593 2604
rect 24627 2601 24639 2635
rect 24581 2595 24639 2601
rect 24946 2592 24952 2644
rect 25004 2592 25010 2644
rect 25038 2592 25044 2644
rect 25096 2592 25102 2644
rect 26326 2592 26332 2644
rect 26384 2632 26390 2644
rect 26605 2635 26663 2641
rect 26605 2632 26617 2635
rect 26384 2604 26617 2632
rect 26384 2592 26390 2604
rect 26605 2601 26617 2604
rect 26651 2601 26663 2635
rect 26605 2595 26663 2601
rect 27154 2592 27160 2644
rect 27212 2632 27218 2644
rect 27249 2635 27307 2641
rect 27249 2632 27261 2635
rect 27212 2604 27261 2632
rect 27212 2592 27218 2604
rect 27249 2601 27261 2604
rect 27295 2601 27307 2635
rect 27249 2595 27307 2601
rect 27338 2592 27344 2644
rect 27396 2632 27402 2644
rect 30926 2632 30932 2644
rect 27396 2604 30932 2632
rect 27396 2592 27402 2604
rect 30926 2592 30932 2604
rect 30984 2592 30990 2644
rect 31018 2592 31024 2644
rect 31076 2632 31082 2644
rect 31389 2635 31447 2641
rect 31389 2632 31401 2635
rect 31076 2604 31401 2632
rect 31076 2592 31082 2604
rect 31389 2601 31401 2604
rect 31435 2601 31447 2635
rect 31389 2595 31447 2601
rect 33502 2592 33508 2644
rect 33560 2592 33566 2644
rect 33778 2592 33784 2644
rect 33836 2632 33842 2644
rect 34146 2632 34152 2644
rect 33836 2604 34152 2632
rect 33836 2592 33842 2604
rect 34146 2592 34152 2604
rect 34204 2592 34210 2644
rect 36354 2592 36360 2644
rect 36412 2592 36418 2644
rect 37366 2592 37372 2644
rect 37424 2632 37430 2644
rect 37737 2635 37795 2641
rect 37737 2632 37749 2635
rect 37424 2604 37749 2632
rect 37424 2592 37430 2604
rect 37737 2601 37749 2604
rect 37783 2601 37795 2635
rect 37737 2595 37795 2601
rect 39485 2635 39543 2641
rect 39485 2601 39497 2635
rect 39531 2632 39543 2635
rect 39942 2632 39948 2644
rect 39531 2604 39948 2632
rect 39531 2601 39543 2604
rect 39485 2595 39543 2601
rect 39942 2592 39948 2604
rect 40000 2592 40006 2644
rect 40678 2592 40684 2644
rect 40736 2592 40742 2644
rect 42245 2635 42303 2641
rect 42245 2601 42257 2635
rect 42291 2632 42303 2635
rect 43254 2632 43260 2644
rect 42291 2604 43260 2632
rect 42291 2601 42303 2604
rect 42245 2595 42303 2601
rect 43254 2592 43260 2604
rect 43312 2592 43318 2644
rect 25222 2564 25228 2576
rect 20303 2536 20392 2564
rect 20456 2536 23980 2564
rect 20303 2533 20315 2536
rect 20257 2527 20315 2533
rect 18690 2456 18696 2508
rect 18748 2496 18754 2508
rect 20364 2496 20392 2536
rect 18748 2468 20300 2496
rect 20364 2468 21404 2496
rect 18748 2456 18754 2468
rect 18782 2388 18788 2440
rect 18840 2388 18846 2440
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2428 18935 2431
rect 19058 2428 19064 2440
rect 18923 2400 19064 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 19058 2388 19064 2400
rect 19116 2388 19122 2440
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 19889 2431 19947 2437
rect 19889 2397 19901 2431
rect 19935 2428 19947 2431
rect 20070 2428 20076 2440
rect 19935 2400 20076 2428
rect 19935 2397 19947 2400
rect 19889 2391 19947 2397
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 20162 2388 20168 2440
rect 20220 2388 20226 2440
rect 20272 2428 20300 2468
rect 20441 2431 20499 2437
rect 20441 2428 20453 2431
rect 20272 2400 20453 2428
rect 20441 2397 20453 2400
rect 20487 2397 20499 2431
rect 20441 2391 20499 2397
rect 20717 2431 20775 2437
rect 20717 2397 20729 2431
rect 20763 2428 20775 2431
rect 20806 2428 20812 2440
rect 20763 2400 20812 2428
rect 20763 2397 20775 2400
rect 20717 2391 20775 2397
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 20990 2388 20996 2440
rect 21048 2388 21054 2440
rect 21266 2388 21272 2440
rect 21324 2388 21330 2440
rect 21376 2437 21404 2468
rect 21361 2431 21419 2437
rect 21361 2397 21373 2431
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 21450 2388 21456 2440
rect 21508 2428 21514 2440
rect 22097 2431 22155 2437
rect 22097 2428 22109 2431
rect 21508 2400 22109 2428
rect 21508 2388 21514 2400
rect 22097 2397 22109 2400
rect 22143 2397 22155 2431
rect 22097 2391 22155 2397
rect 22370 2388 22376 2440
rect 22428 2388 22434 2440
rect 22649 2431 22707 2437
rect 22649 2397 22661 2431
rect 22695 2428 22707 2431
rect 22738 2428 22744 2440
rect 22695 2400 22744 2428
rect 22695 2397 22707 2400
rect 22649 2391 22707 2397
rect 22738 2388 22744 2400
rect 22796 2388 22802 2440
rect 23109 2431 23167 2437
rect 23109 2397 23121 2431
rect 23155 2428 23167 2431
rect 23566 2428 23572 2440
rect 23155 2400 23572 2428
rect 23155 2397 23167 2400
rect 23109 2391 23167 2397
rect 23566 2388 23572 2400
rect 23624 2388 23630 2440
rect 23842 2360 23848 2372
rect 19076 2332 23848 2360
rect 19076 2301 19104 2332
rect 23842 2320 23848 2332
rect 23900 2320 23906 2372
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2261 18659 2295
rect 18601 2255 18659 2261
rect 19061 2295 19119 2301
rect 19061 2261 19073 2295
rect 19107 2261 19119 2295
rect 19061 2255 19119 2261
rect 19705 2295 19763 2301
rect 19705 2261 19717 2295
rect 19751 2292 19763 2295
rect 19886 2292 19892 2304
rect 19751 2264 19892 2292
rect 19751 2261 19763 2264
rect 19705 2255 19763 2261
rect 19886 2252 19892 2264
rect 19944 2252 19950 2304
rect 19981 2295 20039 2301
rect 19981 2261 19993 2295
rect 20027 2292 20039 2295
rect 20438 2292 20444 2304
rect 20027 2264 20444 2292
rect 20027 2261 20039 2264
rect 19981 2255 20039 2261
rect 20438 2252 20444 2264
rect 20496 2252 20502 2304
rect 21085 2295 21143 2301
rect 21085 2261 21097 2295
rect 21131 2292 21143 2295
rect 21266 2292 21272 2304
rect 21131 2264 21272 2292
rect 21131 2261 21143 2264
rect 21085 2255 21143 2261
rect 21266 2252 21272 2264
rect 21324 2252 21330 2304
rect 21542 2252 21548 2304
rect 21600 2252 21606 2304
rect 21913 2295 21971 2301
rect 21913 2261 21925 2295
rect 21959 2292 21971 2295
rect 22002 2292 22008 2304
rect 21959 2264 22008 2292
rect 21959 2261 21971 2264
rect 21913 2255 21971 2261
rect 22002 2252 22008 2264
rect 22060 2252 22066 2304
rect 22186 2252 22192 2304
rect 22244 2252 22250 2304
rect 22465 2295 22523 2301
rect 22465 2261 22477 2295
rect 22511 2292 22523 2295
rect 23198 2292 23204 2304
rect 22511 2264 23204 2292
rect 22511 2261 22523 2264
rect 22465 2255 22523 2261
rect 23198 2252 23204 2264
rect 23256 2252 23262 2304
rect 23952 2292 23980 2536
rect 24780 2536 25228 2564
rect 24780 2437 24808 2536
rect 25222 2524 25228 2536
rect 25280 2524 25286 2576
rect 25317 2567 25375 2573
rect 25317 2533 25329 2567
rect 25363 2533 25375 2567
rect 25317 2527 25375 2533
rect 25332 2496 25360 2527
rect 25590 2524 25596 2576
rect 25648 2524 25654 2576
rect 25866 2524 25872 2576
rect 25924 2524 25930 2576
rect 37642 2564 37648 2576
rect 26528 2536 37648 2564
rect 26528 2496 26556 2536
rect 37642 2524 37648 2536
rect 37700 2524 37706 2576
rect 24872 2468 25360 2496
rect 25700 2468 26556 2496
rect 24397 2431 24455 2437
rect 24397 2397 24409 2431
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 24765 2431 24823 2437
rect 24765 2397 24777 2431
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 24412 2360 24440 2391
rect 24872 2360 24900 2468
rect 25225 2431 25283 2437
rect 25225 2397 25237 2431
rect 25271 2428 25283 2431
rect 25314 2428 25320 2440
rect 25271 2400 25320 2428
rect 25271 2397 25283 2400
rect 25225 2391 25283 2397
rect 25314 2388 25320 2400
rect 25372 2388 25378 2440
rect 25501 2431 25559 2437
rect 25501 2397 25513 2431
rect 25547 2428 25559 2431
rect 25700 2428 25728 2468
rect 26602 2456 26608 2508
rect 26660 2496 26666 2508
rect 34238 2496 34244 2508
rect 26660 2468 30236 2496
rect 26660 2456 26666 2468
rect 25547 2400 25728 2428
rect 25777 2407 25835 2413
rect 25547 2397 25559 2400
rect 25501 2391 25559 2397
rect 25777 2373 25789 2407
rect 25823 2373 25835 2407
rect 25958 2388 25964 2440
rect 26016 2428 26022 2440
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 26016 2400 26065 2428
rect 26016 2388 26022 2400
rect 26053 2397 26065 2400
rect 26099 2397 26111 2431
rect 26053 2391 26111 2397
rect 26326 2388 26332 2440
rect 26384 2388 26390 2440
rect 26418 2388 26424 2440
rect 26476 2388 26482 2440
rect 26786 2388 26792 2440
rect 26844 2428 26850 2440
rect 26881 2431 26939 2437
rect 26881 2428 26893 2431
rect 26844 2400 26893 2428
rect 26844 2388 26850 2400
rect 26881 2397 26893 2400
rect 26927 2397 26939 2431
rect 26881 2391 26939 2397
rect 26970 2388 26976 2440
rect 27028 2428 27034 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27028 2400 27169 2428
rect 27028 2388 27034 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 27430 2388 27436 2440
rect 27488 2388 27494 2440
rect 27709 2431 27767 2437
rect 27709 2397 27721 2431
rect 27755 2428 27767 2431
rect 28074 2428 28080 2440
rect 27755 2400 28080 2428
rect 27755 2397 27767 2400
rect 27709 2391 27767 2397
rect 28074 2388 28080 2400
rect 28132 2388 28138 2440
rect 28166 2388 28172 2440
rect 28224 2388 28230 2440
rect 28353 2431 28411 2437
rect 28353 2397 28365 2431
rect 28399 2397 28411 2431
rect 28353 2391 28411 2397
rect 28721 2431 28779 2437
rect 28721 2397 28733 2431
rect 28767 2428 28779 2431
rect 28994 2428 29000 2440
rect 28767 2400 29000 2428
rect 28767 2397 28779 2400
rect 28721 2391 28779 2397
rect 25777 2367 25835 2373
rect 24412 2332 24900 2360
rect 25792 2292 25820 2367
rect 28368 2360 28396 2391
rect 28994 2388 29000 2400
rect 29052 2388 29058 2440
rect 29178 2388 29184 2440
rect 29236 2388 29242 2440
rect 29733 2431 29791 2437
rect 29733 2397 29745 2431
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 28368 2332 29040 2360
rect 23952 2264 25820 2292
rect 26145 2295 26203 2301
rect 26145 2261 26157 2295
rect 26191 2292 26203 2295
rect 26234 2292 26240 2304
rect 26191 2264 26240 2292
rect 26191 2261 26203 2264
rect 26145 2255 26203 2261
rect 26234 2252 26240 2264
rect 26292 2252 26298 2304
rect 26694 2252 26700 2304
rect 26752 2252 26758 2304
rect 26786 2252 26792 2304
rect 26844 2292 26850 2304
rect 26973 2295 27031 2301
rect 26973 2292 26985 2295
rect 26844 2264 26985 2292
rect 26844 2252 26850 2264
rect 26973 2261 26985 2264
rect 27019 2261 27031 2295
rect 26973 2255 27031 2261
rect 27798 2252 27804 2304
rect 27856 2252 27862 2304
rect 27982 2252 27988 2304
rect 28040 2252 28046 2304
rect 28258 2252 28264 2304
rect 28316 2292 28322 2304
rect 28537 2295 28595 2301
rect 28537 2292 28549 2295
rect 28316 2264 28549 2292
rect 28316 2252 28322 2264
rect 28537 2261 28549 2264
rect 28583 2261 28595 2295
rect 28537 2255 28595 2261
rect 28718 2252 28724 2304
rect 28776 2292 28782 2304
rect 29012 2301 29040 2332
rect 29086 2320 29092 2372
rect 29144 2360 29150 2372
rect 29748 2360 29776 2391
rect 30006 2388 30012 2440
rect 30064 2388 30070 2440
rect 30098 2388 30104 2440
rect 30156 2388 30162 2440
rect 29144 2332 29776 2360
rect 29144 2320 29150 2332
rect 28905 2295 28963 2301
rect 28905 2292 28917 2295
rect 28776 2264 28917 2292
rect 28776 2252 28782 2264
rect 28905 2261 28917 2264
rect 28951 2261 28963 2295
rect 28905 2255 28963 2261
rect 28997 2295 29055 2301
rect 28997 2261 29009 2295
rect 29043 2261 29055 2295
rect 28997 2255 29055 2261
rect 29546 2252 29552 2304
rect 29604 2252 29610 2304
rect 29822 2252 29828 2304
rect 29880 2252 29886 2304
rect 30116 2301 30144 2388
rect 30208 2304 30236 2468
rect 30576 2468 34244 2496
rect 30576 2437 30604 2468
rect 34238 2456 34244 2468
rect 34296 2456 34302 2508
rect 30285 2431 30343 2437
rect 30285 2397 30297 2431
rect 30331 2428 30343 2431
rect 30561 2431 30619 2437
rect 30331 2400 30420 2428
rect 30331 2397 30343 2400
rect 30285 2391 30343 2397
rect 30101 2295 30159 2301
rect 30101 2261 30113 2295
rect 30147 2261 30159 2295
rect 30101 2255 30159 2261
rect 30190 2252 30196 2304
rect 30248 2252 30254 2304
rect 30392 2301 30420 2400
rect 30561 2397 30573 2431
rect 30607 2397 30619 2431
rect 31565 2427 31623 2433
rect 31565 2424 31577 2427
rect 30561 2391 30619 2397
rect 31496 2396 31577 2424
rect 30377 2295 30435 2301
rect 30377 2261 30389 2295
rect 30423 2261 30435 2295
rect 31496 2292 31524 2396
rect 31565 2393 31577 2396
rect 31611 2393 31623 2427
rect 31565 2387 31623 2393
rect 31941 2431 31999 2437
rect 31941 2397 31953 2431
rect 31987 2428 31999 2431
rect 31987 2400 32812 2428
rect 31987 2397 31999 2400
rect 31941 2391 31999 2397
rect 32784 2360 32812 2400
rect 32858 2388 32864 2440
rect 32916 2388 32922 2440
rect 33686 2388 33692 2440
rect 33744 2388 33750 2440
rect 36538 2388 36544 2440
rect 36596 2388 36602 2440
rect 37918 2388 37924 2440
rect 37976 2388 37982 2440
rect 39666 2388 39672 2440
rect 39724 2388 39730 2440
rect 40862 2388 40868 2440
rect 40920 2388 40926 2440
rect 42426 2388 42432 2440
rect 42484 2388 42490 2440
rect 35618 2360 35624 2372
rect 32784 2332 35624 2360
rect 35618 2320 35624 2332
rect 35676 2320 35682 2372
rect 31757 2295 31815 2301
rect 31757 2292 31769 2295
rect 31496 2264 31769 2292
rect 30377 2255 30435 2261
rect 31757 2261 31769 2264
rect 31803 2261 31815 2295
rect 31757 2255 31815 2261
rect 32582 2252 32588 2304
rect 32640 2292 32646 2304
rect 33045 2295 33103 2301
rect 33045 2292 33057 2295
rect 32640 2264 33057 2292
rect 32640 2252 32646 2264
rect 33045 2261 33057 2264
rect 33091 2261 33103 2295
rect 33045 2255 33103 2261
rect 1104 2202 44040 2224
rect 1104 2150 11644 2202
rect 11696 2150 11708 2202
rect 11760 2150 11772 2202
rect 11824 2150 11836 2202
rect 11888 2150 11900 2202
rect 11952 2150 22338 2202
rect 22390 2150 22402 2202
rect 22454 2150 22466 2202
rect 22518 2150 22530 2202
rect 22582 2150 22594 2202
rect 22646 2150 33032 2202
rect 33084 2150 33096 2202
rect 33148 2150 33160 2202
rect 33212 2150 33224 2202
rect 33276 2150 33288 2202
rect 33340 2150 43726 2202
rect 43778 2150 43790 2202
rect 43842 2150 43854 2202
rect 43906 2150 43918 2202
rect 43970 2150 43982 2202
rect 44034 2150 44040 2202
rect 1104 2128 44040 2150
rect 6730 2048 6736 2100
rect 6788 2048 6794 2100
rect 14185 2091 14243 2097
rect 14185 2057 14197 2091
rect 14231 2088 14243 2091
rect 14274 2088 14280 2100
rect 14231 2060 14280 2088
rect 14231 2057 14243 2060
rect 14185 2051 14243 2057
rect 14274 2048 14280 2060
rect 14332 2048 14338 2100
rect 15378 2048 15384 2100
rect 15436 2048 15442 2100
rect 15654 2048 15660 2100
rect 15712 2048 15718 2100
rect 15933 2091 15991 2097
rect 15933 2057 15945 2091
rect 15979 2057 15991 2091
rect 15933 2051 15991 2057
rect 16025 2091 16083 2097
rect 16025 2057 16037 2091
rect 16071 2088 16083 2091
rect 16298 2088 16304 2100
rect 16071 2060 16304 2088
rect 16071 2057 16083 2060
rect 16025 2051 16083 2057
rect 6546 1912 6552 1964
rect 6604 1912 6610 1964
rect 13722 1912 13728 1964
rect 13780 1912 13786 1964
rect 14366 1912 14372 1964
rect 14424 1912 14430 1964
rect 15102 1912 15108 1964
rect 15160 1912 15166 1964
rect 15197 1955 15255 1961
rect 15197 1921 15209 1955
rect 15243 1952 15255 1955
rect 15286 1952 15292 1964
rect 15243 1924 15292 1952
rect 15243 1921 15255 1924
rect 15197 1915 15255 1921
rect 15286 1912 15292 1924
rect 15344 1912 15350 1964
rect 15473 1955 15531 1961
rect 15473 1921 15485 1955
rect 15519 1921 15531 1955
rect 15473 1915 15531 1921
rect 14918 1844 14924 1896
rect 14976 1884 14982 1896
rect 15488 1884 15516 1915
rect 15746 1912 15752 1964
rect 15804 1912 15810 1964
rect 14976 1856 15516 1884
rect 15948 1884 15976 2051
rect 16298 2048 16304 2060
rect 16356 2048 16362 2100
rect 16482 2048 16488 2100
rect 16540 2048 16546 2100
rect 16850 2048 16856 2100
rect 16908 2088 16914 2100
rect 16945 2091 17003 2097
rect 16945 2088 16957 2091
rect 16908 2060 16957 2088
rect 16908 2048 16914 2060
rect 16945 2057 16957 2060
rect 16991 2057 17003 2091
rect 16945 2051 17003 2057
rect 17221 2091 17279 2097
rect 17221 2057 17233 2091
rect 17267 2088 17279 2091
rect 17678 2088 17684 2100
rect 17267 2060 17684 2088
rect 17267 2057 17279 2060
rect 17221 2051 17279 2057
rect 17678 2048 17684 2060
rect 17736 2048 17742 2100
rect 17865 2091 17923 2097
rect 17865 2057 17877 2091
rect 17911 2057 17923 2091
rect 17865 2051 17923 2057
rect 18141 2091 18199 2097
rect 18141 2057 18153 2091
rect 18187 2088 18199 2091
rect 18782 2088 18788 2100
rect 18187 2060 18788 2088
rect 18187 2057 18199 2060
rect 18141 2051 18199 2057
rect 17880 2020 17908 2051
rect 18782 2048 18788 2060
rect 18840 2048 18846 2100
rect 18969 2091 19027 2097
rect 18969 2057 18981 2091
rect 19015 2088 19027 2091
rect 20530 2088 20536 2100
rect 19015 2060 20116 2088
rect 19015 2057 19027 2060
rect 18969 2051 19027 2057
rect 17880 1992 19564 2020
rect 16206 1912 16212 1964
rect 16264 1912 16270 1964
rect 16298 1912 16304 1964
rect 16356 1912 16362 1964
rect 16390 1912 16396 1964
rect 16448 1952 16454 1964
rect 16761 1955 16819 1961
rect 16761 1952 16773 1955
rect 16448 1924 16773 1952
rect 16448 1912 16454 1924
rect 16761 1921 16773 1924
rect 16807 1921 16819 1955
rect 16761 1915 16819 1921
rect 16850 1912 16856 1964
rect 16908 1952 16914 1964
rect 17037 1955 17095 1961
rect 17037 1952 17049 1955
rect 16908 1924 17049 1952
rect 16908 1912 16914 1924
rect 17037 1921 17049 1924
rect 17083 1921 17095 1955
rect 17037 1915 17095 1921
rect 17310 1912 17316 1964
rect 17368 1912 17374 1964
rect 17586 1912 17592 1964
rect 17644 1912 17650 1964
rect 17862 1912 17868 1964
rect 17920 1912 17926 1964
rect 18046 1912 18052 1964
rect 18104 1912 18110 1964
rect 18322 1912 18328 1964
rect 18380 1912 18386 1964
rect 18414 1912 18420 1964
rect 18472 1912 18478 1964
rect 18693 1955 18751 1961
rect 18693 1921 18705 1955
rect 18739 1921 18751 1955
rect 18693 1915 18751 1921
rect 17880 1884 17908 1912
rect 15948 1856 17908 1884
rect 14976 1844 14982 1856
rect 17954 1844 17960 1896
rect 18012 1884 18018 1896
rect 18708 1884 18736 1915
rect 19150 1912 19156 1964
rect 19208 1912 19214 1964
rect 19536 1961 19564 1992
rect 19429 1955 19487 1961
rect 19429 1952 19441 1955
rect 19306 1924 19441 1952
rect 18012 1856 18736 1884
rect 18012 1844 18018 1856
rect 18782 1844 18788 1896
rect 18840 1884 18846 1896
rect 19306 1884 19334 1924
rect 19429 1921 19441 1924
rect 19475 1921 19487 1955
rect 19429 1915 19487 1921
rect 19521 1955 19579 1961
rect 19521 1921 19533 1955
rect 19567 1921 19579 1955
rect 19521 1915 19579 1921
rect 18840 1856 19334 1884
rect 20088 1884 20116 2060
rect 20180 2060 20536 2088
rect 20180 2029 20208 2060
rect 20530 2048 20536 2060
rect 20588 2048 20594 2100
rect 20625 2091 20683 2097
rect 20625 2057 20637 2091
rect 20671 2088 20683 2091
rect 23017 2091 23075 2097
rect 20671 2060 21680 2088
rect 20671 2057 20683 2060
rect 20625 2051 20683 2057
rect 20165 2023 20223 2029
rect 20165 1989 20177 2023
rect 20211 1989 20223 2023
rect 20165 1983 20223 1989
rect 20438 1980 20444 2032
rect 20496 2020 20502 2032
rect 21269 2023 21327 2029
rect 21269 2020 21281 2023
rect 20496 1992 21281 2020
rect 20496 1980 20502 1992
rect 21269 1989 21281 1992
rect 21315 1989 21327 2023
rect 21269 1983 21327 1989
rect 20806 1912 20812 1964
rect 20864 1912 20870 1964
rect 20898 1912 20904 1964
rect 20956 1952 20962 1964
rect 21085 1955 21143 1961
rect 21085 1952 21097 1955
rect 20956 1924 21097 1952
rect 20956 1912 20962 1924
rect 21085 1921 21097 1924
rect 21131 1921 21143 1955
rect 21652 1952 21680 2060
rect 23017 2057 23029 2091
rect 23063 2088 23075 2091
rect 23106 2088 23112 2100
rect 23063 2060 23112 2088
rect 23063 2057 23075 2060
rect 23017 2051 23075 2057
rect 23106 2048 23112 2060
rect 23164 2048 23170 2100
rect 23566 2048 23572 2100
rect 23624 2088 23630 2100
rect 23845 2091 23903 2097
rect 23845 2088 23857 2091
rect 23624 2060 23857 2088
rect 23624 2048 23630 2060
rect 23845 2057 23857 2060
rect 23891 2057 23903 2091
rect 23845 2051 23903 2057
rect 23934 2048 23940 2100
rect 23992 2088 23998 2100
rect 24673 2091 24731 2097
rect 23992 2060 24440 2088
rect 23992 2048 23998 2060
rect 22097 1955 22155 1961
rect 22097 1952 22109 1955
rect 21652 1924 22109 1952
rect 21085 1915 21143 1921
rect 22097 1921 22109 1924
rect 22143 1921 22155 1955
rect 22097 1915 22155 1921
rect 22922 1912 22928 1964
rect 22980 1912 22986 1964
rect 23201 1955 23259 1961
rect 23201 1921 23213 1955
rect 23247 1952 23259 1955
rect 23382 1952 23388 1964
rect 23247 1924 23388 1952
rect 23247 1921 23259 1924
rect 23201 1915 23259 1921
rect 23382 1912 23388 1924
rect 23440 1912 23446 1964
rect 23474 1912 23480 1964
rect 23532 1912 23538 1964
rect 23750 1912 23756 1964
rect 23808 1912 23814 1964
rect 24029 1955 24087 1961
rect 24029 1921 24041 1955
rect 24075 1952 24087 1955
rect 24210 1952 24216 1964
rect 24075 1924 24216 1952
rect 24075 1921 24087 1924
rect 24029 1915 24087 1921
rect 24210 1912 24216 1924
rect 24268 1912 24274 1964
rect 24302 1912 24308 1964
rect 24360 1912 24366 1964
rect 24412 1952 24440 2060
rect 24673 2057 24685 2091
rect 24719 2088 24731 2091
rect 24762 2088 24768 2100
rect 24719 2060 24768 2088
rect 24719 2057 24731 2060
rect 24673 2051 24731 2057
rect 24762 2048 24768 2060
rect 24820 2048 24826 2100
rect 25590 2048 25596 2100
rect 25648 2088 25654 2100
rect 25648 2060 26004 2088
rect 25648 2048 25654 2060
rect 25976 2029 26004 2060
rect 26694 2048 26700 2100
rect 26752 2088 26758 2100
rect 27982 2088 27988 2100
rect 26752 2060 27016 2088
rect 26752 2048 26758 2060
rect 25409 2023 25467 2029
rect 25409 2020 25421 2023
rect 25056 1992 25421 2020
rect 24581 1955 24639 1961
rect 24581 1952 24593 1955
rect 24412 1924 24593 1952
rect 24581 1921 24593 1924
rect 24627 1921 24639 1955
rect 24581 1915 24639 1921
rect 24670 1912 24676 1964
rect 24728 1952 24734 1964
rect 24857 1955 24915 1961
rect 24857 1952 24869 1955
rect 24728 1924 24869 1952
rect 24728 1912 24734 1924
rect 24857 1921 24869 1924
rect 24903 1921 24915 1955
rect 24857 1915 24915 1921
rect 24946 1912 24952 1964
rect 25004 1952 25010 1964
rect 25056 1952 25084 1992
rect 25409 1989 25421 1992
rect 25455 1989 25467 2023
rect 25409 1983 25467 1989
rect 25961 2023 26019 2029
rect 25961 1989 25973 2023
rect 26007 1989 26019 2023
rect 25961 1983 26019 1989
rect 26050 1980 26056 2032
rect 26108 2020 26114 2032
rect 26108 1992 26832 2020
rect 26108 1980 26114 1992
rect 25004 1924 25084 1952
rect 25133 1955 25191 1961
rect 25004 1912 25010 1924
rect 25133 1921 25145 1955
rect 25179 1921 25191 1955
rect 25133 1915 25191 1921
rect 25148 1884 25176 1915
rect 25222 1912 25228 1964
rect 25280 1952 25286 1964
rect 26602 1952 26608 1964
rect 25280 1924 26608 1952
rect 25280 1912 25286 1924
rect 26602 1912 26608 1924
rect 26660 1912 26666 1964
rect 26804 1961 26832 1992
rect 26789 1955 26847 1961
rect 26789 1921 26801 1955
rect 26835 1921 26847 1955
rect 26988 1952 27016 2060
rect 27080 2060 27988 2088
rect 27080 2029 27108 2060
rect 27982 2048 27988 2060
rect 28040 2048 28046 2100
rect 28902 2048 28908 2100
rect 28960 2088 28966 2100
rect 28960 2048 28994 2088
rect 29822 2048 29828 2100
rect 29880 2048 29886 2100
rect 30190 2048 30196 2100
rect 30248 2088 30254 2100
rect 30248 2060 31754 2088
rect 30248 2048 30254 2060
rect 27065 2023 27123 2029
rect 27065 1989 27077 2023
rect 27111 1989 27123 2023
rect 28169 2023 28227 2029
rect 28169 2020 28181 2023
rect 27065 1983 27123 1989
rect 27448 1992 28181 2020
rect 27448 1952 27476 1992
rect 28169 1989 28181 1992
rect 28215 1989 28227 2023
rect 28169 1983 28227 1989
rect 28626 1980 28632 2032
rect 28684 2020 28690 2032
rect 28813 2023 28871 2029
rect 28813 2020 28825 2023
rect 28684 1992 28825 2020
rect 28684 1980 28690 1992
rect 28813 1989 28825 1992
rect 28859 1989 28871 2023
rect 28966 2020 28994 2048
rect 29840 2020 29868 2048
rect 28966 1992 29408 2020
rect 29840 1992 30316 2020
rect 28813 1983 28871 1989
rect 26988 1924 27476 1952
rect 27617 1955 27675 1961
rect 26789 1915 26847 1921
rect 27617 1921 27629 1955
rect 27663 1952 27675 1955
rect 28350 1952 28356 1964
rect 27663 1924 28356 1952
rect 27663 1921 27675 1924
rect 27617 1915 27675 1921
rect 28350 1912 28356 1924
rect 28408 1912 28414 1964
rect 28442 1912 28448 1964
rect 28500 1952 28506 1964
rect 28902 1952 28908 1964
rect 28500 1924 28908 1952
rect 28500 1912 28506 1924
rect 28902 1912 28908 1924
rect 28960 1912 28966 1964
rect 28994 1912 29000 1964
rect 29052 1952 29058 1964
rect 29273 1955 29331 1961
rect 29273 1952 29285 1955
rect 29052 1924 29285 1952
rect 29052 1912 29058 1924
rect 29273 1921 29285 1924
rect 29319 1921 29331 1955
rect 29380 1952 29408 1992
rect 30288 1961 30316 1992
rect 30374 1980 30380 2032
rect 30432 2020 30438 2032
rect 31726 2020 31754 2060
rect 31846 2048 31852 2100
rect 31904 2088 31910 2100
rect 31904 2060 32812 2088
rect 31904 2048 31910 2060
rect 32784 2029 32812 2060
rect 33686 2048 33692 2100
rect 33744 2088 33750 2100
rect 33744 2060 35664 2088
rect 33744 2048 33750 2060
rect 32217 2023 32275 2029
rect 32217 2020 32229 2023
rect 30432 1992 31616 2020
rect 31726 1992 32229 2020
rect 30432 1980 30438 1992
rect 29825 1955 29883 1961
rect 29825 1952 29837 1955
rect 29380 1924 29837 1952
rect 29273 1915 29331 1921
rect 29825 1921 29837 1924
rect 29871 1921 29883 1955
rect 29825 1915 29883 1921
rect 30285 1955 30343 1961
rect 30285 1921 30297 1955
rect 30331 1921 30343 1955
rect 30285 1915 30343 1921
rect 30742 1912 30748 1964
rect 30800 1952 30806 1964
rect 30929 1955 30987 1961
rect 30929 1952 30941 1955
rect 30800 1924 30941 1952
rect 30800 1912 30806 1924
rect 30929 1921 30941 1924
rect 30975 1921 30987 1955
rect 31481 1955 31539 1961
rect 31481 1952 31493 1955
rect 30929 1915 30987 1921
rect 31036 1924 31493 1952
rect 25314 1884 25320 1896
rect 20088 1856 22968 1884
rect 18840 1844 18846 1856
rect 17402 1816 17408 1828
rect 13924 1788 17408 1816
rect 13924 1757 13952 1788
rect 17402 1776 17408 1788
rect 17460 1776 17466 1828
rect 17497 1819 17555 1825
rect 17497 1785 17509 1819
rect 17543 1816 17555 1819
rect 18230 1816 18236 1828
rect 17543 1788 18236 1816
rect 17543 1785 17555 1788
rect 17497 1779 17555 1785
rect 18230 1776 18236 1788
rect 18288 1776 18294 1828
rect 18601 1819 18659 1825
rect 18601 1785 18613 1819
rect 18647 1816 18659 1819
rect 22741 1819 22799 1825
rect 18647 1788 22692 1816
rect 18647 1785 18659 1788
rect 18601 1779 18659 1785
rect 13909 1751 13967 1757
rect 13909 1717 13921 1751
rect 13955 1717 13967 1751
rect 13909 1711 13967 1717
rect 14921 1751 14979 1757
rect 14921 1717 14933 1751
rect 14967 1748 14979 1751
rect 16574 1748 16580 1760
rect 14967 1720 16580 1748
rect 14967 1717 14979 1720
rect 14921 1711 14979 1717
rect 16574 1708 16580 1720
rect 16632 1708 16638 1760
rect 17773 1751 17831 1757
rect 17773 1717 17785 1751
rect 17819 1748 17831 1751
rect 18506 1748 18512 1760
rect 17819 1720 18512 1748
rect 17819 1717 17831 1720
rect 17773 1711 17831 1717
rect 18506 1708 18512 1720
rect 18564 1708 18570 1760
rect 18874 1708 18880 1760
rect 18932 1708 18938 1760
rect 19245 1751 19303 1757
rect 19245 1717 19257 1751
rect 19291 1748 19303 1751
rect 19610 1748 19616 1760
rect 19291 1720 19616 1748
rect 19291 1717 19303 1720
rect 19245 1711 19303 1717
rect 19610 1708 19616 1720
rect 19668 1708 19674 1760
rect 19702 1708 19708 1760
rect 19760 1708 19766 1760
rect 19978 1708 19984 1760
rect 20036 1748 20042 1760
rect 20257 1751 20315 1757
rect 20257 1748 20269 1751
rect 20036 1720 20269 1748
rect 20036 1708 20042 1720
rect 20257 1717 20269 1720
rect 20303 1717 20315 1751
rect 20257 1711 20315 1717
rect 20898 1708 20904 1760
rect 20956 1708 20962 1760
rect 21082 1708 21088 1760
rect 21140 1748 21146 1760
rect 21361 1751 21419 1757
rect 21361 1748 21373 1751
rect 21140 1720 21373 1748
rect 21140 1708 21146 1720
rect 21361 1717 21373 1720
rect 21407 1717 21419 1751
rect 21361 1711 21419 1717
rect 21910 1708 21916 1760
rect 21968 1748 21974 1760
rect 22189 1751 22247 1757
rect 22189 1748 22201 1751
rect 21968 1720 22201 1748
rect 21968 1708 21974 1720
rect 22189 1717 22201 1720
rect 22235 1717 22247 1751
rect 22664 1748 22692 1788
rect 22741 1785 22753 1819
rect 22787 1816 22799 1819
rect 22830 1816 22836 1828
rect 22787 1788 22836 1816
rect 22787 1785 22799 1788
rect 22741 1779 22799 1785
rect 22830 1776 22836 1788
rect 22888 1776 22894 1828
rect 22940 1816 22968 1856
rect 23308 1856 24900 1884
rect 25148 1856 25320 1884
rect 23014 1816 23020 1828
rect 22940 1788 23020 1816
rect 23014 1776 23020 1788
rect 23072 1776 23078 1828
rect 23308 1816 23336 1856
rect 24872 1828 24900 1856
rect 25314 1844 25320 1856
rect 25372 1844 25378 1896
rect 26326 1844 26332 1896
rect 26384 1884 26390 1896
rect 27341 1887 27399 1893
rect 27341 1884 27353 1887
rect 26384 1856 27353 1884
rect 26384 1844 26390 1856
rect 27341 1853 27353 1856
rect 27387 1853 27399 1887
rect 27341 1847 27399 1853
rect 27430 1844 27436 1896
rect 27488 1884 27494 1896
rect 31036 1884 31064 1924
rect 31481 1921 31493 1924
rect 31527 1921 31539 1955
rect 31588 1952 31616 1992
rect 32217 1989 32229 1992
rect 32263 1989 32275 2023
rect 32217 1983 32275 1989
rect 32769 2023 32827 2029
rect 32769 1989 32781 2023
rect 32815 1989 32827 2023
rect 32769 1983 32827 1989
rect 33318 1980 33324 2032
rect 33376 1980 33382 2032
rect 34146 1980 34152 2032
rect 34204 2020 34210 2032
rect 34425 2023 34483 2029
rect 34425 2020 34437 2023
rect 34204 1992 34437 2020
rect 34204 1980 34210 1992
rect 34425 1989 34437 1992
rect 34471 1989 34483 2023
rect 35636 2020 35664 2060
rect 36538 2048 36544 2100
rect 36596 2088 36602 2100
rect 37277 2091 37335 2097
rect 37277 2088 37289 2091
rect 36596 2060 37289 2088
rect 36596 2048 36602 2060
rect 37277 2057 37289 2060
rect 37323 2057 37335 2091
rect 37277 2051 37335 2057
rect 37553 2091 37611 2097
rect 37553 2057 37565 2091
rect 37599 2057 37611 2091
rect 37553 2051 37611 2057
rect 37568 2020 37596 2051
rect 37918 2048 37924 2100
rect 37976 2088 37982 2100
rect 38105 2091 38163 2097
rect 38105 2088 38117 2091
rect 37976 2060 38117 2088
rect 37976 2048 37982 2060
rect 38105 2057 38117 2060
rect 38151 2057 38163 2091
rect 38105 2051 38163 2057
rect 38749 2091 38807 2097
rect 38749 2057 38761 2091
rect 38795 2088 38807 2091
rect 39666 2088 39672 2100
rect 38795 2060 39672 2088
rect 38795 2057 38807 2060
rect 38749 2051 38807 2057
rect 39666 2048 39672 2060
rect 39724 2048 39730 2100
rect 39945 2091 40003 2097
rect 39945 2057 39957 2091
rect 39991 2088 40003 2091
rect 40862 2088 40868 2100
rect 39991 2060 40868 2088
rect 39991 2057 40003 2060
rect 39945 2051 40003 2057
rect 40862 2048 40868 2060
rect 40920 2048 40926 2100
rect 42426 2048 42432 2100
rect 42484 2048 42490 2100
rect 35636 1992 37596 2020
rect 34425 1983 34483 1989
rect 33873 1955 33931 1961
rect 31588 1924 32720 1952
rect 31481 1915 31539 1921
rect 27488 1856 31064 1884
rect 27488 1844 27494 1856
rect 31202 1844 31208 1896
rect 31260 1884 31266 1896
rect 32692 1884 32720 1924
rect 33873 1921 33885 1955
rect 33919 1921 33931 1955
rect 33873 1915 33931 1921
rect 33888 1884 33916 1915
rect 34882 1912 34888 1964
rect 34940 1912 34946 1964
rect 36354 1912 36360 1964
rect 36412 1912 36418 1964
rect 37461 1955 37519 1961
rect 37461 1921 37473 1955
rect 37507 1921 37519 1955
rect 37461 1915 37519 1921
rect 37737 1955 37795 1961
rect 37737 1921 37749 1955
rect 37783 1921 37795 1955
rect 37737 1915 37795 1921
rect 38289 1955 38347 1961
rect 38289 1921 38301 1955
rect 38335 1921 38347 1955
rect 38289 1915 38347 1921
rect 38933 1955 38991 1961
rect 38933 1921 38945 1955
rect 38979 1952 38991 1955
rect 40034 1952 40040 1964
rect 38979 1924 40040 1952
rect 38979 1921 38991 1924
rect 38933 1915 38991 1921
rect 31260 1856 31892 1884
rect 32692 1856 33916 1884
rect 31260 1844 31266 1856
rect 24762 1816 24768 1828
rect 23216 1788 23336 1816
rect 23492 1788 24768 1816
rect 23216 1748 23244 1788
rect 22664 1720 23244 1748
rect 23293 1751 23351 1757
rect 22189 1711 22247 1717
rect 23293 1717 23305 1751
rect 23339 1748 23351 1751
rect 23492 1748 23520 1788
rect 24762 1776 24768 1788
rect 24820 1776 24826 1828
rect 24854 1776 24860 1828
rect 24912 1776 24918 1828
rect 24949 1819 25007 1825
rect 24949 1785 24961 1819
rect 24995 1816 25007 1819
rect 27154 1816 27160 1828
rect 24995 1788 27160 1816
rect 24995 1785 25007 1788
rect 24949 1779 25007 1785
rect 27154 1776 27160 1788
rect 27212 1776 27218 1828
rect 28350 1776 28356 1828
rect 28408 1776 28414 1828
rect 28626 1776 28632 1828
rect 28684 1816 28690 1828
rect 28997 1819 29055 1825
rect 28997 1816 29009 1819
rect 28684 1788 29009 1816
rect 28684 1776 28690 1788
rect 28997 1785 29009 1788
rect 29043 1785 29055 1819
rect 28997 1779 29055 1785
rect 29362 1776 29368 1828
rect 29420 1816 29426 1828
rect 29420 1788 30512 1816
rect 29420 1776 29426 1788
rect 23339 1720 23520 1748
rect 23569 1751 23627 1757
rect 23339 1717 23351 1720
rect 23293 1711 23351 1717
rect 23569 1717 23581 1751
rect 23615 1748 23627 1751
rect 24026 1748 24032 1760
rect 23615 1720 24032 1748
rect 23615 1717 23627 1720
rect 23569 1711 23627 1717
rect 24026 1708 24032 1720
rect 24084 1708 24090 1760
rect 24118 1708 24124 1760
rect 24176 1708 24182 1760
rect 24397 1751 24455 1757
rect 24397 1717 24409 1751
rect 24443 1748 24455 1751
rect 24670 1748 24676 1760
rect 24443 1720 24676 1748
rect 24443 1717 24455 1720
rect 24397 1711 24455 1717
rect 24670 1708 24676 1720
rect 24728 1708 24734 1760
rect 25222 1708 25228 1760
rect 25280 1748 25286 1760
rect 25501 1751 25559 1757
rect 25501 1748 25513 1751
rect 25280 1720 25513 1748
rect 25280 1708 25286 1720
rect 25501 1717 25513 1720
rect 25547 1717 25559 1751
rect 25501 1711 25559 1717
rect 25866 1708 25872 1760
rect 25924 1748 25930 1760
rect 26237 1751 26295 1757
rect 26237 1748 26249 1751
rect 25924 1720 26249 1748
rect 25924 1708 25930 1720
rect 26237 1717 26249 1720
rect 26283 1717 26295 1751
rect 26237 1711 26295 1717
rect 26602 1708 26608 1760
rect 26660 1708 26666 1760
rect 27430 1708 27436 1760
rect 27488 1748 27494 1760
rect 27709 1751 27767 1757
rect 27709 1748 27721 1751
rect 27488 1720 27721 1748
rect 27488 1708 27494 1720
rect 27709 1717 27721 1720
rect 27755 1717 27767 1751
rect 27709 1711 27767 1717
rect 28166 1708 28172 1760
rect 28224 1748 28230 1760
rect 29457 1751 29515 1757
rect 29457 1748 29469 1751
rect 28224 1720 29469 1748
rect 28224 1708 28230 1720
rect 29457 1717 29469 1720
rect 29503 1717 29515 1751
rect 29457 1711 29515 1717
rect 29638 1708 29644 1760
rect 29696 1748 29702 1760
rect 30484 1757 30512 1788
rect 29917 1751 29975 1757
rect 29917 1748 29929 1751
rect 29696 1720 29929 1748
rect 29696 1708 29702 1720
rect 29917 1717 29929 1720
rect 29963 1717 29975 1751
rect 29917 1711 29975 1717
rect 30469 1751 30527 1757
rect 30469 1717 30481 1751
rect 30515 1717 30527 1751
rect 30469 1711 30527 1717
rect 31018 1708 31024 1760
rect 31076 1708 31082 1760
rect 31294 1708 31300 1760
rect 31352 1748 31358 1760
rect 31757 1751 31815 1757
rect 31757 1748 31769 1751
rect 31352 1720 31769 1748
rect 31352 1708 31358 1720
rect 31757 1717 31769 1720
rect 31803 1717 31815 1751
rect 31864 1748 31892 1856
rect 31938 1776 31944 1828
rect 31996 1816 32002 1828
rect 33042 1816 33048 1828
rect 31996 1788 33048 1816
rect 31996 1776 32002 1788
rect 33042 1776 33048 1788
rect 33100 1776 33106 1828
rect 33318 1776 33324 1828
rect 33376 1816 33382 1828
rect 33376 1788 35112 1816
rect 33376 1776 33382 1788
rect 32309 1751 32367 1757
rect 32309 1748 32321 1751
rect 31864 1720 32321 1748
rect 31757 1711 31815 1717
rect 32309 1717 32321 1720
rect 32355 1717 32367 1751
rect 32309 1711 32367 1717
rect 32398 1708 32404 1760
rect 32456 1748 32462 1760
rect 32861 1751 32919 1757
rect 32861 1748 32873 1751
rect 32456 1720 32873 1748
rect 32456 1708 32462 1720
rect 32861 1717 32873 1720
rect 32907 1717 32919 1751
rect 32861 1711 32919 1717
rect 32950 1708 32956 1760
rect 33008 1748 33014 1760
rect 33413 1751 33471 1757
rect 33413 1748 33425 1751
rect 33008 1720 33425 1748
rect 33008 1708 33014 1720
rect 33413 1717 33425 1720
rect 33459 1717 33471 1751
rect 33413 1711 33471 1717
rect 33502 1708 33508 1760
rect 33560 1748 33566 1760
rect 33965 1751 34023 1757
rect 33965 1748 33977 1751
rect 33560 1720 33977 1748
rect 33560 1708 33566 1720
rect 33965 1717 33977 1720
rect 34011 1717 34023 1751
rect 33965 1711 34023 1717
rect 34514 1708 34520 1760
rect 34572 1708 34578 1760
rect 35084 1757 35112 1788
rect 36538 1776 36544 1828
rect 36596 1776 36602 1828
rect 35069 1751 35127 1757
rect 35069 1717 35081 1751
rect 35115 1717 35127 1751
rect 37476 1748 37504 1915
rect 37752 1816 37780 1915
rect 38304 1884 38332 1915
rect 40034 1912 40040 1924
rect 40092 1912 40098 1964
rect 40126 1912 40132 1964
rect 40184 1912 40190 1964
rect 41049 1955 41107 1961
rect 41049 1921 41061 1955
rect 41095 1952 41107 1955
rect 41506 1952 41512 1964
rect 41095 1924 41512 1952
rect 41095 1921 41107 1924
rect 41049 1915 41107 1921
rect 41506 1912 41512 1924
rect 41564 1912 41570 1964
rect 40678 1884 40684 1896
rect 38304 1856 40684 1884
rect 40678 1844 40684 1856
rect 40736 1844 40742 1896
rect 39758 1816 39764 1828
rect 37752 1788 39764 1816
rect 39758 1776 39764 1788
rect 39816 1776 39822 1828
rect 40865 1819 40923 1825
rect 40865 1785 40877 1819
rect 40911 1816 40923 1819
rect 42444 1816 42472 2048
rect 40911 1788 42472 1816
rect 40911 1785 40923 1788
rect 40865 1779 40923 1785
rect 39942 1748 39948 1760
rect 37476 1720 39948 1748
rect 35069 1711 35127 1717
rect 39942 1708 39948 1720
rect 40000 1708 40006 1760
rect 1104 1658 43884 1680
rect 1104 1606 6297 1658
rect 6349 1606 6361 1658
rect 6413 1606 6425 1658
rect 6477 1606 6489 1658
rect 6541 1606 6553 1658
rect 6605 1606 16991 1658
rect 17043 1606 17055 1658
rect 17107 1606 17119 1658
rect 17171 1606 17183 1658
rect 17235 1606 17247 1658
rect 17299 1606 27685 1658
rect 27737 1606 27749 1658
rect 27801 1606 27813 1658
rect 27865 1606 27877 1658
rect 27929 1606 27941 1658
rect 27993 1606 38379 1658
rect 38431 1606 38443 1658
rect 38495 1606 38507 1658
rect 38559 1606 38571 1658
rect 38623 1606 38635 1658
rect 38687 1606 43884 1658
rect 1104 1584 43884 1606
rect 6822 1504 6828 1556
rect 6880 1504 6886 1556
rect 7929 1547 7987 1553
rect 7929 1513 7941 1547
rect 7975 1544 7987 1547
rect 8478 1544 8484 1556
rect 7975 1516 8484 1544
rect 7975 1513 7987 1516
rect 7929 1507 7987 1513
rect 8478 1504 8484 1516
rect 8536 1504 8542 1556
rect 9401 1547 9459 1553
rect 9401 1513 9413 1547
rect 9447 1544 9459 1547
rect 10410 1544 10416 1556
rect 9447 1516 10416 1544
rect 9447 1513 9459 1516
rect 9401 1507 9459 1513
rect 10410 1504 10416 1516
rect 10468 1504 10474 1556
rect 10778 1504 10784 1556
rect 10836 1504 10842 1556
rect 11974 1504 11980 1556
rect 12032 1504 12038 1556
rect 12250 1504 12256 1556
rect 12308 1504 12314 1556
rect 13906 1504 13912 1556
rect 13964 1504 13970 1556
rect 14642 1504 14648 1556
rect 14700 1504 14706 1556
rect 14918 1504 14924 1556
rect 14976 1504 14982 1556
rect 15197 1547 15255 1553
rect 15197 1513 15209 1547
rect 15243 1544 15255 1547
rect 15746 1544 15752 1556
rect 15243 1516 15752 1544
rect 15243 1513 15255 1516
rect 15197 1507 15255 1513
rect 15746 1504 15752 1516
rect 15804 1504 15810 1556
rect 16025 1547 16083 1553
rect 16025 1513 16037 1547
rect 16071 1544 16083 1547
rect 16390 1544 16396 1556
rect 16071 1516 16396 1544
rect 16071 1513 16083 1516
rect 16025 1507 16083 1513
rect 16390 1504 16396 1516
rect 16448 1504 16454 1556
rect 16850 1544 16856 1556
rect 16592 1516 16856 1544
rect 7377 1479 7435 1485
rect 7377 1445 7389 1479
rect 7423 1476 7435 1479
rect 8294 1476 8300 1488
rect 7423 1448 8300 1476
rect 7423 1445 7435 1448
rect 7377 1439 7435 1445
rect 8294 1436 8300 1448
rect 8352 1436 8358 1488
rect 9674 1436 9680 1488
rect 9732 1436 9738 1488
rect 9950 1436 9956 1488
rect 10008 1436 10014 1488
rect 10226 1436 10232 1488
rect 10284 1436 10290 1488
rect 14369 1479 14427 1485
rect 14369 1445 14381 1479
rect 14415 1476 14427 1479
rect 15286 1476 15292 1488
rect 14415 1448 15292 1476
rect 14415 1445 14427 1448
rect 14369 1439 14427 1445
rect 15286 1436 15292 1448
rect 15344 1436 15350 1488
rect 15473 1479 15531 1485
rect 15473 1445 15485 1479
rect 15519 1476 15531 1479
rect 16301 1479 16359 1485
rect 15519 1448 15884 1476
rect 15519 1445 15531 1448
rect 15473 1439 15531 1445
rect 8110 1408 8116 1420
rect 7392 1380 7604 1408
rect 4890 1300 4896 1352
rect 4948 1300 4954 1352
rect 5169 1343 5227 1349
rect 5169 1309 5181 1343
rect 5215 1309 5227 1343
rect 5169 1303 5227 1309
rect 5445 1343 5503 1349
rect 5445 1309 5457 1343
rect 5491 1340 5503 1343
rect 5626 1340 5632 1352
rect 5491 1312 5632 1340
rect 5491 1309 5503 1312
rect 5445 1303 5503 1309
rect 5184 1272 5212 1303
rect 5626 1300 5632 1312
rect 5684 1300 5690 1352
rect 5721 1343 5779 1349
rect 5721 1309 5733 1343
rect 5767 1340 5779 1343
rect 5902 1340 5908 1352
rect 5767 1312 5908 1340
rect 5767 1309 5779 1312
rect 5721 1303 5779 1309
rect 5902 1300 5908 1312
rect 5960 1300 5966 1352
rect 5994 1300 6000 1352
rect 6052 1300 6058 1352
rect 6365 1343 6423 1349
rect 6365 1309 6377 1343
rect 6411 1309 6423 1343
rect 6365 1303 6423 1309
rect 6641 1343 6699 1349
rect 6641 1309 6653 1343
rect 6687 1340 6699 1343
rect 6822 1340 6828 1352
rect 6687 1312 6828 1340
rect 6687 1309 6699 1312
rect 6641 1303 6699 1309
rect 5534 1272 5540 1284
rect 5184 1244 5540 1272
rect 5534 1232 5540 1244
rect 5592 1232 5598 1284
rect 6380 1272 6408 1303
rect 6822 1300 6828 1312
rect 6880 1300 6886 1352
rect 6917 1343 6975 1349
rect 6917 1309 6929 1343
rect 6963 1340 6975 1343
rect 7193 1343 7251 1349
rect 6963 1312 7144 1340
rect 6963 1309 6975 1312
rect 6917 1303 6975 1309
rect 7006 1272 7012 1284
rect 6380 1244 7012 1272
rect 7006 1232 7012 1244
rect 7064 1232 7070 1284
rect 7116 1272 7144 1312
rect 7193 1309 7205 1343
rect 7239 1340 7251 1343
rect 7392 1340 7420 1380
rect 7239 1312 7420 1340
rect 7239 1309 7251 1312
rect 7193 1303 7251 1309
rect 7466 1300 7472 1352
rect 7524 1300 7530 1352
rect 7576 1340 7604 1380
rect 7944 1380 8116 1408
rect 7650 1340 7656 1352
rect 7576 1312 7656 1340
rect 7650 1300 7656 1312
rect 7708 1300 7714 1352
rect 7745 1343 7803 1349
rect 7745 1309 7757 1343
rect 7791 1340 7803 1343
rect 7944 1340 7972 1380
rect 8110 1368 8116 1380
rect 8168 1368 8174 1420
rect 14274 1408 14280 1420
rect 8864 1380 9076 1408
rect 7791 1312 7972 1340
rect 8021 1343 8079 1349
rect 7791 1309 7803 1312
rect 7745 1303 7803 1309
rect 8021 1309 8033 1343
rect 8067 1309 8079 1343
rect 8021 1303 8079 1309
rect 8297 1343 8355 1349
rect 8297 1309 8309 1343
rect 8343 1340 8355 1343
rect 8573 1343 8631 1349
rect 8343 1312 8524 1340
rect 8343 1309 8355 1312
rect 8297 1303 8355 1309
rect 7558 1272 7564 1284
rect 7116 1244 7564 1272
rect 7558 1232 7564 1244
rect 7616 1232 7622 1284
rect 8036 1272 8064 1303
rect 8386 1272 8392 1284
rect 8036 1244 8392 1272
rect 8386 1232 8392 1244
rect 8444 1232 8450 1284
rect 8496 1272 8524 1312
rect 8573 1309 8585 1343
rect 8619 1340 8631 1343
rect 8864 1340 8892 1380
rect 9048 1352 9076 1380
rect 13832 1380 14280 1408
rect 8619 1312 8892 1340
rect 8941 1343 8999 1349
rect 8619 1309 8631 1312
rect 8573 1303 8631 1309
rect 8941 1309 8953 1343
rect 8987 1309 8999 1343
rect 8941 1303 8999 1309
rect 8846 1272 8852 1284
rect 8496 1244 8852 1272
rect 8846 1232 8852 1244
rect 8904 1232 8910 1284
rect 8956 1272 8984 1303
rect 9030 1300 9036 1352
rect 9088 1300 9094 1352
rect 9217 1343 9275 1349
rect 9217 1309 9229 1343
rect 9263 1340 9275 1343
rect 9493 1343 9551 1349
rect 9263 1312 9444 1340
rect 9263 1309 9275 1312
rect 9217 1303 9275 1309
rect 9306 1272 9312 1284
rect 8956 1244 9312 1272
rect 9306 1232 9312 1244
rect 9364 1232 9370 1284
rect 9416 1272 9444 1312
rect 9493 1309 9505 1343
rect 9539 1340 9551 1343
rect 9769 1343 9827 1349
rect 9539 1312 9720 1340
rect 9539 1309 9551 1312
rect 9493 1303 9551 1309
rect 9582 1272 9588 1284
rect 9416 1244 9588 1272
rect 9582 1232 9588 1244
rect 9640 1232 9646 1284
rect 9692 1272 9720 1312
rect 9769 1309 9781 1343
rect 9815 1340 9827 1343
rect 10045 1343 10103 1349
rect 9815 1312 9996 1340
rect 9815 1309 9827 1312
rect 9769 1303 9827 1309
rect 9858 1272 9864 1284
rect 9692 1244 9864 1272
rect 9858 1232 9864 1244
rect 9916 1232 9922 1284
rect 5074 1164 5080 1216
rect 5132 1164 5138 1216
rect 5350 1164 5356 1216
rect 5408 1164 5414 1216
rect 5626 1164 5632 1216
rect 5684 1164 5690 1216
rect 5905 1207 5963 1213
rect 5905 1173 5917 1207
rect 5951 1204 5963 1207
rect 6086 1204 6092 1216
rect 5951 1176 6092 1204
rect 5951 1173 5963 1176
rect 5905 1167 5963 1173
rect 6086 1164 6092 1176
rect 6144 1164 6150 1216
rect 6178 1164 6184 1216
rect 6236 1164 6242 1216
rect 6546 1164 6552 1216
rect 6604 1164 6610 1216
rect 7101 1207 7159 1213
rect 7101 1173 7113 1207
rect 7147 1204 7159 1207
rect 7374 1204 7380 1216
rect 7147 1176 7380 1204
rect 7147 1173 7159 1176
rect 7101 1167 7159 1173
rect 7374 1164 7380 1176
rect 7432 1164 7438 1216
rect 7653 1207 7711 1213
rect 7653 1173 7665 1207
rect 7699 1204 7711 1207
rect 7834 1204 7840 1216
rect 7699 1176 7840 1204
rect 7699 1173 7711 1176
rect 7653 1167 7711 1173
rect 7834 1164 7840 1176
rect 7892 1164 7898 1216
rect 8018 1164 8024 1216
rect 8076 1204 8082 1216
rect 8205 1207 8263 1213
rect 8205 1204 8217 1207
rect 8076 1176 8217 1204
rect 8076 1164 8082 1176
rect 8205 1173 8217 1176
rect 8251 1173 8263 1207
rect 8205 1167 8263 1173
rect 8481 1207 8539 1213
rect 8481 1173 8493 1207
rect 8527 1204 8539 1207
rect 8570 1204 8576 1216
rect 8527 1176 8576 1204
rect 8527 1173 8539 1176
rect 8481 1167 8539 1173
rect 8570 1164 8576 1176
rect 8628 1164 8634 1216
rect 8754 1164 8760 1216
rect 8812 1164 8818 1216
rect 9122 1164 9128 1216
rect 9180 1164 9186 1216
rect 9968 1204 9996 1312
rect 10045 1309 10057 1343
rect 10091 1309 10103 1343
rect 10045 1303 10103 1309
rect 10321 1343 10379 1349
rect 10321 1309 10333 1343
rect 10367 1340 10379 1343
rect 10367 1312 10548 1340
rect 10367 1309 10379 1312
rect 10321 1303 10379 1309
rect 10060 1272 10088 1303
rect 10410 1272 10416 1284
rect 10060 1244 10416 1272
rect 10410 1232 10416 1244
rect 10468 1232 10474 1284
rect 10520 1272 10548 1312
rect 10594 1300 10600 1352
rect 10652 1300 10658 1352
rect 10899 1343 10957 1349
rect 10899 1309 10911 1343
rect 10945 1340 10957 1343
rect 10945 1312 11100 1340
rect 10945 1309 10957 1312
rect 10899 1303 10957 1309
rect 10686 1272 10692 1284
rect 10520 1244 10692 1272
rect 10686 1232 10692 1244
rect 10744 1232 10750 1284
rect 11072 1272 11100 1312
rect 11146 1300 11152 1352
rect 11204 1300 11210 1352
rect 11517 1343 11575 1349
rect 11517 1309 11529 1343
rect 11563 1309 11575 1343
rect 11517 1303 11575 1309
rect 11793 1343 11851 1349
rect 11793 1309 11805 1343
rect 11839 1340 11851 1343
rect 12069 1343 12127 1349
rect 11839 1312 12020 1340
rect 11839 1309 11851 1312
rect 11793 1303 11851 1309
rect 11422 1272 11428 1284
rect 11072 1244 11428 1272
rect 11422 1232 11428 1244
rect 11480 1232 11486 1284
rect 11532 1272 11560 1303
rect 11882 1272 11888 1284
rect 11532 1244 11888 1272
rect 11882 1232 11888 1244
rect 11940 1232 11946 1284
rect 11992 1272 12020 1312
rect 12069 1309 12081 1343
rect 12115 1340 12127 1343
rect 12250 1340 12256 1352
rect 12115 1312 12256 1340
rect 12115 1309 12127 1312
rect 12069 1303 12127 1309
rect 12250 1300 12256 1312
rect 12308 1300 12314 1352
rect 12345 1343 12403 1349
rect 12345 1309 12357 1343
rect 12391 1340 12403 1343
rect 12434 1340 12440 1352
rect 12391 1312 12440 1340
rect 12391 1309 12403 1312
rect 12345 1303 12403 1309
rect 12434 1300 12440 1312
rect 12492 1300 12498 1352
rect 12526 1300 12532 1352
rect 12584 1300 12590 1352
rect 12621 1343 12679 1349
rect 12621 1309 12633 1343
rect 12667 1309 12679 1343
rect 12621 1303 12679 1309
rect 12897 1343 12955 1349
rect 12897 1309 12909 1343
rect 12943 1340 12955 1343
rect 13078 1340 13084 1352
rect 12943 1312 13084 1340
rect 12943 1309 12955 1312
rect 12897 1303 12955 1309
rect 12158 1272 12164 1284
rect 11992 1244 12164 1272
rect 12158 1232 12164 1244
rect 12216 1232 12222 1284
rect 10318 1204 10324 1216
rect 9968 1176 10324 1204
rect 10318 1164 10324 1176
rect 10376 1164 10382 1216
rect 10505 1207 10563 1213
rect 10505 1173 10517 1207
rect 10551 1204 10563 1207
rect 10962 1204 10968 1216
rect 10551 1176 10968 1204
rect 10551 1173 10563 1176
rect 10505 1167 10563 1173
rect 10962 1164 10968 1176
rect 11020 1164 11026 1216
rect 11057 1207 11115 1213
rect 11057 1173 11069 1207
rect 11103 1204 11115 1207
rect 11238 1204 11244 1216
rect 11103 1176 11244 1204
rect 11103 1173 11115 1176
rect 11057 1167 11115 1173
rect 11238 1164 11244 1176
rect 11296 1164 11302 1216
rect 11330 1164 11336 1216
rect 11388 1164 11394 1216
rect 11701 1207 11759 1213
rect 11701 1173 11713 1207
rect 11747 1204 11759 1207
rect 12066 1204 12072 1216
rect 11747 1176 12072 1204
rect 11747 1173 11759 1176
rect 11701 1167 11759 1173
rect 12066 1164 12072 1176
rect 12124 1164 12130 1216
rect 12544 1213 12572 1300
rect 12636 1272 12664 1303
rect 13078 1300 13084 1312
rect 13136 1300 13142 1352
rect 13173 1343 13231 1349
rect 13173 1309 13185 1343
rect 13219 1340 13231 1343
rect 13354 1340 13360 1352
rect 13219 1312 13360 1340
rect 13219 1309 13231 1312
rect 13173 1303 13231 1309
rect 13354 1300 13360 1312
rect 13412 1300 13418 1352
rect 13449 1343 13507 1349
rect 13449 1309 13461 1343
rect 13495 1309 13507 1343
rect 13449 1303 13507 1309
rect 13725 1343 13783 1349
rect 13725 1309 13737 1343
rect 13771 1340 13783 1343
rect 13832 1340 13860 1380
rect 14274 1368 14280 1380
rect 14332 1368 14338 1420
rect 15746 1408 15752 1420
rect 15212 1380 15752 1408
rect 13771 1312 13860 1340
rect 14093 1343 14151 1349
rect 13771 1309 13783 1312
rect 13725 1303 13783 1309
rect 14093 1309 14105 1343
rect 14139 1309 14151 1343
rect 14093 1303 14151 1309
rect 12986 1272 12992 1284
rect 12636 1244 12992 1272
rect 12986 1232 12992 1244
rect 13044 1232 13050 1284
rect 13464 1272 13492 1303
rect 13814 1272 13820 1284
rect 13464 1244 13820 1272
rect 13814 1232 13820 1244
rect 13872 1232 13878 1284
rect 14108 1272 14136 1303
rect 14550 1300 14556 1352
rect 14608 1300 14614 1352
rect 14829 1343 14887 1349
rect 14829 1309 14841 1343
rect 14875 1309 14887 1343
rect 14829 1303 14887 1309
rect 15105 1343 15163 1349
rect 15105 1309 15117 1343
rect 15151 1340 15163 1343
rect 15212 1340 15240 1380
rect 15746 1368 15752 1380
rect 15804 1368 15810 1420
rect 15856 1408 15884 1448
rect 16301 1445 16313 1479
rect 16347 1476 16359 1479
rect 16592 1476 16620 1516
rect 16850 1504 16856 1516
rect 16908 1504 16914 1556
rect 16945 1547 17003 1553
rect 16945 1513 16957 1547
rect 16991 1544 17003 1547
rect 17221 1547 17279 1553
rect 16991 1516 17172 1544
rect 16991 1513 17003 1516
rect 16945 1507 17003 1513
rect 16347 1448 16620 1476
rect 16347 1445 16359 1448
rect 16301 1439 16359 1445
rect 16574 1408 16580 1420
rect 15856 1380 16580 1408
rect 16574 1368 16580 1380
rect 16632 1368 16638 1420
rect 16942 1408 16948 1420
rect 16776 1380 16948 1408
rect 15151 1312 15240 1340
rect 15381 1343 15439 1349
rect 15151 1309 15163 1312
rect 15105 1303 15163 1309
rect 15381 1309 15393 1343
rect 15427 1309 15439 1343
rect 15381 1303 15439 1309
rect 14734 1272 14740 1284
rect 14108 1244 14740 1272
rect 14734 1232 14740 1244
rect 14792 1232 14798 1284
rect 14844 1272 14872 1303
rect 15286 1272 15292 1284
rect 14844 1244 15292 1272
rect 15286 1232 15292 1244
rect 15344 1232 15350 1284
rect 15396 1272 15424 1303
rect 15654 1300 15660 1352
rect 15712 1300 15718 1352
rect 15930 1300 15936 1352
rect 15988 1300 15994 1352
rect 16209 1343 16267 1349
rect 16209 1309 16221 1343
rect 16255 1309 16267 1343
rect 16209 1303 16267 1309
rect 16485 1343 16543 1349
rect 16485 1309 16497 1343
rect 16531 1340 16543 1343
rect 16776 1340 16804 1380
rect 16942 1368 16948 1380
rect 17000 1368 17006 1420
rect 17144 1408 17172 1516
rect 17221 1513 17233 1547
rect 17267 1544 17279 1547
rect 17586 1544 17592 1556
rect 17267 1516 17592 1544
rect 17267 1513 17279 1516
rect 17221 1507 17279 1513
rect 17586 1504 17592 1516
rect 17644 1504 17650 1556
rect 17773 1547 17831 1553
rect 17773 1513 17785 1547
rect 17819 1544 17831 1547
rect 18414 1544 18420 1556
rect 17819 1516 18420 1544
rect 17819 1513 17831 1516
rect 17773 1507 17831 1513
rect 18414 1504 18420 1516
rect 18472 1504 18478 1556
rect 18506 1504 18512 1556
rect 18564 1504 18570 1556
rect 18601 1547 18659 1553
rect 18601 1513 18613 1547
rect 18647 1544 18659 1547
rect 19150 1544 19156 1556
rect 18647 1516 19156 1544
rect 18647 1513 18659 1516
rect 18601 1507 18659 1513
rect 19150 1504 19156 1516
rect 19208 1504 19214 1556
rect 19812 1516 23244 1544
rect 17494 1436 17500 1488
rect 17552 1436 17558 1488
rect 18524 1476 18552 1504
rect 19812 1476 19840 1516
rect 17604 1448 18460 1476
rect 18524 1448 19840 1476
rect 17604 1408 17632 1448
rect 18046 1408 18052 1420
rect 17144 1380 17632 1408
rect 17880 1380 18052 1408
rect 16531 1312 16804 1340
rect 16853 1343 16911 1349
rect 16531 1309 16543 1312
rect 16485 1303 16543 1309
rect 16853 1309 16865 1343
rect 16899 1309 16911 1343
rect 16853 1303 16911 1309
rect 17129 1343 17187 1349
rect 17129 1309 17141 1343
rect 17175 1340 17187 1343
rect 17405 1343 17463 1349
rect 17175 1312 17356 1340
rect 17175 1309 17187 1312
rect 17129 1303 17187 1309
rect 16114 1272 16120 1284
rect 15396 1244 16120 1272
rect 16114 1232 16120 1244
rect 16172 1232 16178 1284
rect 16224 1272 16252 1303
rect 16574 1272 16580 1284
rect 16224 1244 16580 1272
rect 16574 1232 16580 1244
rect 16632 1232 16638 1284
rect 16868 1272 16896 1303
rect 17218 1272 17224 1284
rect 16868 1244 17224 1272
rect 17218 1232 17224 1244
rect 17276 1232 17282 1284
rect 12529 1207 12587 1213
rect 12529 1173 12541 1207
rect 12575 1173 12587 1207
rect 12529 1167 12587 1173
rect 12805 1207 12863 1213
rect 12805 1173 12817 1207
rect 12851 1204 12863 1207
rect 12894 1204 12900 1216
rect 12851 1176 12900 1204
rect 12851 1173 12863 1176
rect 12805 1167 12863 1173
rect 12894 1164 12900 1176
rect 12952 1164 12958 1216
rect 13081 1207 13139 1213
rect 13081 1173 13093 1207
rect 13127 1204 13139 1207
rect 13262 1204 13268 1216
rect 13127 1176 13268 1204
rect 13127 1173 13139 1176
rect 13081 1167 13139 1173
rect 13262 1164 13268 1176
rect 13320 1164 13326 1216
rect 13357 1207 13415 1213
rect 13357 1173 13369 1207
rect 13403 1204 13415 1207
rect 13446 1204 13452 1216
rect 13403 1176 13452 1204
rect 13403 1173 13415 1176
rect 13357 1167 13415 1173
rect 13446 1164 13452 1176
rect 13504 1164 13510 1216
rect 13538 1164 13544 1216
rect 13596 1204 13602 1216
rect 13633 1207 13691 1213
rect 13633 1204 13645 1207
rect 13596 1176 13645 1204
rect 13596 1164 13602 1176
rect 13633 1173 13645 1176
rect 13679 1173 13691 1207
rect 13633 1167 13691 1173
rect 14277 1207 14335 1213
rect 14277 1173 14289 1207
rect 14323 1204 14335 1207
rect 15562 1204 15568 1216
rect 14323 1176 15568 1204
rect 14323 1173 14335 1176
rect 14277 1167 14335 1173
rect 15562 1164 15568 1176
rect 15620 1164 15626 1216
rect 15749 1207 15807 1213
rect 15749 1173 15761 1207
rect 15795 1204 15807 1207
rect 16206 1204 16212 1216
rect 15795 1176 16212 1204
rect 15795 1173 15807 1176
rect 15749 1167 15807 1173
rect 16206 1164 16212 1176
rect 16264 1164 16270 1216
rect 16669 1207 16727 1213
rect 16669 1173 16681 1207
rect 16715 1204 16727 1207
rect 17126 1204 17132 1216
rect 16715 1176 17132 1204
rect 16715 1173 16727 1176
rect 16669 1167 16727 1173
rect 17126 1164 17132 1176
rect 17184 1164 17190 1216
rect 17328 1204 17356 1312
rect 17405 1309 17417 1343
rect 17451 1309 17463 1343
rect 17405 1303 17463 1309
rect 17681 1343 17739 1349
rect 17681 1309 17693 1343
rect 17727 1340 17739 1343
rect 17880 1340 17908 1380
rect 18046 1368 18052 1380
rect 18104 1368 18110 1420
rect 18432 1408 18460 1448
rect 19886 1436 19892 1488
rect 19944 1476 19950 1488
rect 19944 1448 20392 1476
rect 19944 1436 19950 1448
rect 18598 1408 18604 1420
rect 18156 1380 18368 1408
rect 18432 1380 18604 1408
rect 17727 1312 17908 1340
rect 17957 1343 18015 1349
rect 17727 1309 17739 1312
rect 17681 1303 17739 1309
rect 17957 1309 17969 1343
rect 18003 1340 18015 1343
rect 18156 1340 18184 1380
rect 18003 1312 18184 1340
rect 18233 1343 18291 1349
rect 18003 1309 18015 1312
rect 17957 1303 18015 1309
rect 18233 1309 18245 1343
rect 18279 1309 18291 1343
rect 18340 1340 18368 1380
rect 18598 1368 18604 1380
rect 18656 1368 18662 1420
rect 19150 1408 19156 1420
rect 18984 1380 19156 1408
rect 18414 1340 18420 1352
rect 18340 1312 18420 1340
rect 18233 1303 18291 1309
rect 17420 1272 17448 1303
rect 18138 1272 18144 1284
rect 17420 1244 18000 1272
rect 17972 1216 18000 1244
rect 18064 1244 18144 1272
rect 17402 1204 17408 1216
rect 17328 1176 17408 1204
rect 17402 1164 17408 1176
rect 17460 1164 17466 1216
rect 17954 1164 17960 1216
rect 18012 1164 18018 1216
rect 18064 1213 18092 1244
rect 18138 1232 18144 1244
rect 18196 1232 18202 1284
rect 18248 1216 18276 1303
rect 18414 1300 18420 1312
rect 18472 1300 18478 1352
rect 18506 1300 18512 1352
rect 18564 1300 18570 1352
rect 18785 1343 18843 1349
rect 18785 1309 18797 1343
rect 18831 1340 18843 1343
rect 18984 1340 19012 1380
rect 19150 1368 19156 1380
rect 19208 1368 19214 1420
rect 19628 1380 20300 1408
rect 19628 1352 19656 1380
rect 18831 1312 19012 1340
rect 18831 1309 18843 1312
rect 18785 1303 18843 1309
rect 19058 1300 19064 1352
rect 19116 1300 19122 1352
rect 19245 1343 19303 1349
rect 19245 1309 19257 1343
rect 19291 1309 19303 1343
rect 19245 1303 19303 1309
rect 19260 1272 19288 1303
rect 19518 1300 19524 1352
rect 19576 1300 19582 1352
rect 19610 1300 19616 1352
rect 19668 1300 19674 1352
rect 19794 1300 19800 1352
rect 19852 1340 19858 1352
rect 20272 1349 20300 1380
rect 19889 1343 19947 1349
rect 19889 1340 19901 1343
rect 19852 1312 19901 1340
rect 19852 1300 19858 1312
rect 19889 1309 19901 1312
rect 19935 1309 19947 1343
rect 19889 1303 19947 1309
rect 20257 1343 20315 1349
rect 20257 1309 20269 1343
rect 20303 1309 20315 1343
rect 20364 1340 20392 1448
rect 22278 1436 22284 1488
rect 22336 1436 22342 1488
rect 22830 1436 22836 1488
rect 22888 1476 22894 1488
rect 23216 1476 23244 1516
rect 23290 1504 23296 1556
rect 23348 1544 23354 1556
rect 23477 1547 23535 1553
rect 23477 1544 23489 1547
rect 23348 1516 23489 1544
rect 23348 1504 23354 1516
rect 23477 1513 23489 1516
rect 23523 1513 23535 1547
rect 23477 1507 23535 1513
rect 23584 1516 24256 1544
rect 23584 1476 23612 1516
rect 22888 1448 23152 1476
rect 23216 1448 23612 1476
rect 22888 1436 22894 1448
rect 22186 1368 22192 1420
rect 22244 1368 22250 1420
rect 22296 1408 22324 1436
rect 22296 1380 22968 1408
rect 20717 1343 20775 1349
rect 20717 1340 20729 1343
rect 20364 1312 20729 1340
rect 20257 1303 20315 1309
rect 20717 1309 20729 1312
rect 20763 1309 20775 1343
rect 20717 1303 20775 1309
rect 20898 1300 20904 1352
rect 20956 1300 20962 1352
rect 21266 1300 21272 1352
rect 21324 1340 21330 1352
rect 21361 1343 21419 1349
rect 21361 1340 21373 1343
rect 21324 1312 21373 1340
rect 21324 1300 21330 1312
rect 21361 1309 21373 1312
rect 21407 1309 21419 1343
rect 21361 1303 21419 1309
rect 22002 1300 22008 1352
rect 22060 1340 22066 1352
rect 22557 1343 22615 1349
rect 22557 1340 22569 1343
rect 22060 1312 22569 1340
rect 22060 1300 22066 1312
rect 22557 1309 22569 1312
rect 22603 1309 22615 1343
rect 22557 1303 22615 1309
rect 22738 1300 22744 1352
rect 22796 1300 22802 1352
rect 22940 1349 22968 1380
rect 22925 1343 22983 1349
rect 22925 1309 22937 1343
rect 22971 1309 22983 1343
rect 22925 1303 22983 1309
rect 20530 1272 20536 1284
rect 18340 1244 19288 1272
rect 19352 1244 20536 1272
rect 18049 1207 18107 1213
rect 18049 1173 18061 1207
rect 18095 1173 18107 1207
rect 18049 1167 18107 1173
rect 18230 1164 18236 1216
rect 18288 1164 18294 1216
rect 18340 1213 18368 1244
rect 18325 1207 18383 1213
rect 18325 1173 18337 1207
rect 18371 1173 18383 1207
rect 18325 1167 18383 1173
rect 18877 1207 18935 1213
rect 18877 1173 18889 1207
rect 18923 1204 18935 1207
rect 19352 1204 19380 1244
rect 20530 1232 20536 1244
rect 20588 1232 20594 1284
rect 20916 1272 20944 1300
rect 21913 1275 21971 1281
rect 21913 1272 21925 1275
rect 20916 1244 21925 1272
rect 21913 1241 21925 1244
rect 21959 1241 21971 1275
rect 22756 1272 22784 1300
rect 23124 1272 23152 1448
rect 23934 1436 23940 1488
rect 23992 1436 23998 1488
rect 24118 1436 24124 1488
rect 24176 1436 24182 1488
rect 24228 1476 24256 1516
rect 24302 1504 24308 1556
rect 24360 1544 24366 1556
rect 24949 1547 25007 1553
rect 24949 1544 24961 1547
rect 24360 1516 24961 1544
rect 24360 1504 24366 1516
rect 24949 1513 24961 1516
rect 24995 1513 25007 1547
rect 24949 1507 25007 1513
rect 25501 1547 25559 1553
rect 25501 1513 25513 1547
rect 25547 1513 25559 1547
rect 27157 1547 27215 1553
rect 27157 1544 27169 1547
rect 25501 1507 25559 1513
rect 25608 1516 27169 1544
rect 24394 1476 24400 1488
rect 24228 1448 24400 1476
rect 24394 1436 24400 1448
rect 24452 1436 24458 1488
rect 24670 1436 24676 1488
rect 24728 1476 24734 1488
rect 25516 1476 25544 1507
rect 24728 1448 25544 1476
rect 24728 1436 24734 1448
rect 23198 1300 23204 1352
rect 23256 1340 23262 1352
rect 23385 1343 23443 1349
rect 23385 1340 23397 1343
rect 23256 1312 23397 1340
rect 23256 1300 23262 1312
rect 23385 1309 23397 1312
rect 23431 1309 23443 1343
rect 23385 1303 23443 1309
rect 23845 1343 23903 1349
rect 23845 1309 23857 1343
rect 23891 1309 23903 1343
rect 23952 1340 23980 1436
rect 24136 1408 24164 1436
rect 24136 1380 24808 1408
rect 24397 1343 24455 1349
rect 24397 1340 24409 1343
rect 23952 1312 24409 1340
rect 23845 1303 23903 1309
rect 24397 1309 24409 1312
rect 24443 1309 24455 1343
rect 24397 1303 24455 1309
rect 23860 1272 23888 1303
rect 24670 1300 24676 1352
rect 24728 1300 24734 1352
rect 24780 1340 24808 1380
rect 25130 1368 25136 1420
rect 25188 1408 25194 1420
rect 25608 1408 25636 1516
rect 27157 1513 27169 1516
rect 27203 1513 27215 1547
rect 27157 1507 27215 1513
rect 27614 1504 27620 1556
rect 27672 1544 27678 1556
rect 28261 1547 28319 1553
rect 28261 1544 28273 1547
rect 27672 1516 28273 1544
rect 27672 1504 27678 1516
rect 28261 1513 28273 1516
rect 28307 1513 28319 1547
rect 28261 1507 28319 1513
rect 28350 1504 28356 1556
rect 28408 1544 28414 1556
rect 29086 1544 29092 1556
rect 28408 1516 29092 1544
rect 28408 1504 28414 1516
rect 29086 1504 29092 1516
rect 29144 1504 29150 1556
rect 29454 1504 29460 1556
rect 29512 1544 29518 1556
rect 31389 1547 31447 1553
rect 31389 1544 31401 1547
rect 29512 1516 31401 1544
rect 29512 1504 29518 1516
rect 31389 1513 31401 1516
rect 31435 1513 31447 1547
rect 31389 1507 31447 1513
rect 31662 1504 31668 1556
rect 31720 1544 31726 1556
rect 31846 1544 31852 1556
rect 31720 1516 31852 1544
rect 31720 1504 31726 1516
rect 31846 1504 31852 1516
rect 31904 1504 31910 1556
rect 32309 1547 32367 1553
rect 32309 1544 32321 1547
rect 32140 1516 32321 1544
rect 26234 1436 26240 1488
rect 26292 1476 26298 1488
rect 26292 1448 26648 1476
rect 26292 1436 26298 1448
rect 25188 1380 25636 1408
rect 25188 1368 25194 1380
rect 25961 1343 26019 1349
rect 25961 1340 25973 1343
rect 24780 1312 25973 1340
rect 25961 1309 25973 1312
rect 26007 1309 26019 1343
rect 25961 1303 26019 1309
rect 26513 1343 26571 1349
rect 26513 1309 26525 1343
rect 26559 1309 26571 1343
rect 26620 1340 26648 1448
rect 26694 1436 26700 1488
rect 26752 1436 26758 1488
rect 26878 1436 26884 1488
rect 26936 1476 26942 1488
rect 28442 1476 28448 1488
rect 26936 1448 28448 1476
rect 26936 1436 26942 1448
rect 28442 1436 28448 1448
rect 28500 1436 28506 1488
rect 28902 1436 28908 1488
rect 28960 1476 28966 1488
rect 30929 1479 30987 1485
rect 30929 1476 30941 1479
rect 28960 1448 30941 1476
rect 28960 1436 28966 1448
rect 30929 1445 30941 1448
rect 30975 1445 30987 1479
rect 30929 1439 30987 1445
rect 31478 1436 31484 1488
rect 31536 1476 31542 1488
rect 31938 1476 31944 1488
rect 31536 1448 31944 1476
rect 31536 1436 31542 1448
rect 31938 1436 31944 1448
rect 31996 1436 32002 1488
rect 27172 1380 27568 1408
rect 27172 1352 27200 1380
rect 27065 1343 27123 1349
rect 27065 1340 27077 1343
rect 26620 1312 27077 1340
rect 26513 1303 26571 1309
rect 27065 1309 27077 1312
rect 27111 1309 27123 1343
rect 27065 1303 27123 1309
rect 22756 1244 22968 1272
rect 23124 1244 23888 1272
rect 21913 1235 21971 1241
rect 22940 1216 22968 1244
rect 23934 1232 23940 1284
rect 23992 1272 23998 1284
rect 24688 1272 24716 1300
rect 24857 1275 24915 1281
rect 24857 1272 24869 1275
rect 23992 1244 24624 1272
rect 24688 1244 24869 1272
rect 23992 1232 23998 1244
rect 18923 1176 19380 1204
rect 18923 1173 18935 1176
rect 18877 1167 18935 1173
rect 19426 1164 19432 1216
rect 19484 1164 19490 1216
rect 19705 1207 19763 1213
rect 19705 1173 19717 1207
rect 19751 1204 19763 1207
rect 19886 1204 19892 1216
rect 19751 1176 19892 1204
rect 19751 1173 19763 1176
rect 19705 1167 19763 1173
rect 19886 1164 19892 1176
rect 19944 1164 19950 1216
rect 20073 1207 20131 1213
rect 20073 1173 20085 1207
rect 20119 1204 20131 1207
rect 20346 1204 20352 1216
rect 20119 1176 20352 1204
rect 20119 1173 20131 1176
rect 20073 1167 20131 1173
rect 20346 1164 20352 1176
rect 20404 1164 20410 1216
rect 20438 1164 20444 1216
rect 20496 1164 20502 1216
rect 20806 1164 20812 1216
rect 20864 1164 20870 1216
rect 21545 1207 21603 1213
rect 21545 1173 21557 1207
rect 21591 1204 21603 1207
rect 22094 1204 22100 1216
rect 21591 1176 22100 1204
rect 21591 1173 21603 1176
rect 21545 1167 21603 1173
rect 22094 1164 22100 1176
rect 22152 1164 22158 1216
rect 22738 1164 22744 1216
rect 22796 1164 22802 1216
rect 22922 1164 22928 1216
rect 22980 1164 22986 1216
rect 23106 1164 23112 1216
rect 23164 1164 23170 1216
rect 23566 1164 23572 1216
rect 23624 1204 23630 1216
rect 24596 1213 24624 1244
rect 24857 1241 24869 1244
rect 24903 1241 24915 1275
rect 24857 1235 24915 1241
rect 24946 1232 24952 1284
rect 25004 1272 25010 1284
rect 25409 1275 25467 1281
rect 25409 1272 25421 1275
rect 25004 1244 25421 1272
rect 25004 1232 25010 1244
rect 25409 1241 25421 1244
rect 25455 1241 25467 1275
rect 26528 1272 26556 1303
rect 27154 1300 27160 1352
rect 27212 1300 27218 1352
rect 27540 1340 27568 1380
rect 28074 1368 28080 1420
rect 28132 1408 28138 1420
rect 30469 1411 30527 1417
rect 30469 1408 30481 1411
rect 28132 1380 30481 1408
rect 28132 1368 28138 1380
rect 30469 1377 30481 1380
rect 30515 1377 30527 1411
rect 30469 1371 30527 1377
rect 30650 1368 30656 1420
rect 30708 1408 30714 1420
rect 32140 1408 32168 1516
rect 32309 1513 32321 1516
rect 32355 1513 32367 1547
rect 32861 1547 32919 1553
rect 32861 1544 32873 1547
rect 32309 1507 32367 1513
rect 32600 1516 32873 1544
rect 32600 1408 32628 1516
rect 32861 1513 32873 1516
rect 32907 1513 32919 1547
rect 32861 1507 32919 1513
rect 33042 1504 33048 1556
rect 33100 1544 33106 1556
rect 33413 1547 33471 1553
rect 33413 1544 33425 1547
rect 33100 1516 33425 1544
rect 33100 1504 33106 1516
rect 33413 1513 33425 1516
rect 33459 1513 33471 1547
rect 34885 1547 34943 1553
rect 34885 1544 34897 1547
rect 33413 1507 33471 1513
rect 33796 1516 34897 1544
rect 30708 1380 32168 1408
rect 32324 1380 32628 1408
rect 30708 1368 30714 1380
rect 27599 1343 27657 1349
rect 27599 1340 27611 1343
rect 27540 1312 27611 1340
rect 27599 1309 27611 1312
rect 27645 1309 27657 1343
rect 27599 1303 27657 1309
rect 27798 1300 27804 1352
rect 27856 1340 27862 1352
rect 28169 1343 28227 1349
rect 28169 1340 28181 1343
rect 27856 1312 28181 1340
rect 27856 1300 27862 1312
rect 28169 1309 28181 1312
rect 28215 1309 28227 1343
rect 28169 1303 28227 1309
rect 28810 1300 28816 1352
rect 28868 1340 28874 1352
rect 29365 1343 29423 1349
rect 29365 1340 29377 1343
rect 28868 1312 29377 1340
rect 28868 1300 28874 1312
rect 29365 1309 29377 1312
rect 29411 1309 29423 1343
rect 29365 1303 29423 1309
rect 29546 1300 29552 1352
rect 29604 1340 29610 1352
rect 29604 1312 29868 1340
rect 29604 1300 29610 1312
rect 29641 1275 29699 1281
rect 29641 1272 29653 1275
rect 26528 1244 27568 1272
rect 25409 1235 25467 1241
rect 24029 1207 24087 1213
rect 24029 1204 24041 1207
rect 23624 1176 24041 1204
rect 23624 1164 23630 1176
rect 24029 1173 24041 1176
rect 24075 1173 24087 1207
rect 24029 1167 24087 1173
rect 24581 1207 24639 1213
rect 24581 1173 24593 1207
rect 24627 1173 24639 1207
rect 24581 1167 24639 1173
rect 24762 1164 24768 1216
rect 24820 1204 24826 1216
rect 26053 1207 26111 1213
rect 26053 1204 26065 1207
rect 24820 1176 26065 1204
rect 24820 1164 24826 1176
rect 26053 1173 26065 1176
rect 26099 1173 26111 1207
rect 27540 1204 27568 1244
rect 27724 1244 29224 1272
rect 27724 1204 27752 1244
rect 27540 1176 27752 1204
rect 26053 1167 26111 1173
rect 27890 1164 27896 1216
rect 27948 1164 27954 1216
rect 28810 1164 28816 1216
rect 28868 1164 28874 1216
rect 29196 1213 29224 1244
rect 29472 1244 29653 1272
rect 29472 1216 29500 1244
rect 29641 1241 29653 1244
rect 29687 1241 29699 1275
rect 29840 1272 29868 1312
rect 29914 1300 29920 1352
rect 29972 1340 29978 1352
rect 30193 1343 30251 1349
rect 30193 1340 30205 1343
rect 29972 1312 30205 1340
rect 29972 1300 29978 1312
rect 30193 1309 30205 1312
rect 30239 1309 30251 1343
rect 30193 1303 30251 1309
rect 30282 1300 30288 1352
rect 30340 1340 30346 1352
rect 30340 1312 31892 1340
rect 30340 1300 30346 1312
rect 30745 1275 30803 1281
rect 30745 1272 30757 1275
rect 29840 1244 30757 1272
rect 29641 1235 29699 1241
rect 30745 1241 30757 1244
rect 30791 1241 30803 1275
rect 30745 1235 30803 1241
rect 31297 1275 31355 1281
rect 31297 1241 31309 1275
rect 31343 1272 31355 1275
rect 31864 1272 31892 1312
rect 31938 1300 31944 1352
rect 31996 1300 32002 1352
rect 32324 1340 32352 1380
rect 32858 1368 32864 1420
rect 32916 1408 32922 1420
rect 33796 1408 33824 1516
rect 34885 1513 34897 1516
rect 34931 1513 34943 1547
rect 34885 1507 34943 1513
rect 35986 1504 35992 1556
rect 36044 1544 36050 1556
rect 38102 1544 38108 1556
rect 36044 1516 38108 1544
rect 36044 1504 36050 1516
rect 38102 1504 38108 1516
rect 38160 1504 38166 1556
rect 39206 1504 39212 1556
rect 39264 1504 39270 1556
rect 40034 1504 40040 1556
rect 40092 1504 40098 1556
rect 40126 1504 40132 1556
rect 40184 1544 40190 1556
rect 41233 1547 41291 1553
rect 41233 1544 41245 1547
rect 40184 1516 41245 1544
rect 40184 1504 40190 1516
rect 41233 1513 41245 1516
rect 41279 1513 41291 1547
rect 41233 1507 41291 1513
rect 41506 1504 41512 1556
rect 41564 1504 41570 1556
rect 34054 1436 34060 1488
rect 34112 1476 34118 1488
rect 35897 1479 35955 1485
rect 35897 1476 35909 1479
rect 34112 1448 35909 1476
rect 34112 1436 34118 1448
rect 35897 1445 35909 1448
rect 35943 1445 35955 1479
rect 35897 1439 35955 1445
rect 37737 1479 37795 1485
rect 37737 1445 37749 1479
rect 37783 1445 37795 1479
rect 37737 1439 37795 1445
rect 32916 1380 33824 1408
rect 32916 1368 32922 1380
rect 34422 1368 34428 1420
rect 34480 1408 34486 1420
rect 34480 1380 35894 1408
rect 34480 1368 34486 1380
rect 32048 1312 32352 1340
rect 32048 1272 32076 1312
rect 32490 1300 32496 1352
rect 32548 1340 32554 1352
rect 32548 1312 32904 1340
rect 32548 1300 32554 1312
rect 31343 1244 31800 1272
rect 31864 1244 32076 1272
rect 31343 1241 31355 1244
rect 31297 1235 31355 1241
rect 29181 1207 29239 1213
rect 29181 1173 29193 1207
rect 29227 1173 29239 1207
rect 29181 1167 29239 1173
rect 29454 1164 29460 1216
rect 29512 1164 29518 1216
rect 29730 1164 29736 1216
rect 29788 1164 29794 1216
rect 31772 1213 31800 1244
rect 32214 1232 32220 1284
rect 32272 1232 32278 1284
rect 32766 1232 32772 1284
rect 32824 1232 32830 1284
rect 32876 1272 32904 1312
rect 33134 1300 33140 1352
rect 33192 1340 33198 1352
rect 33321 1343 33379 1349
rect 33321 1340 33333 1343
rect 33192 1312 33333 1340
rect 33192 1300 33198 1312
rect 33321 1309 33333 1312
rect 33367 1309 33379 1343
rect 33321 1303 33379 1309
rect 33870 1300 33876 1352
rect 33928 1300 33934 1352
rect 34054 1300 34060 1352
rect 34112 1340 34118 1352
rect 34333 1343 34391 1349
rect 34333 1340 34345 1343
rect 34112 1312 34345 1340
rect 34112 1300 34118 1312
rect 34333 1309 34345 1312
rect 34379 1309 34391 1343
rect 34333 1303 34391 1309
rect 34514 1300 34520 1352
rect 34572 1300 34578 1352
rect 35066 1300 35072 1352
rect 35124 1340 35130 1352
rect 35713 1343 35771 1349
rect 35713 1340 35725 1343
rect 35124 1312 35725 1340
rect 35124 1300 35130 1312
rect 35713 1309 35725 1312
rect 35759 1309 35771 1343
rect 35866 1340 35894 1380
rect 37200 1380 37412 1408
rect 36357 1343 36415 1349
rect 36357 1340 36369 1343
rect 35866 1312 36369 1340
rect 35713 1303 35771 1309
rect 36357 1309 36369 1312
rect 36403 1309 36415 1343
rect 36357 1303 36415 1309
rect 36449 1343 36507 1349
rect 36449 1309 36461 1343
rect 36495 1309 36507 1343
rect 36449 1303 36507 1309
rect 34532 1272 34560 1300
rect 32876 1244 34560 1272
rect 34606 1232 34612 1284
rect 34664 1272 34670 1284
rect 34793 1275 34851 1281
rect 34793 1272 34805 1275
rect 34664 1244 34805 1272
rect 34664 1232 34670 1244
rect 34793 1241 34805 1244
rect 34839 1241 34851 1275
rect 34793 1235 34851 1241
rect 31757 1207 31815 1213
rect 31757 1173 31769 1207
rect 31803 1173 31815 1207
rect 31757 1167 31815 1173
rect 31846 1164 31852 1216
rect 31904 1204 31910 1216
rect 33965 1207 34023 1213
rect 33965 1204 33977 1207
rect 31904 1176 33977 1204
rect 31904 1164 31910 1176
rect 33965 1173 33977 1176
rect 34011 1173 34023 1207
rect 33965 1167 34023 1173
rect 34514 1164 34520 1216
rect 34572 1164 34578 1216
rect 34808 1204 34836 1235
rect 34974 1232 34980 1284
rect 35032 1272 35038 1284
rect 36464 1272 36492 1303
rect 36722 1300 36728 1352
rect 36780 1300 36786 1352
rect 35032 1244 36492 1272
rect 35032 1232 35038 1244
rect 36538 1232 36544 1284
rect 36596 1272 36602 1284
rect 37200 1272 37228 1380
rect 37274 1300 37280 1352
rect 37332 1300 37338 1352
rect 36596 1244 37228 1272
rect 36596 1232 36602 1244
rect 35437 1207 35495 1213
rect 35437 1204 35449 1207
rect 34808 1176 35449 1204
rect 35437 1173 35449 1176
rect 35483 1173 35495 1207
rect 35437 1167 35495 1173
rect 36170 1164 36176 1216
rect 36228 1164 36234 1216
rect 36630 1164 36636 1216
rect 36688 1164 36694 1216
rect 36906 1164 36912 1216
rect 36964 1164 36970 1216
rect 37292 1213 37320 1300
rect 37384 1272 37412 1380
rect 37458 1300 37464 1352
rect 37516 1300 37522 1352
rect 37550 1300 37556 1352
rect 37608 1300 37614 1352
rect 37642 1300 37648 1352
rect 37700 1340 37706 1352
rect 37752 1340 37780 1439
rect 39850 1436 39856 1488
rect 39908 1436 39914 1488
rect 40052 1476 40080 1504
rect 40957 1479 41015 1485
rect 40957 1476 40969 1479
rect 40052 1448 40969 1476
rect 40957 1445 40969 1448
rect 41003 1445 41015 1479
rect 40957 1439 41015 1445
rect 39298 1368 39304 1420
rect 39356 1408 39362 1420
rect 39356 1380 41460 1408
rect 39356 1368 39362 1380
rect 37700 1312 37780 1340
rect 37700 1300 37706 1312
rect 37826 1300 37832 1352
rect 37884 1300 37890 1352
rect 38102 1300 38108 1352
rect 38160 1300 38166 1352
rect 38381 1343 38439 1349
rect 38381 1309 38393 1343
rect 38427 1309 38439 1343
rect 38381 1303 38439 1309
rect 38396 1272 38424 1303
rect 38654 1300 38660 1352
rect 38712 1300 38718 1352
rect 38930 1300 38936 1352
rect 38988 1300 38994 1352
rect 39390 1300 39396 1352
rect 39448 1300 39454 1352
rect 39485 1343 39543 1349
rect 39485 1309 39497 1343
rect 39531 1309 39543 1343
rect 39485 1303 39543 1309
rect 37384 1244 38424 1272
rect 38470 1232 38476 1284
rect 38528 1272 38534 1284
rect 39500 1272 39528 1303
rect 40034 1300 40040 1352
rect 40092 1300 40098 1352
rect 40310 1300 40316 1352
rect 40368 1300 40374 1352
rect 40586 1300 40592 1352
rect 40644 1300 40650 1352
rect 40862 1300 40868 1352
rect 40920 1300 40926 1352
rect 41138 1300 41144 1352
rect 41196 1300 41202 1352
rect 41432 1349 41460 1380
rect 41417 1343 41475 1349
rect 41417 1309 41429 1343
rect 41463 1309 41475 1343
rect 41417 1303 41475 1309
rect 41693 1343 41751 1349
rect 41693 1309 41705 1343
rect 41739 1309 41751 1343
rect 41693 1303 41751 1309
rect 38528 1244 39528 1272
rect 38528 1232 38534 1244
rect 39942 1232 39948 1284
rect 40000 1272 40006 1284
rect 41708 1272 41736 1303
rect 40000 1244 41736 1272
rect 40000 1232 40006 1244
rect 37277 1207 37335 1213
rect 37277 1173 37289 1207
rect 37323 1173 37335 1207
rect 37277 1167 37335 1173
rect 37366 1164 37372 1216
rect 37424 1204 37430 1216
rect 38013 1207 38071 1213
rect 38013 1204 38025 1207
rect 37424 1176 38025 1204
rect 37424 1164 37430 1176
rect 38013 1173 38025 1176
rect 38059 1173 38071 1207
rect 38013 1167 38071 1173
rect 38286 1164 38292 1216
rect 38344 1164 38350 1216
rect 38562 1164 38568 1216
rect 38620 1164 38626 1216
rect 38838 1164 38844 1216
rect 38896 1164 38902 1216
rect 39114 1164 39120 1216
rect 39172 1164 39178 1216
rect 39206 1164 39212 1216
rect 39264 1204 39270 1216
rect 39669 1207 39727 1213
rect 39669 1204 39681 1207
rect 39264 1176 39681 1204
rect 39264 1164 39270 1176
rect 39669 1173 39681 1176
rect 39715 1173 39727 1207
rect 39669 1167 39727 1173
rect 39758 1164 39764 1216
rect 39816 1204 39822 1216
rect 40129 1207 40187 1213
rect 40129 1204 40141 1207
rect 39816 1176 40141 1204
rect 39816 1164 39822 1176
rect 40129 1173 40141 1176
rect 40175 1173 40187 1207
rect 40129 1167 40187 1173
rect 40218 1164 40224 1216
rect 40276 1204 40282 1216
rect 40405 1207 40463 1213
rect 40405 1204 40417 1207
rect 40276 1176 40417 1204
rect 40276 1164 40282 1176
rect 40405 1173 40417 1176
rect 40451 1173 40463 1207
rect 40405 1167 40463 1173
rect 40678 1164 40684 1216
rect 40736 1164 40742 1216
rect 1104 1114 44040 1136
rect 1104 1062 11644 1114
rect 11696 1062 11708 1114
rect 11760 1062 11772 1114
rect 11824 1062 11836 1114
rect 11888 1062 11900 1114
rect 11952 1062 22338 1114
rect 22390 1062 22402 1114
rect 22454 1062 22466 1114
rect 22518 1062 22530 1114
rect 22582 1062 22594 1114
rect 22646 1062 33032 1114
rect 33084 1062 33096 1114
rect 33148 1062 33160 1114
rect 33212 1062 33224 1114
rect 33276 1062 33288 1114
rect 33340 1062 43726 1114
rect 43778 1062 43790 1114
rect 43842 1062 43854 1114
rect 43906 1062 43918 1114
rect 43970 1062 43982 1114
rect 44034 1062 44040 1114
rect 1104 1040 44040 1062
rect 5074 960 5080 1012
rect 5132 960 5138 1012
rect 5626 960 5632 1012
rect 5684 1000 5690 1012
rect 5684 972 15700 1000
rect 5684 960 5690 972
rect 5092 864 5120 960
rect 9950 892 9956 944
rect 10008 892 10014 944
rect 10226 892 10232 944
rect 10284 932 10290 944
rect 15672 932 15700 972
rect 19058 960 19064 1012
rect 19116 960 19122 1012
rect 19426 960 19432 1012
rect 19484 1000 19490 1012
rect 19484 972 25820 1000
rect 19484 960 19490 972
rect 19076 932 19104 960
rect 10284 904 15516 932
rect 15672 904 19104 932
rect 10284 892 10290 904
rect 5092 836 6914 864
rect 6886 796 6914 836
rect 7374 824 7380 876
rect 7432 864 7438 876
rect 9968 864 9996 892
rect 7432 836 9904 864
rect 9968 836 15424 864
rect 7432 824 7438 836
rect 9876 796 9904 836
rect 6886 768 8708 796
rect 9876 768 12434 796
rect 5994 688 6000 740
rect 6052 728 6058 740
rect 6730 728 6736 740
rect 6052 700 6736 728
rect 6052 688 6058 700
rect 6730 688 6736 700
rect 6788 688 6794 740
rect 7466 688 7472 740
rect 7524 728 7530 740
rect 8110 728 8116 740
rect 7524 700 8116 728
rect 7524 688 7530 700
rect 8110 688 8116 700
rect 8168 688 8174 740
rect 8570 688 8576 740
rect 8628 688 8634 740
rect 6086 620 6092 672
rect 6144 620 6150 672
rect 7834 620 7840 672
rect 7892 620 7898 672
rect 6104 320 6132 620
rect 7852 524 7880 620
rect 8588 592 8616 688
rect 8680 660 8708 768
rect 10410 688 10416 740
rect 10468 728 10474 740
rect 10594 728 10600 740
rect 10468 700 10600 728
rect 10468 688 10474 700
rect 10594 688 10600 700
rect 10652 688 10658 740
rect 11146 688 11152 740
rect 11204 728 11210 740
rect 11698 728 11704 740
rect 11204 700 11704 728
rect 11204 688 11210 700
rect 11698 688 11704 700
rect 11756 688 11762 740
rect 11514 660 11520 672
rect 8680 632 11520 660
rect 11514 620 11520 632
rect 11572 620 11578 672
rect 12406 660 12434 768
rect 13354 688 13360 740
rect 13412 728 13418 740
rect 13814 728 13820 740
rect 13412 700 13820 728
rect 13412 688 13418 700
rect 13814 688 13820 700
rect 13872 688 13878 740
rect 14550 688 14556 740
rect 14608 728 14614 740
rect 15194 728 15200 740
rect 14608 700 15200 728
rect 14608 688 14614 700
rect 15194 688 15200 700
rect 15252 688 15258 740
rect 12406 632 15240 660
rect 14458 592 14464 604
rect 8588 564 14464 592
rect 14458 552 14464 564
rect 14516 552 14522 604
rect 12710 524 12716 536
rect 7852 496 12716 524
rect 12710 484 12716 496
rect 12768 484 12774 536
rect 15212 524 15240 632
rect 15396 592 15424 836
rect 15488 796 15516 904
rect 22094 892 22100 944
rect 22152 932 22158 944
rect 22462 932 22468 944
rect 22152 904 22468 932
rect 22152 892 22158 904
rect 22462 892 22468 904
rect 22520 892 22526 944
rect 24026 892 24032 944
rect 24084 932 24090 944
rect 24946 932 24952 944
rect 24084 904 24952 932
rect 24084 892 24090 904
rect 24946 892 24952 904
rect 25004 892 25010 944
rect 15562 824 15568 876
rect 15620 864 15626 876
rect 25314 864 25320 876
rect 15620 836 25320 864
rect 15620 824 15626 836
rect 25314 824 25320 836
rect 25372 824 25378 876
rect 16206 796 16212 808
rect 15488 768 16212 796
rect 16206 756 16212 768
rect 16264 756 16270 808
rect 18874 756 18880 808
rect 18932 796 18938 808
rect 25792 796 25820 972
rect 27338 960 27344 1012
rect 27396 1000 27402 1012
rect 29730 1000 29736 1012
rect 27396 972 29736 1000
rect 27396 960 27402 972
rect 29730 960 29736 972
rect 29788 960 29794 1012
rect 36170 1000 36176 1012
rect 31726 972 36176 1000
rect 26050 892 26056 944
rect 26108 932 26114 944
rect 27614 932 27620 944
rect 26108 904 27620 932
rect 26108 892 26114 904
rect 27614 892 27620 904
rect 27672 892 27678 944
rect 28994 892 29000 944
rect 29052 932 29058 944
rect 31726 932 31754 972
rect 36170 960 36176 972
rect 36228 960 36234 1012
rect 37182 960 37188 1012
rect 37240 1000 37246 1012
rect 38930 1000 38936 1012
rect 37240 972 38936 1000
rect 37240 960 37246 972
rect 38930 960 38936 972
rect 38988 960 38994 1012
rect 39114 960 39120 1012
rect 39172 960 39178 1012
rect 29052 904 31754 932
rect 29052 892 29058 904
rect 34698 892 34704 944
rect 34756 932 34762 944
rect 39132 932 39160 960
rect 34756 904 39160 932
rect 34756 892 34762 904
rect 25866 824 25872 876
rect 25924 864 25930 876
rect 36630 864 36636 876
rect 25924 836 36636 864
rect 25924 824 25930 836
rect 36630 824 36636 836
rect 36688 824 36694 876
rect 38838 864 38844 876
rect 37660 836 38844 864
rect 32214 796 32220 808
rect 18932 768 22094 796
rect 25792 768 32220 796
rect 18932 756 18938 768
rect 15654 688 15660 740
rect 15712 728 15718 740
rect 16390 728 16396 740
rect 15712 700 16396 728
rect 15712 688 15718 700
rect 16390 688 16396 700
rect 16448 688 16454 740
rect 18506 688 18512 740
rect 18564 728 18570 740
rect 19150 728 19156 740
rect 18564 700 19156 728
rect 18564 688 18570 700
rect 19150 688 19156 700
rect 19208 688 19214 740
rect 20162 688 20168 740
rect 20220 688 20226 740
rect 15930 620 15936 672
rect 15988 660 15994 672
rect 16666 660 16672 672
rect 15988 632 16672 660
rect 15988 620 15994 632
rect 16666 620 16672 632
rect 16724 620 16730 672
rect 18230 620 18236 672
rect 18288 660 18294 672
rect 18874 660 18880 672
rect 18288 632 18880 660
rect 18288 620 18294 632
rect 18874 620 18880 632
rect 18932 620 18938 672
rect 20180 592 20208 688
rect 20438 620 20444 672
rect 20496 660 20502 672
rect 21174 660 21180 672
rect 20496 632 21180 660
rect 20496 620 20502 632
rect 21174 620 21180 632
rect 21232 620 21238 672
rect 15396 564 20208 592
rect 22066 592 22094 768
rect 32214 756 32220 768
rect 32272 756 32278 808
rect 35434 756 35440 808
rect 35492 796 35498 808
rect 37458 796 37464 808
rect 35492 768 37464 796
rect 35492 756 35498 768
rect 37458 756 37464 768
rect 37516 756 37522 808
rect 23658 688 23664 740
rect 23716 688 23722 740
rect 26786 688 26792 740
rect 26844 728 26850 740
rect 29454 728 29460 740
rect 26844 700 29460 728
rect 26844 688 26850 700
rect 29454 688 29460 700
rect 29512 688 29518 740
rect 29546 688 29552 740
rect 29604 728 29610 740
rect 29604 700 32904 728
rect 29604 688 29610 700
rect 23676 660 23704 688
rect 28810 660 28816 672
rect 23676 632 28816 660
rect 28810 620 28816 632
rect 28868 620 28874 672
rect 28920 632 29592 660
rect 28920 592 28948 632
rect 22066 564 28948 592
rect 29564 592 29592 632
rect 32766 620 32772 672
rect 32824 620 32830 672
rect 32784 592 32812 620
rect 29564 564 32812 592
rect 32876 592 32904 700
rect 35158 688 35164 740
rect 35216 728 35222 740
rect 36722 728 36728 740
rect 35216 700 36728 728
rect 35216 688 35222 700
rect 36722 688 36728 700
rect 36780 688 36786 740
rect 35434 620 35440 672
rect 35492 660 35498 672
rect 37550 660 37556 672
rect 35492 632 37556 660
rect 35492 620 35498 632
rect 37550 620 37556 632
rect 37608 620 37614 672
rect 37660 592 37688 836
rect 38838 824 38844 836
rect 38896 824 38902 876
rect 39114 824 39120 876
rect 39172 864 39178 876
rect 40862 864 40868 876
rect 39172 836 40868 864
rect 39172 824 39178 836
rect 40862 824 40868 836
rect 40920 824 40926 876
rect 37734 756 37740 808
rect 37792 796 37798 808
rect 39390 796 39396 808
rect 37792 768 39396 796
rect 37792 756 37798 768
rect 39390 756 39396 768
rect 39448 756 39454 808
rect 38286 688 38292 740
rect 38344 688 38350 740
rect 39114 688 39120 740
rect 39172 728 39178 740
rect 41138 728 41144 740
rect 39172 700 41144 728
rect 39172 688 39178 700
rect 41138 688 41144 700
rect 41196 688 41202 740
rect 32876 564 37688 592
rect 23382 524 23388 536
rect 15212 496 23388 524
rect 23382 484 23388 496
rect 23440 484 23446 536
rect 24486 484 24492 536
rect 24544 524 24550 536
rect 29546 524 29552 536
rect 24544 496 29552 524
rect 24544 484 24550 496
rect 29546 484 29552 496
rect 29604 484 29610 536
rect 29730 484 29736 536
rect 29788 524 29794 536
rect 34698 524 34704 536
rect 29788 496 34704 524
rect 29788 484 29794 496
rect 34698 484 34704 496
rect 34756 484 34762 536
rect 8754 416 8760 468
rect 8812 416 8818 468
rect 13446 416 13452 468
rect 13504 456 13510 468
rect 15010 456 15016 468
rect 13504 428 15016 456
rect 13504 416 13510 428
rect 15010 416 15016 428
rect 15068 416 15074 468
rect 19886 416 19892 468
rect 19944 456 19950 468
rect 20254 456 20260 468
rect 19944 428 20260 456
rect 19944 416 19950 428
rect 20254 416 20260 428
rect 20312 416 20318 468
rect 20714 416 20720 468
rect 20772 416 20778 468
rect 38304 456 38332 688
rect 38562 620 38568 672
rect 38620 660 38626 672
rect 40586 660 40592 672
rect 38620 632 40592 660
rect 38620 620 38626 632
rect 40586 620 40592 632
rect 40644 620 40650 672
rect 39850 456 39856 468
rect 22066 428 26648 456
rect 6104 292 6914 320
rect 6886 48 6914 292
rect 8772 184 8800 416
rect 20732 388 20760 416
rect 12636 360 20760 388
rect 12636 184 12664 360
rect 21726 348 21732 400
rect 21784 388 21790 400
rect 22066 388 22094 428
rect 21784 360 22094 388
rect 21784 348 21790 360
rect 13262 280 13268 332
rect 13320 320 13326 332
rect 26510 320 26516 332
rect 13320 292 26516 320
rect 13320 280 13326 292
rect 26510 280 26516 292
rect 26568 280 26574 332
rect 26620 320 26648 428
rect 29656 428 38332 456
rect 38396 428 39856 456
rect 29656 320 29684 428
rect 37366 388 37372 400
rect 26620 292 29684 320
rect 29748 360 37372 388
rect 14458 212 14464 264
rect 14516 252 14522 264
rect 21450 252 21456 264
rect 14516 224 21456 252
rect 14516 212 14522 224
rect 21450 212 21456 224
rect 21508 212 21514 264
rect 26142 212 26148 264
rect 26200 252 26206 264
rect 29748 252 29776 360
rect 37366 348 37372 360
rect 37424 348 37430 400
rect 38396 388 38424 428
rect 39850 416 39856 428
rect 39908 416 39914 468
rect 37844 360 38424 388
rect 34514 320 34520 332
rect 26200 224 29776 252
rect 31726 292 34520 320
rect 26200 212 26206 224
rect 8772 156 12664 184
rect 12710 144 12716 196
rect 12768 184 12774 196
rect 22922 184 22928 196
rect 12768 156 22928 184
rect 12768 144 12774 156
rect 22922 144 22928 156
rect 22980 144 22986 196
rect 25406 144 25412 196
rect 25464 184 25470 196
rect 31726 184 31754 292
rect 34514 280 34520 292
rect 34572 280 34578 332
rect 35618 280 35624 332
rect 35676 320 35682 332
rect 37844 320 37872 360
rect 38470 348 38476 400
rect 38528 388 38534 400
rect 40310 388 40316 400
rect 38528 360 40316 388
rect 38528 348 38534 360
rect 40310 348 40316 360
rect 40368 348 40374 400
rect 35676 292 37872 320
rect 35676 280 35682 292
rect 37918 280 37924 332
rect 37976 320 37982 332
rect 40034 320 40040 332
rect 37976 292 40040 320
rect 37976 280 37982 292
rect 40034 280 40040 292
rect 40092 280 40098 332
rect 36814 212 36820 264
rect 36872 252 36878 264
rect 38654 252 38660 264
rect 36872 224 38660 252
rect 36872 212 36878 224
rect 38654 212 38660 224
rect 38712 212 38718 264
rect 25464 156 31754 184
rect 25464 144 25470 156
rect 35802 144 35808 196
rect 35860 184 35866 196
rect 37458 184 37464 196
rect 35860 156 37464 184
rect 35860 144 35866 156
rect 37458 144 37464 156
rect 37516 144 37522 196
rect 9122 76 9128 128
rect 9180 116 9186 128
rect 13446 116 13452 128
rect 9180 88 13452 116
rect 9180 76 9186 88
rect 13446 76 13452 88
rect 13504 76 13510 128
rect 13538 76 13544 128
rect 13596 116 13602 128
rect 25958 116 25964 128
rect 13596 88 25964 116
rect 13596 76 13602 88
rect 25958 76 25964 88
rect 26016 76 26022 128
rect 26418 76 26424 128
rect 26476 116 26482 128
rect 29730 116 29736 128
rect 26476 88 29736 116
rect 26476 76 26482 88
rect 29730 76 29736 88
rect 29788 76 29794 128
rect 31754 76 31760 128
rect 31812 116 31818 128
rect 36906 116 36912 128
rect 31812 88 36912 116
rect 31812 76 31818 88
rect 36906 76 36912 88
rect 36964 76 36970 128
rect 10502 48 10508 60
rect 6886 20 10508 48
rect 10502 8 10508 20
rect 10560 8 10566 60
rect 12894 8 12900 60
rect 12952 48 12958 60
rect 26970 48 26976 60
rect 12952 20 26976 48
rect 12952 8 12958 20
rect 26970 8 26976 20
rect 27028 8 27034 60
rect 34238 8 34244 60
rect 34296 48 34302 60
rect 39206 48 39212 60
rect 34296 20 39212 48
rect 34296 8 34302 20
rect 39206 8 39212 20
rect 39264 8 39270 60
<< via1 >>
rect 13912 8780 13964 8832
rect 23572 8780 23624 8832
rect 11644 8678 11696 8730
rect 11708 8678 11760 8730
rect 11772 8678 11824 8730
rect 11836 8678 11888 8730
rect 11900 8678 11952 8730
rect 22338 8678 22390 8730
rect 22402 8678 22454 8730
rect 22466 8678 22518 8730
rect 22530 8678 22582 8730
rect 22594 8678 22646 8730
rect 33032 8678 33084 8730
rect 33096 8678 33148 8730
rect 33160 8678 33212 8730
rect 33224 8678 33276 8730
rect 33288 8678 33340 8730
rect 43726 8678 43778 8730
rect 43790 8678 43842 8730
rect 43854 8678 43906 8730
rect 43918 8678 43970 8730
rect 43982 8678 44034 8730
rect 1400 8576 1452 8628
rect 3424 8576 3476 8628
rect 5632 8619 5684 8628
rect 5632 8585 5641 8619
rect 5641 8585 5675 8619
rect 5675 8585 5684 8619
rect 5632 8576 5684 8585
rect 7656 8576 7708 8628
rect 10048 8619 10100 8628
rect 10048 8585 10057 8619
rect 10057 8585 10091 8619
rect 10091 8585 10100 8619
rect 10048 8576 10100 8585
rect 11980 8576 12032 8628
rect 14004 8576 14056 8628
rect 16120 8576 16172 8628
rect 18236 8576 18288 8628
rect 20352 8576 20404 8628
rect 22744 8619 22796 8628
rect 22744 8585 22753 8619
rect 22753 8585 22787 8619
rect 22787 8585 22796 8619
rect 22744 8576 22796 8585
rect 24676 8619 24728 8628
rect 24676 8585 24685 8619
rect 24685 8585 24719 8619
rect 24719 8585 24728 8619
rect 24676 8576 24728 8585
rect 26700 8576 26752 8628
rect 28908 8619 28960 8628
rect 28908 8585 28917 8619
rect 28917 8585 28951 8619
rect 28951 8585 28960 8619
rect 28908 8576 28960 8585
rect 30932 8576 30984 8628
rect 32956 8576 33008 8628
rect 35164 8576 35216 8628
rect 37464 8619 37516 8628
rect 37464 8585 37473 8619
rect 37473 8585 37507 8619
rect 37507 8585 37516 8619
rect 37464 8576 37516 8585
rect 39396 8576 39448 8628
rect 41512 8576 41564 8628
rect 43628 8576 43680 8628
rect 22100 8508 22152 8560
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 9772 8483 9824 8492
rect 9772 8449 9797 8483
rect 9797 8449 9824 8483
rect 9772 8440 9824 8449
rect 13912 8440 13964 8492
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 16212 8483 16264 8492
rect 16212 8449 16221 8483
rect 16221 8449 16255 8483
rect 16255 8449 16264 8483
rect 16212 8440 16264 8449
rect 18604 8440 18656 8492
rect 20444 8483 20496 8492
rect 20444 8449 20453 8483
rect 20453 8449 20487 8483
rect 20487 8449 20496 8483
rect 20444 8440 20496 8449
rect 22928 8440 22980 8492
rect 25044 8440 25096 8492
rect 26976 8483 27028 8492
rect 26976 8449 26985 8483
rect 26985 8449 27019 8483
rect 27019 8449 27028 8483
rect 26976 8440 27028 8449
rect 30104 8440 30156 8492
rect 31024 8483 31076 8492
rect 31024 8449 31033 8483
rect 31033 8449 31067 8483
rect 31067 8449 31076 8483
rect 31024 8440 31076 8449
rect 33508 8440 33560 8492
rect 26332 8372 26384 8424
rect 4436 8347 4488 8356
rect 4436 8313 4445 8347
rect 4445 8313 4479 8347
rect 4479 8313 4488 8347
rect 4436 8304 4488 8313
rect 9772 8304 9824 8356
rect 23296 8304 23348 8356
rect 37372 8483 37424 8492
rect 37372 8449 37381 8483
rect 37381 8449 37415 8483
rect 37415 8449 37424 8483
rect 37372 8440 37424 8449
rect 39948 8483 40000 8492
rect 39948 8449 39957 8483
rect 39957 8449 39991 8483
rect 39991 8449 40000 8483
rect 39948 8440 40000 8449
rect 40684 8440 40736 8492
rect 43260 8483 43312 8492
rect 43260 8449 43269 8483
rect 43269 8449 43303 8483
rect 43303 8449 43312 8483
rect 43260 8440 43312 8449
rect 36360 8304 36412 8356
rect 6297 8134 6349 8186
rect 6361 8134 6413 8186
rect 6425 8134 6477 8186
rect 6489 8134 6541 8186
rect 6553 8134 6605 8186
rect 16991 8134 17043 8186
rect 17055 8134 17107 8186
rect 17119 8134 17171 8186
rect 17183 8134 17235 8186
rect 17247 8134 17299 8186
rect 27685 8134 27737 8186
rect 27749 8134 27801 8186
rect 27813 8134 27865 8186
rect 27877 8134 27929 8186
rect 27941 8134 27993 8186
rect 38379 8134 38431 8186
rect 38443 8134 38495 8186
rect 38507 8134 38559 8186
rect 38571 8134 38623 8186
rect 38635 8134 38687 8186
rect 11644 7590 11696 7642
rect 11708 7590 11760 7642
rect 11772 7590 11824 7642
rect 11836 7590 11888 7642
rect 11900 7590 11952 7642
rect 22338 7590 22390 7642
rect 22402 7590 22454 7642
rect 22466 7590 22518 7642
rect 22530 7590 22582 7642
rect 22594 7590 22646 7642
rect 33032 7590 33084 7642
rect 33096 7590 33148 7642
rect 33160 7590 33212 7642
rect 33224 7590 33276 7642
rect 33288 7590 33340 7642
rect 43726 7590 43778 7642
rect 43790 7590 43842 7642
rect 43854 7590 43906 7642
rect 43918 7590 43970 7642
rect 43982 7590 44034 7642
rect 6297 7046 6349 7098
rect 6361 7046 6413 7098
rect 6425 7046 6477 7098
rect 6489 7046 6541 7098
rect 6553 7046 6605 7098
rect 16991 7046 17043 7098
rect 17055 7046 17107 7098
rect 17119 7046 17171 7098
rect 17183 7046 17235 7098
rect 17247 7046 17299 7098
rect 27685 7046 27737 7098
rect 27749 7046 27801 7098
rect 27813 7046 27865 7098
rect 27877 7046 27929 7098
rect 27941 7046 27993 7098
rect 38379 7046 38431 7098
rect 38443 7046 38495 7098
rect 38507 7046 38559 7098
rect 38571 7046 38623 7098
rect 38635 7046 38687 7098
rect 11644 6502 11696 6554
rect 11708 6502 11760 6554
rect 11772 6502 11824 6554
rect 11836 6502 11888 6554
rect 11900 6502 11952 6554
rect 22338 6502 22390 6554
rect 22402 6502 22454 6554
rect 22466 6502 22518 6554
rect 22530 6502 22582 6554
rect 22594 6502 22646 6554
rect 33032 6502 33084 6554
rect 33096 6502 33148 6554
rect 33160 6502 33212 6554
rect 33224 6502 33276 6554
rect 33288 6502 33340 6554
rect 43726 6502 43778 6554
rect 43790 6502 43842 6554
rect 43854 6502 43906 6554
rect 43918 6502 43970 6554
rect 43982 6502 44034 6554
rect 6297 5958 6349 6010
rect 6361 5958 6413 6010
rect 6425 5958 6477 6010
rect 6489 5958 6541 6010
rect 6553 5958 6605 6010
rect 16991 5958 17043 6010
rect 17055 5958 17107 6010
rect 17119 5958 17171 6010
rect 17183 5958 17235 6010
rect 17247 5958 17299 6010
rect 27685 5958 27737 6010
rect 27749 5958 27801 6010
rect 27813 5958 27865 6010
rect 27877 5958 27929 6010
rect 27941 5958 27993 6010
rect 38379 5958 38431 6010
rect 38443 5958 38495 6010
rect 38507 5958 38559 6010
rect 38571 5958 38623 6010
rect 38635 5958 38687 6010
rect 11644 5414 11696 5466
rect 11708 5414 11760 5466
rect 11772 5414 11824 5466
rect 11836 5414 11888 5466
rect 11900 5414 11952 5466
rect 22338 5414 22390 5466
rect 22402 5414 22454 5466
rect 22466 5414 22518 5466
rect 22530 5414 22582 5466
rect 22594 5414 22646 5466
rect 33032 5414 33084 5466
rect 33096 5414 33148 5466
rect 33160 5414 33212 5466
rect 33224 5414 33276 5466
rect 33288 5414 33340 5466
rect 43726 5414 43778 5466
rect 43790 5414 43842 5466
rect 43854 5414 43906 5466
rect 43918 5414 43970 5466
rect 43982 5414 44034 5466
rect 6297 4870 6349 4922
rect 6361 4870 6413 4922
rect 6425 4870 6477 4922
rect 6489 4870 6541 4922
rect 6553 4870 6605 4922
rect 16991 4870 17043 4922
rect 17055 4870 17107 4922
rect 17119 4870 17171 4922
rect 17183 4870 17235 4922
rect 17247 4870 17299 4922
rect 27685 4870 27737 4922
rect 27749 4870 27801 4922
rect 27813 4870 27865 4922
rect 27877 4870 27929 4922
rect 27941 4870 27993 4922
rect 38379 4870 38431 4922
rect 38443 4870 38495 4922
rect 38507 4870 38559 4922
rect 38571 4870 38623 4922
rect 38635 4870 38687 4922
rect 6828 4632 6880 4684
rect 23480 4632 23532 4684
rect 6736 4564 6788 4616
rect 23940 4564 23992 4616
rect 11980 4496 12032 4548
rect 28080 4496 28132 4548
rect 11336 4428 11388 4480
rect 28816 4428 28868 4480
rect 11644 4326 11696 4378
rect 11708 4326 11760 4378
rect 11772 4326 11824 4378
rect 11836 4326 11888 4378
rect 11900 4326 11952 4378
rect 22338 4326 22390 4378
rect 22402 4326 22454 4378
rect 22466 4326 22518 4378
rect 22530 4326 22582 4378
rect 22594 4326 22646 4378
rect 33032 4326 33084 4378
rect 33096 4326 33148 4378
rect 33160 4326 33212 4378
rect 33224 4326 33276 4378
rect 33288 4326 33340 4378
rect 43726 4326 43778 4378
rect 43790 4326 43842 4378
rect 43854 4326 43906 4378
rect 43918 4326 43970 4378
rect 43982 4326 44034 4378
rect 16488 4224 16540 4276
rect 33784 4224 33836 4276
rect 15660 4156 15712 4208
rect 34888 4156 34940 4208
rect 6297 3782 6349 3834
rect 6361 3782 6413 3834
rect 6425 3782 6477 3834
rect 6489 3782 6541 3834
rect 6553 3782 6605 3834
rect 16991 3782 17043 3834
rect 17055 3782 17107 3834
rect 17119 3782 17171 3834
rect 17183 3782 17235 3834
rect 17247 3782 17299 3834
rect 27685 3782 27737 3834
rect 27749 3782 27801 3834
rect 27813 3782 27865 3834
rect 27877 3782 27929 3834
rect 27941 3782 27993 3834
rect 38379 3782 38431 3834
rect 38443 3782 38495 3834
rect 38507 3782 38559 3834
rect 38571 3782 38623 3834
rect 38635 3782 38687 3834
rect 16304 3408 16356 3460
rect 30380 3408 30432 3460
rect 8024 3340 8076 3392
rect 21456 3340 21508 3392
rect 11644 3238 11696 3290
rect 11708 3238 11760 3290
rect 11772 3238 11824 3290
rect 11836 3238 11888 3290
rect 11900 3238 11952 3290
rect 22338 3238 22390 3290
rect 22402 3238 22454 3290
rect 22466 3238 22518 3290
rect 22530 3238 22582 3290
rect 22594 3238 22646 3290
rect 33032 3238 33084 3290
rect 33096 3238 33148 3290
rect 33160 3238 33212 3290
rect 33224 3238 33276 3290
rect 33288 3238 33340 3290
rect 43726 3238 43778 3290
rect 43790 3238 43842 3290
rect 43854 3238 43906 3290
rect 43918 3238 43970 3290
rect 43982 3238 44034 3290
rect 17960 3136 18012 3188
rect 26148 3136 26200 3188
rect 29920 3136 29972 3188
rect 17684 3068 17736 3120
rect 5356 3000 5408 3052
rect 25412 3000 25464 3052
rect 26056 3000 26108 3052
rect 12256 2932 12308 2984
rect 28080 3000 28132 3052
rect 28264 3043 28316 3052
rect 28264 3009 28273 3043
rect 28273 3009 28307 3043
rect 28307 3009 28316 3043
rect 28264 3000 28316 3009
rect 27620 2932 27672 2984
rect 28816 3043 28868 3052
rect 28816 3009 28825 3043
rect 28825 3009 28859 3043
rect 28859 3009 28868 3043
rect 28816 3000 28868 3009
rect 16580 2864 16632 2916
rect 11520 2796 11572 2848
rect 19340 2796 19392 2848
rect 19432 2839 19484 2848
rect 19432 2805 19441 2839
rect 19441 2805 19475 2839
rect 19475 2805 19484 2839
rect 19432 2796 19484 2805
rect 22100 2907 22152 2916
rect 22100 2873 22109 2907
rect 22109 2873 22143 2907
rect 22143 2873 22152 2907
rect 22100 2864 22152 2873
rect 24676 2864 24728 2916
rect 25228 2864 25280 2916
rect 25872 2864 25924 2916
rect 27436 2864 27488 2916
rect 37280 3068 37332 3120
rect 39212 3000 39264 3052
rect 25320 2796 25372 2848
rect 26240 2796 26292 2848
rect 26424 2796 26476 2848
rect 27252 2839 27304 2848
rect 27252 2805 27261 2839
rect 27261 2805 27295 2839
rect 27295 2805 27304 2839
rect 27252 2796 27304 2805
rect 28080 2839 28132 2848
rect 28080 2805 28089 2839
rect 28089 2805 28123 2839
rect 28123 2805 28132 2839
rect 28080 2796 28132 2805
rect 28356 2839 28408 2848
rect 28356 2805 28365 2839
rect 28365 2805 28399 2839
rect 28399 2805 28408 2839
rect 28356 2796 28408 2805
rect 28632 2839 28684 2848
rect 28632 2805 28641 2839
rect 28641 2805 28675 2839
rect 28675 2805 28684 2839
rect 28632 2796 28684 2805
rect 31760 2864 31812 2916
rect 29368 2839 29420 2848
rect 29368 2805 29377 2839
rect 29377 2805 29411 2839
rect 29411 2805 29420 2839
rect 29368 2796 29420 2805
rect 31116 2796 31168 2848
rect 32956 2796 33008 2848
rect 6297 2694 6349 2746
rect 6361 2694 6413 2746
rect 6425 2694 6477 2746
rect 6489 2694 6541 2746
rect 6553 2694 6605 2746
rect 16991 2694 17043 2746
rect 17055 2694 17107 2746
rect 17119 2694 17171 2746
rect 17183 2694 17235 2746
rect 17247 2694 17299 2746
rect 27685 2694 27737 2746
rect 27749 2694 27801 2746
rect 27813 2694 27865 2746
rect 27877 2694 27929 2746
rect 27941 2694 27993 2746
rect 38379 2694 38431 2746
rect 38443 2694 38495 2746
rect 38507 2694 38559 2746
rect 38571 2694 38623 2746
rect 38635 2694 38687 2746
rect 14096 2635 14148 2644
rect 14096 2601 14105 2635
rect 14105 2601 14139 2635
rect 14139 2601 14148 2635
rect 14096 2592 14148 2601
rect 16304 2635 16356 2644
rect 16304 2601 16313 2635
rect 16313 2601 16347 2635
rect 16347 2601 16356 2635
rect 16304 2592 16356 2601
rect 16396 2592 16448 2644
rect 18512 2635 18564 2644
rect 18512 2601 18521 2635
rect 18521 2601 18555 2635
rect 18555 2601 18564 2635
rect 18512 2592 18564 2601
rect 18604 2592 18656 2644
rect 18972 2592 19024 2644
rect 17776 2524 17828 2576
rect 14280 2431 14332 2440
rect 14280 2397 14289 2431
rect 14289 2397 14323 2431
rect 14323 2397 14332 2431
rect 14280 2388 14332 2397
rect 14648 2388 14700 2440
rect 16304 2388 16356 2440
rect 16764 2388 16816 2440
rect 18420 2388 18472 2440
rect 18512 2388 18564 2440
rect 10416 2320 10468 2372
rect 9680 2252 9732 2304
rect 18512 2252 18564 2304
rect 19800 2524 19852 2576
rect 20536 2635 20588 2644
rect 20536 2601 20545 2635
rect 20545 2601 20579 2635
rect 20579 2601 20588 2635
rect 20536 2592 20588 2601
rect 20812 2635 20864 2644
rect 20812 2601 20821 2635
rect 20821 2601 20855 2635
rect 20855 2601 20864 2635
rect 20812 2592 20864 2601
rect 22928 2635 22980 2644
rect 22928 2601 22937 2635
rect 22937 2601 22971 2635
rect 22971 2601 22980 2635
rect 22928 2592 22980 2601
rect 23572 2592 23624 2644
rect 24952 2635 25004 2644
rect 24952 2601 24961 2635
rect 24961 2601 24995 2635
rect 24995 2601 25004 2635
rect 24952 2592 25004 2601
rect 25044 2635 25096 2644
rect 25044 2601 25053 2635
rect 25053 2601 25087 2635
rect 25087 2601 25096 2635
rect 25044 2592 25096 2601
rect 26332 2592 26384 2644
rect 27160 2592 27212 2644
rect 27344 2592 27396 2644
rect 30932 2592 30984 2644
rect 31024 2592 31076 2644
rect 33508 2635 33560 2644
rect 33508 2601 33517 2635
rect 33517 2601 33551 2635
rect 33551 2601 33560 2635
rect 33508 2592 33560 2601
rect 33784 2592 33836 2644
rect 34152 2592 34204 2644
rect 36360 2635 36412 2644
rect 36360 2601 36369 2635
rect 36369 2601 36403 2635
rect 36403 2601 36412 2635
rect 36360 2592 36412 2601
rect 37372 2592 37424 2644
rect 39948 2592 40000 2644
rect 40684 2635 40736 2644
rect 40684 2601 40693 2635
rect 40693 2601 40727 2635
rect 40727 2601 40736 2635
rect 40684 2592 40736 2601
rect 43260 2592 43312 2644
rect 18696 2456 18748 2508
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 19064 2388 19116 2440
rect 19340 2388 19392 2440
rect 20076 2388 20128 2440
rect 20168 2431 20220 2440
rect 20168 2397 20177 2431
rect 20177 2397 20211 2431
rect 20211 2397 20220 2431
rect 20168 2388 20220 2397
rect 20812 2388 20864 2440
rect 20996 2431 21048 2440
rect 20996 2397 21005 2431
rect 21005 2397 21039 2431
rect 21039 2397 21048 2431
rect 20996 2388 21048 2397
rect 21272 2431 21324 2440
rect 21272 2397 21281 2431
rect 21281 2397 21315 2431
rect 21315 2397 21324 2431
rect 21272 2388 21324 2397
rect 21456 2388 21508 2440
rect 22376 2431 22428 2440
rect 22376 2397 22385 2431
rect 22385 2397 22419 2431
rect 22419 2397 22428 2431
rect 22376 2388 22428 2397
rect 22744 2388 22796 2440
rect 23572 2388 23624 2440
rect 23848 2320 23900 2372
rect 19892 2252 19944 2304
rect 20444 2252 20496 2304
rect 21272 2252 21324 2304
rect 21548 2295 21600 2304
rect 21548 2261 21557 2295
rect 21557 2261 21591 2295
rect 21591 2261 21600 2295
rect 21548 2252 21600 2261
rect 22008 2252 22060 2304
rect 22192 2295 22244 2304
rect 22192 2261 22201 2295
rect 22201 2261 22235 2295
rect 22235 2261 22244 2295
rect 22192 2252 22244 2261
rect 23204 2252 23256 2304
rect 25228 2524 25280 2576
rect 25596 2567 25648 2576
rect 25596 2533 25605 2567
rect 25605 2533 25639 2567
rect 25639 2533 25648 2567
rect 25596 2524 25648 2533
rect 25872 2567 25924 2576
rect 25872 2533 25881 2567
rect 25881 2533 25915 2567
rect 25915 2533 25924 2567
rect 25872 2524 25924 2533
rect 37648 2524 37700 2576
rect 25320 2388 25372 2440
rect 26608 2456 26660 2508
rect 25964 2388 26016 2440
rect 26332 2431 26384 2440
rect 26332 2397 26341 2431
rect 26341 2397 26375 2431
rect 26375 2397 26384 2431
rect 26332 2388 26384 2397
rect 26424 2431 26476 2440
rect 26424 2397 26433 2431
rect 26433 2397 26467 2431
rect 26467 2397 26476 2431
rect 26424 2388 26476 2397
rect 26792 2388 26844 2440
rect 26976 2388 27028 2440
rect 27436 2431 27488 2440
rect 27436 2397 27445 2431
rect 27445 2397 27479 2431
rect 27479 2397 27488 2431
rect 27436 2388 27488 2397
rect 28080 2388 28132 2440
rect 28172 2431 28224 2440
rect 28172 2397 28181 2431
rect 28181 2397 28215 2431
rect 28215 2397 28224 2431
rect 28172 2388 28224 2397
rect 29000 2388 29052 2440
rect 29184 2431 29236 2440
rect 29184 2397 29193 2431
rect 29193 2397 29227 2431
rect 29227 2397 29236 2431
rect 29184 2388 29236 2397
rect 26240 2252 26292 2304
rect 26700 2295 26752 2304
rect 26700 2261 26709 2295
rect 26709 2261 26743 2295
rect 26743 2261 26752 2295
rect 26700 2252 26752 2261
rect 26792 2252 26844 2304
rect 27804 2295 27856 2304
rect 27804 2261 27813 2295
rect 27813 2261 27847 2295
rect 27847 2261 27856 2295
rect 27804 2252 27856 2261
rect 27988 2295 28040 2304
rect 27988 2261 27997 2295
rect 27997 2261 28031 2295
rect 28031 2261 28040 2295
rect 27988 2252 28040 2261
rect 28264 2252 28316 2304
rect 28724 2252 28776 2304
rect 29092 2320 29144 2372
rect 30012 2431 30064 2440
rect 30012 2397 30021 2431
rect 30021 2397 30055 2431
rect 30055 2397 30064 2431
rect 30012 2388 30064 2397
rect 30104 2388 30156 2440
rect 29552 2295 29604 2304
rect 29552 2261 29561 2295
rect 29561 2261 29595 2295
rect 29595 2261 29604 2295
rect 29552 2252 29604 2261
rect 29828 2295 29880 2304
rect 29828 2261 29837 2295
rect 29837 2261 29871 2295
rect 29871 2261 29880 2295
rect 29828 2252 29880 2261
rect 34244 2456 34296 2508
rect 30196 2252 30248 2304
rect 32864 2431 32916 2440
rect 32864 2397 32873 2431
rect 32873 2397 32907 2431
rect 32907 2397 32916 2431
rect 32864 2388 32916 2397
rect 33692 2431 33744 2440
rect 33692 2397 33701 2431
rect 33701 2397 33735 2431
rect 33735 2397 33744 2431
rect 33692 2388 33744 2397
rect 36544 2431 36596 2440
rect 36544 2397 36553 2431
rect 36553 2397 36587 2431
rect 36587 2397 36596 2431
rect 36544 2388 36596 2397
rect 37924 2431 37976 2440
rect 37924 2397 37933 2431
rect 37933 2397 37967 2431
rect 37967 2397 37976 2431
rect 37924 2388 37976 2397
rect 39672 2431 39724 2440
rect 39672 2397 39681 2431
rect 39681 2397 39715 2431
rect 39715 2397 39724 2431
rect 39672 2388 39724 2397
rect 40868 2431 40920 2440
rect 40868 2397 40877 2431
rect 40877 2397 40911 2431
rect 40911 2397 40920 2431
rect 40868 2388 40920 2397
rect 42432 2431 42484 2440
rect 42432 2397 42441 2431
rect 42441 2397 42475 2431
rect 42475 2397 42484 2431
rect 42432 2388 42484 2397
rect 35624 2320 35676 2372
rect 32588 2252 32640 2304
rect 11644 2150 11696 2202
rect 11708 2150 11760 2202
rect 11772 2150 11824 2202
rect 11836 2150 11888 2202
rect 11900 2150 11952 2202
rect 22338 2150 22390 2202
rect 22402 2150 22454 2202
rect 22466 2150 22518 2202
rect 22530 2150 22582 2202
rect 22594 2150 22646 2202
rect 33032 2150 33084 2202
rect 33096 2150 33148 2202
rect 33160 2150 33212 2202
rect 33224 2150 33276 2202
rect 33288 2150 33340 2202
rect 43726 2150 43778 2202
rect 43790 2150 43842 2202
rect 43854 2150 43906 2202
rect 43918 2150 43970 2202
rect 43982 2150 44034 2202
rect 6736 2091 6788 2100
rect 6736 2057 6745 2091
rect 6745 2057 6779 2091
rect 6779 2057 6788 2091
rect 6736 2048 6788 2057
rect 14280 2048 14332 2100
rect 15384 2091 15436 2100
rect 15384 2057 15393 2091
rect 15393 2057 15427 2091
rect 15427 2057 15436 2091
rect 15384 2048 15436 2057
rect 15660 2091 15712 2100
rect 15660 2057 15669 2091
rect 15669 2057 15703 2091
rect 15703 2057 15712 2091
rect 15660 2048 15712 2057
rect 6552 1955 6604 1964
rect 6552 1921 6561 1955
rect 6561 1921 6595 1955
rect 6595 1921 6604 1955
rect 6552 1912 6604 1921
rect 13728 1955 13780 1964
rect 13728 1921 13737 1955
rect 13737 1921 13771 1955
rect 13771 1921 13780 1955
rect 13728 1912 13780 1921
rect 14372 1955 14424 1964
rect 14372 1921 14381 1955
rect 14381 1921 14415 1955
rect 14415 1921 14424 1955
rect 14372 1912 14424 1921
rect 15108 1955 15160 1964
rect 15108 1921 15117 1955
rect 15117 1921 15151 1955
rect 15151 1921 15160 1955
rect 15108 1912 15160 1921
rect 15292 1912 15344 1964
rect 14924 1844 14976 1896
rect 15752 1955 15804 1964
rect 15752 1921 15761 1955
rect 15761 1921 15795 1955
rect 15795 1921 15804 1955
rect 15752 1912 15804 1921
rect 16304 2048 16356 2100
rect 16488 2091 16540 2100
rect 16488 2057 16497 2091
rect 16497 2057 16531 2091
rect 16531 2057 16540 2091
rect 16488 2048 16540 2057
rect 16856 2048 16908 2100
rect 17684 2048 17736 2100
rect 18788 2048 18840 2100
rect 16212 1955 16264 1964
rect 16212 1921 16221 1955
rect 16221 1921 16255 1955
rect 16255 1921 16264 1955
rect 16212 1912 16264 1921
rect 16304 1955 16356 1964
rect 16304 1921 16313 1955
rect 16313 1921 16347 1955
rect 16347 1921 16356 1955
rect 16304 1912 16356 1921
rect 16396 1912 16448 1964
rect 16856 1912 16908 1964
rect 17316 1955 17368 1964
rect 17316 1921 17325 1955
rect 17325 1921 17359 1955
rect 17359 1921 17368 1955
rect 17316 1912 17368 1921
rect 17592 1955 17644 1964
rect 17592 1921 17601 1955
rect 17601 1921 17635 1955
rect 17635 1921 17644 1955
rect 17592 1912 17644 1921
rect 17868 1912 17920 1964
rect 18052 1955 18104 1964
rect 18052 1921 18061 1955
rect 18061 1921 18095 1955
rect 18095 1921 18104 1955
rect 18052 1912 18104 1921
rect 18328 1955 18380 1964
rect 18328 1921 18337 1955
rect 18337 1921 18371 1955
rect 18371 1921 18380 1955
rect 18328 1912 18380 1921
rect 18420 1955 18472 1964
rect 18420 1921 18429 1955
rect 18429 1921 18463 1955
rect 18463 1921 18472 1955
rect 18420 1912 18472 1921
rect 17960 1844 18012 1896
rect 19156 1955 19208 1964
rect 19156 1921 19165 1955
rect 19165 1921 19199 1955
rect 19199 1921 19208 1955
rect 19156 1912 19208 1921
rect 18788 1844 18840 1896
rect 20536 2048 20588 2100
rect 20444 1980 20496 2032
rect 20812 1955 20864 1964
rect 20812 1921 20821 1955
rect 20821 1921 20855 1955
rect 20855 1921 20864 1955
rect 20812 1912 20864 1921
rect 20904 1912 20956 1964
rect 23112 2048 23164 2100
rect 23572 2048 23624 2100
rect 23940 2048 23992 2100
rect 22928 1955 22980 1964
rect 22928 1921 22937 1955
rect 22937 1921 22971 1955
rect 22971 1921 22980 1955
rect 22928 1912 22980 1921
rect 23388 1912 23440 1964
rect 23480 1955 23532 1964
rect 23480 1921 23489 1955
rect 23489 1921 23523 1955
rect 23523 1921 23532 1955
rect 23480 1912 23532 1921
rect 23756 1955 23808 1964
rect 23756 1921 23765 1955
rect 23765 1921 23799 1955
rect 23799 1921 23808 1955
rect 23756 1912 23808 1921
rect 24216 1912 24268 1964
rect 24308 1955 24360 1964
rect 24308 1921 24317 1955
rect 24317 1921 24351 1955
rect 24351 1921 24360 1955
rect 24308 1912 24360 1921
rect 24768 2048 24820 2100
rect 25596 2048 25648 2100
rect 26700 2048 26752 2100
rect 24676 1912 24728 1964
rect 24952 1912 25004 1964
rect 26056 1980 26108 2032
rect 25228 1912 25280 1964
rect 26608 1912 26660 1964
rect 27988 2048 28040 2100
rect 28908 2048 28960 2100
rect 29828 2048 29880 2100
rect 30196 2048 30248 2100
rect 28632 1980 28684 2032
rect 28356 1912 28408 1964
rect 28448 1912 28500 1964
rect 28908 1912 28960 1964
rect 29000 1912 29052 1964
rect 30380 1980 30432 2032
rect 31852 2048 31904 2100
rect 33692 2048 33744 2100
rect 30748 1912 30800 1964
rect 17408 1776 17460 1828
rect 18236 1776 18288 1828
rect 16580 1708 16632 1760
rect 18512 1708 18564 1760
rect 18880 1751 18932 1760
rect 18880 1717 18889 1751
rect 18889 1717 18923 1751
rect 18923 1717 18932 1751
rect 18880 1708 18932 1717
rect 19616 1708 19668 1760
rect 19708 1751 19760 1760
rect 19708 1717 19717 1751
rect 19717 1717 19751 1751
rect 19751 1717 19760 1751
rect 19708 1708 19760 1717
rect 19984 1708 20036 1760
rect 20904 1751 20956 1760
rect 20904 1717 20913 1751
rect 20913 1717 20947 1751
rect 20947 1717 20956 1751
rect 20904 1708 20956 1717
rect 21088 1708 21140 1760
rect 21916 1708 21968 1760
rect 22836 1776 22888 1828
rect 23020 1776 23072 1828
rect 25320 1844 25372 1896
rect 26332 1844 26384 1896
rect 27436 1844 27488 1896
rect 33324 2023 33376 2032
rect 33324 1989 33333 2023
rect 33333 1989 33367 2023
rect 33367 1989 33376 2023
rect 33324 1980 33376 1989
rect 34152 1980 34204 2032
rect 36544 2048 36596 2100
rect 37924 2048 37976 2100
rect 39672 2048 39724 2100
rect 40868 2048 40920 2100
rect 42432 2048 42484 2100
rect 31208 1844 31260 1896
rect 34888 1955 34940 1964
rect 34888 1921 34897 1955
rect 34897 1921 34931 1955
rect 34931 1921 34940 1955
rect 34888 1912 34940 1921
rect 36360 1955 36412 1964
rect 36360 1921 36369 1955
rect 36369 1921 36403 1955
rect 36403 1921 36412 1955
rect 36360 1912 36412 1921
rect 24768 1776 24820 1828
rect 24860 1776 24912 1828
rect 27160 1776 27212 1828
rect 28356 1819 28408 1828
rect 28356 1785 28365 1819
rect 28365 1785 28399 1819
rect 28399 1785 28408 1819
rect 28356 1776 28408 1785
rect 28632 1776 28684 1828
rect 29368 1776 29420 1828
rect 24032 1708 24084 1760
rect 24124 1751 24176 1760
rect 24124 1717 24133 1751
rect 24133 1717 24167 1751
rect 24167 1717 24176 1751
rect 24124 1708 24176 1717
rect 24676 1708 24728 1760
rect 25228 1708 25280 1760
rect 25872 1708 25924 1760
rect 26608 1751 26660 1760
rect 26608 1717 26617 1751
rect 26617 1717 26651 1751
rect 26651 1717 26660 1751
rect 26608 1708 26660 1717
rect 27436 1708 27488 1760
rect 28172 1708 28224 1760
rect 29644 1708 29696 1760
rect 31024 1751 31076 1760
rect 31024 1717 31033 1751
rect 31033 1717 31067 1751
rect 31067 1717 31076 1751
rect 31024 1708 31076 1717
rect 31300 1708 31352 1760
rect 31944 1776 31996 1828
rect 33048 1776 33100 1828
rect 33324 1776 33376 1828
rect 32404 1708 32456 1760
rect 32956 1708 33008 1760
rect 33508 1708 33560 1760
rect 34520 1751 34572 1760
rect 34520 1717 34529 1751
rect 34529 1717 34563 1751
rect 34563 1717 34572 1751
rect 34520 1708 34572 1717
rect 36544 1819 36596 1828
rect 36544 1785 36553 1819
rect 36553 1785 36587 1819
rect 36587 1785 36596 1819
rect 36544 1776 36596 1785
rect 40040 1912 40092 1964
rect 40132 1955 40184 1964
rect 40132 1921 40141 1955
rect 40141 1921 40175 1955
rect 40175 1921 40184 1955
rect 40132 1912 40184 1921
rect 41512 1912 41564 1964
rect 40684 1844 40736 1896
rect 39764 1776 39816 1828
rect 39948 1708 40000 1760
rect 6297 1606 6349 1658
rect 6361 1606 6413 1658
rect 6425 1606 6477 1658
rect 6489 1606 6541 1658
rect 6553 1606 6605 1658
rect 16991 1606 17043 1658
rect 17055 1606 17107 1658
rect 17119 1606 17171 1658
rect 17183 1606 17235 1658
rect 17247 1606 17299 1658
rect 27685 1606 27737 1658
rect 27749 1606 27801 1658
rect 27813 1606 27865 1658
rect 27877 1606 27929 1658
rect 27941 1606 27993 1658
rect 38379 1606 38431 1658
rect 38443 1606 38495 1658
rect 38507 1606 38559 1658
rect 38571 1606 38623 1658
rect 38635 1606 38687 1658
rect 6828 1547 6880 1556
rect 6828 1513 6837 1547
rect 6837 1513 6871 1547
rect 6871 1513 6880 1547
rect 6828 1504 6880 1513
rect 8484 1504 8536 1556
rect 10416 1504 10468 1556
rect 10784 1547 10836 1556
rect 10784 1513 10793 1547
rect 10793 1513 10827 1547
rect 10827 1513 10836 1547
rect 10784 1504 10836 1513
rect 11980 1547 12032 1556
rect 11980 1513 11989 1547
rect 11989 1513 12023 1547
rect 12023 1513 12032 1547
rect 11980 1504 12032 1513
rect 12256 1547 12308 1556
rect 12256 1513 12265 1547
rect 12265 1513 12299 1547
rect 12299 1513 12308 1547
rect 12256 1504 12308 1513
rect 13912 1547 13964 1556
rect 13912 1513 13921 1547
rect 13921 1513 13955 1547
rect 13955 1513 13964 1547
rect 13912 1504 13964 1513
rect 14648 1547 14700 1556
rect 14648 1513 14657 1547
rect 14657 1513 14691 1547
rect 14691 1513 14700 1547
rect 14648 1504 14700 1513
rect 14924 1547 14976 1556
rect 14924 1513 14933 1547
rect 14933 1513 14967 1547
rect 14967 1513 14976 1547
rect 14924 1504 14976 1513
rect 15752 1504 15804 1556
rect 16396 1504 16448 1556
rect 8300 1436 8352 1488
rect 9680 1479 9732 1488
rect 9680 1445 9689 1479
rect 9689 1445 9723 1479
rect 9723 1445 9732 1479
rect 9680 1436 9732 1445
rect 9956 1479 10008 1488
rect 9956 1445 9965 1479
rect 9965 1445 9999 1479
rect 9999 1445 10008 1479
rect 9956 1436 10008 1445
rect 10232 1479 10284 1488
rect 10232 1445 10241 1479
rect 10241 1445 10275 1479
rect 10275 1445 10284 1479
rect 10232 1436 10284 1445
rect 15292 1436 15344 1488
rect 4896 1343 4948 1352
rect 4896 1309 4905 1343
rect 4905 1309 4939 1343
rect 4939 1309 4948 1343
rect 4896 1300 4948 1309
rect 5632 1300 5684 1352
rect 5908 1300 5960 1352
rect 6000 1343 6052 1352
rect 6000 1309 6009 1343
rect 6009 1309 6043 1343
rect 6043 1309 6052 1343
rect 6000 1300 6052 1309
rect 5540 1232 5592 1284
rect 6828 1300 6880 1352
rect 7012 1232 7064 1284
rect 7472 1343 7524 1352
rect 7472 1309 7481 1343
rect 7481 1309 7515 1343
rect 7515 1309 7524 1343
rect 7472 1300 7524 1309
rect 7656 1300 7708 1352
rect 8116 1368 8168 1420
rect 7564 1232 7616 1284
rect 8392 1232 8444 1284
rect 8852 1232 8904 1284
rect 9036 1300 9088 1352
rect 9312 1232 9364 1284
rect 9588 1232 9640 1284
rect 9864 1232 9916 1284
rect 5080 1207 5132 1216
rect 5080 1173 5089 1207
rect 5089 1173 5123 1207
rect 5123 1173 5132 1207
rect 5080 1164 5132 1173
rect 5356 1207 5408 1216
rect 5356 1173 5365 1207
rect 5365 1173 5399 1207
rect 5399 1173 5408 1207
rect 5356 1164 5408 1173
rect 5632 1207 5684 1216
rect 5632 1173 5641 1207
rect 5641 1173 5675 1207
rect 5675 1173 5684 1207
rect 5632 1164 5684 1173
rect 6092 1164 6144 1216
rect 6184 1207 6236 1216
rect 6184 1173 6193 1207
rect 6193 1173 6227 1207
rect 6227 1173 6236 1207
rect 6184 1164 6236 1173
rect 6552 1207 6604 1216
rect 6552 1173 6561 1207
rect 6561 1173 6595 1207
rect 6595 1173 6604 1207
rect 6552 1164 6604 1173
rect 7380 1164 7432 1216
rect 7840 1164 7892 1216
rect 8024 1164 8076 1216
rect 8576 1164 8628 1216
rect 8760 1207 8812 1216
rect 8760 1173 8769 1207
rect 8769 1173 8803 1207
rect 8803 1173 8812 1207
rect 8760 1164 8812 1173
rect 9128 1207 9180 1216
rect 9128 1173 9137 1207
rect 9137 1173 9171 1207
rect 9171 1173 9180 1207
rect 9128 1164 9180 1173
rect 10416 1232 10468 1284
rect 10600 1343 10652 1352
rect 10600 1309 10609 1343
rect 10609 1309 10643 1343
rect 10643 1309 10652 1343
rect 10600 1300 10652 1309
rect 10692 1232 10744 1284
rect 11152 1343 11204 1352
rect 11152 1309 11161 1343
rect 11161 1309 11195 1343
rect 11195 1309 11204 1343
rect 11152 1300 11204 1309
rect 11428 1232 11480 1284
rect 11888 1232 11940 1284
rect 12256 1300 12308 1352
rect 12440 1300 12492 1352
rect 12532 1300 12584 1352
rect 12164 1232 12216 1284
rect 10324 1164 10376 1216
rect 10968 1164 11020 1216
rect 11244 1164 11296 1216
rect 11336 1207 11388 1216
rect 11336 1173 11345 1207
rect 11345 1173 11379 1207
rect 11379 1173 11388 1207
rect 11336 1164 11388 1173
rect 12072 1164 12124 1216
rect 13084 1300 13136 1352
rect 13360 1300 13412 1352
rect 14280 1368 14332 1420
rect 12992 1232 13044 1284
rect 13820 1232 13872 1284
rect 14556 1343 14608 1352
rect 14556 1309 14565 1343
rect 14565 1309 14599 1343
rect 14599 1309 14608 1343
rect 14556 1300 14608 1309
rect 15752 1368 15804 1420
rect 16856 1504 16908 1556
rect 16580 1368 16632 1420
rect 14740 1232 14792 1284
rect 15292 1232 15344 1284
rect 15660 1343 15712 1352
rect 15660 1309 15669 1343
rect 15669 1309 15703 1343
rect 15703 1309 15712 1343
rect 15660 1300 15712 1309
rect 15936 1343 15988 1352
rect 15936 1309 15945 1343
rect 15945 1309 15979 1343
rect 15979 1309 15988 1343
rect 15936 1300 15988 1309
rect 16948 1368 17000 1420
rect 17592 1504 17644 1556
rect 18420 1504 18472 1556
rect 18512 1504 18564 1556
rect 19156 1504 19208 1556
rect 17500 1479 17552 1488
rect 17500 1445 17509 1479
rect 17509 1445 17543 1479
rect 17543 1445 17552 1479
rect 17500 1436 17552 1445
rect 16120 1232 16172 1284
rect 16580 1232 16632 1284
rect 17224 1232 17276 1284
rect 12900 1164 12952 1216
rect 13268 1164 13320 1216
rect 13452 1164 13504 1216
rect 13544 1164 13596 1216
rect 15568 1164 15620 1216
rect 16212 1164 16264 1216
rect 17132 1164 17184 1216
rect 18052 1368 18104 1420
rect 19892 1436 19944 1488
rect 18604 1368 18656 1420
rect 17408 1164 17460 1216
rect 17960 1164 18012 1216
rect 18144 1232 18196 1284
rect 18420 1300 18472 1352
rect 18512 1343 18564 1352
rect 18512 1309 18521 1343
rect 18521 1309 18555 1343
rect 18555 1309 18564 1343
rect 18512 1300 18564 1309
rect 19156 1368 19208 1420
rect 19064 1343 19116 1352
rect 19064 1309 19073 1343
rect 19073 1309 19107 1343
rect 19107 1309 19116 1343
rect 19064 1300 19116 1309
rect 19524 1343 19576 1352
rect 19524 1309 19533 1343
rect 19533 1309 19567 1343
rect 19567 1309 19576 1343
rect 19524 1300 19576 1309
rect 19616 1300 19668 1352
rect 19800 1300 19852 1352
rect 22284 1436 22336 1488
rect 22836 1436 22888 1488
rect 23296 1504 23348 1556
rect 22192 1411 22244 1420
rect 22192 1377 22201 1411
rect 22201 1377 22235 1411
rect 22235 1377 22244 1411
rect 22192 1368 22244 1377
rect 20904 1300 20956 1352
rect 21272 1300 21324 1352
rect 22008 1300 22060 1352
rect 22744 1300 22796 1352
rect 18236 1164 18288 1216
rect 20536 1232 20588 1284
rect 23940 1436 23992 1488
rect 24124 1436 24176 1488
rect 24308 1504 24360 1556
rect 24400 1436 24452 1488
rect 24676 1436 24728 1488
rect 23204 1300 23256 1352
rect 24676 1300 24728 1352
rect 25136 1368 25188 1420
rect 27620 1504 27672 1556
rect 28356 1504 28408 1556
rect 29092 1504 29144 1556
rect 29460 1504 29512 1556
rect 31668 1504 31720 1556
rect 31852 1504 31904 1556
rect 26240 1436 26292 1488
rect 26700 1479 26752 1488
rect 26700 1445 26709 1479
rect 26709 1445 26743 1479
rect 26743 1445 26752 1479
rect 26700 1436 26752 1445
rect 26884 1436 26936 1488
rect 28448 1436 28500 1488
rect 28908 1436 28960 1488
rect 31484 1436 31536 1488
rect 31944 1436 31996 1488
rect 23940 1232 23992 1284
rect 19432 1207 19484 1216
rect 19432 1173 19441 1207
rect 19441 1173 19475 1207
rect 19475 1173 19484 1207
rect 19432 1164 19484 1173
rect 19892 1164 19944 1216
rect 20352 1164 20404 1216
rect 20444 1207 20496 1216
rect 20444 1173 20453 1207
rect 20453 1173 20487 1207
rect 20487 1173 20496 1207
rect 20444 1164 20496 1173
rect 20812 1207 20864 1216
rect 20812 1173 20821 1207
rect 20821 1173 20855 1207
rect 20855 1173 20864 1207
rect 20812 1164 20864 1173
rect 22100 1164 22152 1216
rect 22744 1207 22796 1216
rect 22744 1173 22753 1207
rect 22753 1173 22787 1207
rect 22787 1173 22796 1207
rect 22744 1164 22796 1173
rect 22928 1164 22980 1216
rect 23112 1207 23164 1216
rect 23112 1173 23121 1207
rect 23121 1173 23155 1207
rect 23155 1173 23164 1207
rect 23112 1164 23164 1173
rect 23572 1164 23624 1216
rect 24952 1232 25004 1284
rect 27160 1300 27212 1352
rect 28080 1368 28132 1420
rect 30656 1368 30708 1420
rect 33048 1504 33100 1556
rect 27804 1300 27856 1352
rect 28816 1300 28868 1352
rect 29552 1300 29604 1352
rect 24768 1164 24820 1216
rect 27896 1207 27948 1216
rect 27896 1173 27905 1207
rect 27905 1173 27939 1207
rect 27939 1173 27948 1207
rect 27896 1164 27948 1173
rect 28816 1207 28868 1216
rect 28816 1173 28825 1207
rect 28825 1173 28859 1207
rect 28859 1173 28868 1207
rect 28816 1164 28868 1173
rect 29920 1300 29972 1352
rect 30288 1300 30340 1352
rect 31944 1343 31996 1352
rect 31944 1309 31953 1343
rect 31953 1309 31987 1343
rect 31987 1309 31996 1343
rect 31944 1300 31996 1309
rect 32864 1368 32916 1420
rect 35992 1504 36044 1556
rect 38108 1504 38160 1556
rect 39212 1547 39264 1556
rect 39212 1513 39221 1547
rect 39221 1513 39255 1547
rect 39255 1513 39264 1547
rect 39212 1504 39264 1513
rect 40040 1504 40092 1556
rect 40132 1504 40184 1556
rect 41512 1547 41564 1556
rect 41512 1513 41521 1547
rect 41521 1513 41555 1547
rect 41555 1513 41564 1547
rect 41512 1504 41564 1513
rect 34060 1436 34112 1488
rect 34428 1368 34480 1420
rect 32496 1300 32548 1352
rect 29460 1164 29512 1216
rect 29736 1207 29788 1216
rect 29736 1173 29745 1207
rect 29745 1173 29779 1207
rect 29779 1173 29788 1207
rect 29736 1164 29788 1173
rect 32220 1275 32272 1284
rect 32220 1241 32229 1275
rect 32229 1241 32263 1275
rect 32263 1241 32272 1275
rect 32220 1232 32272 1241
rect 32772 1275 32824 1284
rect 32772 1241 32781 1275
rect 32781 1241 32815 1275
rect 32815 1241 32824 1275
rect 32772 1232 32824 1241
rect 33140 1300 33192 1352
rect 33876 1343 33928 1352
rect 33876 1309 33885 1343
rect 33885 1309 33919 1343
rect 33919 1309 33928 1343
rect 33876 1300 33928 1309
rect 34060 1300 34112 1352
rect 34520 1300 34572 1352
rect 35072 1300 35124 1352
rect 34612 1232 34664 1284
rect 31852 1164 31904 1216
rect 34520 1207 34572 1216
rect 34520 1173 34529 1207
rect 34529 1173 34563 1207
rect 34563 1173 34572 1207
rect 34520 1164 34572 1173
rect 34980 1232 35032 1284
rect 36728 1343 36780 1352
rect 36728 1309 36737 1343
rect 36737 1309 36771 1343
rect 36771 1309 36780 1343
rect 36728 1300 36780 1309
rect 36544 1232 36596 1284
rect 37280 1300 37332 1352
rect 36176 1207 36228 1216
rect 36176 1173 36185 1207
rect 36185 1173 36219 1207
rect 36219 1173 36228 1207
rect 36176 1164 36228 1173
rect 36636 1207 36688 1216
rect 36636 1173 36645 1207
rect 36645 1173 36679 1207
rect 36679 1173 36688 1207
rect 36636 1164 36688 1173
rect 36912 1207 36964 1216
rect 36912 1173 36921 1207
rect 36921 1173 36955 1207
rect 36955 1173 36964 1207
rect 36912 1164 36964 1173
rect 37464 1343 37516 1352
rect 37464 1309 37473 1343
rect 37473 1309 37507 1343
rect 37507 1309 37516 1343
rect 37464 1300 37516 1309
rect 37556 1343 37608 1352
rect 37556 1309 37565 1343
rect 37565 1309 37599 1343
rect 37599 1309 37608 1343
rect 37556 1300 37608 1309
rect 37648 1300 37700 1352
rect 39856 1479 39908 1488
rect 39856 1445 39865 1479
rect 39865 1445 39899 1479
rect 39899 1445 39908 1479
rect 39856 1436 39908 1445
rect 39304 1368 39356 1420
rect 37832 1343 37884 1352
rect 37832 1309 37841 1343
rect 37841 1309 37875 1343
rect 37875 1309 37884 1343
rect 37832 1300 37884 1309
rect 38108 1343 38160 1352
rect 38108 1309 38117 1343
rect 38117 1309 38151 1343
rect 38151 1309 38160 1343
rect 38108 1300 38160 1309
rect 38660 1343 38712 1352
rect 38660 1309 38669 1343
rect 38669 1309 38703 1343
rect 38703 1309 38712 1343
rect 38660 1300 38712 1309
rect 38936 1343 38988 1352
rect 38936 1309 38945 1343
rect 38945 1309 38979 1343
rect 38979 1309 38988 1343
rect 38936 1300 38988 1309
rect 39396 1343 39448 1352
rect 39396 1309 39405 1343
rect 39405 1309 39439 1343
rect 39439 1309 39448 1343
rect 39396 1300 39448 1309
rect 38476 1232 38528 1284
rect 40040 1343 40092 1352
rect 40040 1309 40049 1343
rect 40049 1309 40083 1343
rect 40083 1309 40092 1343
rect 40040 1300 40092 1309
rect 40316 1343 40368 1352
rect 40316 1309 40325 1343
rect 40325 1309 40359 1343
rect 40359 1309 40368 1343
rect 40316 1300 40368 1309
rect 40592 1343 40644 1352
rect 40592 1309 40601 1343
rect 40601 1309 40635 1343
rect 40635 1309 40644 1343
rect 40592 1300 40644 1309
rect 40868 1343 40920 1352
rect 40868 1309 40877 1343
rect 40877 1309 40911 1343
rect 40911 1309 40920 1343
rect 40868 1300 40920 1309
rect 41144 1343 41196 1352
rect 41144 1309 41153 1343
rect 41153 1309 41187 1343
rect 41187 1309 41196 1343
rect 41144 1300 41196 1309
rect 39948 1232 40000 1284
rect 37372 1164 37424 1216
rect 38292 1207 38344 1216
rect 38292 1173 38301 1207
rect 38301 1173 38335 1207
rect 38335 1173 38344 1207
rect 38292 1164 38344 1173
rect 38568 1207 38620 1216
rect 38568 1173 38577 1207
rect 38577 1173 38611 1207
rect 38611 1173 38620 1207
rect 38568 1164 38620 1173
rect 38844 1207 38896 1216
rect 38844 1173 38853 1207
rect 38853 1173 38887 1207
rect 38887 1173 38896 1207
rect 38844 1164 38896 1173
rect 39120 1207 39172 1216
rect 39120 1173 39129 1207
rect 39129 1173 39163 1207
rect 39163 1173 39172 1207
rect 39120 1164 39172 1173
rect 39212 1164 39264 1216
rect 39764 1164 39816 1216
rect 40224 1164 40276 1216
rect 40684 1207 40736 1216
rect 40684 1173 40693 1207
rect 40693 1173 40727 1207
rect 40727 1173 40736 1207
rect 40684 1164 40736 1173
rect 11644 1062 11696 1114
rect 11708 1062 11760 1114
rect 11772 1062 11824 1114
rect 11836 1062 11888 1114
rect 11900 1062 11952 1114
rect 22338 1062 22390 1114
rect 22402 1062 22454 1114
rect 22466 1062 22518 1114
rect 22530 1062 22582 1114
rect 22594 1062 22646 1114
rect 33032 1062 33084 1114
rect 33096 1062 33148 1114
rect 33160 1062 33212 1114
rect 33224 1062 33276 1114
rect 33288 1062 33340 1114
rect 43726 1062 43778 1114
rect 43790 1062 43842 1114
rect 43854 1062 43906 1114
rect 43918 1062 43970 1114
rect 43982 1062 44034 1114
rect 5080 960 5132 1012
rect 5632 960 5684 1012
rect 9956 892 10008 944
rect 10232 892 10284 944
rect 19064 960 19116 1012
rect 19432 960 19484 1012
rect 7380 824 7432 876
rect 6000 688 6052 740
rect 6736 688 6788 740
rect 7472 688 7524 740
rect 8116 688 8168 740
rect 8576 688 8628 740
rect 6092 620 6144 672
rect 7840 620 7892 672
rect 10416 688 10468 740
rect 10600 688 10652 740
rect 11152 688 11204 740
rect 11704 688 11756 740
rect 11520 620 11572 672
rect 13360 688 13412 740
rect 13820 688 13872 740
rect 14556 688 14608 740
rect 15200 688 15252 740
rect 14464 552 14516 604
rect 12716 484 12768 536
rect 22100 892 22152 944
rect 22468 892 22520 944
rect 24032 892 24084 944
rect 24952 892 25004 944
rect 15568 824 15620 876
rect 25320 824 25372 876
rect 16212 756 16264 808
rect 18880 756 18932 808
rect 27344 960 27396 1012
rect 29736 960 29788 1012
rect 26056 892 26108 944
rect 27620 892 27672 944
rect 29000 892 29052 944
rect 36176 960 36228 1012
rect 37188 960 37240 1012
rect 38936 960 38988 1012
rect 39120 960 39172 1012
rect 34704 892 34756 944
rect 25872 824 25924 876
rect 36636 824 36688 876
rect 15660 688 15712 740
rect 16396 688 16448 740
rect 18512 688 18564 740
rect 19156 688 19208 740
rect 20168 688 20220 740
rect 15936 620 15988 672
rect 16672 620 16724 672
rect 18236 620 18288 672
rect 18880 620 18932 672
rect 20444 620 20496 672
rect 21180 620 21232 672
rect 32220 756 32272 808
rect 35440 756 35492 808
rect 37464 756 37516 808
rect 23664 688 23716 740
rect 26792 688 26844 740
rect 29460 688 29512 740
rect 29552 688 29604 740
rect 28816 620 28868 672
rect 32772 620 32824 672
rect 35164 688 35216 740
rect 36728 688 36780 740
rect 35440 620 35492 672
rect 37556 620 37608 672
rect 38844 824 38896 876
rect 39120 824 39172 876
rect 40868 824 40920 876
rect 37740 756 37792 808
rect 39396 756 39448 808
rect 38292 688 38344 740
rect 39120 688 39172 740
rect 41144 688 41196 740
rect 23388 484 23440 536
rect 24492 484 24544 536
rect 29552 484 29604 536
rect 29736 484 29788 536
rect 34704 484 34756 536
rect 8760 416 8812 468
rect 13452 416 13504 468
rect 15016 416 15068 468
rect 19892 416 19944 468
rect 20260 416 20312 468
rect 20720 416 20772 468
rect 38568 620 38620 672
rect 40592 620 40644 672
rect 21732 348 21784 400
rect 13268 280 13320 332
rect 26516 280 26568 332
rect 14464 212 14516 264
rect 21456 212 21508 264
rect 26148 212 26200 264
rect 37372 348 37424 400
rect 39856 416 39908 468
rect 12716 144 12768 196
rect 22928 144 22980 196
rect 25412 144 25464 196
rect 34520 280 34572 332
rect 35624 280 35676 332
rect 38476 348 38528 400
rect 40316 348 40368 400
rect 37924 280 37976 332
rect 40040 280 40092 332
rect 36820 212 36872 264
rect 38660 212 38712 264
rect 35808 144 35860 196
rect 37464 144 37516 196
rect 9128 76 9180 128
rect 13452 76 13504 128
rect 13544 76 13596 128
rect 25964 76 26016 128
rect 26424 76 26476 128
rect 29736 76 29788 128
rect 31760 76 31812 128
rect 36912 76 36964 128
rect 10508 8 10560 60
rect 12900 8 12952 60
rect 26976 8 27028 60
rect 34244 8 34296 60
rect 39212 8 39264 60
<< metal2 >>
rect 1306 9840 1362 10000
rect 3422 9840 3478 10000
rect 5538 9840 5594 10000
rect 7654 9840 7710 10000
rect 9770 9840 9826 10000
rect 9876 9846 10088 9874
rect 1320 8514 1348 9840
rect 3436 8634 3464 9840
rect 5552 9058 5580 9840
rect 5552 9030 5672 9058
rect 5644 8634 5672 9030
rect 7668 8634 7696 9840
rect 9784 9738 9812 9840
rect 9876 9738 9904 9846
rect 9784 9710 9904 9738
rect 10060 8634 10088 9846
rect 11886 9840 11942 10000
rect 14002 9840 14058 10000
rect 16118 9840 16174 10000
rect 18234 9840 18290 10000
rect 20350 9840 20406 10000
rect 22466 9840 22522 10000
rect 22572 9846 22784 9874
rect 11900 8922 11928 9840
rect 11900 8894 12020 8922
rect 11644 8732 11952 8741
rect 11644 8730 11650 8732
rect 11706 8730 11730 8732
rect 11786 8730 11810 8732
rect 11866 8730 11890 8732
rect 11946 8730 11952 8732
rect 11706 8678 11708 8730
rect 11888 8678 11890 8730
rect 11644 8676 11650 8678
rect 11706 8676 11730 8678
rect 11786 8676 11810 8678
rect 11866 8676 11890 8678
rect 11946 8676 11952 8678
rect 11644 8667 11952 8676
rect 11992 8634 12020 8894
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 1412 8514 1440 8570
rect 1320 8486 1440 8514
rect 5538 8528 5594 8537
rect 13924 8498 13952 8774
rect 14016 8634 14044 9840
rect 16132 8634 16160 9840
rect 18248 8634 18276 9840
rect 20364 8634 20392 9840
rect 22480 9738 22508 9840
rect 22572 9738 22600 9846
rect 22480 9710 22600 9738
rect 22338 8732 22646 8741
rect 22338 8730 22344 8732
rect 22400 8730 22424 8732
rect 22480 8730 22504 8732
rect 22560 8730 22584 8732
rect 22640 8730 22646 8732
rect 22400 8678 22402 8730
rect 22582 8678 22584 8730
rect 22338 8676 22344 8678
rect 22400 8676 22424 8678
rect 22480 8676 22504 8678
rect 22560 8676 22584 8678
rect 22640 8676 22646 8678
rect 22338 8667 22646 8676
rect 22756 8634 22784 9846
rect 24582 9840 24638 10000
rect 26698 9840 26754 10000
rect 28814 9840 28870 10000
rect 30930 9840 30986 10000
rect 33046 9840 33102 10000
rect 35162 9840 35218 10000
rect 37278 9840 37334 10000
rect 39394 9840 39450 10000
rect 41510 9840 41566 10000
rect 43626 9840 43682 10000
rect 24596 9058 24624 9840
rect 24596 9030 24716 9058
rect 23572 8832 23624 8838
rect 23572 8774 23624 8780
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22100 8560 22152 8566
rect 22100 8502 22152 8508
rect 5538 8463 5540 8472
rect 5592 8463 5594 8472
rect 9772 8492 9824 8498
rect 5540 8434 5592 8440
rect 9772 8434 9824 8440
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 4434 8392 4490 8401
rect 9784 8362 9812 8434
rect 4434 8327 4436 8336
rect 4488 8327 4490 8336
rect 9772 8356 9824 8362
rect 4436 8298 4488 8304
rect 9772 8298 9824 8304
rect 6297 8188 6605 8197
rect 6297 8186 6303 8188
rect 6359 8186 6383 8188
rect 6439 8186 6463 8188
rect 6519 8186 6543 8188
rect 6599 8186 6605 8188
rect 6359 8134 6361 8186
rect 6541 8134 6543 8186
rect 6297 8132 6303 8134
rect 6359 8132 6383 8134
rect 6439 8132 6463 8134
rect 6519 8132 6543 8134
rect 6599 8132 6605 8134
rect 6297 8123 6605 8132
rect 11644 7644 11952 7653
rect 11644 7642 11650 7644
rect 11706 7642 11730 7644
rect 11786 7642 11810 7644
rect 11866 7642 11890 7644
rect 11946 7642 11952 7644
rect 11706 7590 11708 7642
rect 11888 7590 11890 7642
rect 11644 7588 11650 7590
rect 11706 7588 11730 7590
rect 11786 7588 11810 7590
rect 11866 7588 11890 7590
rect 11946 7588 11952 7590
rect 11644 7579 11952 7588
rect 6297 7100 6605 7109
rect 6297 7098 6303 7100
rect 6359 7098 6383 7100
rect 6439 7098 6463 7100
rect 6519 7098 6543 7100
rect 6599 7098 6605 7100
rect 6359 7046 6361 7098
rect 6541 7046 6543 7098
rect 6297 7044 6303 7046
rect 6359 7044 6383 7046
rect 6439 7044 6463 7046
rect 6519 7044 6543 7046
rect 6599 7044 6605 7046
rect 6297 7035 6605 7044
rect 11644 6556 11952 6565
rect 11644 6554 11650 6556
rect 11706 6554 11730 6556
rect 11786 6554 11810 6556
rect 11866 6554 11890 6556
rect 11946 6554 11952 6556
rect 11706 6502 11708 6554
rect 11888 6502 11890 6554
rect 11644 6500 11650 6502
rect 11706 6500 11730 6502
rect 11786 6500 11810 6502
rect 11866 6500 11890 6502
rect 11946 6500 11952 6502
rect 11644 6491 11952 6500
rect 6297 6012 6605 6021
rect 6297 6010 6303 6012
rect 6359 6010 6383 6012
rect 6439 6010 6463 6012
rect 6519 6010 6543 6012
rect 6599 6010 6605 6012
rect 6359 5958 6361 6010
rect 6541 5958 6543 6010
rect 6297 5956 6303 5958
rect 6359 5956 6383 5958
rect 6439 5956 6463 5958
rect 6519 5956 6543 5958
rect 6599 5956 6605 5958
rect 6297 5947 6605 5956
rect 11644 5468 11952 5477
rect 11644 5466 11650 5468
rect 11706 5466 11730 5468
rect 11786 5466 11810 5468
rect 11866 5466 11890 5468
rect 11946 5466 11952 5468
rect 11706 5414 11708 5466
rect 11888 5414 11890 5466
rect 11644 5412 11650 5414
rect 11706 5412 11730 5414
rect 11786 5412 11810 5414
rect 11866 5412 11890 5414
rect 11946 5412 11952 5414
rect 11644 5403 11952 5412
rect 6297 4924 6605 4933
rect 6297 4922 6303 4924
rect 6359 4922 6383 4924
rect 6439 4922 6463 4924
rect 6519 4922 6543 4924
rect 6599 4922 6605 4924
rect 6359 4870 6361 4922
rect 6541 4870 6543 4922
rect 6297 4868 6303 4870
rect 6359 4868 6383 4870
rect 6439 4868 6463 4870
rect 6519 4868 6543 4870
rect 6599 4868 6605 4870
rect 6297 4859 6605 4868
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6297 3836 6605 3845
rect 6297 3834 6303 3836
rect 6359 3834 6383 3836
rect 6439 3834 6463 3836
rect 6519 3834 6543 3836
rect 6599 3834 6605 3836
rect 6359 3782 6361 3834
rect 6541 3782 6543 3834
rect 6297 3780 6303 3782
rect 6359 3780 6383 3782
rect 6439 3780 6463 3782
rect 6519 3780 6543 3782
rect 6599 3780 6605 3782
rect 6297 3771 6605 3780
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 4896 1352 4948 1358
rect 4896 1294 4948 1300
rect 4908 82 4936 1294
rect 5368 1222 5396 2994
rect 6297 2748 6605 2757
rect 6297 2746 6303 2748
rect 6359 2746 6383 2748
rect 6439 2746 6463 2748
rect 6519 2746 6543 2748
rect 6599 2746 6605 2748
rect 6359 2694 6361 2746
rect 6541 2694 6543 2746
rect 6297 2692 6303 2694
rect 6359 2692 6383 2694
rect 6439 2692 6463 2694
rect 6519 2692 6543 2694
rect 6599 2692 6605 2694
rect 6297 2683 6605 2692
rect 6748 2106 6776 4558
rect 6736 2100 6788 2106
rect 6736 2042 6788 2048
rect 6552 1964 6604 1970
rect 6552 1906 6604 1912
rect 6564 1850 6592 1906
rect 6564 1822 6684 1850
rect 6297 1660 6605 1669
rect 6297 1658 6303 1660
rect 6359 1658 6383 1660
rect 6439 1658 6463 1660
rect 6519 1658 6543 1660
rect 6599 1658 6605 1660
rect 6359 1606 6361 1658
rect 6541 1606 6543 1658
rect 6297 1604 6303 1606
rect 6359 1604 6383 1606
rect 6439 1604 6463 1606
rect 6519 1604 6543 1606
rect 6599 1604 6605 1606
rect 6297 1595 6605 1604
rect 5632 1352 5684 1358
rect 5908 1352 5960 1358
rect 5684 1300 5764 1306
rect 5632 1294 5764 1300
rect 5908 1294 5960 1300
rect 6000 1352 6052 1358
rect 6000 1294 6052 1300
rect 5540 1284 5592 1290
rect 5644 1278 5764 1294
rect 5540 1226 5592 1232
rect 5080 1216 5132 1222
rect 5080 1158 5132 1164
rect 5356 1216 5408 1222
rect 5356 1158 5408 1164
rect 5092 1018 5120 1158
rect 5080 1012 5132 1018
rect 5080 954 5132 960
rect 5552 762 5580 1226
rect 5632 1216 5684 1222
rect 5632 1158 5684 1164
rect 5644 1018 5672 1158
rect 5632 1012 5684 1018
rect 5632 954 5684 960
rect 5552 734 5672 762
rect 5644 160 5672 734
rect 5354 82 5410 160
rect 4908 54 5410 82
rect 5354 0 5410 54
rect 5630 0 5686 160
rect 5736 82 5764 1278
rect 5920 490 5948 1294
rect 6012 746 6040 1294
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 6184 1216 6236 1222
rect 6184 1158 6236 1164
rect 6552 1216 6604 1222
rect 6552 1158 6604 1164
rect 6000 740 6052 746
rect 6000 682 6052 688
rect 6104 678 6132 1158
rect 6092 672 6144 678
rect 6196 649 6224 1158
rect 6092 614 6144 620
rect 6182 640 6238 649
rect 6182 575 6238 584
rect 5920 462 6040 490
rect 5906 82 5962 160
rect 5736 54 5962 82
rect 6012 82 6040 462
rect 6564 377 6592 1158
rect 6550 368 6606 377
rect 6550 303 6606 312
rect 6182 82 6238 160
rect 6012 54 6238 82
rect 5906 0 5962 54
rect 6182 0 6238 54
rect 6458 82 6514 160
rect 6656 82 6684 1822
rect 6840 1562 6868 4626
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 6828 1556 6880 1562
rect 6828 1498 6880 1504
rect 6840 1414 7144 1442
rect 6840 1358 6868 1414
rect 6828 1352 6880 1358
rect 6828 1294 6880 1300
rect 7012 1284 7064 1290
rect 7012 1226 7064 1232
rect 6736 740 6788 746
rect 6736 682 6788 688
rect 6748 160 6776 682
rect 7024 160 7052 1226
rect 6458 54 6684 82
rect 6458 0 6514 54
rect 6734 0 6790 160
rect 7010 0 7066 160
rect 7116 82 7144 1414
rect 7472 1352 7524 1358
rect 7472 1294 7524 1300
rect 7656 1352 7708 1358
rect 7656 1294 7708 1300
rect 7380 1216 7432 1222
rect 7380 1158 7432 1164
rect 7392 882 7420 1158
rect 7380 876 7432 882
rect 7380 818 7432 824
rect 7484 746 7512 1294
rect 7564 1284 7616 1290
rect 7564 1226 7616 1232
rect 7472 740 7524 746
rect 7472 682 7524 688
rect 7576 160 7604 1226
rect 7286 82 7342 160
rect 7116 54 7342 82
rect 7286 0 7342 54
rect 7562 0 7618 160
rect 7668 82 7696 1294
rect 8036 1222 8064 3334
rect 8482 2544 8538 2553
rect 8482 2479 8538 2488
rect 8496 1562 8524 2479
rect 10416 2372 10468 2378
rect 10416 2314 10468 2320
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 9692 1494 9720 2246
rect 10428 1562 10456 2314
rect 10782 2000 10838 2009
rect 10782 1935 10838 1944
rect 10690 1864 10746 1873
rect 10520 1822 10690 1850
rect 10416 1556 10468 1562
rect 10416 1498 10468 1504
rect 8300 1488 8352 1494
rect 8298 1456 8300 1465
rect 9680 1488 9732 1494
rect 8352 1456 8354 1465
rect 8116 1420 8168 1426
rect 8168 1380 8248 1408
rect 9680 1430 9732 1436
rect 9956 1488 10008 1494
rect 9956 1430 10008 1436
rect 10232 1488 10284 1494
rect 10232 1430 10284 1436
rect 8298 1391 8354 1400
rect 8116 1362 8168 1368
rect 7840 1216 7892 1222
rect 7840 1158 7892 1164
rect 8024 1216 8076 1222
rect 8024 1158 8076 1164
rect 7852 678 7880 1158
rect 8116 740 8168 746
rect 8116 682 8168 688
rect 7840 672 7892 678
rect 7840 614 7892 620
rect 8128 160 8156 682
rect 7838 82 7894 160
rect 7668 54 7894 82
rect 7838 0 7894 54
rect 8114 0 8170 160
rect 8220 82 8248 1380
rect 9036 1352 9088 1358
rect 9088 1312 9260 1340
rect 9036 1294 9088 1300
rect 8392 1284 8444 1290
rect 8852 1284 8904 1290
rect 8444 1244 8524 1272
rect 8392 1226 8444 1232
rect 8390 82 8446 160
rect 8220 54 8446 82
rect 8496 82 8524 1244
rect 8904 1244 8984 1272
rect 8852 1226 8904 1232
rect 8576 1216 8628 1222
rect 8576 1158 8628 1164
rect 8760 1216 8812 1222
rect 8760 1158 8812 1164
rect 8588 746 8616 1158
rect 8576 740 8628 746
rect 8576 682 8628 688
rect 8772 474 8800 1158
rect 8760 468 8812 474
rect 8760 410 8812 416
rect 8956 160 8984 1244
rect 9128 1216 9180 1222
rect 9128 1158 9180 1164
rect 8666 82 8722 160
rect 8496 54 8722 82
rect 8390 0 8446 54
rect 8666 0 8722 54
rect 8942 0 8998 160
rect 9140 134 9168 1158
rect 9232 160 9260 1312
rect 9312 1284 9364 1290
rect 9588 1284 9640 1290
rect 9364 1244 9536 1272
rect 9312 1226 9364 1232
rect 9508 160 9536 1244
rect 9864 1284 9916 1290
rect 9640 1244 9812 1272
rect 9588 1226 9640 1232
rect 9784 160 9812 1244
rect 9864 1226 9916 1232
rect 9876 728 9904 1226
rect 9968 950 9996 1430
rect 10244 950 10272 1430
rect 10416 1284 10468 1290
rect 10416 1226 10468 1232
rect 10324 1216 10376 1222
rect 10324 1158 10376 1164
rect 9956 944 10008 950
rect 9956 886 10008 892
rect 10232 944 10284 950
rect 10232 886 10284 892
rect 9876 700 10088 728
rect 10060 160 10088 700
rect 10336 160 10364 1158
rect 10428 746 10456 1226
rect 10416 740 10468 746
rect 10416 682 10468 688
rect 9128 128 9180 134
rect 9128 70 9180 76
rect 9218 0 9274 160
rect 9494 0 9550 160
rect 9770 0 9826 160
rect 10046 0 10102 160
rect 10322 0 10378 160
rect 10520 66 10548 1822
rect 10690 1799 10746 1808
rect 10796 1562 10824 1935
rect 10784 1556 10836 1562
rect 10784 1498 10836 1504
rect 10612 1414 11100 1442
rect 10612 1358 10640 1414
rect 10600 1352 10652 1358
rect 10600 1294 10652 1300
rect 10692 1284 10744 1290
rect 10744 1244 10916 1272
rect 10692 1226 10744 1232
rect 10600 740 10652 746
rect 10600 682 10652 688
rect 10612 160 10640 682
rect 10888 160 10916 1244
rect 10968 1216 11020 1222
rect 10968 1158 11020 1164
rect 10980 785 11008 1158
rect 10966 776 11022 785
rect 10966 711 11022 720
rect 11072 626 11100 1414
rect 11152 1352 11204 1358
rect 11152 1294 11204 1300
rect 11164 746 11192 1294
rect 11348 1222 11376 4422
rect 11644 4380 11952 4389
rect 11644 4378 11650 4380
rect 11706 4378 11730 4380
rect 11786 4378 11810 4380
rect 11866 4378 11890 4380
rect 11946 4378 11952 4380
rect 11706 4326 11708 4378
rect 11888 4326 11890 4378
rect 11644 4324 11650 4326
rect 11706 4324 11730 4326
rect 11786 4324 11810 4326
rect 11866 4324 11890 4326
rect 11946 4324 11952 4326
rect 11644 4315 11952 4324
rect 11644 3292 11952 3301
rect 11644 3290 11650 3292
rect 11706 3290 11730 3292
rect 11786 3290 11810 3292
rect 11866 3290 11890 3292
rect 11946 3290 11952 3292
rect 11706 3238 11708 3290
rect 11888 3238 11890 3290
rect 11644 3236 11650 3238
rect 11706 3236 11730 3238
rect 11786 3236 11810 3238
rect 11866 3236 11890 3238
rect 11946 3236 11952 3238
rect 11644 3227 11952 3236
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11428 1284 11480 1290
rect 11428 1226 11480 1232
rect 11244 1216 11296 1222
rect 11244 1158 11296 1164
rect 11336 1216 11388 1222
rect 11336 1158 11388 1164
rect 11256 921 11284 1158
rect 11242 912 11298 921
rect 11242 847 11298 856
rect 11152 740 11204 746
rect 11152 682 11204 688
rect 11072 598 11192 626
rect 11164 160 11192 598
rect 11440 160 11468 1226
rect 11532 678 11560 2790
rect 11644 2204 11952 2213
rect 11644 2202 11650 2204
rect 11706 2202 11730 2204
rect 11786 2202 11810 2204
rect 11866 2202 11890 2204
rect 11946 2202 11952 2204
rect 11706 2150 11708 2202
rect 11888 2150 11890 2202
rect 11644 2148 11650 2150
rect 11706 2148 11730 2150
rect 11786 2148 11810 2150
rect 11866 2148 11890 2150
rect 11946 2148 11952 2150
rect 11644 2139 11952 2148
rect 11992 1562 12020 4490
rect 12530 4040 12586 4049
rect 12530 3975 12586 3984
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 12070 2408 12126 2417
rect 12070 2343 12126 2352
rect 11980 1556 12032 1562
rect 11980 1498 12032 1504
rect 11888 1284 11940 1290
rect 11940 1244 12020 1272
rect 11888 1226 11940 1232
rect 11644 1116 11952 1125
rect 11644 1114 11650 1116
rect 11706 1114 11730 1116
rect 11786 1114 11810 1116
rect 11866 1114 11890 1116
rect 11946 1114 11952 1116
rect 11706 1062 11708 1114
rect 11888 1062 11890 1114
rect 11644 1060 11650 1062
rect 11706 1060 11730 1062
rect 11786 1060 11810 1062
rect 11866 1060 11890 1062
rect 11946 1060 11952 1062
rect 11644 1051 11952 1060
rect 11704 740 11756 746
rect 11704 682 11756 688
rect 11520 672 11572 678
rect 11520 614 11572 620
rect 11716 160 11744 682
rect 11992 160 12020 1244
rect 12084 1222 12112 2343
rect 12268 1562 12296 2926
rect 12256 1556 12308 1562
rect 12256 1498 12308 1504
rect 12544 1358 12572 3975
rect 14108 2650 14136 8434
rect 16224 5658 16252 8434
rect 16991 8188 17299 8197
rect 16991 8186 16997 8188
rect 17053 8186 17077 8188
rect 17133 8186 17157 8188
rect 17213 8186 17237 8188
rect 17293 8186 17299 8188
rect 17053 8134 17055 8186
rect 17235 8134 17237 8186
rect 16991 8132 16997 8134
rect 17053 8132 17077 8134
rect 17133 8132 17157 8134
rect 17213 8132 17237 8134
rect 17293 8132 17299 8134
rect 16991 8123 17299 8132
rect 16991 7100 17299 7109
rect 16991 7098 16997 7100
rect 17053 7098 17077 7100
rect 17133 7098 17157 7100
rect 17213 7098 17237 7100
rect 17293 7098 17299 7100
rect 17053 7046 17055 7098
rect 17235 7046 17237 7098
rect 16991 7044 16997 7046
rect 17053 7044 17077 7046
rect 17133 7044 17157 7046
rect 17213 7044 17237 7046
rect 17293 7044 17299 7046
rect 16991 7035 17299 7044
rect 16991 6012 17299 6021
rect 16991 6010 16997 6012
rect 17053 6010 17077 6012
rect 17133 6010 17157 6012
rect 17213 6010 17237 6012
rect 17293 6010 17299 6012
rect 17053 5958 17055 6010
rect 17235 5958 17237 6010
rect 16991 5956 16997 5958
rect 17053 5956 17077 5958
rect 17133 5956 17157 5958
rect 17213 5956 17237 5958
rect 17293 5956 17299 5958
rect 16991 5947 17299 5956
rect 16224 5630 16436 5658
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15382 3632 15438 3641
rect 15382 3567 15438 3576
rect 14370 3224 14426 3233
rect 14370 3159 14426 3168
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 13910 2136 13966 2145
rect 14292 2106 14320 2382
rect 13910 2071 13966 2080
rect 14280 2100 14332 2106
rect 13542 2000 13598 2009
rect 13542 1935 13598 1944
rect 13728 1964 13780 1970
rect 12256 1352 12308 1358
rect 12440 1352 12492 1358
rect 12308 1312 12388 1340
rect 12256 1294 12308 1300
rect 12164 1284 12216 1290
rect 12164 1226 12216 1232
rect 12072 1216 12124 1222
rect 12072 1158 12124 1164
rect 10508 60 10560 66
rect 10508 2 10560 8
rect 10598 0 10654 160
rect 10874 0 10930 160
rect 11150 0 11206 160
rect 11426 0 11482 160
rect 11702 0 11758 160
rect 11978 0 12034 160
rect 12176 82 12204 1226
rect 12254 82 12310 160
rect 12176 54 12310 82
rect 12360 82 12388 1312
rect 12440 1294 12492 1300
rect 12532 1352 12584 1358
rect 12532 1294 12584 1300
rect 13084 1352 13136 1358
rect 13360 1352 13412 1358
rect 13136 1312 13216 1340
rect 13084 1294 13136 1300
rect 12452 218 12480 1294
rect 12992 1284 13044 1290
rect 12992 1226 13044 1232
rect 12900 1216 12952 1222
rect 12900 1158 12952 1164
rect 12716 536 12768 542
rect 12716 478 12768 484
rect 12452 190 12664 218
rect 12728 202 12756 478
rect 12530 82 12586 160
rect 12360 54 12586 82
rect 12636 82 12664 190
rect 12716 196 12768 202
rect 12716 138 12768 144
rect 12806 82 12862 160
rect 12636 54 12862 82
rect 12912 66 12940 1158
rect 13004 82 13032 1226
rect 13082 82 13138 160
rect 12254 0 12310 54
rect 12530 0 12586 54
rect 12806 0 12862 54
rect 12900 60 12952 66
rect 13004 54 13138 82
rect 13188 82 13216 1312
rect 13556 1306 13584 1935
rect 13728 1906 13780 1912
rect 13360 1294 13412 1300
rect 13268 1216 13320 1222
rect 13268 1158 13320 1164
rect 13280 338 13308 1158
rect 13372 746 13400 1294
rect 13464 1278 13584 1306
rect 13464 1222 13492 1278
rect 13452 1216 13504 1222
rect 13452 1158 13504 1164
rect 13544 1216 13596 1222
rect 13544 1158 13596 1164
rect 13360 740 13412 746
rect 13360 682 13412 688
rect 13452 468 13504 474
rect 13452 410 13504 416
rect 13268 332 13320 338
rect 13268 274 13320 280
rect 13358 82 13414 160
rect 13464 134 13492 410
rect 13556 134 13584 1158
rect 13188 54 13414 82
rect 13452 128 13504 134
rect 13452 70 13504 76
rect 13544 128 13596 134
rect 13544 70 13596 76
rect 13634 82 13690 160
rect 13740 82 13768 1906
rect 13924 1562 13952 2071
rect 14280 2042 14332 2048
rect 14384 1970 14412 3159
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14372 1964 14424 1970
rect 14372 1906 14424 1912
rect 14660 1562 14688 2382
rect 15396 2106 15424 3567
rect 15672 2106 15700 4150
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16210 2952 16266 2961
rect 16210 2887 16266 2896
rect 15384 2100 15436 2106
rect 15384 2042 15436 2048
rect 15660 2100 15712 2106
rect 15660 2042 15712 2048
rect 16224 1970 16252 2887
rect 16316 2650 16344 3402
rect 16408 2650 16436 5630
rect 16991 4924 17299 4933
rect 16991 4922 16997 4924
rect 17053 4922 17077 4924
rect 17133 4922 17157 4924
rect 17213 4922 17237 4924
rect 17293 4922 17299 4924
rect 17053 4870 17055 4922
rect 17235 4870 17237 4922
rect 16991 4868 16997 4870
rect 17053 4868 17077 4870
rect 17133 4868 17157 4870
rect 17213 4868 17237 4870
rect 17293 4868 17299 4870
rect 16991 4859 17299 4868
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16316 2106 16344 2382
rect 16500 2106 16528 4218
rect 18234 4040 18290 4049
rect 18234 3975 18290 3984
rect 16991 3836 17299 3845
rect 16991 3834 16997 3836
rect 17053 3834 17077 3836
rect 17133 3834 17157 3836
rect 17213 3834 17237 3836
rect 17293 3834 17299 3836
rect 17053 3782 17055 3834
rect 17235 3782 17237 3834
rect 16991 3780 16997 3782
rect 17053 3780 17077 3782
rect 17133 3780 17157 3782
rect 17213 3780 17237 3782
rect 17293 3780 17299 3782
rect 16991 3771 17299 3780
rect 16854 3496 16910 3505
rect 16854 3431 16910 3440
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 16304 2100 16356 2106
rect 16304 2042 16356 2048
rect 16488 2100 16540 2106
rect 16488 2042 16540 2048
rect 15108 1964 15160 1970
rect 15108 1906 15160 1912
rect 15292 1964 15344 1970
rect 15292 1906 15344 1912
rect 15752 1964 15804 1970
rect 15752 1906 15804 1912
rect 16212 1964 16264 1970
rect 16212 1906 16264 1912
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 16396 1964 16448 1970
rect 16396 1906 16448 1912
rect 14924 1896 14976 1902
rect 14924 1838 14976 1844
rect 14936 1562 14964 1838
rect 13912 1556 13964 1562
rect 13912 1498 13964 1504
rect 14648 1556 14700 1562
rect 14648 1498 14700 1504
rect 14924 1556 14976 1562
rect 14924 1498 14976 1504
rect 14280 1420 14332 1426
rect 14280 1362 14332 1368
rect 13820 1284 13872 1290
rect 13872 1244 14044 1272
rect 13820 1226 13872 1232
rect 13820 740 13872 746
rect 13820 682 13872 688
rect 12900 2 12952 8
rect 13082 0 13138 54
rect 13358 0 13414 54
rect 13634 54 13768 82
rect 13832 82 13860 682
rect 13910 82 13966 160
rect 13832 54 13966 82
rect 14016 82 14044 1244
rect 14186 82 14242 160
rect 14016 54 14242 82
rect 14292 82 14320 1362
rect 14556 1352 14608 1358
rect 14556 1294 14608 1300
rect 15014 1320 15070 1329
rect 14568 746 14596 1294
rect 14740 1284 14792 1290
rect 15014 1255 15070 1264
rect 14740 1226 14792 1232
rect 14556 740 14608 746
rect 14556 682 14608 688
rect 14464 604 14516 610
rect 14464 546 14516 552
rect 14476 270 14504 546
rect 14464 264 14516 270
rect 14464 206 14516 212
rect 14752 160 14780 1226
rect 15028 474 15056 1255
rect 15016 468 15068 474
rect 15016 410 15068 416
rect 14462 82 14518 160
rect 14292 54 14518 82
rect 13634 0 13690 54
rect 13910 0 13966 54
rect 14186 0 14242 54
rect 14462 0 14518 54
rect 14738 0 14794 160
rect 15014 82 15070 160
rect 15120 82 15148 1906
rect 15304 1494 15332 1906
rect 15764 1562 15792 1906
rect 15752 1556 15804 1562
rect 15752 1498 15804 1504
rect 15292 1488 15344 1494
rect 15292 1430 15344 1436
rect 15752 1420 15804 1426
rect 15804 1380 15884 1408
rect 15752 1362 15804 1368
rect 15660 1352 15712 1358
rect 15660 1294 15712 1300
rect 15292 1284 15344 1290
rect 15344 1244 15424 1272
rect 15292 1226 15344 1232
rect 15200 740 15252 746
rect 15200 682 15252 688
rect 15014 54 15148 82
rect 15212 82 15240 682
rect 15290 82 15346 160
rect 15212 54 15346 82
rect 15396 82 15424 1244
rect 15568 1216 15620 1222
rect 15568 1158 15620 1164
rect 15580 882 15608 1158
rect 15568 876 15620 882
rect 15568 818 15620 824
rect 15672 746 15700 1294
rect 15660 740 15712 746
rect 15660 682 15712 688
rect 15856 160 15884 1380
rect 15936 1352 15988 1358
rect 15936 1294 15988 1300
rect 15948 678 15976 1294
rect 16120 1284 16172 1290
rect 16120 1226 16172 1232
rect 15936 672 15988 678
rect 15936 614 15988 620
rect 16132 160 16160 1226
rect 16212 1216 16264 1222
rect 16316 1204 16344 1906
rect 16408 1562 16436 1906
rect 16592 1766 16620 2858
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16580 1760 16632 1766
rect 16580 1702 16632 1708
rect 16396 1556 16448 1562
rect 16776 1544 16804 2382
rect 16868 2106 16896 3431
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 16991 2748 17299 2757
rect 16991 2746 16997 2748
rect 17053 2746 17077 2748
rect 17133 2746 17157 2748
rect 17213 2746 17237 2748
rect 17293 2746 17299 2748
rect 17053 2694 17055 2746
rect 17235 2694 17237 2746
rect 16991 2692 16997 2694
rect 17053 2692 17077 2694
rect 17133 2692 17157 2694
rect 17213 2692 17237 2694
rect 17293 2692 17299 2694
rect 16991 2683 17299 2692
rect 17406 2680 17462 2689
rect 17406 2615 17462 2624
rect 17420 2281 17448 2615
rect 17406 2272 17462 2281
rect 17406 2207 17462 2216
rect 17696 2106 17724 3062
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 16856 2100 16908 2106
rect 16856 2042 16908 2048
rect 17684 2100 17736 2106
rect 17684 2042 17736 2048
rect 16856 1964 16908 1970
rect 16856 1906 16908 1912
rect 17316 1964 17368 1970
rect 17316 1906 17368 1912
rect 17592 1964 17644 1970
rect 17592 1906 17644 1912
rect 16868 1562 16896 1906
rect 16991 1660 17299 1669
rect 16991 1658 16997 1660
rect 17053 1658 17077 1660
rect 17133 1658 17157 1660
rect 17213 1658 17237 1660
rect 17293 1658 17299 1660
rect 17053 1606 17055 1658
rect 17235 1606 17237 1658
rect 16991 1604 16997 1606
rect 17053 1604 17077 1606
rect 17133 1604 17157 1606
rect 17213 1604 17237 1606
rect 17293 1604 17299 1606
rect 16991 1595 17299 1604
rect 16396 1498 16448 1504
rect 16592 1516 16804 1544
rect 16856 1556 16908 1562
rect 16592 1426 16620 1516
rect 16856 1498 16908 1504
rect 17328 1476 17356 1906
rect 17408 1828 17460 1834
rect 17408 1770 17460 1776
rect 17420 1737 17448 1770
rect 17406 1728 17462 1737
rect 17406 1663 17462 1672
rect 17498 1592 17554 1601
rect 17604 1562 17632 1906
rect 17498 1527 17554 1536
rect 17592 1556 17644 1562
rect 17512 1494 17540 1527
rect 17592 1498 17644 1504
rect 17236 1448 17356 1476
rect 17500 1488 17552 1494
rect 16580 1420 16632 1426
rect 16580 1362 16632 1368
rect 16948 1420 17000 1426
rect 17236 1408 17264 1448
rect 17500 1430 17552 1436
rect 17788 1442 17816 2518
rect 17972 1986 18000 3130
rect 17880 1970 18000 1986
rect 17868 1964 18000 1970
rect 17920 1958 18000 1964
rect 18052 1964 18104 1970
rect 17868 1906 17920 1912
rect 18052 1906 18104 1912
rect 17960 1896 18012 1902
rect 18064 1873 18092 1906
rect 17960 1838 18012 1844
rect 18050 1864 18106 1873
rect 17788 1414 17908 1442
rect 17000 1380 17080 1408
rect 16948 1362 17000 1368
rect 16580 1284 16632 1290
rect 16632 1244 16988 1272
rect 16580 1226 16632 1232
rect 16264 1176 16344 1204
rect 16854 1184 16910 1193
rect 16212 1158 16264 1164
rect 16854 1119 16910 1128
rect 16212 808 16264 814
rect 16212 750 16264 756
rect 16224 241 16252 750
rect 16396 740 16448 746
rect 16396 682 16448 688
rect 16210 232 16266 241
rect 16210 167 16266 176
rect 16408 160 16436 682
rect 16672 672 16724 678
rect 16868 649 16896 1119
rect 16672 614 16724 620
rect 16854 640 16910 649
rect 16684 160 16712 614
rect 16854 575 16910 584
rect 16960 160 16988 1244
rect 15566 82 15622 160
rect 15396 54 15622 82
rect 15014 0 15070 54
rect 15290 0 15346 54
rect 15566 0 15622 54
rect 15842 0 15898 160
rect 16118 0 16174 160
rect 16394 0 16450 160
rect 16670 0 16726 160
rect 16946 0 17002 160
rect 17052 82 17080 1380
rect 17144 1380 17264 1408
rect 17144 1222 17172 1380
rect 17224 1284 17276 1290
rect 17276 1244 17356 1272
rect 17224 1226 17276 1232
rect 17132 1216 17184 1222
rect 17132 1158 17184 1164
rect 17222 82 17278 160
rect 17052 54 17278 82
rect 17328 82 17356 1244
rect 17408 1216 17460 1222
rect 17460 1176 17632 1204
rect 17408 1158 17460 1164
rect 17498 82 17554 160
rect 17328 54 17554 82
rect 17604 82 17632 1176
rect 17880 1034 17908 1414
rect 17972 1306 18000 1838
rect 18248 1834 18276 3975
rect 18510 3088 18566 3097
rect 18510 3023 18566 3032
rect 18524 2650 18552 3023
rect 18616 2650 18644 8434
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19432 2848 19484 2854
rect 19484 2796 19564 2802
rect 19432 2790 19564 2796
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 18524 2514 18736 2530
rect 18524 2508 18748 2514
rect 18524 2502 18696 2508
rect 18524 2446 18552 2502
rect 18696 2450 18748 2456
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 18326 2136 18382 2145
rect 18326 2071 18382 2080
rect 18432 2088 18460 2382
rect 18512 2304 18564 2310
rect 18564 2264 18736 2292
rect 18512 2246 18564 2252
rect 18340 1970 18368 2071
rect 18432 2060 18644 2088
rect 18328 1964 18380 1970
rect 18328 1906 18380 1912
rect 18420 1964 18472 1970
rect 18420 1906 18472 1912
rect 18050 1799 18106 1808
rect 18236 1828 18288 1834
rect 18236 1770 18288 1776
rect 18432 1562 18460 1906
rect 18512 1760 18564 1766
rect 18512 1702 18564 1708
rect 18524 1562 18552 1702
rect 18420 1556 18472 1562
rect 18420 1498 18472 1504
rect 18512 1556 18564 1562
rect 18512 1498 18564 1504
rect 18616 1426 18644 2060
rect 18708 1986 18736 2264
rect 18800 2106 18828 2382
rect 18984 2281 19012 2586
rect 19352 2446 19380 2790
rect 19444 2774 19564 2790
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 18970 2272 19026 2281
rect 18970 2207 19026 2216
rect 18788 2100 18840 2106
rect 18788 2042 18840 2048
rect 18708 1958 18828 1986
rect 18800 1902 18828 1958
rect 18788 1896 18840 1902
rect 18788 1838 18840 1844
rect 18880 1760 18932 1766
rect 18880 1702 18932 1708
rect 18052 1420 18104 1426
rect 18604 1420 18656 1426
rect 18104 1380 18368 1408
rect 18052 1362 18104 1368
rect 17972 1290 18184 1306
rect 17972 1284 18196 1290
rect 17972 1278 18144 1284
rect 18144 1226 18196 1232
rect 17960 1216 18012 1222
rect 18236 1216 18288 1222
rect 18012 1176 18092 1204
rect 17960 1158 18012 1164
rect 17958 1048 18014 1057
rect 17880 1006 17958 1034
rect 17958 983 18014 992
rect 18064 160 18092 1176
rect 18236 1158 18288 1164
rect 18248 678 18276 1158
rect 18236 672 18288 678
rect 18236 614 18288 620
rect 18340 160 18368 1380
rect 18604 1362 18656 1368
rect 18420 1352 18472 1358
rect 18420 1294 18472 1300
rect 18512 1352 18564 1358
rect 18512 1294 18564 1300
rect 17774 82 17830 160
rect 17604 54 17830 82
rect 17222 0 17278 54
rect 17498 0 17554 54
rect 17774 0 17830 54
rect 18050 0 18106 160
rect 18326 0 18382 160
rect 18432 82 18460 1294
rect 18524 746 18552 1294
rect 18892 814 18920 1702
rect 19076 1601 19104 2382
rect 19156 1964 19208 1970
rect 19156 1906 19208 1912
rect 19062 1592 19118 1601
rect 19168 1562 19196 1906
rect 19062 1527 19118 1536
rect 19156 1556 19208 1562
rect 19156 1498 19208 1504
rect 19156 1420 19208 1426
rect 19208 1380 19380 1408
rect 19156 1362 19208 1368
rect 19064 1352 19116 1358
rect 19064 1294 19116 1300
rect 19076 1018 19104 1294
rect 19064 1012 19116 1018
rect 19064 954 19116 960
rect 18880 808 18932 814
rect 18880 750 18932 756
rect 18512 740 18564 746
rect 18512 682 18564 688
rect 19156 740 19208 746
rect 19156 682 19208 688
rect 18880 672 18932 678
rect 18880 614 18932 620
rect 18892 160 18920 614
rect 19168 160 19196 682
rect 19352 660 19380 1380
rect 19536 1358 19564 2774
rect 20456 2774 20484 8434
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 20456 2746 20576 2774
rect 20548 2650 20576 2746
rect 20536 2644 20588 2650
rect 20536 2586 20588 2592
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 19800 2576 19852 2582
rect 19800 2518 19852 2524
rect 19616 1760 19668 1766
rect 19616 1702 19668 1708
rect 19708 1760 19760 1766
rect 19708 1702 19760 1708
rect 19628 1358 19656 1702
rect 19524 1352 19576 1358
rect 19524 1294 19576 1300
rect 19616 1352 19668 1358
rect 19616 1294 19668 1300
rect 19432 1216 19484 1222
rect 19432 1158 19484 1164
rect 19444 1018 19472 1158
rect 19432 1012 19484 1018
rect 19432 954 19484 960
rect 19352 632 19472 660
rect 19444 160 19472 632
rect 19720 160 19748 1702
rect 19812 1358 19840 2518
rect 20824 2446 20852 2586
rect 21468 2446 21496 3334
rect 21546 3224 21602 3233
rect 21546 3159 21602 3168
rect 21560 2961 21588 3159
rect 21546 2952 21602 2961
rect 22112 2922 22140 8502
rect 22928 8492 22980 8498
rect 22928 8434 22980 8440
rect 22338 7644 22646 7653
rect 22338 7642 22344 7644
rect 22400 7642 22424 7644
rect 22480 7642 22504 7644
rect 22560 7642 22584 7644
rect 22640 7642 22646 7644
rect 22400 7590 22402 7642
rect 22582 7590 22584 7642
rect 22338 7588 22344 7590
rect 22400 7588 22424 7590
rect 22480 7588 22504 7590
rect 22560 7588 22584 7590
rect 22640 7588 22646 7590
rect 22338 7579 22646 7588
rect 22338 6556 22646 6565
rect 22338 6554 22344 6556
rect 22400 6554 22424 6556
rect 22480 6554 22504 6556
rect 22560 6554 22584 6556
rect 22640 6554 22646 6556
rect 22400 6502 22402 6554
rect 22582 6502 22584 6554
rect 22338 6500 22344 6502
rect 22400 6500 22424 6502
rect 22480 6500 22504 6502
rect 22560 6500 22584 6502
rect 22640 6500 22646 6502
rect 22338 6491 22646 6500
rect 22338 5468 22646 5477
rect 22338 5466 22344 5468
rect 22400 5466 22424 5468
rect 22480 5466 22504 5468
rect 22560 5466 22584 5468
rect 22640 5466 22646 5468
rect 22400 5414 22402 5466
rect 22582 5414 22584 5466
rect 22338 5412 22344 5414
rect 22400 5412 22424 5414
rect 22480 5412 22504 5414
rect 22560 5412 22584 5414
rect 22640 5412 22646 5414
rect 22338 5403 22646 5412
rect 22338 4380 22646 4389
rect 22338 4378 22344 4380
rect 22400 4378 22424 4380
rect 22480 4378 22504 4380
rect 22560 4378 22584 4380
rect 22640 4378 22646 4380
rect 22400 4326 22402 4378
rect 22582 4326 22584 4378
rect 22338 4324 22344 4326
rect 22400 4324 22424 4326
rect 22480 4324 22504 4326
rect 22560 4324 22584 4326
rect 22640 4324 22646 4326
rect 22338 4315 22646 4324
rect 22338 3292 22646 3301
rect 22338 3290 22344 3292
rect 22400 3290 22424 3292
rect 22480 3290 22504 3292
rect 22560 3290 22584 3292
rect 22640 3290 22646 3292
rect 22400 3238 22402 3290
rect 22582 3238 22584 3290
rect 22338 3236 22344 3238
rect 22400 3236 22424 3238
rect 22480 3236 22504 3238
rect 22560 3236 22584 3238
rect 22640 3236 22646 3238
rect 22338 3227 22646 3236
rect 21546 2887 21602 2896
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 22940 2650 22968 8434
rect 23296 8356 23348 8362
rect 23296 8298 23348 8304
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 22374 2544 22430 2553
rect 22374 2479 22430 2488
rect 22388 2446 22416 2479
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 21272 2440 21324 2446
rect 21456 2440 21508 2446
rect 21324 2400 21404 2428
rect 21272 2382 21324 2388
rect 19892 2304 19944 2310
rect 19892 2246 19944 2252
rect 19904 1494 19932 2246
rect 19984 1760 20036 1766
rect 19984 1702 20036 1708
rect 19892 1488 19944 1494
rect 19892 1430 19944 1436
rect 19800 1352 19852 1358
rect 19800 1294 19852 1300
rect 19892 1216 19944 1222
rect 19892 1158 19944 1164
rect 19904 474 19932 1158
rect 19892 468 19944 474
rect 19892 410 19944 416
rect 19996 160 20024 1702
rect 20088 241 20116 2382
rect 20180 746 20208 2382
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 20456 2038 20484 2246
rect 20536 2100 20588 2106
rect 20536 2042 20588 2048
rect 20732 2094 20944 2122
rect 20444 2032 20496 2038
rect 20444 1974 20496 1980
rect 20548 1290 20576 2042
rect 20536 1284 20588 1290
rect 20536 1226 20588 1232
rect 20352 1216 20404 1222
rect 20352 1158 20404 1164
rect 20444 1216 20496 1222
rect 20444 1158 20496 1164
rect 20168 740 20220 746
rect 20168 682 20220 688
rect 20260 468 20312 474
rect 20260 410 20312 416
rect 20074 232 20130 241
rect 20074 167 20130 176
rect 20272 160 20300 410
rect 18602 82 18658 160
rect 18432 54 18658 82
rect 18602 0 18658 54
rect 18878 0 18934 160
rect 19154 0 19210 160
rect 19430 0 19486 160
rect 19706 0 19762 160
rect 19982 0 20038 160
rect 20258 0 20314 160
rect 20364 82 20392 1158
rect 20456 678 20484 1158
rect 20444 672 20496 678
rect 20444 614 20496 620
rect 20732 474 20760 2094
rect 20916 1970 20944 2094
rect 20812 1964 20864 1970
rect 20812 1906 20864 1912
rect 20904 1964 20956 1970
rect 20904 1906 20956 1912
rect 20824 1329 20852 1906
rect 20904 1760 20956 1766
rect 20904 1702 20956 1708
rect 20916 1358 20944 1702
rect 20904 1352 20956 1358
rect 20810 1320 20866 1329
rect 20904 1294 20956 1300
rect 20810 1255 20866 1264
rect 20812 1216 20864 1222
rect 20812 1158 20864 1164
rect 20720 468 20772 474
rect 20720 410 20772 416
rect 20824 160 20852 1158
rect 21008 513 21036 2382
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 21088 1760 21140 1766
rect 21088 1702 21140 1708
rect 20994 504 21050 513
rect 20994 439 21050 448
rect 21100 160 21128 1702
rect 21284 1358 21312 2246
rect 21272 1352 21324 1358
rect 21272 1294 21324 1300
rect 21376 762 21404 2400
rect 21456 2382 21508 2388
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 22744 2440 22796 2446
rect 22744 2382 22796 2388
rect 21548 2304 21600 2310
rect 21548 2246 21600 2252
rect 22008 2304 22060 2310
rect 22008 2246 22060 2252
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 21376 734 21496 762
rect 21180 672 21232 678
rect 21232 632 21404 660
rect 21180 614 21232 620
rect 21376 160 21404 632
rect 21468 270 21496 734
rect 21456 264 21508 270
rect 21456 206 21508 212
rect 20534 82 20590 160
rect 20364 54 20590 82
rect 20534 0 20590 54
rect 20810 0 20866 160
rect 21086 0 21142 160
rect 21362 0 21418 160
rect 21560 82 21588 2246
rect 21916 1760 21968 1766
rect 21916 1702 21968 1708
rect 21730 1320 21786 1329
rect 21730 1255 21786 1264
rect 21744 406 21772 1255
rect 21822 1048 21878 1057
rect 21822 983 21878 992
rect 21836 513 21864 983
rect 21822 504 21878 513
rect 21822 439 21878 448
rect 21732 400 21784 406
rect 21732 342 21784 348
rect 21928 160 21956 1702
rect 22020 1358 22048 2246
rect 22204 1578 22232 2246
rect 22338 2204 22646 2213
rect 22338 2202 22344 2204
rect 22400 2202 22424 2204
rect 22480 2202 22504 2204
rect 22560 2202 22584 2204
rect 22640 2202 22646 2204
rect 22400 2150 22402 2202
rect 22582 2150 22584 2202
rect 22338 2148 22344 2150
rect 22400 2148 22424 2150
rect 22480 2148 22504 2150
rect 22560 2148 22584 2150
rect 22640 2148 22646 2150
rect 22338 2139 22646 2148
rect 22204 1550 22324 1578
rect 22296 1494 22324 1550
rect 22284 1488 22336 1494
rect 22284 1430 22336 1436
rect 22192 1420 22244 1426
rect 22192 1362 22244 1368
rect 22008 1352 22060 1358
rect 22008 1294 22060 1300
rect 22100 1216 22152 1222
rect 22100 1158 22152 1164
rect 22112 950 22140 1158
rect 22100 944 22152 950
rect 22100 886 22152 892
rect 22204 160 22232 1362
rect 22756 1358 22784 2382
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 23112 2100 23164 2106
rect 23112 2042 23164 2048
rect 22928 1964 22980 1970
rect 22928 1906 22980 1912
rect 22836 1828 22888 1834
rect 22836 1770 22888 1776
rect 22848 1494 22876 1770
rect 22836 1488 22888 1494
rect 22940 1465 22968 1906
rect 23020 1828 23072 1834
rect 23020 1770 23072 1776
rect 22836 1430 22888 1436
rect 22926 1456 22982 1465
rect 22926 1391 22982 1400
rect 22744 1352 22796 1358
rect 22744 1294 22796 1300
rect 22744 1216 22796 1222
rect 22744 1158 22796 1164
rect 22928 1216 22980 1222
rect 23032 1193 23060 1770
rect 23124 1601 23152 2042
rect 23110 1592 23166 1601
rect 23110 1527 23166 1536
rect 23216 1358 23244 2246
rect 23308 2145 23336 8298
rect 23480 4684 23532 4690
rect 23480 4626 23532 4632
rect 23294 2136 23350 2145
rect 23294 2071 23350 2080
rect 23492 1970 23520 4626
rect 23584 2650 23612 8774
rect 24688 8634 24716 9030
rect 26712 8634 26740 9840
rect 28828 9058 28856 9840
rect 28828 9030 28948 9058
rect 28920 8634 28948 9030
rect 30944 8634 30972 9840
rect 33060 9058 33088 9840
rect 32968 9030 33088 9058
rect 32968 8634 32996 9030
rect 33032 8732 33340 8741
rect 33032 8730 33038 8732
rect 33094 8730 33118 8732
rect 33174 8730 33198 8732
rect 33254 8730 33278 8732
rect 33334 8730 33340 8732
rect 33094 8678 33096 8730
rect 33276 8678 33278 8730
rect 33032 8676 33038 8678
rect 33094 8676 33118 8678
rect 33174 8676 33198 8678
rect 33254 8676 33278 8678
rect 33334 8676 33340 8678
rect 33032 8667 33340 8676
rect 35176 8634 35204 9840
rect 37292 9058 37320 9840
rect 37292 9030 37504 9058
rect 37476 8634 37504 9030
rect 39408 8634 39436 9840
rect 41524 8634 41552 9840
rect 43640 8634 43668 9840
rect 43726 8732 44034 8741
rect 43726 8730 43732 8732
rect 43788 8730 43812 8732
rect 43868 8730 43892 8732
rect 43948 8730 43972 8732
rect 44028 8730 44034 8732
rect 43788 8678 43790 8730
rect 43970 8678 43972 8730
rect 43726 8676 43732 8678
rect 43788 8676 43812 8678
rect 43868 8676 43892 8678
rect 43948 8676 43972 8678
rect 44028 8676 44034 8678
rect 43726 8667 44034 8676
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 26700 8628 26752 8634
rect 26700 8570 26752 8576
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 30932 8628 30984 8634
rect 30932 8570 30984 8576
rect 32956 8628 33008 8634
rect 32956 8570 33008 8576
rect 35164 8628 35216 8634
rect 35164 8570 35216 8576
rect 37464 8628 37516 8634
rect 37464 8570 37516 8576
rect 39396 8628 39448 8634
rect 39396 8570 39448 8576
rect 41512 8628 41564 8634
rect 41512 8570 41564 8576
rect 43628 8628 43680 8634
rect 43628 8570 43680 8576
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 26976 8492 27028 8498
rect 26976 8434 27028 8440
rect 30104 8492 30156 8498
rect 30104 8434 30156 8440
rect 31024 8492 31076 8498
rect 31024 8434 31076 8440
rect 33508 8492 33560 8498
rect 33508 8434 33560 8440
rect 37372 8492 37424 8498
rect 37372 8434 37424 8440
rect 39948 8492 40000 8498
rect 39948 8434 40000 8440
rect 40684 8492 40736 8498
rect 40684 8434 40736 8440
rect 43260 8492 43312 8498
rect 43260 8434 43312 8440
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 23572 2644 23624 2650
rect 23572 2586 23624 2592
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 23584 2106 23612 2382
rect 23848 2372 23900 2378
rect 23848 2314 23900 2320
rect 23572 2100 23624 2106
rect 23572 2042 23624 2048
rect 23388 1964 23440 1970
rect 23388 1906 23440 1912
rect 23480 1964 23532 1970
rect 23480 1906 23532 1912
rect 23756 1964 23808 1970
rect 23756 1906 23808 1912
rect 23296 1556 23348 1562
rect 23296 1498 23348 1504
rect 23204 1352 23256 1358
rect 23204 1294 23256 1300
rect 23112 1216 23164 1222
rect 22928 1158 22980 1164
rect 23018 1184 23074 1193
rect 22338 1116 22646 1125
rect 22338 1114 22344 1116
rect 22400 1114 22424 1116
rect 22480 1114 22504 1116
rect 22560 1114 22584 1116
rect 22640 1114 22646 1116
rect 22400 1062 22402 1114
rect 22582 1062 22584 1114
rect 22338 1060 22344 1062
rect 22400 1060 22424 1062
rect 22480 1060 22504 1062
rect 22560 1060 22584 1062
rect 22640 1060 22646 1062
rect 22338 1051 22646 1060
rect 22468 944 22520 950
rect 22468 886 22520 892
rect 22480 160 22508 886
rect 22756 160 22784 1158
rect 22940 202 22968 1158
rect 23112 1158 23164 1164
rect 23018 1119 23074 1128
rect 22928 196 22980 202
rect 21638 82 21694 160
rect 21560 54 21694 82
rect 21638 0 21694 54
rect 21914 0 21970 160
rect 22190 0 22246 160
rect 22466 0 22522 160
rect 22742 0 22798 160
rect 22928 138 22980 144
rect 23018 82 23074 160
rect 23124 82 23152 1158
rect 23308 160 23336 1498
rect 23400 542 23428 1906
rect 23662 1728 23718 1737
rect 23662 1663 23718 1672
rect 23572 1216 23624 1222
rect 23572 1158 23624 1164
rect 23388 536 23440 542
rect 23388 478 23440 484
rect 23584 160 23612 1158
rect 23676 746 23704 1663
rect 23664 740 23716 746
rect 23664 682 23716 688
rect 23768 649 23796 1906
rect 23860 1465 23888 2314
rect 23952 2106 23980 4558
rect 24676 2916 24728 2922
rect 24676 2858 24728 2864
rect 23940 2100 23992 2106
rect 23940 2042 23992 2048
rect 24228 2094 24532 2122
rect 24228 1970 24256 2094
rect 24216 1964 24268 1970
rect 24216 1906 24268 1912
rect 24308 1964 24360 1970
rect 24308 1906 24360 1912
rect 24032 1760 24084 1766
rect 24032 1702 24084 1708
rect 24124 1760 24176 1766
rect 24320 1714 24348 1906
rect 24398 1864 24454 1873
rect 24398 1799 24454 1808
rect 24124 1702 24176 1708
rect 23938 1592 23994 1601
rect 23938 1527 23994 1536
rect 23952 1494 23980 1527
rect 23940 1488 23992 1494
rect 23846 1456 23902 1465
rect 23940 1430 23992 1436
rect 23846 1391 23902 1400
rect 23860 1290 23980 1306
rect 23860 1284 23992 1290
rect 23860 1278 23940 1284
rect 23754 640 23810 649
rect 23754 575 23810 584
rect 23860 160 23888 1278
rect 23940 1226 23992 1232
rect 24044 950 24072 1702
rect 24136 1494 24164 1702
rect 24228 1686 24348 1714
rect 24124 1488 24176 1494
rect 24124 1430 24176 1436
rect 24228 1329 24256 1686
rect 24308 1556 24360 1562
rect 24308 1498 24360 1504
rect 24214 1320 24270 1329
rect 24214 1255 24270 1264
rect 24032 944 24084 950
rect 24032 886 24084 892
rect 23018 54 23152 82
rect 23018 0 23074 54
rect 23294 0 23350 160
rect 23570 0 23626 160
rect 23846 0 23902 160
rect 24122 82 24178 160
rect 24320 82 24348 1498
rect 24412 1494 24440 1799
rect 24400 1488 24452 1494
rect 24400 1430 24452 1436
rect 24504 542 24532 2094
rect 24688 1970 24716 2858
rect 24950 2680 25006 2689
rect 25056 2650 25084 8434
rect 26332 8424 26384 8430
rect 26332 8366 26384 8372
rect 26148 3188 26200 3194
rect 26148 3130 26200 3136
rect 26160 3097 26188 3130
rect 26146 3088 26202 3097
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 26056 3052 26108 3058
rect 26146 3023 26202 3032
rect 26056 2994 26108 3000
rect 25228 2916 25280 2922
rect 25228 2858 25280 2864
rect 24950 2615 24952 2624
rect 25004 2615 25006 2624
rect 25044 2644 25096 2650
rect 24952 2586 25004 2592
rect 25044 2586 25096 2592
rect 25240 2582 25268 2858
rect 25320 2848 25372 2854
rect 25320 2790 25372 2796
rect 25228 2576 25280 2582
rect 25228 2518 25280 2524
rect 25332 2446 25360 2790
rect 25320 2440 25372 2446
rect 25320 2382 25372 2388
rect 24768 2100 24820 2106
rect 24820 2060 24992 2088
rect 24768 2042 24820 2048
rect 24964 1970 24992 2060
rect 24676 1964 24728 1970
rect 24676 1906 24728 1912
rect 24952 1964 25004 1970
rect 24952 1906 25004 1912
rect 25228 1964 25280 1970
rect 25228 1906 25280 1912
rect 25240 1850 25268 1906
rect 24768 1828 24820 1834
rect 24768 1770 24820 1776
rect 24860 1828 24912 1834
rect 24964 1822 25268 1850
rect 25320 1896 25372 1902
rect 25320 1838 25372 1844
rect 24964 1816 24992 1822
rect 24912 1788 24992 1816
rect 24860 1770 24912 1776
rect 24676 1760 24728 1766
rect 24676 1702 24728 1708
rect 24688 1601 24716 1702
rect 24674 1592 24730 1601
rect 24674 1527 24730 1536
rect 24676 1488 24728 1494
rect 24596 1448 24676 1476
rect 24492 536 24544 542
rect 24492 478 24544 484
rect 24596 388 24624 1448
rect 24676 1430 24728 1436
rect 24676 1352 24728 1358
rect 24780 1340 24808 1770
rect 25228 1760 25280 1766
rect 25228 1702 25280 1708
rect 25136 1420 25188 1426
rect 25136 1362 25188 1368
rect 24728 1312 24808 1340
rect 24676 1294 24728 1300
rect 24952 1284 25004 1290
rect 24952 1226 25004 1232
rect 24768 1216 24820 1222
rect 24768 1158 24820 1164
rect 24412 360 24624 388
rect 24412 160 24440 360
rect 24122 54 24348 82
rect 24122 0 24178 54
rect 24398 0 24454 160
rect 24674 82 24730 160
rect 24780 82 24808 1158
rect 24964 950 24992 1226
rect 24952 944 25004 950
rect 24952 886 25004 892
rect 24674 54 24808 82
rect 24950 82 25006 160
rect 25148 82 25176 1362
rect 25240 160 25268 1702
rect 25332 882 25360 1838
rect 25320 876 25372 882
rect 25320 818 25372 824
rect 25424 202 25452 2994
rect 25872 2916 25924 2922
rect 25872 2858 25924 2864
rect 25884 2582 25912 2858
rect 26068 2689 26096 2994
rect 26146 2952 26202 2961
rect 26146 2887 26202 2896
rect 26054 2680 26110 2689
rect 26054 2615 26110 2624
rect 25596 2576 25648 2582
rect 25596 2518 25648 2524
rect 25872 2576 25924 2582
rect 25872 2518 25924 2524
rect 25608 2106 25636 2518
rect 25964 2440 26016 2446
rect 25964 2382 26016 2388
rect 25596 2100 25648 2106
rect 25596 2042 25648 2048
rect 25872 1760 25924 1766
rect 25792 1720 25872 1748
rect 25502 640 25558 649
rect 25502 575 25558 584
rect 25412 196 25464 202
rect 24950 54 25176 82
rect 24674 0 24730 54
rect 24950 0 25006 54
rect 25226 0 25282 160
rect 25516 160 25544 575
rect 25792 160 25820 1720
rect 25872 1702 25924 1708
rect 25976 1544 26004 2382
rect 26056 2032 26108 2038
rect 26056 1974 26108 1980
rect 25884 1516 26004 1544
rect 25884 882 25912 1516
rect 26068 1442 26096 1974
rect 25976 1414 26096 1442
rect 25872 876 25924 882
rect 25872 818 25924 824
rect 25412 138 25464 144
rect 25502 0 25558 160
rect 25778 0 25834 160
rect 25976 134 26004 1414
rect 26056 944 26108 950
rect 26056 886 26108 892
rect 26068 160 26096 886
rect 26160 270 26188 2887
rect 26240 2848 26292 2854
rect 26240 2790 26292 2796
rect 26252 2310 26280 2790
rect 26344 2650 26372 8366
rect 26424 2848 26476 2854
rect 26424 2790 26476 2796
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 26436 2446 26464 2790
rect 26988 2774 27016 8434
rect 27685 8188 27993 8197
rect 27685 8186 27691 8188
rect 27747 8186 27771 8188
rect 27827 8186 27851 8188
rect 27907 8186 27931 8188
rect 27987 8186 27993 8188
rect 27747 8134 27749 8186
rect 27929 8134 27931 8186
rect 27685 8132 27691 8134
rect 27747 8132 27771 8134
rect 27827 8132 27851 8134
rect 27907 8132 27931 8134
rect 27987 8132 27993 8134
rect 27685 8123 27993 8132
rect 27685 7100 27993 7109
rect 27685 7098 27691 7100
rect 27747 7098 27771 7100
rect 27827 7098 27851 7100
rect 27907 7098 27931 7100
rect 27987 7098 27993 7100
rect 27747 7046 27749 7098
rect 27929 7046 27931 7098
rect 27685 7044 27691 7046
rect 27747 7044 27771 7046
rect 27827 7044 27851 7046
rect 27907 7044 27931 7046
rect 27987 7044 27993 7046
rect 27685 7035 27993 7044
rect 27685 6012 27993 6021
rect 27685 6010 27691 6012
rect 27747 6010 27771 6012
rect 27827 6010 27851 6012
rect 27907 6010 27931 6012
rect 27987 6010 27993 6012
rect 27747 5958 27749 6010
rect 27929 5958 27931 6010
rect 27685 5956 27691 5958
rect 27747 5956 27771 5958
rect 27827 5956 27851 5958
rect 27907 5956 27931 5958
rect 27987 5956 27993 5958
rect 27685 5947 27993 5956
rect 27685 4924 27993 4933
rect 27685 4922 27691 4924
rect 27747 4922 27771 4924
rect 27827 4922 27851 4924
rect 27907 4922 27931 4924
rect 27987 4922 27993 4924
rect 27747 4870 27749 4922
rect 27929 4870 27931 4922
rect 27685 4868 27691 4870
rect 27747 4868 27771 4870
rect 27827 4868 27851 4870
rect 27907 4868 27931 4870
rect 27987 4868 27993 4870
rect 27685 4859 27993 4868
rect 28080 4548 28132 4554
rect 28080 4490 28132 4496
rect 27685 3836 27993 3845
rect 27685 3834 27691 3836
rect 27747 3834 27771 3836
rect 27827 3834 27851 3836
rect 27907 3834 27931 3836
rect 27987 3834 27993 3836
rect 27747 3782 27749 3834
rect 27929 3782 27931 3834
rect 27685 3780 27691 3782
rect 27747 3780 27771 3782
rect 27827 3780 27851 3782
rect 27907 3780 27931 3782
rect 27987 3780 27993 3782
rect 27526 3768 27582 3777
rect 27685 3771 27993 3780
rect 27582 3726 27660 3754
rect 27526 3703 27582 3712
rect 27632 2990 27660 3726
rect 28092 3058 28120 4490
rect 28816 4480 28868 4486
rect 28816 4422 28868 4428
rect 28828 3058 28856 4422
rect 29920 3188 29972 3194
rect 29920 3130 29972 3136
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 28264 3052 28316 3058
rect 28264 2994 28316 3000
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 27620 2984 27672 2990
rect 27250 2952 27306 2961
rect 27620 2926 27672 2932
rect 28276 2938 28304 2994
rect 28906 2952 28962 2961
rect 27250 2887 27306 2896
rect 27436 2916 27488 2922
rect 27264 2854 27292 2887
rect 28276 2910 28488 2938
rect 27436 2858 27488 2864
rect 27252 2848 27304 2854
rect 27252 2790 27304 2796
rect 26988 2746 27200 2774
rect 26528 2638 26832 2666
rect 27172 2650 27200 2746
rect 27342 2680 27398 2689
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 26240 2304 26292 2310
rect 26240 2246 26292 2252
rect 26344 1986 26372 2382
rect 26344 1958 26464 1986
rect 26332 1896 26384 1902
rect 26332 1838 26384 1844
rect 26238 1592 26294 1601
rect 26238 1527 26294 1536
rect 26252 1494 26280 1527
rect 26240 1488 26292 1494
rect 26240 1430 26292 1436
rect 26148 264 26200 270
rect 26148 206 26200 212
rect 26344 160 26372 1838
rect 25964 128 26016 134
rect 25964 70 26016 76
rect 26054 0 26110 160
rect 26330 0 26386 160
rect 26436 134 26464 1958
rect 26528 338 26556 2638
rect 26608 2508 26660 2514
rect 26608 2450 26660 2456
rect 26620 1970 26648 2450
rect 26804 2446 26832 2638
rect 27160 2644 27212 2650
rect 27342 2615 27344 2624
rect 27160 2586 27212 2592
rect 27396 2615 27398 2624
rect 27344 2586 27396 2592
rect 27448 2446 27476 2858
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 27685 2748 27993 2757
rect 27685 2746 27691 2748
rect 27747 2746 27771 2748
rect 27827 2746 27851 2748
rect 27907 2746 27931 2748
rect 27987 2746 27993 2748
rect 27747 2694 27749 2746
rect 27929 2694 27931 2746
rect 27685 2692 27691 2694
rect 27747 2692 27771 2694
rect 27827 2692 27851 2694
rect 27907 2692 27931 2694
rect 27987 2692 27993 2694
rect 27685 2683 27993 2692
rect 28092 2446 28120 2790
rect 26792 2440 26844 2446
rect 26792 2382 26844 2388
rect 26976 2440 27028 2446
rect 26976 2382 27028 2388
rect 27436 2440 27488 2446
rect 27436 2382 27488 2388
rect 28080 2440 28132 2446
rect 28080 2382 28132 2388
rect 28172 2440 28224 2446
rect 28172 2382 28224 2388
rect 26700 2304 26752 2310
rect 26700 2246 26752 2252
rect 26792 2304 26844 2310
rect 26792 2246 26844 2252
rect 26712 2106 26740 2246
rect 26700 2100 26752 2106
rect 26700 2042 26752 2048
rect 26608 1964 26660 1970
rect 26608 1906 26660 1912
rect 26608 1760 26660 1766
rect 26608 1702 26660 1708
rect 26620 1329 26648 1702
rect 26700 1488 26752 1494
rect 26700 1430 26752 1436
rect 26606 1320 26662 1329
rect 26606 1255 26662 1264
rect 26516 332 26568 338
rect 26516 274 26568 280
rect 26424 128 26476 134
rect 26424 70 26476 76
rect 26606 82 26662 160
rect 26712 82 26740 1430
rect 26804 746 26832 2246
rect 26884 1488 26936 1494
rect 26884 1430 26936 1436
rect 26792 740 26844 746
rect 26792 682 26844 688
rect 26896 160 26924 1430
rect 26606 54 26740 82
rect 26606 0 26662 54
rect 26882 0 26938 160
rect 26988 66 27016 2382
rect 27804 2304 27856 2310
rect 27802 2272 27804 2281
rect 27988 2304 28040 2310
rect 27856 2272 27858 2281
rect 27988 2246 28040 2252
rect 27802 2207 27858 2216
rect 28000 2106 28028 2246
rect 27988 2100 28040 2106
rect 27988 2042 28040 2048
rect 28184 1986 28212 2382
rect 28264 2304 28316 2310
rect 28264 2246 28316 2252
rect 27356 1958 28212 1986
rect 27160 1828 27212 1834
rect 27160 1770 27212 1776
rect 27172 1358 27200 1770
rect 27356 1737 27384 1958
rect 27436 1896 27488 1902
rect 27434 1864 27436 1873
rect 27488 1864 27490 1873
rect 27434 1799 27490 1808
rect 27436 1760 27488 1766
rect 27342 1728 27398 1737
rect 27436 1702 27488 1708
rect 28172 1760 28224 1766
rect 28172 1702 28224 1708
rect 27342 1663 27398 1672
rect 27160 1352 27212 1358
rect 27160 1294 27212 1300
rect 27344 1012 27396 1018
rect 27344 954 27396 960
rect 27356 626 27384 954
rect 27172 598 27384 626
rect 27172 160 27200 598
rect 27448 160 27476 1702
rect 27685 1660 27993 1669
rect 27685 1658 27691 1660
rect 27747 1658 27771 1660
rect 27827 1658 27851 1660
rect 27907 1658 27931 1660
rect 27987 1658 27993 1660
rect 27747 1606 27749 1658
rect 27929 1606 27931 1658
rect 27685 1604 27691 1606
rect 27747 1604 27771 1606
rect 27827 1604 27851 1606
rect 27907 1604 27931 1606
rect 27987 1604 27993 1606
rect 27685 1595 27993 1604
rect 27620 1556 27672 1562
rect 28184 1544 28212 1702
rect 27620 1498 27672 1504
rect 27724 1516 28212 1544
rect 27632 950 27660 1498
rect 27620 944 27672 950
rect 27620 886 27672 892
rect 27724 160 27752 1516
rect 28080 1420 28132 1426
rect 28080 1362 28132 1368
rect 27804 1352 27856 1358
rect 27802 1320 27804 1329
rect 27856 1320 27858 1329
rect 27802 1255 27858 1264
rect 27896 1216 27948 1222
rect 27896 1158 27948 1164
rect 27908 649 27936 1158
rect 27894 640 27950 649
rect 27894 575 27950 584
rect 26976 60 27028 66
rect 26976 2 27028 8
rect 27158 0 27214 160
rect 27434 0 27490 160
rect 27710 0 27766 160
rect 27986 82 28042 160
rect 28092 82 28120 1362
rect 28276 160 28304 2246
rect 28368 1970 28396 2790
rect 28460 1970 28488 2910
rect 28906 2887 28962 2896
rect 28632 2848 28684 2854
rect 28632 2790 28684 2796
rect 28644 2038 28672 2790
rect 28724 2304 28776 2310
rect 28920 2292 28948 2887
rect 29368 2848 29420 2854
rect 29196 2796 29368 2802
rect 29196 2790 29420 2796
rect 29196 2774 29408 2790
rect 29196 2666 29224 2774
rect 29012 2638 29224 2666
rect 29012 2446 29040 2638
rect 29000 2440 29052 2446
rect 29184 2440 29236 2446
rect 29000 2382 29052 2388
rect 29182 2408 29184 2417
rect 29236 2408 29238 2417
rect 29092 2372 29144 2378
rect 29182 2343 29238 2352
rect 29092 2314 29144 2320
rect 28920 2264 29040 2292
rect 28724 2246 28776 2252
rect 28736 2145 28764 2246
rect 28722 2136 28778 2145
rect 28908 2100 28960 2106
rect 28722 2071 28778 2080
rect 28828 2060 28908 2088
rect 28632 2032 28684 2038
rect 28632 1974 28684 1980
rect 28356 1964 28408 1970
rect 28356 1906 28408 1912
rect 28448 1964 28500 1970
rect 28448 1906 28500 1912
rect 28356 1828 28408 1834
rect 28632 1828 28684 1834
rect 28408 1788 28488 1816
rect 28356 1770 28408 1776
rect 28356 1556 28408 1562
rect 28356 1498 28408 1504
rect 28368 921 28396 1498
rect 28460 1494 28488 1788
rect 28552 1788 28632 1816
rect 28448 1488 28500 1494
rect 28448 1430 28500 1436
rect 28354 912 28410 921
rect 28354 847 28410 856
rect 28552 160 28580 1788
rect 28632 1770 28684 1776
rect 28828 1442 28856 2060
rect 28908 2042 28960 2048
rect 29012 1970 29040 2264
rect 28908 1964 28960 1970
rect 28908 1906 28960 1912
rect 29000 1964 29052 1970
rect 29000 1906 29052 1912
rect 28920 1714 28948 1906
rect 28920 1686 29040 1714
rect 28736 1414 28856 1442
rect 28908 1488 28960 1494
rect 28908 1430 28960 1436
rect 28736 1193 28764 1414
rect 28816 1352 28868 1358
rect 28816 1294 28868 1300
rect 28828 1222 28856 1294
rect 28816 1216 28868 1222
rect 28722 1184 28778 1193
rect 28816 1158 28868 1164
rect 28722 1119 28778 1128
rect 28828 678 28856 1158
rect 28816 672 28868 678
rect 28816 614 28868 620
rect 27986 54 28120 82
rect 27986 0 28042 54
rect 28262 0 28318 160
rect 28538 0 28594 160
rect 28814 82 28870 160
rect 28920 82 28948 1430
rect 29012 950 29040 1686
rect 29104 1562 29132 2314
rect 29552 2304 29604 2310
rect 29552 2246 29604 2252
rect 29828 2304 29880 2310
rect 29828 2246 29880 2252
rect 29368 1828 29420 1834
rect 29288 1788 29368 1816
rect 29092 1556 29144 1562
rect 29092 1498 29144 1504
rect 29000 944 29052 950
rect 29000 886 29052 892
rect 28814 54 28948 82
rect 29090 82 29146 160
rect 29288 82 29316 1788
rect 29368 1770 29420 1776
rect 29460 1556 29512 1562
rect 29380 1516 29460 1544
rect 29380 160 29408 1516
rect 29460 1498 29512 1504
rect 29564 1358 29592 2246
rect 29840 2106 29868 2246
rect 29828 2100 29880 2106
rect 29828 2042 29880 2048
rect 29644 1760 29696 1766
rect 29644 1702 29696 1708
rect 29552 1352 29604 1358
rect 29552 1294 29604 1300
rect 29460 1216 29512 1222
rect 29460 1158 29512 1164
rect 29472 746 29500 1158
rect 29460 740 29512 746
rect 29460 682 29512 688
rect 29552 740 29604 746
rect 29552 682 29604 688
rect 29564 542 29592 682
rect 29552 536 29604 542
rect 29552 478 29604 484
rect 29656 160 29684 1702
rect 29932 1358 29960 3130
rect 30010 2544 30066 2553
rect 30010 2479 30066 2488
rect 30024 2446 30052 2479
rect 30116 2446 30144 8434
rect 30380 3460 30432 3466
rect 30380 3402 30432 3408
rect 30012 2440 30064 2446
rect 30012 2382 30064 2388
rect 30104 2440 30156 2446
rect 30104 2382 30156 2388
rect 30196 2304 30248 2310
rect 30196 2246 30248 2252
rect 30208 2106 30236 2246
rect 30196 2100 30248 2106
rect 30196 2042 30248 2048
rect 30392 2038 30420 3402
rect 31036 2650 31064 8434
rect 33032 7644 33340 7653
rect 33032 7642 33038 7644
rect 33094 7642 33118 7644
rect 33174 7642 33198 7644
rect 33254 7642 33278 7644
rect 33334 7642 33340 7644
rect 33094 7590 33096 7642
rect 33276 7590 33278 7642
rect 33032 7588 33038 7590
rect 33094 7588 33118 7590
rect 33174 7588 33198 7590
rect 33254 7588 33278 7590
rect 33334 7588 33340 7590
rect 33032 7579 33340 7588
rect 33032 6556 33340 6565
rect 33032 6554 33038 6556
rect 33094 6554 33118 6556
rect 33174 6554 33198 6556
rect 33254 6554 33278 6556
rect 33334 6554 33340 6556
rect 33094 6502 33096 6554
rect 33276 6502 33278 6554
rect 33032 6500 33038 6502
rect 33094 6500 33118 6502
rect 33174 6500 33198 6502
rect 33254 6500 33278 6502
rect 33334 6500 33340 6502
rect 33032 6491 33340 6500
rect 33032 5468 33340 5477
rect 33032 5466 33038 5468
rect 33094 5466 33118 5468
rect 33174 5466 33198 5468
rect 33254 5466 33278 5468
rect 33334 5466 33340 5468
rect 33094 5414 33096 5466
rect 33276 5414 33278 5466
rect 33032 5412 33038 5414
rect 33094 5412 33118 5414
rect 33174 5412 33198 5414
rect 33254 5412 33278 5414
rect 33334 5412 33340 5414
rect 33032 5403 33340 5412
rect 33032 4380 33340 4389
rect 33032 4378 33038 4380
rect 33094 4378 33118 4380
rect 33174 4378 33198 4380
rect 33254 4378 33278 4380
rect 33334 4378 33340 4380
rect 33094 4326 33096 4378
rect 33276 4326 33278 4378
rect 33032 4324 33038 4326
rect 33094 4324 33118 4326
rect 33174 4324 33198 4326
rect 33254 4324 33278 4326
rect 33334 4324 33340 4326
rect 33032 4315 33340 4324
rect 32862 3496 32918 3505
rect 32862 3431 32918 3440
rect 31114 3360 31170 3369
rect 31114 3295 31170 3304
rect 31128 2854 31156 3295
rect 31760 2916 31812 2922
rect 31760 2858 31812 2864
rect 31116 2848 31168 2854
rect 31116 2790 31168 2796
rect 30932 2644 30984 2650
rect 30932 2586 30984 2592
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 30944 2281 30972 2586
rect 30930 2272 30986 2281
rect 30930 2207 30986 2216
rect 30380 2032 30432 2038
rect 30380 1974 30432 1980
rect 30748 1964 30800 1970
rect 30748 1906 30800 1912
rect 30852 1958 31248 1986
rect 30760 1465 30788 1906
rect 30746 1456 30802 1465
rect 30116 1426 30696 1442
rect 30116 1420 30708 1426
rect 30116 1414 30656 1420
rect 29920 1352 29972 1358
rect 29920 1294 29972 1300
rect 29736 1216 29788 1222
rect 29736 1158 29788 1164
rect 29748 1018 29776 1158
rect 29736 1012 29788 1018
rect 29736 954 29788 960
rect 29736 536 29788 542
rect 29736 478 29788 484
rect 29090 54 29316 82
rect 28814 0 28870 54
rect 29090 0 29146 54
rect 29366 0 29422 160
rect 29642 0 29698 160
rect 29748 134 29776 478
rect 29736 128 29788 134
rect 29736 70 29788 76
rect 29918 82 29974 160
rect 30116 82 30144 1414
rect 30746 1391 30802 1400
rect 30656 1362 30708 1368
rect 30288 1352 30340 1358
rect 30288 1294 30340 1300
rect 29918 54 30144 82
rect 30194 82 30250 160
rect 30300 82 30328 1294
rect 30852 218 30880 1958
rect 31220 1902 31248 1958
rect 31208 1896 31260 1902
rect 31208 1838 31260 1844
rect 31024 1760 31076 1766
rect 31300 1760 31352 1766
rect 31024 1702 31076 1708
rect 31220 1720 31300 1748
rect 31036 388 31064 1702
rect 30668 190 30880 218
rect 30944 360 31064 388
rect 30194 54 30328 82
rect 30470 82 30526 160
rect 30668 82 30696 190
rect 30470 54 30696 82
rect 30746 82 30802 160
rect 30944 82 30972 360
rect 30746 54 30972 82
rect 31022 82 31078 160
rect 31220 82 31248 1720
rect 31300 1702 31352 1708
rect 31668 1556 31720 1562
rect 31588 1516 31668 1544
rect 31484 1488 31536 1494
rect 31484 1430 31536 1436
rect 31022 54 31248 82
rect 31298 82 31354 160
rect 31496 82 31524 1430
rect 31588 160 31616 1516
rect 31668 1498 31720 1504
rect 31298 54 31524 82
rect 29918 0 29974 54
rect 30194 0 30250 54
rect 30470 0 30526 54
rect 30746 0 30802 54
rect 31022 0 31078 54
rect 31298 0 31354 54
rect 31574 0 31630 160
rect 31772 134 31800 2858
rect 32876 2446 32904 3431
rect 33032 3292 33340 3301
rect 33032 3290 33038 3292
rect 33094 3290 33118 3292
rect 33174 3290 33198 3292
rect 33254 3290 33278 3292
rect 33334 3290 33340 3292
rect 33094 3238 33096 3290
rect 33276 3238 33278 3290
rect 33032 3236 33038 3238
rect 33094 3236 33118 3238
rect 33174 3236 33198 3238
rect 33254 3236 33278 3238
rect 33334 3236 33340 3238
rect 33032 3227 33340 3236
rect 33414 3088 33470 3097
rect 33414 3023 33470 3032
rect 32956 2848 33008 2854
rect 32956 2790 33008 2796
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 32588 2304 32640 2310
rect 31850 2272 31906 2281
rect 32588 2246 32640 2252
rect 31850 2207 31906 2216
rect 31864 2106 31892 2207
rect 31852 2100 31904 2106
rect 31852 2042 31904 2048
rect 31944 1828 31996 1834
rect 31944 1770 31996 1776
rect 31852 1556 31904 1562
rect 31852 1498 31904 1504
rect 31864 1222 31892 1498
rect 31956 1494 31984 1770
rect 32404 1760 32456 1766
rect 32048 1720 32404 1748
rect 31944 1488 31996 1494
rect 31944 1430 31996 1436
rect 31944 1352 31996 1358
rect 31944 1294 31996 1300
rect 31852 1216 31904 1222
rect 31852 1158 31904 1164
rect 31956 785 31984 1294
rect 31942 776 31998 785
rect 31942 711 31998 720
rect 31760 128 31812 134
rect 31760 70 31812 76
rect 31850 82 31906 160
rect 32048 82 32076 1720
rect 32404 1702 32456 1708
rect 32600 1578 32628 2246
rect 32968 1952 32996 2790
rect 33032 2204 33340 2213
rect 33032 2202 33038 2204
rect 33094 2202 33118 2204
rect 33174 2202 33198 2204
rect 33254 2202 33278 2204
rect 33334 2202 33340 2204
rect 33094 2150 33096 2202
rect 33276 2150 33278 2202
rect 33032 2148 33038 2150
rect 33094 2148 33118 2150
rect 33174 2148 33198 2150
rect 33254 2148 33278 2150
rect 33334 2148 33340 2150
rect 33032 2139 33340 2148
rect 33324 2032 33376 2038
rect 33428 1986 33456 3023
rect 33520 2650 33548 8434
rect 36360 8356 36412 8362
rect 36360 8298 36412 8304
rect 33784 4276 33836 4282
rect 33784 4218 33836 4224
rect 33796 2650 33824 4218
rect 34888 4208 34940 4214
rect 34888 4150 34940 4156
rect 33874 4040 33930 4049
rect 33930 3998 34008 4026
rect 33874 3975 33930 3984
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 33784 2644 33836 2650
rect 33784 2586 33836 2592
rect 33692 2440 33744 2446
rect 33692 2382 33744 2388
rect 33704 2106 33732 2382
rect 33692 2100 33744 2106
rect 33692 2042 33744 2048
rect 33980 1986 34008 3998
rect 34152 2644 34204 2650
rect 34152 2586 34204 2592
rect 34164 2038 34192 2586
rect 34244 2508 34296 2514
rect 34244 2450 34296 2456
rect 33376 1980 33456 1986
rect 33324 1974 33456 1980
rect 33336 1958 33456 1974
rect 33888 1958 34008 1986
rect 34152 2032 34204 2038
rect 34152 1974 34204 1980
rect 32968 1924 33180 1952
rect 33048 1828 33100 1834
rect 33048 1770 33100 1776
rect 32956 1760 33008 1766
rect 32956 1702 33008 1708
rect 32324 1550 32628 1578
rect 32220 1284 32272 1290
rect 32220 1226 32272 1232
rect 32232 814 32260 1226
rect 32220 808 32272 814
rect 32220 750 32272 756
rect 31850 54 32076 82
rect 32126 82 32182 160
rect 32324 82 32352 1550
rect 32864 1420 32916 1426
rect 32864 1362 32916 1368
rect 32496 1352 32548 1358
rect 32496 1294 32548 1300
rect 32126 54 32352 82
rect 32402 82 32458 160
rect 32508 82 32536 1294
rect 32772 1284 32824 1290
rect 32772 1226 32824 1232
rect 32784 678 32812 1226
rect 32772 672 32824 678
rect 32772 614 32824 620
rect 32402 54 32536 82
rect 32678 82 32734 160
rect 32876 82 32904 1362
rect 32968 160 32996 1702
rect 33060 1562 33088 1770
rect 33048 1556 33100 1562
rect 33048 1498 33100 1504
rect 33152 1358 33180 1924
rect 33324 1828 33376 1834
rect 33324 1770 33376 1776
rect 33140 1352 33192 1358
rect 33140 1294 33192 1300
rect 33336 1306 33364 1770
rect 33508 1760 33560 1766
rect 33508 1702 33560 1708
rect 33336 1278 33456 1306
rect 33032 1116 33340 1125
rect 33032 1114 33038 1116
rect 33094 1114 33118 1116
rect 33174 1114 33198 1116
rect 33254 1114 33278 1116
rect 33334 1114 33340 1116
rect 33094 1062 33096 1114
rect 33276 1062 33278 1114
rect 33032 1060 33038 1062
rect 33094 1060 33118 1062
rect 33174 1060 33198 1062
rect 33254 1060 33278 1062
rect 33334 1060 33340 1062
rect 33032 1051 33340 1060
rect 32678 54 32904 82
rect 31850 0 31906 54
rect 32126 0 32182 54
rect 32402 0 32458 54
rect 32678 0 32734 54
rect 32954 0 33010 160
rect 33230 82 33286 160
rect 33428 82 33456 1278
rect 33520 160 33548 1702
rect 33888 1358 33916 1958
rect 34060 1488 34112 1494
rect 33980 1448 34060 1476
rect 33876 1352 33928 1358
rect 33876 1294 33928 1300
rect 33230 54 33456 82
rect 33230 0 33286 54
rect 33506 0 33562 160
rect 33782 82 33838 160
rect 33980 82 34008 1448
rect 34060 1430 34112 1436
rect 34060 1352 34112 1358
rect 34060 1294 34112 1300
rect 34072 160 34100 1294
rect 33782 54 34008 82
rect 33782 0 33838 54
rect 34058 0 34114 160
rect 34256 66 34284 2450
rect 34900 1970 34928 4150
rect 36372 2650 36400 8298
rect 37280 3120 37332 3126
rect 37280 3062 37332 3068
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 36544 2440 36596 2446
rect 36544 2382 36596 2388
rect 35624 2372 35676 2378
rect 35624 2314 35676 2320
rect 34888 1964 34940 1970
rect 34888 1906 34940 1912
rect 34520 1760 34572 1766
rect 34520 1702 34572 1708
rect 34428 1420 34480 1426
rect 34428 1362 34480 1368
rect 34440 762 34468 1362
rect 34532 1358 34560 1702
rect 34520 1352 34572 1358
rect 35072 1352 35124 1358
rect 35070 1320 35072 1329
rect 35124 1320 35126 1329
rect 34520 1294 34572 1300
rect 34808 1290 35020 1306
rect 34612 1284 34664 1290
rect 34612 1226 34664 1232
rect 34808 1284 35032 1290
rect 34808 1278 34980 1284
rect 34520 1216 34572 1222
rect 34520 1158 34572 1164
rect 34348 734 34468 762
rect 34348 160 34376 734
rect 34532 338 34560 1158
rect 34624 513 34652 1226
rect 34704 944 34756 950
rect 34704 886 34756 892
rect 34716 542 34744 886
rect 34704 536 34756 542
rect 34610 504 34666 513
rect 34704 478 34756 484
rect 34610 439 34666 448
rect 34520 332 34572 338
rect 34520 274 34572 280
rect 34244 60 34296 66
rect 34244 2 34296 8
rect 34334 0 34390 160
rect 34610 82 34666 160
rect 34808 82 34836 1278
rect 35070 1255 35126 1264
rect 34980 1226 35032 1232
rect 35440 808 35492 814
rect 35360 756 35440 762
rect 35360 750 35492 756
rect 35164 740 35216 746
rect 35164 682 35216 688
rect 35360 734 35480 750
rect 35176 626 35204 682
rect 34900 598 35204 626
rect 34900 160 34928 598
rect 34610 54 34836 82
rect 34610 0 34666 54
rect 34886 0 34942 160
rect 35162 82 35218 160
rect 35360 82 35388 734
rect 35440 672 35492 678
rect 35440 614 35492 620
rect 35452 160 35480 614
rect 35636 338 35664 2314
rect 36556 2106 36584 2382
rect 36544 2100 36596 2106
rect 36544 2042 36596 2048
rect 36542 2000 36598 2009
rect 36360 1964 36412 1970
rect 36542 1935 36598 1944
rect 36360 1906 36412 1912
rect 35992 1556 36044 1562
rect 35992 1498 36044 1504
rect 35624 332 35676 338
rect 35624 274 35676 280
rect 35808 196 35860 202
rect 35162 54 35388 82
rect 35162 0 35218 54
rect 35438 0 35494 160
rect 35714 82 35770 160
rect 36004 160 36032 1498
rect 36176 1216 36228 1222
rect 36176 1158 36228 1164
rect 36188 1018 36216 1158
rect 36176 1012 36228 1018
rect 36176 954 36228 960
rect 35808 138 35860 144
rect 35820 82 35848 138
rect 35714 54 35848 82
rect 35714 0 35770 54
rect 35990 0 36046 160
rect 36266 82 36322 160
rect 36372 82 36400 1906
rect 36556 1834 36584 1935
rect 36544 1828 36596 1834
rect 36544 1770 36596 1776
rect 37292 1358 37320 3062
rect 37384 2650 37412 8434
rect 38379 8188 38687 8197
rect 38379 8186 38385 8188
rect 38441 8186 38465 8188
rect 38521 8186 38545 8188
rect 38601 8186 38625 8188
rect 38681 8186 38687 8188
rect 38441 8134 38443 8186
rect 38623 8134 38625 8186
rect 38379 8132 38385 8134
rect 38441 8132 38465 8134
rect 38521 8132 38545 8134
rect 38601 8132 38625 8134
rect 38681 8132 38687 8134
rect 38379 8123 38687 8132
rect 38379 7100 38687 7109
rect 38379 7098 38385 7100
rect 38441 7098 38465 7100
rect 38521 7098 38545 7100
rect 38601 7098 38625 7100
rect 38681 7098 38687 7100
rect 38441 7046 38443 7098
rect 38623 7046 38625 7098
rect 38379 7044 38385 7046
rect 38441 7044 38465 7046
rect 38521 7044 38545 7046
rect 38601 7044 38625 7046
rect 38681 7044 38687 7046
rect 38379 7035 38687 7044
rect 38379 6012 38687 6021
rect 38379 6010 38385 6012
rect 38441 6010 38465 6012
rect 38521 6010 38545 6012
rect 38601 6010 38625 6012
rect 38681 6010 38687 6012
rect 38441 5958 38443 6010
rect 38623 5958 38625 6010
rect 38379 5956 38385 5958
rect 38441 5956 38465 5958
rect 38521 5956 38545 5958
rect 38601 5956 38625 5958
rect 38681 5956 38687 5958
rect 38379 5947 38687 5956
rect 38379 4924 38687 4933
rect 38379 4922 38385 4924
rect 38441 4922 38465 4924
rect 38521 4922 38545 4924
rect 38601 4922 38625 4924
rect 38681 4922 38687 4924
rect 38441 4870 38443 4922
rect 38623 4870 38625 4922
rect 38379 4868 38385 4870
rect 38441 4868 38465 4870
rect 38521 4868 38545 4870
rect 38601 4868 38625 4870
rect 38681 4868 38687 4870
rect 38379 4859 38687 4868
rect 38379 3836 38687 3845
rect 38379 3834 38385 3836
rect 38441 3834 38465 3836
rect 38521 3834 38545 3836
rect 38601 3834 38625 3836
rect 38681 3834 38687 3836
rect 38441 3782 38443 3834
rect 38623 3782 38625 3834
rect 38379 3780 38385 3782
rect 38441 3780 38465 3782
rect 38521 3780 38545 3782
rect 38601 3780 38625 3782
rect 38681 3780 38687 3782
rect 38379 3771 38687 3780
rect 39212 3052 39264 3058
rect 39212 2994 39264 3000
rect 38379 2748 38687 2757
rect 38379 2746 38385 2748
rect 38441 2746 38465 2748
rect 38521 2746 38545 2748
rect 38601 2746 38625 2748
rect 38681 2746 38687 2748
rect 38441 2694 38443 2746
rect 38623 2694 38625 2746
rect 38379 2692 38385 2694
rect 38441 2692 38465 2694
rect 38521 2692 38545 2694
rect 38601 2692 38625 2694
rect 38681 2692 38687 2694
rect 38379 2683 38687 2692
rect 37372 2644 37424 2650
rect 37372 2586 37424 2592
rect 37648 2576 37700 2582
rect 37648 2518 37700 2524
rect 37660 1358 37688 2518
rect 37924 2440 37976 2446
rect 37924 2382 37976 2388
rect 37936 2106 37964 2382
rect 37924 2100 37976 2106
rect 37924 2042 37976 2048
rect 38379 1660 38687 1669
rect 38379 1658 38385 1660
rect 38441 1658 38465 1660
rect 38521 1658 38545 1660
rect 38601 1658 38625 1660
rect 38681 1658 38687 1660
rect 38441 1606 38443 1658
rect 38623 1606 38625 1658
rect 38379 1604 38385 1606
rect 38441 1604 38465 1606
rect 38521 1604 38545 1606
rect 38601 1604 38625 1606
rect 38681 1604 38687 1606
rect 38379 1595 38687 1604
rect 39224 1562 39252 2994
rect 39960 2650 39988 8434
rect 40696 2650 40724 8434
rect 43272 2650 43300 8434
rect 43726 7644 44034 7653
rect 43726 7642 43732 7644
rect 43788 7642 43812 7644
rect 43868 7642 43892 7644
rect 43948 7642 43972 7644
rect 44028 7642 44034 7644
rect 43788 7590 43790 7642
rect 43970 7590 43972 7642
rect 43726 7588 43732 7590
rect 43788 7588 43812 7590
rect 43868 7588 43892 7590
rect 43948 7588 43972 7590
rect 44028 7588 44034 7590
rect 43726 7579 44034 7588
rect 43726 6556 44034 6565
rect 43726 6554 43732 6556
rect 43788 6554 43812 6556
rect 43868 6554 43892 6556
rect 43948 6554 43972 6556
rect 44028 6554 44034 6556
rect 43788 6502 43790 6554
rect 43970 6502 43972 6554
rect 43726 6500 43732 6502
rect 43788 6500 43812 6502
rect 43868 6500 43892 6502
rect 43948 6500 43972 6502
rect 44028 6500 44034 6502
rect 43726 6491 44034 6500
rect 43726 5468 44034 5477
rect 43726 5466 43732 5468
rect 43788 5466 43812 5468
rect 43868 5466 43892 5468
rect 43948 5466 43972 5468
rect 44028 5466 44034 5468
rect 43788 5414 43790 5466
rect 43970 5414 43972 5466
rect 43726 5412 43732 5414
rect 43788 5412 43812 5414
rect 43868 5412 43892 5414
rect 43948 5412 43972 5414
rect 44028 5412 44034 5414
rect 43726 5403 44034 5412
rect 43726 4380 44034 4389
rect 43726 4378 43732 4380
rect 43788 4378 43812 4380
rect 43868 4378 43892 4380
rect 43948 4378 43972 4380
rect 44028 4378 44034 4380
rect 43788 4326 43790 4378
rect 43970 4326 43972 4378
rect 43726 4324 43732 4326
rect 43788 4324 43812 4326
rect 43868 4324 43892 4326
rect 43948 4324 43972 4326
rect 44028 4324 44034 4326
rect 43726 4315 44034 4324
rect 43726 3292 44034 3301
rect 43726 3290 43732 3292
rect 43788 3290 43812 3292
rect 43868 3290 43892 3292
rect 43948 3290 43972 3292
rect 44028 3290 44034 3292
rect 43788 3238 43790 3290
rect 43970 3238 43972 3290
rect 43726 3236 43732 3238
rect 43788 3236 43812 3238
rect 43868 3236 43892 3238
rect 43948 3236 43972 3238
rect 44028 3236 44034 3238
rect 43726 3227 44034 3236
rect 39948 2644 40000 2650
rect 39948 2586 40000 2592
rect 40684 2644 40736 2650
rect 40684 2586 40736 2592
rect 43260 2644 43312 2650
rect 43260 2586 43312 2592
rect 39672 2440 39724 2446
rect 39672 2382 39724 2388
rect 40868 2440 40920 2446
rect 40868 2382 40920 2388
rect 42432 2440 42484 2446
rect 42432 2382 42484 2388
rect 39684 2106 39712 2382
rect 40880 2106 40908 2382
rect 42444 2106 42472 2382
rect 43726 2204 44034 2213
rect 43726 2202 43732 2204
rect 43788 2202 43812 2204
rect 43868 2202 43892 2204
rect 43948 2202 43972 2204
rect 44028 2202 44034 2204
rect 43788 2150 43790 2202
rect 43970 2150 43972 2202
rect 43726 2148 43732 2150
rect 43788 2148 43812 2150
rect 43868 2148 43892 2150
rect 43948 2148 43972 2150
rect 44028 2148 44034 2150
rect 43726 2139 44034 2148
rect 39672 2100 39724 2106
rect 39672 2042 39724 2048
rect 40868 2100 40920 2106
rect 40868 2042 40920 2048
rect 42432 2100 42484 2106
rect 42432 2042 42484 2048
rect 40040 1964 40092 1970
rect 40040 1906 40092 1912
rect 40132 1964 40184 1970
rect 40132 1906 40184 1912
rect 41512 1964 41564 1970
rect 41512 1906 41564 1912
rect 39764 1828 39816 1834
rect 39764 1770 39816 1776
rect 38108 1556 38160 1562
rect 38108 1498 38160 1504
rect 39212 1556 39264 1562
rect 39212 1498 39264 1504
rect 38120 1358 38148 1498
rect 39304 1420 39356 1426
rect 39304 1362 39356 1368
rect 36728 1352 36780 1358
rect 36728 1294 36780 1300
rect 37280 1352 37332 1358
rect 37280 1294 37332 1300
rect 37464 1352 37516 1358
rect 37464 1294 37516 1300
rect 37556 1352 37608 1358
rect 37556 1294 37608 1300
rect 37648 1352 37700 1358
rect 37648 1294 37700 1300
rect 37832 1352 37884 1358
rect 37832 1294 37884 1300
rect 38108 1352 38160 1358
rect 38108 1294 38160 1300
rect 38660 1352 38712 1358
rect 38660 1294 38712 1300
rect 38936 1352 38988 1358
rect 38936 1294 38988 1300
rect 36544 1284 36596 1290
rect 36544 1226 36596 1232
rect 36556 160 36584 1226
rect 36636 1216 36688 1222
rect 36636 1158 36688 1164
rect 36648 882 36676 1158
rect 36636 876 36688 882
rect 36636 818 36688 824
rect 36740 746 36768 1294
rect 36912 1216 36964 1222
rect 36912 1158 36964 1164
rect 37372 1216 37424 1222
rect 37372 1158 37424 1164
rect 36728 740 36780 746
rect 36728 682 36780 688
rect 36820 264 36872 270
rect 36820 206 36872 212
rect 36832 160 36860 206
rect 36266 54 36400 82
rect 36266 0 36322 54
rect 36542 0 36598 160
rect 36818 0 36874 160
rect 36924 134 36952 1158
rect 37188 1012 37240 1018
rect 37188 954 37240 960
rect 36912 128 36964 134
rect 36912 70 36964 76
rect 37094 82 37150 160
rect 37200 82 37228 954
rect 37384 406 37412 1158
rect 37476 814 37504 1294
rect 37464 808 37516 814
rect 37464 750 37516 756
rect 37568 678 37596 1294
rect 37844 898 37872 1294
rect 38476 1284 38528 1290
rect 38476 1226 38528 1232
rect 38292 1216 38344 1222
rect 38292 1158 38344 1164
rect 37660 870 37872 898
rect 37556 672 37608 678
rect 37556 614 37608 620
rect 37660 490 37688 870
rect 37740 808 37792 814
rect 37740 750 37792 756
rect 37476 462 37688 490
rect 37372 400 37424 406
rect 37372 342 37424 348
rect 37476 202 37504 462
rect 37752 218 37780 750
rect 38304 746 38332 1158
rect 38292 740 38344 746
rect 38292 682 38344 688
rect 38488 490 38516 1226
rect 38568 1216 38620 1222
rect 38568 1158 38620 1164
rect 38580 785 38608 1158
rect 38566 776 38622 785
rect 38566 711 38622 720
rect 38568 672 38620 678
rect 38568 614 38620 620
rect 37464 196 37516 202
rect 37094 54 37228 82
rect 37370 82 37426 160
rect 37464 138 37516 144
rect 37568 190 37780 218
rect 37844 462 38516 490
rect 37568 82 37596 190
rect 37370 54 37596 82
rect 37646 82 37702 160
rect 37844 82 37872 462
rect 38476 400 38528 406
rect 38396 348 38476 354
rect 38396 342 38528 348
rect 37924 332 37976 338
rect 37924 274 37976 280
rect 38396 326 38516 342
rect 37936 160 37964 274
rect 37646 54 37872 82
rect 37094 0 37150 54
rect 37370 0 37426 54
rect 37646 0 37702 54
rect 37922 0 37978 160
rect 38198 82 38254 160
rect 38396 82 38424 326
rect 38198 54 38424 82
rect 38474 82 38530 160
rect 38580 82 38608 614
rect 38672 270 38700 1294
rect 38844 1216 38896 1222
rect 38844 1158 38896 1164
rect 38856 882 38884 1158
rect 38948 1018 38976 1294
rect 39120 1216 39172 1222
rect 39120 1158 39172 1164
rect 39212 1216 39264 1222
rect 39212 1158 39264 1164
rect 39132 1018 39160 1158
rect 38936 1012 38988 1018
rect 38936 954 38988 960
rect 39120 1012 39172 1018
rect 39120 954 39172 960
rect 38948 882 39160 898
rect 38844 876 38896 882
rect 38844 818 38896 824
rect 38948 876 39172 882
rect 38948 870 39120 876
rect 38660 264 38712 270
rect 38660 206 38712 212
rect 38474 54 38608 82
rect 38750 82 38806 160
rect 38948 82 38976 870
rect 39120 818 39172 824
rect 39120 740 39172 746
rect 39120 682 39172 688
rect 39132 626 39160 682
rect 39040 598 39160 626
rect 39040 160 39068 598
rect 38750 54 38976 82
rect 38198 0 38254 54
rect 38474 0 38530 54
rect 38750 0 38806 54
rect 39026 0 39082 160
rect 39224 66 39252 1158
rect 39316 160 39344 1362
rect 39396 1352 39448 1358
rect 39396 1294 39448 1300
rect 39408 814 39436 1294
rect 39776 1222 39804 1770
rect 39948 1760 40000 1766
rect 39948 1702 40000 1708
rect 39856 1488 39908 1494
rect 39856 1430 39908 1436
rect 39960 1442 39988 1702
rect 40052 1562 40080 1906
rect 40144 1562 40172 1906
rect 40684 1896 40736 1902
rect 40684 1838 40736 1844
rect 40040 1556 40092 1562
rect 40040 1498 40092 1504
rect 40132 1556 40184 1562
rect 40132 1498 40184 1504
rect 39764 1216 39816 1222
rect 39764 1158 39816 1164
rect 39396 808 39448 814
rect 39396 750 39448 756
rect 39868 474 39896 1430
rect 39960 1414 40264 1442
rect 40040 1352 40092 1358
rect 40040 1294 40092 1300
rect 39948 1284 40000 1290
rect 39948 1226 40000 1232
rect 39856 468 39908 474
rect 39856 410 39908 416
rect 39212 60 39264 66
rect 39212 2 39264 8
rect 39302 0 39358 160
rect 39578 82 39634 160
rect 39960 82 39988 1226
rect 40052 338 40080 1294
rect 40236 1222 40264 1414
rect 40316 1352 40368 1358
rect 40316 1294 40368 1300
rect 40592 1352 40644 1358
rect 40592 1294 40644 1300
rect 40224 1216 40276 1222
rect 40224 1158 40276 1164
rect 40328 406 40356 1294
rect 40604 678 40632 1294
rect 40696 1222 40724 1838
rect 41524 1562 41552 1906
rect 41512 1556 41564 1562
rect 41512 1498 41564 1504
rect 40868 1352 40920 1358
rect 40868 1294 40920 1300
rect 41144 1352 41196 1358
rect 41144 1294 41196 1300
rect 40684 1216 40736 1222
rect 40684 1158 40736 1164
rect 40880 882 40908 1294
rect 40868 876 40920 882
rect 40868 818 40920 824
rect 41156 746 41184 1294
rect 43726 1116 44034 1125
rect 43726 1114 43732 1116
rect 43788 1114 43812 1116
rect 43868 1114 43892 1116
rect 43948 1114 43972 1116
rect 44028 1114 44034 1116
rect 43788 1062 43790 1114
rect 43970 1062 43972 1114
rect 43726 1060 43732 1062
rect 43788 1060 43812 1062
rect 43868 1060 43892 1062
rect 43948 1060 43972 1062
rect 44028 1060 44034 1062
rect 43726 1051 44034 1060
rect 41144 740 41196 746
rect 41144 682 41196 688
rect 40592 672 40644 678
rect 40592 614 40644 620
rect 40316 400 40368 406
rect 40316 342 40368 348
rect 40040 332 40092 338
rect 40040 274 40092 280
rect 39578 54 39988 82
rect 39578 0 39634 54
<< via2 >>
rect 11650 8730 11706 8732
rect 11730 8730 11786 8732
rect 11810 8730 11866 8732
rect 11890 8730 11946 8732
rect 11650 8678 11696 8730
rect 11696 8678 11706 8730
rect 11730 8678 11760 8730
rect 11760 8678 11772 8730
rect 11772 8678 11786 8730
rect 11810 8678 11824 8730
rect 11824 8678 11836 8730
rect 11836 8678 11866 8730
rect 11890 8678 11900 8730
rect 11900 8678 11946 8730
rect 11650 8676 11706 8678
rect 11730 8676 11786 8678
rect 11810 8676 11866 8678
rect 11890 8676 11946 8678
rect 5538 8492 5594 8528
rect 22344 8730 22400 8732
rect 22424 8730 22480 8732
rect 22504 8730 22560 8732
rect 22584 8730 22640 8732
rect 22344 8678 22390 8730
rect 22390 8678 22400 8730
rect 22424 8678 22454 8730
rect 22454 8678 22466 8730
rect 22466 8678 22480 8730
rect 22504 8678 22518 8730
rect 22518 8678 22530 8730
rect 22530 8678 22560 8730
rect 22584 8678 22594 8730
rect 22594 8678 22640 8730
rect 22344 8676 22400 8678
rect 22424 8676 22480 8678
rect 22504 8676 22560 8678
rect 22584 8676 22640 8678
rect 5538 8472 5540 8492
rect 5540 8472 5592 8492
rect 5592 8472 5594 8492
rect 4434 8356 4490 8392
rect 4434 8336 4436 8356
rect 4436 8336 4488 8356
rect 4488 8336 4490 8356
rect 6303 8186 6359 8188
rect 6383 8186 6439 8188
rect 6463 8186 6519 8188
rect 6543 8186 6599 8188
rect 6303 8134 6349 8186
rect 6349 8134 6359 8186
rect 6383 8134 6413 8186
rect 6413 8134 6425 8186
rect 6425 8134 6439 8186
rect 6463 8134 6477 8186
rect 6477 8134 6489 8186
rect 6489 8134 6519 8186
rect 6543 8134 6553 8186
rect 6553 8134 6599 8186
rect 6303 8132 6359 8134
rect 6383 8132 6439 8134
rect 6463 8132 6519 8134
rect 6543 8132 6599 8134
rect 11650 7642 11706 7644
rect 11730 7642 11786 7644
rect 11810 7642 11866 7644
rect 11890 7642 11946 7644
rect 11650 7590 11696 7642
rect 11696 7590 11706 7642
rect 11730 7590 11760 7642
rect 11760 7590 11772 7642
rect 11772 7590 11786 7642
rect 11810 7590 11824 7642
rect 11824 7590 11836 7642
rect 11836 7590 11866 7642
rect 11890 7590 11900 7642
rect 11900 7590 11946 7642
rect 11650 7588 11706 7590
rect 11730 7588 11786 7590
rect 11810 7588 11866 7590
rect 11890 7588 11946 7590
rect 6303 7098 6359 7100
rect 6383 7098 6439 7100
rect 6463 7098 6519 7100
rect 6543 7098 6599 7100
rect 6303 7046 6349 7098
rect 6349 7046 6359 7098
rect 6383 7046 6413 7098
rect 6413 7046 6425 7098
rect 6425 7046 6439 7098
rect 6463 7046 6477 7098
rect 6477 7046 6489 7098
rect 6489 7046 6519 7098
rect 6543 7046 6553 7098
rect 6553 7046 6599 7098
rect 6303 7044 6359 7046
rect 6383 7044 6439 7046
rect 6463 7044 6519 7046
rect 6543 7044 6599 7046
rect 11650 6554 11706 6556
rect 11730 6554 11786 6556
rect 11810 6554 11866 6556
rect 11890 6554 11946 6556
rect 11650 6502 11696 6554
rect 11696 6502 11706 6554
rect 11730 6502 11760 6554
rect 11760 6502 11772 6554
rect 11772 6502 11786 6554
rect 11810 6502 11824 6554
rect 11824 6502 11836 6554
rect 11836 6502 11866 6554
rect 11890 6502 11900 6554
rect 11900 6502 11946 6554
rect 11650 6500 11706 6502
rect 11730 6500 11786 6502
rect 11810 6500 11866 6502
rect 11890 6500 11946 6502
rect 6303 6010 6359 6012
rect 6383 6010 6439 6012
rect 6463 6010 6519 6012
rect 6543 6010 6599 6012
rect 6303 5958 6349 6010
rect 6349 5958 6359 6010
rect 6383 5958 6413 6010
rect 6413 5958 6425 6010
rect 6425 5958 6439 6010
rect 6463 5958 6477 6010
rect 6477 5958 6489 6010
rect 6489 5958 6519 6010
rect 6543 5958 6553 6010
rect 6553 5958 6599 6010
rect 6303 5956 6359 5958
rect 6383 5956 6439 5958
rect 6463 5956 6519 5958
rect 6543 5956 6599 5958
rect 11650 5466 11706 5468
rect 11730 5466 11786 5468
rect 11810 5466 11866 5468
rect 11890 5466 11946 5468
rect 11650 5414 11696 5466
rect 11696 5414 11706 5466
rect 11730 5414 11760 5466
rect 11760 5414 11772 5466
rect 11772 5414 11786 5466
rect 11810 5414 11824 5466
rect 11824 5414 11836 5466
rect 11836 5414 11866 5466
rect 11890 5414 11900 5466
rect 11900 5414 11946 5466
rect 11650 5412 11706 5414
rect 11730 5412 11786 5414
rect 11810 5412 11866 5414
rect 11890 5412 11946 5414
rect 6303 4922 6359 4924
rect 6383 4922 6439 4924
rect 6463 4922 6519 4924
rect 6543 4922 6599 4924
rect 6303 4870 6349 4922
rect 6349 4870 6359 4922
rect 6383 4870 6413 4922
rect 6413 4870 6425 4922
rect 6425 4870 6439 4922
rect 6463 4870 6477 4922
rect 6477 4870 6489 4922
rect 6489 4870 6519 4922
rect 6543 4870 6553 4922
rect 6553 4870 6599 4922
rect 6303 4868 6359 4870
rect 6383 4868 6439 4870
rect 6463 4868 6519 4870
rect 6543 4868 6599 4870
rect 6303 3834 6359 3836
rect 6383 3834 6439 3836
rect 6463 3834 6519 3836
rect 6543 3834 6599 3836
rect 6303 3782 6349 3834
rect 6349 3782 6359 3834
rect 6383 3782 6413 3834
rect 6413 3782 6425 3834
rect 6425 3782 6439 3834
rect 6463 3782 6477 3834
rect 6477 3782 6489 3834
rect 6489 3782 6519 3834
rect 6543 3782 6553 3834
rect 6553 3782 6599 3834
rect 6303 3780 6359 3782
rect 6383 3780 6439 3782
rect 6463 3780 6519 3782
rect 6543 3780 6599 3782
rect 6303 2746 6359 2748
rect 6383 2746 6439 2748
rect 6463 2746 6519 2748
rect 6543 2746 6599 2748
rect 6303 2694 6349 2746
rect 6349 2694 6359 2746
rect 6383 2694 6413 2746
rect 6413 2694 6425 2746
rect 6425 2694 6439 2746
rect 6463 2694 6477 2746
rect 6477 2694 6489 2746
rect 6489 2694 6519 2746
rect 6543 2694 6553 2746
rect 6553 2694 6599 2746
rect 6303 2692 6359 2694
rect 6383 2692 6439 2694
rect 6463 2692 6519 2694
rect 6543 2692 6599 2694
rect 6303 1658 6359 1660
rect 6383 1658 6439 1660
rect 6463 1658 6519 1660
rect 6543 1658 6599 1660
rect 6303 1606 6349 1658
rect 6349 1606 6359 1658
rect 6383 1606 6413 1658
rect 6413 1606 6425 1658
rect 6425 1606 6439 1658
rect 6463 1606 6477 1658
rect 6477 1606 6489 1658
rect 6489 1606 6519 1658
rect 6543 1606 6553 1658
rect 6553 1606 6599 1658
rect 6303 1604 6359 1606
rect 6383 1604 6439 1606
rect 6463 1604 6519 1606
rect 6543 1604 6599 1606
rect 6182 584 6238 640
rect 6550 312 6606 368
rect 8482 2488 8538 2544
rect 10782 1944 10838 2000
rect 8298 1436 8300 1456
rect 8300 1436 8352 1456
rect 8352 1436 8354 1456
rect 8298 1400 8354 1436
rect 10690 1808 10746 1864
rect 10966 720 11022 776
rect 11650 4378 11706 4380
rect 11730 4378 11786 4380
rect 11810 4378 11866 4380
rect 11890 4378 11946 4380
rect 11650 4326 11696 4378
rect 11696 4326 11706 4378
rect 11730 4326 11760 4378
rect 11760 4326 11772 4378
rect 11772 4326 11786 4378
rect 11810 4326 11824 4378
rect 11824 4326 11836 4378
rect 11836 4326 11866 4378
rect 11890 4326 11900 4378
rect 11900 4326 11946 4378
rect 11650 4324 11706 4326
rect 11730 4324 11786 4326
rect 11810 4324 11866 4326
rect 11890 4324 11946 4326
rect 11650 3290 11706 3292
rect 11730 3290 11786 3292
rect 11810 3290 11866 3292
rect 11890 3290 11946 3292
rect 11650 3238 11696 3290
rect 11696 3238 11706 3290
rect 11730 3238 11760 3290
rect 11760 3238 11772 3290
rect 11772 3238 11786 3290
rect 11810 3238 11824 3290
rect 11824 3238 11836 3290
rect 11836 3238 11866 3290
rect 11890 3238 11900 3290
rect 11900 3238 11946 3290
rect 11650 3236 11706 3238
rect 11730 3236 11786 3238
rect 11810 3236 11866 3238
rect 11890 3236 11946 3238
rect 11242 856 11298 912
rect 11650 2202 11706 2204
rect 11730 2202 11786 2204
rect 11810 2202 11866 2204
rect 11890 2202 11946 2204
rect 11650 2150 11696 2202
rect 11696 2150 11706 2202
rect 11730 2150 11760 2202
rect 11760 2150 11772 2202
rect 11772 2150 11786 2202
rect 11810 2150 11824 2202
rect 11824 2150 11836 2202
rect 11836 2150 11866 2202
rect 11890 2150 11900 2202
rect 11900 2150 11946 2202
rect 11650 2148 11706 2150
rect 11730 2148 11786 2150
rect 11810 2148 11866 2150
rect 11890 2148 11946 2150
rect 12530 3984 12586 4040
rect 12070 2352 12126 2408
rect 11650 1114 11706 1116
rect 11730 1114 11786 1116
rect 11810 1114 11866 1116
rect 11890 1114 11946 1116
rect 11650 1062 11696 1114
rect 11696 1062 11706 1114
rect 11730 1062 11760 1114
rect 11760 1062 11772 1114
rect 11772 1062 11786 1114
rect 11810 1062 11824 1114
rect 11824 1062 11836 1114
rect 11836 1062 11866 1114
rect 11890 1062 11900 1114
rect 11900 1062 11946 1114
rect 11650 1060 11706 1062
rect 11730 1060 11786 1062
rect 11810 1060 11866 1062
rect 11890 1060 11946 1062
rect 16997 8186 17053 8188
rect 17077 8186 17133 8188
rect 17157 8186 17213 8188
rect 17237 8186 17293 8188
rect 16997 8134 17043 8186
rect 17043 8134 17053 8186
rect 17077 8134 17107 8186
rect 17107 8134 17119 8186
rect 17119 8134 17133 8186
rect 17157 8134 17171 8186
rect 17171 8134 17183 8186
rect 17183 8134 17213 8186
rect 17237 8134 17247 8186
rect 17247 8134 17293 8186
rect 16997 8132 17053 8134
rect 17077 8132 17133 8134
rect 17157 8132 17213 8134
rect 17237 8132 17293 8134
rect 16997 7098 17053 7100
rect 17077 7098 17133 7100
rect 17157 7098 17213 7100
rect 17237 7098 17293 7100
rect 16997 7046 17043 7098
rect 17043 7046 17053 7098
rect 17077 7046 17107 7098
rect 17107 7046 17119 7098
rect 17119 7046 17133 7098
rect 17157 7046 17171 7098
rect 17171 7046 17183 7098
rect 17183 7046 17213 7098
rect 17237 7046 17247 7098
rect 17247 7046 17293 7098
rect 16997 7044 17053 7046
rect 17077 7044 17133 7046
rect 17157 7044 17213 7046
rect 17237 7044 17293 7046
rect 16997 6010 17053 6012
rect 17077 6010 17133 6012
rect 17157 6010 17213 6012
rect 17237 6010 17293 6012
rect 16997 5958 17043 6010
rect 17043 5958 17053 6010
rect 17077 5958 17107 6010
rect 17107 5958 17119 6010
rect 17119 5958 17133 6010
rect 17157 5958 17171 6010
rect 17171 5958 17183 6010
rect 17183 5958 17213 6010
rect 17237 5958 17247 6010
rect 17247 5958 17293 6010
rect 16997 5956 17053 5958
rect 17077 5956 17133 5958
rect 17157 5956 17213 5958
rect 17237 5956 17293 5958
rect 15382 3576 15438 3632
rect 14370 3168 14426 3224
rect 13910 2080 13966 2136
rect 13542 1944 13598 2000
rect 16210 2896 16266 2952
rect 16997 4922 17053 4924
rect 17077 4922 17133 4924
rect 17157 4922 17213 4924
rect 17237 4922 17293 4924
rect 16997 4870 17043 4922
rect 17043 4870 17053 4922
rect 17077 4870 17107 4922
rect 17107 4870 17119 4922
rect 17119 4870 17133 4922
rect 17157 4870 17171 4922
rect 17171 4870 17183 4922
rect 17183 4870 17213 4922
rect 17237 4870 17247 4922
rect 17247 4870 17293 4922
rect 16997 4868 17053 4870
rect 17077 4868 17133 4870
rect 17157 4868 17213 4870
rect 17237 4868 17293 4870
rect 18234 3984 18290 4040
rect 16997 3834 17053 3836
rect 17077 3834 17133 3836
rect 17157 3834 17213 3836
rect 17237 3834 17293 3836
rect 16997 3782 17043 3834
rect 17043 3782 17053 3834
rect 17077 3782 17107 3834
rect 17107 3782 17119 3834
rect 17119 3782 17133 3834
rect 17157 3782 17171 3834
rect 17171 3782 17183 3834
rect 17183 3782 17213 3834
rect 17237 3782 17247 3834
rect 17247 3782 17293 3834
rect 16997 3780 17053 3782
rect 17077 3780 17133 3782
rect 17157 3780 17213 3782
rect 17237 3780 17293 3782
rect 16854 3440 16910 3496
rect 15014 1264 15070 1320
rect 16997 2746 17053 2748
rect 17077 2746 17133 2748
rect 17157 2746 17213 2748
rect 17237 2746 17293 2748
rect 16997 2694 17043 2746
rect 17043 2694 17053 2746
rect 17077 2694 17107 2746
rect 17107 2694 17119 2746
rect 17119 2694 17133 2746
rect 17157 2694 17171 2746
rect 17171 2694 17183 2746
rect 17183 2694 17213 2746
rect 17237 2694 17247 2746
rect 17247 2694 17293 2746
rect 16997 2692 17053 2694
rect 17077 2692 17133 2694
rect 17157 2692 17213 2694
rect 17237 2692 17293 2694
rect 17406 2624 17462 2680
rect 17406 2216 17462 2272
rect 16997 1658 17053 1660
rect 17077 1658 17133 1660
rect 17157 1658 17213 1660
rect 17237 1658 17293 1660
rect 16997 1606 17043 1658
rect 17043 1606 17053 1658
rect 17077 1606 17107 1658
rect 17107 1606 17119 1658
rect 17119 1606 17133 1658
rect 17157 1606 17171 1658
rect 17171 1606 17183 1658
rect 17183 1606 17213 1658
rect 17237 1606 17247 1658
rect 17247 1606 17293 1658
rect 16997 1604 17053 1606
rect 17077 1604 17133 1606
rect 17157 1604 17213 1606
rect 17237 1604 17293 1606
rect 17406 1672 17462 1728
rect 17498 1536 17554 1592
rect 16854 1128 16910 1184
rect 16210 176 16266 232
rect 16854 584 16910 640
rect 18050 1808 18106 1864
rect 18510 3032 18566 3088
rect 18326 2080 18382 2136
rect 18970 2216 19026 2272
rect 17958 992 18014 1048
rect 19062 1536 19118 1592
rect 21546 3168 21602 3224
rect 21546 2896 21602 2952
rect 22344 7642 22400 7644
rect 22424 7642 22480 7644
rect 22504 7642 22560 7644
rect 22584 7642 22640 7644
rect 22344 7590 22390 7642
rect 22390 7590 22400 7642
rect 22424 7590 22454 7642
rect 22454 7590 22466 7642
rect 22466 7590 22480 7642
rect 22504 7590 22518 7642
rect 22518 7590 22530 7642
rect 22530 7590 22560 7642
rect 22584 7590 22594 7642
rect 22594 7590 22640 7642
rect 22344 7588 22400 7590
rect 22424 7588 22480 7590
rect 22504 7588 22560 7590
rect 22584 7588 22640 7590
rect 22344 6554 22400 6556
rect 22424 6554 22480 6556
rect 22504 6554 22560 6556
rect 22584 6554 22640 6556
rect 22344 6502 22390 6554
rect 22390 6502 22400 6554
rect 22424 6502 22454 6554
rect 22454 6502 22466 6554
rect 22466 6502 22480 6554
rect 22504 6502 22518 6554
rect 22518 6502 22530 6554
rect 22530 6502 22560 6554
rect 22584 6502 22594 6554
rect 22594 6502 22640 6554
rect 22344 6500 22400 6502
rect 22424 6500 22480 6502
rect 22504 6500 22560 6502
rect 22584 6500 22640 6502
rect 22344 5466 22400 5468
rect 22424 5466 22480 5468
rect 22504 5466 22560 5468
rect 22584 5466 22640 5468
rect 22344 5414 22390 5466
rect 22390 5414 22400 5466
rect 22424 5414 22454 5466
rect 22454 5414 22466 5466
rect 22466 5414 22480 5466
rect 22504 5414 22518 5466
rect 22518 5414 22530 5466
rect 22530 5414 22560 5466
rect 22584 5414 22594 5466
rect 22594 5414 22640 5466
rect 22344 5412 22400 5414
rect 22424 5412 22480 5414
rect 22504 5412 22560 5414
rect 22584 5412 22640 5414
rect 22344 4378 22400 4380
rect 22424 4378 22480 4380
rect 22504 4378 22560 4380
rect 22584 4378 22640 4380
rect 22344 4326 22390 4378
rect 22390 4326 22400 4378
rect 22424 4326 22454 4378
rect 22454 4326 22466 4378
rect 22466 4326 22480 4378
rect 22504 4326 22518 4378
rect 22518 4326 22530 4378
rect 22530 4326 22560 4378
rect 22584 4326 22594 4378
rect 22594 4326 22640 4378
rect 22344 4324 22400 4326
rect 22424 4324 22480 4326
rect 22504 4324 22560 4326
rect 22584 4324 22640 4326
rect 22344 3290 22400 3292
rect 22424 3290 22480 3292
rect 22504 3290 22560 3292
rect 22584 3290 22640 3292
rect 22344 3238 22390 3290
rect 22390 3238 22400 3290
rect 22424 3238 22454 3290
rect 22454 3238 22466 3290
rect 22466 3238 22480 3290
rect 22504 3238 22518 3290
rect 22518 3238 22530 3290
rect 22530 3238 22560 3290
rect 22584 3238 22594 3290
rect 22594 3238 22640 3290
rect 22344 3236 22400 3238
rect 22424 3236 22480 3238
rect 22504 3236 22560 3238
rect 22584 3236 22640 3238
rect 22374 2488 22430 2544
rect 20074 176 20130 232
rect 20810 1264 20866 1320
rect 20994 448 21050 504
rect 21730 1264 21786 1320
rect 21822 992 21878 1048
rect 21822 448 21878 504
rect 22344 2202 22400 2204
rect 22424 2202 22480 2204
rect 22504 2202 22560 2204
rect 22584 2202 22640 2204
rect 22344 2150 22390 2202
rect 22390 2150 22400 2202
rect 22424 2150 22454 2202
rect 22454 2150 22466 2202
rect 22466 2150 22480 2202
rect 22504 2150 22518 2202
rect 22518 2150 22530 2202
rect 22530 2150 22560 2202
rect 22584 2150 22594 2202
rect 22594 2150 22640 2202
rect 22344 2148 22400 2150
rect 22424 2148 22480 2150
rect 22504 2148 22560 2150
rect 22584 2148 22640 2150
rect 22926 1400 22982 1456
rect 23110 1536 23166 1592
rect 23294 2080 23350 2136
rect 33038 8730 33094 8732
rect 33118 8730 33174 8732
rect 33198 8730 33254 8732
rect 33278 8730 33334 8732
rect 33038 8678 33084 8730
rect 33084 8678 33094 8730
rect 33118 8678 33148 8730
rect 33148 8678 33160 8730
rect 33160 8678 33174 8730
rect 33198 8678 33212 8730
rect 33212 8678 33224 8730
rect 33224 8678 33254 8730
rect 33278 8678 33288 8730
rect 33288 8678 33334 8730
rect 33038 8676 33094 8678
rect 33118 8676 33174 8678
rect 33198 8676 33254 8678
rect 33278 8676 33334 8678
rect 43732 8730 43788 8732
rect 43812 8730 43868 8732
rect 43892 8730 43948 8732
rect 43972 8730 44028 8732
rect 43732 8678 43778 8730
rect 43778 8678 43788 8730
rect 43812 8678 43842 8730
rect 43842 8678 43854 8730
rect 43854 8678 43868 8730
rect 43892 8678 43906 8730
rect 43906 8678 43918 8730
rect 43918 8678 43948 8730
rect 43972 8678 43982 8730
rect 43982 8678 44028 8730
rect 43732 8676 43788 8678
rect 43812 8676 43868 8678
rect 43892 8676 43948 8678
rect 43972 8676 44028 8678
rect 22344 1114 22400 1116
rect 22424 1114 22480 1116
rect 22504 1114 22560 1116
rect 22584 1114 22640 1116
rect 22344 1062 22390 1114
rect 22390 1062 22400 1114
rect 22424 1062 22454 1114
rect 22454 1062 22466 1114
rect 22466 1062 22480 1114
rect 22504 1062 22518 1114
rect 22518 1062 22530 1114
rect 22530 1062 22560 1114
rect 22584 1062 22594 1114
rect 22594 1062 22640 1114
rect 22344 1060 22400 1062
rect 22424 1060 22480 1062
rect 22504 1060 22560 1062
rect 22584 1060 22640 1062
rect 23018 1128 23074 1184
rect 23662 1672 23718 1728
rect 24398 1808 24454 1864
rect 23938 1536 23994 1592
rect 23846 1400 23902 1456
rect 23754 584 23810 640
rect 24214 1264 24270 1320
rect 24950 2644 25006 2680
rect 26146 3032 26202 3088
rect 24950 2624 24952 2644
rect 24952 2624 25004 2644
rect 25004 2624 25006 2644
rect 24674 1536 24730 1592
rect 26146 2896 26202 2952
rect 26054 2624 26110 2680
rect 25502 584 25558 640
rect 27691 8186 27747 8188
rect 27771 8186 27827 8188
rect 27851 8186 27907 8188
rect 27931 8186 27987 8188
rect 27691 8134 27737 8186
rect 27737 8134 27747 8186
rect 27771 8134 27801 8186
rect 27801 8134 27813 8186
rect 27813 8134 27827 8186
rect 27851 8134 27865 8186
rect 27865 8134 27877 8186
rect 27877 8134 27907 8186
rect 27931 8134 27941 8186
rect 27941 8134 27987 8186
rect 27691 8132 27747 8134
rect 27771 8132 27827 8134
rect 27851 8132 27907 8134
rect 27931 8132 27987 8134
rect 27691 7098 27747 7100
rect 27771 7098 27827 7100
rect 27851 7098 27907 7100
rect 27931 7098 27987 7100
rect 27691 7046 27737 7098
rect 27737 7046 27747 7098
rect 27771 7046 27801 7098
rect 27801 7046 27813 7098
rect 27813 7046 27827 7098
rect 27851 7046 27865 7098
rect 27865 7046 27877 7098
rect 27877 7046 27907 7098
rect 27931 7046 27941 7098
rect 27941 7046 27987 7098
rect 27691 7044 27747 7046
rect 27771 7044 27827 7046
rect 27851 7044 27907 7046
rect 27931 7044 27987 7046
rect 27691 6010 27747 6012
rect 27771 6010 27827 6012
rect 27851 6010 27907 6012
rect 27931 6010 27987 6012
rect 27691 5958 27737 6010
rect 27737 5958 27747 6010
rect 27771 5958 27801 6010
rect 27801 5958 27813 6010
rect 27813 5958 27827 6010
rect 27851 5958 27865 6010
rect 27865 5958 27877 6010
rect 27877 5958 27907 6010
rect 27931 5958 27941 6010
rect 27941 5958 27987 6010
rect 27691 5956 27747 5958
rect 27771 5956 27827 5958
rect 27851 5956 27907 5958
rect 27931 5956 27987 5958
rect 27691 4922 27747 4924
rect 27771 4922 27827 4924
rect 27851 4922 27907 4924
rect 27931 4922 27987 4924
rect 27691 4870 27737 4922
rect 27737 4870 27747 4922
rect 27771 4870 27801 4922
rect 27801 4870 27813 4922
rect 27813 4870 27827 4922
rect 27851 4870 27865 4922
rect 27865 4870 27877 4922
rect 27877 4870 27907 4922
rect 27931 4870 27941 4922
rect 27941 4870 27987 4922
rect 27691 4868 27747 4870
rect 27771 4868 27827 4870
rect 27851 4868 27907 4870
rect 27931 4868 27987 4870
rect 27691 3834 27747 3836
rect 27771 3834 27827 3836
rect 27851 3834 27907 3836
rect 27931 3834 27987 3836
rect 27691 3782 27737 3834
rect 27737 3782 27747 3834
rect 27771 3782 27801 3834
rect 27801 3782 27813 3834
rect 27813 3782 27827 3834
rect 27851 3782 27865 3834
rect 27865 3782 27877 3834
rect 27877 3782 27907 3834
rect 27931 3782 27941 3834
rect 27941 3782 27987 3834
rect 27691 3780 27747 3782
rect 27771 3780 27827 3782
rect 27851 3780 27907 3782
rect 27931 3780 27987 3782
rect 27526 3712 27582 3768
rect 27250 2896 27306 2952
rect 26238 1536 26294 1592
rect 27342 2644 27398 2680
rect 27342 2624 27344 2644
rect 27344 2624 27396 2644
rect 27396 2624 27398 2644
rect 27691 2746 27747 2748
rect 27771 2746 27827 2748
rect 27851 2746 27907 2748
rect 27931 2746 27987 2748
rect 27691 2694 27737 2746
rect 27737 2694 27747 2746
rect 27771 2694 27801 2746
rect 27801 2694 27813 2746
rect 27813 2694 27827 2746
rect 27851 2694 27865 2746
rect 27865 2694 27877 2746
rect 27877 2694 27907 2746
rect 27931 2694 27941 2746
rect 27941 2694 27987 2746
rect 27691 2692 27747 2694
rect 27771 2692 27827 2694
rect 27851 2692 27907 2694
rect 27931 2692 27987 2694
rect 26606 1264 26662 1320
rect 27802 2252 27804 2272
rect 27804 2252 27856 2272
rect 27856 2252 27858 2272
rect 27802 2216 27858 2252
rect 27434 1844 27436 1864
rect 27436 1844 27488 1864
rect 27488 1844 27490 1864
rect 27434 1808 27490 1844
rect 27342 1672 27398 1728
rect 27691 1658 27747 1660
rect 27771 1658 27827 1660
rect 27851 1658 27907 1660
rect 27931 1658 27987 1660
rect 27691 1606 27737 1658
rect 27737 1606 27747 1658
rect 27771 1606 27801 1658
rect 27801 1606 27813 1658
rect 27813 1606 27827 1658
rect 27851 1606 27865 1658
rect 27865 1606 27877 1658
rect 27877 1606 27907 1658
rect 27931 1606 27941 1658
rect 27941 1606 27987 1658
rect 27691 1604 27747 1606
rect 27771 1604 27827 1606
rect 27851 1604 27907 1606
rect 27931 1604 27987 1606
rect 27802 1300 27804 1320
rect 27804 1300 27856 1320
rect 27856 1300 27858 1320
rect 27802 1264 27858 1300
rect 27894 584 27950 640
rect 28906 2896 28962 2952
rect 29182 2388 29184 2408
rect 29184 2388 29236 2408
rect 29236 2388 29238 2408
rect 29182 2352 29238 2388
rect 28722 2080 28778 2136
rect 28354 856 28410 912
rect 28722 1128 28778 1184
rect 30010 2488 30066 2544
rect 33038 7642 33094 7644
rect 33118 7642 33174 7644
rect 33198 7642 33254 7644
rect 33278 7642 33334 7644
rect 33038 7590 33084 7642
rect 33084 7590 33094 7642
rect 33118 7590 33148 7642
rect 33148 7590 33160 7642
rect 33160 7590 33174 7642
rect 33198 7590 33212 7642
rect 33212 7590 33224 7642
rect 33224 7590 33254 7642
rect 33278 7590 33288 7642
rect 33288 7590 33334 7642
rect 33038 7588 33094 7590
rect 33118 7588 33174 7590
rect 33198 7588 33254 7590
rect 33278 7588 33334 7590
rect 33038 6554 33094 6556
rect 33118 6554 33174 6556
rect 33198 6554 33254 6556
rect 33278 6554 33334 6556
rect 33038 6502 33084 6554
rect 33084 6502 33094 6554
rect 33118 6502 33148 6554
rect 33148 6502 33160 6554
rect 33160 6502 33174 6554
rect 33198 6502 33212 6554
rect 33212 6502 33224 6554
rect 33224 6502 33254 6554
rect 33278 6502 33288 6554
rect 33288 6502 33334 6554
rect 33038 6500 33094 6502
rect 33118 6500 33174 6502
rect 33198 6500 33254 6502
rect 33278 6500 33334 6502
rect 33038 5466 33094 5468
rect 33118 5466 33174 5468
rect 33198 5466 33254 5468
rect 33278 5466 33334 5468
rect 33038 5414 33084 5466
rect 33084 5414 33094 5466
rect 33118 5414 33148 5466
rect 33148 5414 33160 5466
rect 33160 5414 33174 5466
rect 33198 5414 33212 5466
rect 33212 5414 33224 5466
rect 33224 5414 33254 5466
rect 33278 5414 33288 5466
rect 33288 5414 33334 5466
rect 33038 5412 33094 5414
rect 33118 5412 33174 5414
rect 33198 5412 33254 5414
rect 33278 5412 33334 5414
rect 33038 4378 33094 4380
rect 33118 4378 33174 4380
rect 33198 4378 33254 4380
rect 33278 4378 33334 4380
rect 33038 4326 33084 4378
rect 33084 4326 33094 4378
rect 33118 4326 33148 4378
rect 33148 4326 33160 4378
rect 33160 4326 33174 4378
rect 33198 4326 33212 4378
rect 33212 4326 33224 4378
rect 33224 4326 33254 4378
rect 33278 4326 33288 4378
rect 33288 4326 33334 4378
rect 33038 4324 33094 4326
rect 33118 4324 33174 4326
rect 33198 4324 33254 4326
rect 33278 4324 33334 4326
rect 32862 3440 32918 3496
rect 31114 3304 31170 3360
rect 30930 2216 30986 2272
rect 30746 1400 30802 1456
rect 33038 3290 33094 3292
rect 33118 3290 33174 3292
rect 33198 3290 33254 3292
rect 33278 3290 33334 3292
rect 33038 3238 33084 3290
rect 33084 3238 33094 3290
rect 33118 3238 33148 3290
rect 33148 3238 33160 3290
rect 33160 3238 33174 3290
rect 33198 3238 33212 3290
rect 33212 3238 33224 3290
rect 33224 3238 33254 3290
rect 33278 3238 33288 3290
rect 33288 3238 33334 3290
rect 33038 3236 33094 3238
rect 33118 3236 33174 3238
rect 33198 3236 33254 3238
rect 33278 3236 33334 3238
rect 33414 3032 33470 3088
rect 31850 2216 31906 2272
rect 31942 720 31998 776
rect 33038 2202 33094 2204
rect 33118 2202 33174 2204
rect 33198 2202 33254 2204
rect 33278 2202 33334 2204
rect 33038 2150 33084 2202
rect 33084 2150 33094 2202
rect 33118 2150 33148 2202
rect 33148 2150 33160 2202
rect 33160 2150 33174 2202
rect 33198 2150 33212 2202
rect 33212 2150 33224 2202
rect 33224 2150 33254 2202
rect 33278 2150 33288 2202
rect 33288 2150 33334 2202
rect 33038 2148 33094 2150
rect 33118 2148 33174 2150
rect 33198 2148 33254 2150
rect 33278 2148 33334 2150
rect 33874 3984 33930 4040
rect 33038 1114 33094 1116
rect 33118 1114 33174 1116
rect 33198 1114 33254 1116
rect 33278 1114 33334 1116
rect 33038 1062 33084 1114
rect 33084 1062 33094 1114
rect 33118 1062 33148 1114
rect 33148 1062 33160 1114
rect 33160 1062 33174 1114
rect 33198 1062 33212 1114
rect 33212 1062 33224 1114
rect 33224 1062 33254 1114
rect 33278 1062 33288 1114
rect 33288 1062 33334 1114
rect 33038 1060 33094 1062
rect 33118 1060 33174 1062
rect 33198 1060 33254 1062
rect 33278 1060 33334 1062
rect 35070 1300 35072 1320
rect 35072 1300 35124 1320
rect 35124 1300 35126 1320
rect 34610 448 34666 504
rect 35070 1264 35126 1300
rect 36542 1944 36598 2000
rect 38385 8186 38441 8188
rect 38465 8186 38521 8188
rect 38545 8186 38601 8188
rect 38625 8186 38681 8188
rect 38385 8134 38431 8186
rect 38431 8134 38441 8186
rect 38465 8134 38495 8186
rect 38495 8134 38507 8186
rect 38507 8134 38521 8186
rect 38545 8134 38559 8186
rect 38559 8134 38571 8186
rect 38571 8134 38601 8186
rect 38625 8134 38635 8186
rect 38635 8134 38681 8186
rect 38385 8132 38441 8134
rect 38465 8132 38521 8134
rect 38545 8132 38601 8134
rect 38625 8132 38681 8134
rect 38385 7098 38441 7100
rect 38465 7098 38521 7100
rect 38545 7098 38601 7100
rect 38625 7098 38681 7100
rect 38385 7046 38431 7098
rect 38431 7046 38441 7098
rect 38465 7046 38495 7098
rect 38495 7046 38507 7098
rect 38507 7046 38521 7098
rect 38545 7046 38559 7098
rect 38559 7046 38571 7098
rect 38571 7046 38601 7098
rect 38625 7046 38635 7098
rect 38635 7046 38681 7098
rect 38385 7044 38441 7046
rect 38465 7044 38521 7046
rect 38545 7044 38601 7046
rect 38625 7044 38681 7046
rect 38385 6010 38441 6012
rect 38465 6010 38521 6012
rect 38545 6010 38601 6012
rect 38625 6010 38681 6012
rect 38385 5958 38431 6010
rect 38431 5958 38441 6010
rect 38465 5958 38495 6010
rect 38495 5958 38507 6010
rect 38507 5958 38521 6010
rect 38545 5958 38559 6010
rect 38559 5958 38571 6010
rect 38571 5958 38601 6010
rect 38625 5958 38635 6010
rect 38635 5958 38681 6010
rect 38385 5956 38441 5958
rect 38465 5956 38521 5958
rect 38545 5956 38601 5958
rect 38625 5956 38681 5958
rect 38385 4922 38441 4924
rect 38465 4922 38521 4924
rect 38545 4922 38601 4924
rect 38625 4922 38681 4924
rect 38385 4870 38431 4922
rect 38431 4870 38441 4922
rect 38465 4870 38495 4922
rect 38495 4870 38507 4922
rect 38507 4870 38521 4922
rect 38545 4870 38559 4922
rect 38559 4870 38571 4922
rect 38571 4870 38601 4922
rect 38625 4870 38635 4922
rect 38635 4870 38681 4922
rect 38385 4868 38441 4870
rect 38465 4868 38521 4870
rect 38545 4868 38601 4870
rect 38625 4868 38681 4870
rect 38385 3834 38441 3836
rect 38465 3834 38521 3836
rect 38545 3834 38601 3836
rect 38625 3834 38681 3836
rect 38385 3782 38431 3834
rect 38431 3782 38441 3834
rect 38465 3782 38495 3834
rect 38495 3782 38507 3834
rect 38507 3782 38521 3834
rect 38545 3782 38559 3834
rect 38559 3782 38571 3834
rect 38571 3782 38601 3834
rect 38625 3782 38635 3834
rect 38635 3782 38681 3834
rect 38385 3780 38441 3782
rect 38465 3780 38521 3782
rect 38545 3780 38601 3782
rect 38625 3780 38681 3782
rect 38385 2746 38441 2748
rect 38465 2746 38521 2748
rect 38545 2746 38601 2748
rect 38625 2746 38681 2748
rect 38385 2694 38431 2746
rect 38431 2694 38441 2746
rect 38465 2694 38495 2746
rect 38495 2694 38507 2746
rect 38507 2694 38521 2746
rect 38545 2694 38559 2746
rect 38559 2694 38571 2746
rect 38571 2694 38601 2746
rect 38625 2694 38635 2746
rect 38635 2694 38681 2746
rect 38385 2692 38441 2694
rect 38465 2692 38521 2694
rect 38545 2692 38601 2694
rect 38625 2692 38681 2694
rect 38385 1658 38441 1660
rect 38465 1658 38521 1660
rect 38545 1658 38601 1660
rect 38625 1658 38681 1660
rect 38385 1606 38431 1658
rect 38431 1606 38441 1658
rect 38465 1606 38495 1658
rect 38495 1606 38507 1658
rect 38507 1606 38521 1658
rect 38545 1606 38559 1658
rect 38559 1606 38571 1658
rect 38571 1606 38601 1658
rect 38625 1606 38635 1658
rect 38635 1606 38681 1658
rect 38385 1604 38441 1606
rect 38465 1604 38521 1606
rect 38545 1604 38601 1606
rect 38625 1604 38681 1606
rect 43732 7642 43788 7644
rect 43812 7642 43868 7644
rect 43892 7642 43948 7644
rect 43972 7642 44028 7644
rect 43732 7590 43778 7642
rect 43778 7590 43788 7642
rect 43812 7590 43842 7642
rect 43842 7590 43854 7642
rect 43854 7590 43868 7642
rect 43892 7590 43906 7642
rect 43906 7590 43918 7642
rect 43918 7590 43948 7642
rect 43972 7590 43982 7642
rect 43982 7590 44028 7642
rect 43732 7588 43788 7590
rect 43812 7588 43868 7590
rect 43892 7588 43948 7590
rect 43972 7588 44028 7590
rect 43732 6554 43788 6556
rect 43812 6554 43868 6556
rect 43892 6554 43948 6556
rect 43972 6554 44028 6556
rect 43732 6502 43778 6554
rect 43778 6502 43788 6554
rect 43812 6502 43842 6554
rect 43842 6502 43854 6554
rect 43854 6502 43868 6554
rect 43892 6502 43906 6554
rect 43906 6502 43918 6554
rect 43918 6502 43948 6554
rect 43972 6502 43982 6554
rect 43982 6502 44028 6554
rect 43732 6500 43788 6502
rect 43812 6500 43868 6502
rect 43892 6500 43948 6502
rect 43972 6500 44028 6502
rect 43732 5466 43788 5468
rect 43812 5466 43868 5468
rect 43892 5466 43948 5468
rect 43972 5466 44028 5468
rect 43732 5414 43778 5466
rect 43778 5414 43788 5466
rect 43812 5414 43842 5466
rect 43842 5414 43854 5466
rect 43854 5414 43868 5466
rect 43892 5414 43906 5466
rect 43906 5414 43918 5466
rect 43918 5414 43948 5466
rect 43972 5414 43982 5466
rect 43982 5414 44028 5466
rect 43732 5412 43788 5414
rect 43812 5412 43868 5414
rect 43892 5412 43948 5414
rect 43972 5412 44028 5414
rect 43732 4378 43788 4380
rect 43812 4378 43868 4380
rect 43892 4378 43948 4380
rect 43972 4378 44028 4380
rect 43732 4326 43778 4378
rect 43778 4326 43788 4378
rect 43812 4326 43842 4378
rect 43842 4326 43854 4378
rect 43854 4326 43868 4378
rect 43892 4326 43906 4378
rect 43906 4326 43918 4378
rect 43918 4326 43948 4378
rect 43972 4326 43982 4378
rect 43982 4326 44028 4378
rect 43732 4324 43788 4326
rect 43812 4324 43868 4326
rect 43892 4324 43948 4326
rect 43972 4324 44028 4326
rect 43732 3290 43788 3292
rect 43812 3290 43868 3292
rect 43892 3290 43948 3292
rect 43972 3290 44028 3292
rect 43732 3238 43778 3290
rect 43778 3238 43788 3290
rect 43812 3238 43842 3290
rect 43842 3238 43854 3290
rect 43854 3238 43868 3290
rect 43892 3238 43906 3290
rect 43906 3238 43918 3290
rect 43918 3238 43948 3290
rect 43972 3238 43982 3290
rect 43982 3238 44028 3290
rect 43732 3236 43788 3238
rect 43812 3236 43868 3238
rect 43892 3236 43948 3238
rect 43972 3236 44028 3238
rect 43732 2202 43788 2204
rect 43812 2202 43868 2204
rect 43892 2202 43948 2204
rect 43972 2202 44028 2204
rect 43732 2150 43778 2202
rect 43778 2150 43788 2202
rect 43812 2150 43842 2202
rect 43842 2150 43854 2202
rect 43854 2150 43868 2202
rect 43892 2150 43906 2202
rect 43906 2150 43918 2202
rect 43918 2150 43948 2202
rect 43972 2150 43982 2202
rect 43982 2150 44028 2202
rect 43732 2148 43788 2150
rect 43812 2148 43868 2150
rect 43892 2148 43948 2150
rect 43972 2148 44028 2150
rect 38566 720 38622 776
rect 43732 1114 43788 1116
rect 43812 1114 43868 1116
rect 43892 1114 43948 1116
rect 43972 1114 44028 1116
rect 43732 1062 43778 1114
rect 43778 1062 43788 1114
rect 43812 1062 43842 1114
rect 43842 1062 43854 1114
rect 43854 1062 43868 1114
rect 43892 1062 43906 1114
rect 43906 1062 43918 1114
rect 43918 1062 43948 1114
rect 43972 1062 43982 1114
rect 43982 1062 44028 1114
rect 43732 1060 43788 1062
rect 43812 1060 43868 1062
rect 43892 1060 43948 1062
rect 43972 1060 44028 1062
<< metal3 >>
rect 11640 8736 11956 8737
rect 11640 8672 11646 8736
rect 11710 8672 11726 8736
rect 11790 8672 11806 8736
rect 11870 8672 11886 8736
rect 11950 8672 11956 8736
rect 11640 8671 11956 8672
rect 22334 8736 22650 8737
rect 22334 8672 22340 8736
rect 22404 8672 22420 8736
rect 22484 8672 22500 8736
rect 22564 8672 22580 8736
rect 22644 8672 22650 8736
rect 22334 8671 22650 8672
rect 33028 8736 33344 8737
rect 33028 8672 33034 8736
rect 33098 8672 33114 8736
rect 33178 8672 33194 8736
rect 33258 8672 33274 8736
rect 33338 8672 33344 8736
rect 33028 8671 33344 8672
rect 43722 8736 44038 8737
rect 43722 8672 43728 8736
rect 43792 8672 43808 8736
rect 43872 8672 43888 8736
rect 43952 8672 43968 8736
rect 44032 8672 44038 8736
rect 43722 8671 44038 8672
rect 5533 8530 5599 8533
rect 24894 8530 24900 8532
rect 5533 8528 24900 8530
rect 5533 8472 5538 8528
rect 5594 8472 24900 8528
rect 5533 8470 24900 8472
rect 5533 8467 5599 8470
rect 24894 8468 24900 8470
rect 24964 8468 24970 8532
rect 4429 8394 4495 8397
rect 25078 8394 25084 8396
rect 4429 8392 25084 8394
rect 4429 8336 4434 8392
rect 4490 8336 25084 8392
rect 4429 8334 25084 8336
rect 4429 8331 4495 8334
rect 25078 8332 25084 8334
rect 25148 8332 25154 8396
rect 6293 8192 6609 8193
rect 6293 8128 6299 8192
rect 6363 8128 6379 8192
rect 6443 8128 6459 8192
rect 6523 8128 6539 8192
rect 6603 8128 6609 8192
rect 6293 8127 6609 8128
rect 16987 8192 17303 8193
rect 16987 8128 16993 8192
rect 17057 8128 17073 8192
rect 17137 8128 17153 8192
rect 17217 8128 17233 8192
rect 17297 8128 17303 8192
rect 16987 8127 17303 8128
rect 27681 8192 27997 8193
rect 27681 8128 27687 8192
rect 27751 8128 27767 8192
rect 27831 8128 27847 8192
rect 27911 8128 27927 8192
rect 27991 8128 27997 8192
rect 27681 8127 27997 8128
rect 38375 8192 38691 8193
rect 38375 8128 38381 8192
rect 38445 8128 38461 8192
rect 38525 8128 38541 8192
rect 38605 8128 38621 8192
rect 38685 8128 38691 8192
rect 38375 8127 38691 8128
rect 11640 7648 11956 7649
rect 11640 7584 11646 7648
rect 11710 7584 11726 7648
rect 11790 7584 11806 7648
rect 11870 7584 11886 7648
rect 11950 7584 11956 7648
rect 11640 7583 11956 7584
rect 22334 7648 22650 7649
rect 22334 7584 22340 7648
rect 22404 7584 22420 7648
rect 22484 7584 22500 7648
rect 22564 7584 22580 7648
rect 22644 7584 22650 7648
rect 22334 7583 22650 7584
rect 33028 7648 33344 7649
rect 33028 7584 33034 7648
rect 33098 7584 33114 7648
rect 33178 7584 33194 7648
rect 33258 7584 33274 7648
rect 33338 7584 33344 7648
rect 33028 7583 33344 7584
rect 43722 7648 44038 7649
rect 43722 7584 43728 7648
rect 43792 7584 43808 7648
rect 43872 7584 43888 7648
rect 43952 7584 43968 7648
rect 44032 7584 44038 7648
rect 43722 7583 44038 7584
rect 6293 7104 6609 7105
rect 6293 7040 6299 7104
rect 6363 7040 6379 7104
rect 6443 7040 6459 7104
rect 6523 7040 6539 7104
rect 6603 7040 6609 7104
rect 6293 7039 6609 7040
rect 16987 7104 17303 7105
rect 16987 7040 16993 7104
rect 17057 7040 17073 7104
rect 17137 7040 17153 7104
rect 17217 7040 17233 7104
rect 17297 7040 17303 7104
rect 16987 7039 17303 7040
rect 27681 7104 27997 7105
rect 27681 7040 27687 7104
rect 27751 7040 27767 7104
rect 27831 7040 27847 7104
rect 27911 7040 27927 7104
rect 27991 7040 27997 7104
rect 27681 7039 27997 7040
rect 38375 7104 38691 7105
rect 38375 7040 38381 7104
rect 38445 7040 38461 7104
rect 38525 7040 38541 7104
rect 38605 7040 38621 7104
rect 38685 7040 38691 7104
rect 38375 7039 38691 7040
rect 11640 6560 11956 6561
rect 11640 6496 11646 6560
rect 11710 6496 11726 6560
rect 11790 6496 11806 6560
rect 11870 6496 11886 6560
rect 11950 6496 11956 6560
rect 11640 6495 11956 6496
rect 22334 6560 22650 6561
rect 22334 6496 22340 6560
rect 22404 6496 22420 6560
rect 22484 6496 22500 6560
rect 22564 6496 22580 6560
rect 22644 6496 22650 6560
rect 22334 6495 22650 6496
rect 33028 6560 33344 6561
rect 33028 6496 33034 6560
rect 33098 6496 33114 6560
rect 33178 6496 33194 6560
rect 33258 6496 33274 6560
rect 33338 6496 33344 6560
rect 33028 6495 33344 6496
rect 43722 6560 44038 6561
rect 43722 6496 43728 6560
rect 43792 6496 43808 6560
rect 43872 6496 43888 6560
rect 43952 6496 43968 6560
rect 44032 6496 44038 6560
rect 43722 6495 44038 6496
rect 6293 6016 6609 6017
rect 6293 5952 6299 6016
rect 6363 5952 6379 6016
rect 6443 5952 6459 6016
rect 6523 5952 6539 6016
rect 6603 5952 6609 6016
rect 6293 5951 6609 5952
rect 16987 6016 17303 6017
rect 16987 5952 16993 6016
rect 17057 5952 17073 6016
rect 17137 5952 17153 6016
rect 17217 5952 17233 6016
rect 17297 5952 17303 6016
rect 16987 5951 17303 5952
rect 27681 6016 27997 6017
rect 27681 5952 27687 6016
rect 27751 5952 27767 6016
rect 27831 5952 27847 6016
rect 27911 5952 27927 6016
rect 27991 5952 27997 6016
rect 27681 5951 27997 5952
rect 38375 6016 38691 6017
rect 38375 5952 38381 6016
rect 38445 5952 38461 6016
rect 38525 5952 38541 6016
rect 38605 5952 38621 6016
rect 38685 5952 38691 6016
rect 38375 5951 38691 5952
rect 11640 5472 11956 5473
rect 11640 5408 11646 5472
rect 11710 5408 11726 5472
rect 11790 5408 11806 5472
rect 11870 5408 11886 5472
rect 11950 5408 11956 5472
rect 11640 5407 11956 5408
rect 22334 5472 22650 5473
rect 22334 5408 22340 5472
rect 22404 5408 22420 5472
rect 22484 5408 22500 5472
rect 22564 5408 22580 5472
rect 22644 5408 22650 5472
rect 22334 5407 22650 5408
rect 33028 5472 33344 5473
rect 33028 5408 33034 5472
rect 33098 5408 33114 5472
rect 33178 5408 33194 5472
rect 33258 5408 33274 5472
rect 33338 5408 33344 5472
rect 33028 5407 33344 5408
rect 43722 5472 44038 5473
rect 43722 5408 43728 5472
rect 43792 5408 43808 5472
rect 43872 5408 43888 5472
rect 43952 5408 43968 5472
rect 44032 5408 44038 5472
rect 43722 5407 44038 5408
rect 6293 4928 6609 4929
rect 6293 4864 6299 4928
rect 6363 4864 6379 4928
rect 6443 4864 6459 4928
rect 6523 4864 6539 4928
rect 6603 4864 6609 4928
rect 6293 4863 6609 4864
rect 16987 4928 17303 4929
rect 16987 4864 16993 4928
rect 17057 4864 17073 4928
rect 17137 4864 17153 4928
rect 17217 4864 17233 4928
rect 17297 4864 17303 4928
rect 16987 4863 17303 4864
rect 27681 4928 27997 4929
rect 27681 4864 27687 4928
rect 27751 4864 27767 4928
rect 27831 4864 27847 4928
rect 27911 4864 27927 4928
rect 27991 4864 27997 4928
rect 27681 4863 27997 4864
rect 38375 4928 38691 4929
rect 38375 4864 38381 4928
rect 38445 4864 38461 4928
rect 38525 4864 38541 4928
rect 38605 4864 38621 4928
rect 38685 4864 38691 4928
rect 38375 4863 38691 4864
rect 11640 4384 11956 4385
rect 11640 4320 11646 4384
rect 11710 4320 11726 4384
rect 11790 4320 11806 4384
rect 11870 4320 11886 4384
rect 11950 4320 11956 4384
rect 11640 4319 11956 4320
rect 22334 4384 22650 4385
rect 22334 4320 22340 4384
rect 22404 4320 22420 4384
rect 22484 4320 22500 4384
rect 22564 4320 22580 4384
rect 22644 4320 22650 4384
rect 22334 4319 22650 4320
rect 33028 4384 33344 4385
rect 33028 4320 33034 4384
rect 33098 4320 33114 4384
rect 33178 4320 33194 4384
rect 33258 4320 33274 4384
rect 33338 4320 33344 4384
rect 33028 4319 33344 4320
rect 43722 4384 44038 4385
rect 43722 4320 43728 4384
rect 43792 4320 43808 4384
rect 43872 4320 43888 4384
rect 43952 4320 43968 4384
rect 44032 4320 44038 4384
rect 43722 4319 44038 4320
rect 12525 4042 12591 4045
rect 18229 4042 18295 4045
rect 33869 4042 33935 4045
rect 12525 4040 17464 4042
rect 12525 3984 12530 4040
rect 12586 3984 17464 4040
rect 12525 3982 17464 3984
rect 12525 3979 12591 3982
rect 17404 3906 17464 3982
rect 18229 4040 33935 4042
rect 18229 3984 18234 4040
rect 18290 3984 33874 4040
rect 33930 3984 33935 4040
rect 18229 3982 33935 3984
rect 18229 3979 18295 3982
rect 33869 3979 33935 3982
rect 17404 3846 22110 3906
rect 6293 3840 6609 3841
rect 6293 3776 6299 3840
rect 6363 3776 6379 3840
rect 6443 3776 6459 3840
rect 6523 3776 6539 3840
rect 6603 3776 6609 3840
rect 6293 3775 6609 3776
rect 16987 3840 17303 3841
rect 16987 3776 16993 3840
rect 17057 3776 17073 3840
rect 17137 3776 17153 3840
rect 17217 3776 17233 3840
rect 17297 3776 17303 3840
rect 16987 3775 17303 3776
rect 22050 3770 22110 3846
rect 27681 3840 27997 3841
rect 27681 3776 27687 3840
rect 27751 3776 27767 3840
rect 27831 3776 27847 3840
rect 27911 3776 27927 3840
rect 27991 3776 27997 3840
rect 27681 3775 27997 3776
rect 38375 3840 38691 3841
rect 38375 3776 38381 3840
rect 38445 3776 38461 3840
rect 38525 3776 38541 3840
rect 38605 3776 38621 3840
rect 38685 3776 38691 3840
rect 38375 3775 38691 3776
rect 27521 3770 27587 3773
rect 22050 3768 27587 3770
rect 22050 3712 27526 3768
rect 27582 3712 27587 3768
rect 22050 3710 27587 3712
rect 27521 3707 27587 3710
rect 15377 3634 15443 3637
rect 34462 3634 34468 3636
rect 15377 3632 34468 3634
rect 15377 3576 15382 3632
rect 15438 3576 34468 3632
rect 15377 3574 34468 3576
rect 15377 3571 15443 3574
rect 34462 3572 34468 3574
rect 34532 3572 34538 3636
rect 16849 3498 16915 3501
rect 32857 3498 32923 3501
rect 16849 3496 32923 3498
rect 16849 3440 16854 3496
rect 16910 3440 32862 3496
rect 32918 3440 32923 3496
rect 16849 3438 32923 3440
rect 16849 3435 16915 3438
rect 32857 3435 32923 3438
rect 31109 3362 31175 3365
rect 26052 3360 31175 3362
rect 26052 3304 31114 3360
rect 31170 3304 31175 3360
rect 26052 3302 31175 3304
rect 11640 3296 11956 3297
rect 11640 3232 11646 3296
rect 11710 3232 11726 3296
rect 11790 3232 11806 3296
rect 11870 3232 11886 3296
rect 11950 3232 11956 3296
rect 11640 3231 11956 3232
rect 22334 3296 22650 3297
rect 22334 3232 22340 3296
rect 22404 3232 22420 3296
rect 22484 3232 22500 3296
rect 22564 3232 22580 3296
rect 22644 3232 22650 3296
rect 22334 3231 22650 3232
rect 14365 3226 14431 3229
rect 21541 3226 21607 3229
rect 26052 3226 26112 3302
rect 31109 3299 31175 3302
rect 33028 3296 33344 3297
rect 33028 3232 33034 3296
rect 33098 3232 33114 3296
rect 33178 3232 33194 3296
rect 33258 3232 33274 3296
rect 33338 3232 33344 3296
rect 33028 3231 33344 3232
rect 43722 3296 44038 3297
rect 43722 3232 43728 3296
rect 43792 3232 43808 3296
rect 43872 3232 43888 3296
rect 43952 3232 43968 3296
rect 44032 3232 44038 3296
rect 43722 3231 44038 3232
rect 14365 3224 21607 3226
rect 14365 3168 14370 3224
rect 14426 3168 21546 3224
rect 21602 3168 21607 3224
rect 14365 3166 21607 3168
rect 14365 3163 14431 3166
rect 21541 3163 21607 3166
rect 26006 3166 26112 3226
rect 18505 3090 18571 3093
rect 26006 3090 26066 3166
rect 18505 3088 26066 3090
rect 18505 3032 18510 3088
rect 18566 3032 26066 3088
rect 18505 3030 26066 3032
rect 26141 3090 26207 3093
rect 33409 3090 33475 3093
rect 26141 3088 33475 3090
rect 26141 3032 26146 3088
rect 26202 3032 33414 3088
rect 33470 3032 33475 3088
rect 26141 3030 33475 3032
rect 18505 3027 18571 3030
rect 26141 3027 26207 3030
rect 33409 3027 33475 3030
rect 16205 2954 16271 2957
rect 21541 2954 21607 2957
rect 26141 2954 26207 2957
rect 16205 2952 21466 2954
rect 16205 2896 16210 2952
rect 16266 2896 21466 2952
rect 16205 2894 21466 2896
rect 16205 2891 16271 2894
rect 21406 2820 21466 2894
rect 21541 2952 26207 2954
rect 21541 2896 21546 2952
rect 21602 2896 26146 2952
rect 26202 2896 26207 2952
rect 21541 2894 26207 2896
rect 21541 2891 21607 2894
rect 26141 2891 26207 2894
rect 27245 2954 27311 2957
rect 28901 2954 28967 2957
rect 27245 2952 28967 2954
rect 27245 2896 27250 2952
rect 27306 2896 28906 2952
rect 28962 2896 28967 2952
rect 27245 2894 28967 2896
rect 27245 2891 27311 2894
rect 28901 2891 28967 2894
rect 21398 2756 21404 2820
rect 21468 2756 21474 2820
rect 6293 2752 6609 2753
rect 6293 2688 6299 2752
rect 6363 2688 6379 2752
rect 6443 2688 6459 2752
rect 6523 2688 6539 2752
rect 6603 2688 6609 2752
rect 6293 2687 6609 2688
rect 16987 2752 17303 2753
rect 16987 2688 16993 2752
rect 17057 2688 17073 2752
rect 17137 2688 17153 2752
rect 17217 2688 17233 2752
rect 17297 2688 17303 2752
rect 16987 2687 17303 2688
rect 27681 2752 27997 2753
rect 27681 2688 27687 2752
rect 27751 2688 27767 2752
rect 27831 2688 27847 2752
rect 27911 2688 27927 2752
rect 27991 2688 27997 2752
rect 27681 2687 27997 2688
rect 38375 2752 38691 2753
rect 38375 2688 38381 2752
rect 38445 2688 38461 2752
rect 38525 2688 38541 2752
rect 38605 2688 38621 2752
rect 38685 2688 38691 2752
rect 38375 2687 38691 2688
rect 17401 2682 17467 2685
rect 24945 2684 25011 2685
rect 17401 2680 24778 2682
rect 17401 2624 17406 2680
rect 17462 2624 24778 2680
rect 17401 2622 24778 2624
rect 17401 2619 17467 2622
rect 8477 2546 8543 2549
rect 22369 2546 22435 2549
rect 8477 2544 22435 2546
rect 8477 2488 8482 2544
rect 8538 2488 22374 2544
rect 22430 2488 22435 2544
rect 8477 2486 22435 2488
rect 24718 2546 24778 2622
rect 24894 2620 24900 2684
rect 24964 2682 25011 2684
rect 26049 2682 26115 2685
rect 27337 2682 27403 2685
rect 24964 2680 25056 2682
rect 25006 2624 25056 2680
rect 24964 2622 25056 2624
rect 26049 2680 27403 2682
rect 26049 2624 26054 2680
rect 26110 2624 27342 2680
rect 27398 2624 27403 2680
rect 26049 2622 27403 2624
rect 24964 2620 25011 2622
rect 24945 2619 25011 2620
rect 26049 2619 26115 2622
rect 27337 2619 27403 2622
rect 30005 2546 30071 2549
rect 24718 2544 30071 2546
rect 24718 2488 30010 2544
rect 30066 2488 30071 2544
rect 24718 2486 30071 2488
rect 8477 2483 8543 2486
rect 22369 2483 22435 2486
rect 30005 2483 30071 2486
rect 12065 2410 12131 2413
rect 29177 2410 29243 2413
rect 12065 2408 29243 2410
rect 12065 2352 12070 2408
rect 12126 2352 29182 2408
rect 29238 2352 29243 2408
rect 12065 2350 29243 2352
rect 12065 2347 12131 2350
rect 29177 2347 29243 2350
rect 17401 2274 17467 2277
rect 18965 2274 19031 2277
rect 12022 2272 17467 2274
rect 12022 2216 17406 2272
rect 17462 2216 17467 2272
rect 12022 2214 17467 2216
rect 11640 2208 11956 2209
rect 11640 2144 11646 2208
rect 11710 2144 11726 2208
rect 11790 2144 11806 2208
rect 11870 2144 11886 2208
rect 11950 2144 11956 2208
rect 11640 2143 11956 2144
rect 10777 2002 10843 2005
rect 12022 2002 12082 2214
rect 17401 2211 17467 2214
rect 17542 2272 19031 2274
rect 17542 2216 18970 2272
rect 19026 2216 19031 2272
rect 17542 2214 19031 2216
rect 13905 2138 13971 2141
rect 17542 2138 17602 2214
rect 18965 2211 19031 2214
rect 25078 2212 25084 2276
rect 25148 2274 25154 2276
rect 27797 2274 27863 2277
rect 25148 2272 27863 2274
rect 25148 2216 27802 2272
rect 27858 2216 27863 2272
rect 25148 2214 27863 2216
rect 25148 2212 25154 2214
rect 27797 2211 27863 2214
rect 30925 2274 30991 2277
rect 31845 2274 31911 2277
rect 30925 2272 31911 2274
rect 30925 2216 30930 2272
rect 30986 2216 31850 2272
rect 31906 2216 31911 2272
rect 30925 2214 31911 2216
rect 30925 2211 30991 2214
rect 31845 2211 31911 2214
rect 22334 2208 22650 2209
rect 22334 2144 22340 2208
rect 22404 2144 22420 2208
rect 22484 2144 22500 2208
rect 22564 2144 22580 2208
rect 22644 2144 22650 2208
rect 22334 2143 22650 2144
rect 33028 2208 33344 2209
rect 33028 2144 33034 2208
rect 33098 2144 33114 2208
rect 33178 2144 33194 2208
rect 33258 2144 33274 2208
rect 33338 2144 33344 2208
rect 33028 2143 33344 2144
rect 43722 2208 44038 2209
rect 43722 2144 43728 2208
rect 43792 2144 43808 2208
rect 43872 2144 43888 2208
rect 43952 2144 43968 2208
rect 44032 2144 44038 2208
rect 43722 2143 44038 2144
rect 13905 2136 17602 2138
rect 13905 2080 13910 2136
rect 13966 2080 17602 2136
rect 13905 2078 17602 2080
rect 18321 2138 18387 2141
rect 23289 2138 23355 2141
rect 28717 2138 28783 2141
rect 18321 2136 22110 2138
rect 18321 2080 18326 2136
rect 18382 2080 22110 2136
rect 18321 2078 22110 2080
rect 13905 2075 13971 2078
rect 18321 2075 18387 2078
rect 10777 2000 12082 2002
rect 10777 1944 10782 2000
rect 10838 1944 12082 2000
rect 10777 1942 12082 1944
rect 13537 2002 13603 2005
rect 22050 2002 22110 2078
rect 23289 2136 28783 2138
rect 23289 2080 23294 2136
rect 23350 2080 28722 2136
rect 28778 2080 28783 2136
rect 23289 2078 28783 2080
rect 23289 2075 23355 2078
rect 28717 2075 28783 2078
rect 36537 2002 36603 2005
rect 13537 2000 18338 2002
rect 13537 1944 13542 2000
rect 13598 1944 18338 2000
rect 13537 1942 18338 1944
rect 22050 2000 36603 2002
rect 22050 1944 36542 2000
rect 36598 1944 36603 2000
rect 22050 1942 36603 1944
rect 10777 1939 10843 1942
rect 13537 1939 13603 1942
rect 10685 1866 10751 1869
rect 18045 1866 18111 1869
rect 10685 1864 18111 1866
rect 10685 1808 10690 1864
rect 10746 1808 18050 1864
rect 18106 1808 18111 1864
rect 10685 1806 18111 1808
rect 18278 1866 18338 1942
rect 36537 1939 36603 1942
rect 24393 1866 24459 1869
rect 27429 1866 27495 1869
rect 18278 1806 23858 1866
rect 10685 1803 10751 1806
rect 18045 1803 18111 1806
rect 17401 1730 17467 1733
rect 23657 1730 23723 1733
rect 17401 1728 23723 1730
rect 17401 1672 17406 1728
rect 17462 1672 23662 1728
rect 23718 1672 23723 1728
rect 17401 1670 23723 1672
rect 23798 1730 23858 1806
rect 24393 1864 27495 1866
rect 24393 1808 24398 1864
rect 24454 1808 27434 1864
rect 27490 1808 27495 1864
rect 24393 1806 27495 1808
rect 24393 1803 24459 1806
rect 27429 1803 27495 1806
rect 27337 1730 27403 1733
rect 23798 1728 27403 1730
rect 23798 1672 27342 1728
rect 27398 1672 27403 1728
rect 23798 1670 27403 1672
rect 17401 1667 17467 1670
rect 23657 1667 23723 1670
rect 27337 1667 27403 1670
rect 6293 1664 6609 1665
rect 6293 1600 6299 1664
rect 6363 1600 6379 1664
rect 6443 1600 6459 1664
rect 6523 1600 6539 1664
rect 6603 1600 6609 1664
rect 6293 1599 6609 1600
rect 16987 1664 17303 1665
rect 16987 1600 16993 1664
rect 17057 1600 17073 1664
rect 17137 1600 17153 1664
rect 17217 1600 17233 1664
rect 17297 1600 17303 1664
rect 16987 1599 17303 1600
rect 27681 1664 27997 1665
rect 27681 1600 27687 1664
rect 27751 1600 27767 1664
rect 27831 1600 27847 1664
rect 27911 1600 27927 1664
rect 27991 1600 27997 1664
rect 27681 1599 27997 1600
rect 38375 1664 38691 1665
rect 38375 1600 38381 1664
rect 38445 1600 38461 1664
rect 38525 1600 38541 1664
rect 38605 1600 38621 1664
rect 38685 1600 38691 1664
rect 38375 1599 38691 1600
rect 17493 1594 17559 1597
rect 19057 1594 19123 1597
rect 17493 1592 19123 1594
rect 17493 1536 17498 1592
rect 17554 1536 19062 1592
rect 19118 1536 19123 1592
rect 17493 1534 19123 1536
rect 17493 1531 17559 1534
rect 19057 1531 19123 1534
rect 23105 1594 23171 1597
rect 23933 1594 23999 1597
rect 23105 1592 23999 1594
rect 23105 1536 23110 1592
rect 23166 1536 23938 1592
rect 23994 1536 23999 1592
rect 23105 1534 23999 1536
rect 23105 1531 23171 1534
rect 23933 1531 23999 1534
rect 24669 1594 24735 1597
rect 26233 1594 26299 1597
rect 24669 1592 26299 1594
rect 24669 1536 24674 1592
rect 24730 1536 26238 1592
rect 26294 1536 26299 1592
rect 24669 1534 26299 1536
rect 24669 1531 24735 1534
rect 26233 1531 26299 1534
rect 8293 1458 8359 1461
rect 22921 1458 22987 1461
rect 8293 1456 22987 1458
rect 8293 1400 8298 1456
rect 8354 1400 22926 1456
rect 22982 1400 22987 1456
rect 8293 1398 22987 1400
rect 8293 1395 8359 1398
rect 22921 1395 22987 1398
rect 23841 1458 23907 1461
rect 30741 1458 30807 1461
rect 23841 1456 30807 1458
rect 23841 1400 23846 1456
rect 23902 1400 30746 1456
rect 30802 1400 30807 1456
rect 23841 1398 30807 1400
rect 23841 1395 23907 1398
rect 30741 1395 30807 1398
rect 15009 1322 15075 1325
rect 20805 1322 20871 1325
rect 15009 1320 20871 1322
rect 15009 1264 15014 1320
rect 15070 1264 20810 1320
rect 20866 1264 20871 1320
rect 15009 1262 20871 1264
rect 15009 1259 15075 1262
rect 20805 1259 20871 1262
rect 21398 1260 21404 1324
rect 21468 1322 21474 1324
rect 21725 1322 21791 1325
rect 24209 1322 24275 1325
rect 21468 1320 21791 1322
rect 21468 1264 21730 1320
rect 21786 1264 21791 1320
rect 21468 1262 21791 1264
rect 21468 1260 21474 1262
rect 21725 1259 21791 1262
rect 22050 1320 24275 1322
rect 22050 1264 24214 1320
rect 24270 1264 24275 1320
rect 22050 1262 24275 1264
rect 16849 1186 16915 1189
rect 22050 1186 22110 1262
rect 24209 1259 24275 1262
rect 26601 1322 26667 1325
rect 27797 1322 27863 1325
rect 26601 1320 27863 1322
rect 26601 1264 26606 1320
rect 26662 1264 27802 1320
rect 27858 1264 27863 1320
rect 26601 1262 27863 1264
rect 26601 1259 26667 1262
rect 27797 1259 27863 1262
rect 34462 1260 34468 1324
rect 34532 1322 34538 1324
rect 35065 1322 35131 1325
rect 34532 1320 35131 1322
rect 34532 1264 35070 1320
rect 35126 1264 35131 1320
rect 34532 1262 35131 1264
rect 34532 1260 34538 1262
rect 35065 1259 35131 1262
rect 16849 1184 22110 1186
rect 16849 1128 16854 1184
rect 16910 1128 22110 1184
rect 16849 1126 22110 1128
rect 23013 1186 23079 1189
rect 28717 1186 28783 1189
rect 23013 1184 28783 1186
rect 23013 1128 23018 1184
rect 23074 1128 28722 1184
rect 28778 1128 28783 1184
rect 23013 1126 28783 1128
rect 16849 1123 16915 1126
rect 23013 1123 23079 1126
rect 28717 1123 28783 1126
rect 11640 1120 11956 1121
rect 11640 1056 11646 1120
rect 11710 1056 11726 1120
rect 11790 1056 11806 1120
rect 11870 1056 11886 1120
rect 11950 1056 11956 1120
rect 11640 1055 11956 1056
rect 22334 1120 22650 1121
rect 22334 1056 22340 1120
rect 22404 1056 22420 1120
rect 22484 1056 22500 1120
rect 22564 1056 22580 1120
rect 22644 1056 22650 1120
rect 22334 1055 22650 1056
rect 33028 1120 33344 1121
rect 33028 1056 33034 1120
rect 33098 1056 33114 1120
rect 33178 1056 33194 1120
rect 33258 1056 33274 1120
rect 33338 1056 33344 1120
rect 33028 1055 33344 1056
rect 43722 1120 44038 1121
rect 43722 1056 43728 1120
rect 43792 1056 43808 1120
rect 43872 1056 43888 1120
rect 43952 1056 43968 1120
rect 44032 1056 44038 1120
rect 43722 1055 44038 1056
rect 17953 1050 18019 1053
rect 21817 1050 21883 1053
rect 17953 1048 21883 1050
rect 17953 992 17958 1048
rect 18014 992 21822 1048
rect 21878 992 21883 1048
rect 17953 990 21883 992
rect 17953 987 18019 990
rect 21817 987 21883 990
rect 11237 914 11303 917
rect 28349 914 28415 917
rect 11237 912 28415 914
rect 11237 856 11242 912
rect 11298 856 28354 912
rect 28410 856 28415 912
rect 11237 854 28415 856
rect 11237 851 11303 854
rect 28349 851 28415 854
rect 10961 778 11027 781
rect 31937 778 32003 781
rect 38561 778 38627 781
rect 10961 776 32003 778
rect 10961 720 10966 776
rect 11022 720 31942 776
rect 31998 720 32003 776
rect 10961 718 32003 720
rect 10961 715 11027 718
rect 31937 715 32003 718
rect 35206 776 38627 778
rect 35206 720 38566 776
rect 38622 720 38627 776
rect 35206 718 38627 720
rect 6177 642 6243 645
rect 16849 642 16915 645
rect 23749 642 23815 645
rect 6177 640 16915 642
rect 6177 584 6182 640
rect 6238 584 16854 640
rect 16910 584 16915 640
rect 6177 582 16915 584
rect 6177 579 6243 582
rect 16849 579 16915 582
rect 17174 640 23815 642
rect 17174 584 23754 640
rect 23810 584 23815 640
rect 17174 582 23815 584
rect 6545 370 6611 373
rect 17174 370 17234 582
rect 23749 579 23815 582
rect 25497 642 25563 645
rect 27889 642 27955 645
rect 25497 640 27955 642
rect 25497 584 25502 640
rect 25558 584 27894 640
rect 27950 584 27955 640
rect 25497 582 27955 584
rect 25497 579 25563 582
rect 27889 579 27955 582
rect 20989 506 21055 509
rect 21817 506 21883 509
rect 34605 506 34671 509
rect 20989 504 21650 506
rect 20989 448 20994 504
rect 21050 448 21650 504
rect 20989 446 21650 448
rect 20989 443 21055 446
rect 6545 368 17234 370
rect 6545 312 6550 368
rect 6606 312 17234 368
rect 6545 310 17234 312
rect 6545 307 6611 310
rect 16205 234 16271 237
rect 20069 234 20135 237
rect 16205 232 20135 234
rect 16205 176 16210 232
rect 16266 176 20074 232
rect 20130 176 20135 232
rect 16205 174 20135 176
rect 21590 234 21650 446
rect 21817 504 34671 506
rect 21817 448 21822 504
rect 21878 448 34610 504
rect 34666 448 34671 504
rect 21817 446 34671 448
rect 21817 443 21883 446
rect 34605 443 34671 446
rect 35206 234 35266 718
rect 38561 715 38627 718
rect 21590 174 35266 234
rect 16205 171 16271 174
rect 20069 171 20135 174
<< via3 >>
rect 11646 8732 11710 8736
rect 11646 8676 11650 8732
rect 11650 8676 11706 8732
rect 11706 8676 11710 8732
rect 11646 8672 11710 8676
rect 11726 8732 11790 8736
rect 11726 8676 11730 8732
rect 11730 8676 11786 8732
rect 11786 8676 11790 8732
rect 11726 8672 11790 8676
rect 11806 8732 11870 8736
rect 11806 8676 11810 8732
rect 11810 8676 11866 8732
rect 11866 8676 11870 8732
rect 11806 8672 11870 8676
rect 11886 8732 11950 8736
rect 11886 8676 11890 8732
rect 11890 8676 11946 8732
rect 11946 8676 11950 8732
rect 11886 8672 11950 8676
rect 22340 8732 22404 8736
rect 22340 8676 22344 8732
rect 22344 8676 22400 8732
rect 22400 8676 22404 8732
rect 22340 8672 22404 8676
rect 22420 8732 22484 8736
rect 22420 8676 22424 8732
rect 22424 8676 22480 8732
rect 22480 8676 22484 8732
rect 22420 8672 22484 8676
rect 22500 8732 22564 8736
rect 22500 8676 22504 8732
rect 22504 8676 22560 8732
rect 22560 8676 22564 8732
rect 22500 8672 22564 8676
rect 22580 8732 22644 8736
rect 22580 8676 22584 8732
rect 22584 8676 22640 8732
rect 22640 8676 22644 8732
rect 22580 8672 22644 8676
rect 33034 8732 33098 8736
rect 33034 8676 33038 8732
rect 33038 8676 33094 8732
rect 33094 8676 33098 8732
rect 33034 8672 33098 8676
rect 33114 8732 33178 8736
rect 33114 8676 33118 8732
rect 33118 8676 33174 8732
rect 33174 8676 33178 8732
rect 33114 8672 33178 8676
rect 33194 8732 33258 8736
rect 33194 8676 33198 8732
rect 33198 8676 33254 8732
rect 33254 8676 33258 8732
rect 33194 8672 33258 8676
rect 33274 8732 33338 8736
rect 33274 8676 33278 8732
rect 33278 8676 33334 8732
rect 33334 8676 33338 8732
rect 33274 8672 33338 8676
rect 43728 8732 43792 8736
rect 43728 8676 43732 8732
rect 43732 8676 43788 8732
rect 43788 8676 43792 8732
rect 43728 8672 43792 8676
rect 43808 8732 43872 8736
rect 43808 8676 43812 8732
rect 43812 8676 43868 8732
rect 43868 8676 43872 8732
rect 43808 8672 43872 8676
rect 43888 8732 43952 8736
rect 43888 8676 43892 8732
rect 43892 8676 43948 8732
rect 43948 8676 43952 8732
rect 43888 8672 43952 8676
rect 43968 8732 44032 8736
rect 43968 8676 43972 8732
rect 43972 8676 44028 8732
rect 44028 8676 44032 8732
rect 43968 8672 44032 8676
rect 24900 8468 24964 8532
rect 25084 8332 25148 8396
rect 6299 8188 6363 8192
rect 6299 8132 6303 8188
rect 6303 8132 6359 8188
rect 6359 8132 6363 8188
rect 6299 8128 6363 8132
rect 6379 8188 6443 8192
rect 6379 8132 6383 8188
rect 6383 8132 6439 8188
rect 6439 8132 6443 8188
rect 6379 8128 6443 8132
rect 6459 8188 6523 8192
rect 6459 8132 6463 8188
rect 6463 8132 6519 8188
rect 6519 8132 6523 8188
rect 6459 8128 6523 8132
rect 6539 8188 6603 8192
rect 6539 8132 6543 8188
rect 6543 8132 6599 8188
rect 6599 8132 6603 8188
rect 6539 8128 6603 8132
rect 16993 8188 17057 8192
rect 16993 8132 16997 8188
rect 16997 8132 17053 8188
rect 17053 8132 17057 8188
rect 16993 8128 17057 8132
rect 17073 8188 17137 8192
rect 17073 8132 17077 8188
rect 17077 8132 17133 8188
rect 17133 8132 17137 8188
rect 17073 8128 17137 8132
rect 17153 8188 17217 8192
rect 17153 8132 17157 8188
rect 17157 8132 17213 8188
rect 17213 8132 17217 8188
rect 17153 8128 17217 8132
rect 17233 8188 17297 8192
rect 17233 8132 17237 8188
rect 17237 8132 17293 8188
rect 17293 8132 17297 8188
rect 17233 8128 17297 8132
rect 27687 8188 27751 8192
rect 27687 8132 27691 8188
rect 27691 8132 27747 8188
rect 27747 8132 27751 8188
rect 27687 8128 27751 8132
rect 27767 8188 27831 8192
rect 27767 8132 27771 8188
rect 27771 8132 27827 8188
rect 27827 8132 27831 8188
rect 27767 8128 27831 8132
rect 27847 8188 27911 8192
rect 27847 8132 27851 8188
rect 27851 8132 27907 8188
rect 27907 8132 27911 8188
rect 27847 8128 27911 8132
rect 27927 8188 27991 8192
rect 27927 8132 27931 8188
rect 27931 8132 27987 8188
rect 27987 8132 27991 8188
rect 27927 8128 27991 8132
rect 38381 8188 38445 8192
rect 38381 8132 38385 8188
rect 38385 8132 38441 8188
rect 38441 8132 38445 8188
rect 38381 8128 38445 8132
rect 38461 8188 38525 8192
rect 38461 8132 38465 8188
rect 38465 8132 38521 8188
rect 38521 8132 38525 8188
rect 38461 8128 38525 8132
rect 38541 8188 38605 8192
rect 38541 8132 38545 8188
rect 38545 8132 38601 8188
rect 38601 8132 38605 8188
rect 38541 8128 38605 8132
rect 38621 8188 38685 8192
rect 38621 8132 38625 8188
rect 38625 8132 38681 8188
rect 38681 8132 38685 8188
rect 38621 8128 38685 8132
rect 11646 7644 11710 7648
rect 11646 7588 11650 7644
rect 11650 7588 11706 7644
rect 11706 7588 11710 7644
rect 11646 7584 11710 7588
rect 11726 7644 11790 7648
rect 11726 7588 11730 7644
rect 11730 7588 11786 7644
rect 11786 7588 11790 7644
rect 11726 7584 11790 7588
rect 11806 7644 11870 7648
rect 11806 7588 11810 7644
rect 11810 7588 11866 7644
rect 11866 7588 11870 7644
rect 11806 7584 11870 7588
rect 11886 7644 11950 7648
rect 11886 7588 11890 7644
rect 11890 7588 11946 7644
rect 11946 7588 11950 7644
rect 11886 7584 11950 7588
rect 22340 7644 22404 7648
rect 22340 7588 22344 7644
rect 22344 7588 22400 7644
rect 22400 7588 22404 7644
rect 22340 7584 22404 7588
rect 22420 7644 22484 7648
rect 22420 7588 22424 7644
rect 22424 7588 22480 7644
rect 22480 7588 22484 7644
rect 22420 7584 22484 7588
rect 22500 7644 22564 7648
rect 22500 7588 22504 7644
rect 22504 7588 22560 7644
rect 22560 7588 22564 7644
rect 22500 7584 22564 7588
rect 22580 7644 22644 7648
rect 22580 7588 22584 7644
rect 22584 7588 22640 7644
rect 22640 7588 22644 7644
rect 22580 7584 22644 7588
rect 33034 7644 33098 7648
rect 33034 7588 33038 7644
rect 33038 7588 33094 7644
rect 33094 7588 33098 7644
rect 33034 7584 33098 7588
rect 33114 7644 33178 7648
rect 33114 7588 33118 7644
rect 33118 7588 33174 7644
rect 33174 7588 33178 7644
rect 33114 7584 33178 7588
rect 33194 7644 33258 7648
rect 33194 7588 33198 7644
rect 33198 7588 33254 7644
rect 33254 7588 33258 7644
rect 33194 7584 33258 7588
rect 33274 7644 33338 7648
rect 33274 7588 33278 7644
rect 33278 7588 33334 7644
rect 33334 7588 33338 7644
rect 33274 7584 33338 7588
rect 43728 7644 43792 7648
rect 43728 7588 43732 7644
rect 43732 7588 43788 7644
rect 43788 7588 43792 7644
rect 43728 7584 43792 7588
rect 43808 7644 43872 7648
rect 43808 7588 43812 7644
rect 43812 7588 43868 7644
rect 43868 7588 43872 7644
rect 43808 7584 43872 7588
rect 43888 7644 43952 7648
rect 43888 7588 43892 7644
rect 43892 7588 43948 7644
rect 43948 7588 43952 7644
rect 43888 7584 43952 7588
rect 43968 7644 44032 7648
rect 43968 7588 43972 7644
rect 43972 7588 44028 7644
rect 44028 7588 44032 7644
rect 43968 7584 44032 7588
rect 6299 7100 6363 7104
rect 6299 7044 6303 7100
rect 6303 7044 6359 7100
rect 6359 7044 6363 7100
rect 6299 7040 6363 7044
rect 6379 7100 6443 7104
rect 6379 7044 6383 7100
rect 6383 7044 6439 7100
rect 6439 7044 6443 7100
rect 6379 7040 6443 7044
rect 6459 7100 6523 7104
rect 6459 7044 6463 7100
rect 6463 7044 6519 7100
rect 6519 7044 6523 7100
rect 6459 7040 6523 7044
rect 6539 7100 6603 7104
rect 6539 7044 6543 7100
rect 6543 7044 6599 7100
rect 6599 7044 6603 7100
rect 6539 7040 6603 7044
rect 16993 7100 17057 7104
rect 16993 7044 16997 7100
rect 16997 7044 17053 7100
rect 17053 7044 17057 7100
rect 16993 7040 17057 7044
rect 17073 7100 17137 7104
rect 17073 7044 17077 7100
rect 17077 7044 17133 7100
rect 17133 7044 17137 7100
rect 17073 7040 17137 7044
rect 17153 7100 17217 7104
rect 17153 7044 17157 7100
rect 17157 7044 17213 7100
rect 17213 7044 17217 7100
rect 17153 7040 17217 7044
rect 17233 7100 17297 7104
rect 17233 7044 17237 7100
rect 17237 7044 17293 7100
rect 17293 7044 17297 7100
rect 17233 7040 17297 7044
rect 27687 7100 27751 7104
rect 27687 7044 27691 7100
rect 27691 7044 27747 7100
rect 27747 7044 27751 7100
rect 27687 7040 27751 7044
rect 27767 7100 27831 7104
rect 27767 7044 27771 7100
rect 27771 7044 27827 7100
rect 27827 7044 27831 7100
rect 27767 7040 27831 7044
rect 27847 7100 27911 7104
rect 27847 7044 27851 7100
rect 27851 7044 27907 7100
rect 27907 7044 27911 7100
rect 27847 7040 27911 7044
rect 27927 7100 27991 7104
rect 27927 7044 27931 7100
rect 27931 7044 27987 7100
rect 27987 7044 27991 7100
rect 27927 7040 27991 7044
rect 38381 7100 38445 7104
rect 38381 7044 38385 7100
rect 38385 7044 38441 7100
rect 38441 7044 38445 7100
rect 38381 7040 38445 7044
rect 38461 7100 38525 7104
rect 38461 7044 38465 7100
rect 38465 7044 38521 7100
rect 38521 7044 38525 7100
rect 38461 7040 38525 7044
rect 38541 7100 38605 7104
rect 38541 7044 38545 7100
rect 38545 7044 38601 7100
rect 38601 7044 38605 7100
rect 38541 7040 38605 7044
rect 38621 7100 38685 7104
rect 38621 7044 38625 7100
rect 38625 7044 38681 7100
rect 38681 7044 38685 7100
rect 38621 7040 38685 7044
rect 11646 6556 11710 6560
rect 11646 6500 11650 6556
rect 11650 6500 11706 6556
rect 11706 6500 11710 6556
rect 11646 6496 11710 6500
rect 11726 6556 11790 6560
rect 11726 6500 11730 6556
rect 11730 6500 11786 6556
rect 11786 6500 11790 6556
rect 11726 6496 11790 6500
rect 11806 6556 11870 6560
rect 11806 6500 11810 6556
rect 11810 6500 11866 6556
rect 11866 6500 11870 6556
rect 11806 6496 11870 6500
rect 11886 6556 11950 6560
rect 11886 6500 11890 6556
rect 11890 6500 11946 6556
rect 11946 6500 11950 6556
rect 11886 6496 11950 6500
rect 22340 6556 22404 6560
rect 22340 6500 22344 6556
rect 22344 6500 22400 6556
rect 22400 6500 22404 6556
rect 22340 6496 22404 6500
rect 22420 6556 22484 6560
rect 22420 6500 22424 6556
rect 22424 6500 22480 6556
rect 22480 6500 22484 6556
rect 22420 6496 22484 6500
rect 22500 6556 22564 6560
rect 22500 6500 22504 6556
rect 22504 6500 22560 6556
rect 22560 6500 22564 6556
rect 22500 6496 22564 6500
rect 22580 6556 22644 6560
rect 22580 6500 22584 6556
rect 22584 6500 22640 6556
rect 22640 6500 22644 6556
rect 22580 6496 22644 6500
rect 33034 6556 33098 6560
rect 33034 6500 33038 6556
rect 33038 6500 33094 6556
rect 33094 6500 33098 6556
rect 33034 6496 33098 6500
rect 33114 6556 33178 6560
rect 33114 6500 33118 6556
rect 33118 6500 33174 6556
rect 33174 6500 33178 6556
rect 33114 6496 33178 6500
rect 33194 6556 33258 6560
rect 33194 6500 33198 6556
rect 33198 6500 33254 6556
rect 33254 6500 33258 6556
rect 33194 6496 33258 6500
rect 33274 6556 33338 6560
rect 33274 6500 33278 6556
rect 33278 6500 33334 6556
rect 33334 6500 33338 6556
rect 33274 6496 33338 6500
rect 43728 6556 43792 6560
rect 43728 6500 43732 6556
rect 43732 6500 43788 6556
rect 43788 6500 43792 6556
rect 43728 6496 43792 6500
rect 43808 6556 43872 6560
rect 43808 6500 43812 6556
rect 43812 6500 43868 6556
rect 43868 6500 43872 6556
rect 43808 6496 43872 6500
rect 43888 6556 43952 6560
rect 43888 6500 43892 6556
rect 43892 6500 43948 6556
rect 43948 6500 43952 6556
rect 43888 6496 43952 6500
rect 43968 6556 44032 6560
rect 43968 6500 43972 6556
rect 43972 6500 44028 6556
rect 44028 6500 44032 6556
rect 43968 6496 44032 6500
rect 6299 6012 6363 6016
rect 6299 5956 6303 6012
rect 6303 5956 6359 6012
rect 6359 5956 6363 6012
rect 6299 5952 6363 5956
rect 6379 6012 6443 6016
rect 6379 5956 6383 6012
rect 6383 5956 6439 6012
rect 6439 5956 6443 6012
rect 6379 5952 6443 5956
rect 6459 6012 6523 6016
rect 6459 5956 6463 6012
rect 6463 5956 6519 6012
rect 6519 5956 6523 6012
rect 6459 5952 6523 5956
rect 6539 6012 6603 6016
rect 6539 5956 6543 6012
rect 6543 5956 6599 6012
rect 6599 5956 6603 6012
rect 6539 5952 6603 5956
rect 16993 6012 17057 6016
rect 16993 5956 16997 6012
rect 16997 5956 17053 6012
rect 17053 5956 17057 6012
rect 16993 5952 17057 5956
rect 17073 6012 17137 6016
rect 17073 5956 17077 6012
rect 17077 5956 17133 6012
rect 17133 5956 17137 6012
rect 17073 5952 17137 5956
rect 17153 6012 17217 6016
rect 17153 5956 17157 6012
rect 17157 5956 17213 6012
rect 17213 5956 17217 6012
rect 17153 5952 17217 5956
rect 17233 6012 17297 6016
rect 17233 5956 17237 6012
rect 17237 5956 17293 6012
rect 17293 5956 17297 6012
rect 17233 5952 17297 5956
rect 27687 6012 27751 6016
rect 27687 5956 27691 6012
rect 27691 5956 27747 6012
rect 27747 5956 27751 6012
rect 27687 5952 27751 5956
rect 27767 6012 27831 6016
rect 27767 5956 27771 6012
rect 27771 5956 27827 6012
rect 27827 5956 27831 6012
rect 27767 5952 27831 5956
rect 27847 6012 27911 6016
rect 27847 5956 27851 6012
rect 27851 5956 27907 6012
rect 27907 5956 27911 6012
rect 27847 5952 27911 5956
rect 27927 6012 27991 6016
rect 27927 5956 27931 6012
rect 27931 5956 27987 6012
rect 27987 5956 27991 6012
rect 27927 5952 27991 5956
rect 38381 6012 38445 6016
rect 38381 5956 38385 6012
rect 38385 5956 38441 6012
rect 38441 5956 38445 6012
rect 38381 5952 38445 5956
rect 38461 6012 38525 6016
rect 38461 5956 38465 6012
rect 38465 5956 38521 6012
rect 38521 5956 38525 6012
rect 38461 5952 38525 5956
rect 38541 6012 38605 6016
rect 38541 5956 38545 6012
rect 38545 5956 38601 6012
rect 38601 5956 38605 6012
rect 38541 5952 38605 5956
rect 38621 6012 38685 6016
rect 38621 5956 38625 6012
rect 38625 5956 38681 6012
rect 38681 5956 38685 6012
rect 38621 5952 38685 5956
rect 11646 5468 11710 5472
rect 11646 5412 11650 5468
rect 11650 5412 11706 5468
rect 11706 5412 11710 5468
rect 11646 5408 11710 5412
rect 11726 5468 11790 5472
rect 11726 5412 11730 5468
rect 11730 5412 11786 5468
rect 11786 5412 11790 5468
rect 11726 5408 11790 5412
rect 11806 5468 11870 5472
rect 11806 5412 11810 5468
rect 11810 5412 11866 5468
rect 11866 5412 11870 5468
rect 11806 5408 11870 5412
rect 11886 5468 11950 5472
rect 11886 5412 11890 5468
rect 11890 5412 11946 5468
rect 11946 5412 11950 5468
rect 11886 5408 11950 5412
rect 22340 5468 22404 5472
rect 22340 5412 22344 5468
rect 22344 5412 22400 5468
rect 22400 5412 22404 5468
rect 22340 5408 22404 5412
rect 22420 5468 22484 5472
rect 22420 5412 22424 5468
rect 22424 5412 22480 5468
rect 22480 5412 22484 5468
rect 22420 5408 22484 5412
rect 22500 5468 22564 5472
rect 22500 5412 22504 5468
rect 22504 5412 22560 5468
rect 22560 5412 22564 5468
rect 22500 5408 22564 5412
rect 22580 5468 22644 5472
rect 22580 5412 22584 5468
rect 22584 5412 22640 5468
rect 22640 5412 22644 5468
rect 22580 5408 22644 5412
rect 33034 5468 33098 5472
rect 33034 5412 33038 5468
rect 33038 5412 33094 5468
rect 33094 5412 33098 5468
rect 33034 5408 33098 5412
rect 33114 5468 33178 5472
rect 33114 5412 33118 5468
rect 33118 5412 33174 5468
rect 33174 5412 33178 5468
rect 33114 5408 33178 5412
rect 33194 5468 33258 5472
rect 33194 5412 33198 5468
rect 33198 5412 33254 5468
rect 33254 5412 33258 5468
rect 33194 5408 33258 5412
rect 33274 5468 33338 5472
rect 33274 5412 33278 5468
rect 33278 5412 33334 5468
rect 33334 5412 33338 5468
rect 33274 5408 33338 5412
rect 43728 5468 43792 5472
rect 43728 5412 43732 5468
rect 43732 5412 43788 5468
rect 43788 5412 43792 5468
rect 43728 5408 43792 5412
rect 43808 5468 43872 5472
rect 43808 5412 43812 5468
rect 43812 5412 43868 5468
rect 43868 5412 43872 5468
rect 43808 5408 43872 5412
rect 43888 5468 43952 5472
rect 43888 5412 43892 5468
rect 43892 5412 43948 5468
rect 43948 5412 43952 5468
rect 43888 5408 43952 5412
rect 43968 5468 44032 5472
rect 43968 5412 43972 5468
rect 43972 5412 44028 5468
rect 44028 5412 44032 5468
rect 43968 5408 44032 5412
rect 6299 4924 6363 4928
rect 6299 4868 6303 4924
rect 6303 4868 6359 4924
rect 6359 4868 6363 4924
rect 6299 4864 6363 4868
rect 6379 4924 6443 4928
rect 6379 4868 6383 4924
rect 6383 4868 6439 4924
rect 6439 4868 6443 4924
rect 6379 4864 6443 4868
rect 6459 4924 6523 4928
rect 6459 4868 6463 4924
rect 6463 4868 6519 4924
rect 6519 4868 6523 4924
rect 6459 4864 6523 4868
rect 6539 4924 6603 4928
rect 6539 4868 6543 4924
rect 6543 4868 6599 4924
rect 6599 4868 6603 4924
rect 6539 4864 6603 4868
rect 16993 4924 17057 4928
rect 16993 4868 16997 4924
rect 16997 4868 17053 4924
rect 17053 4868 17057 4924
rect 16993 4864 17057 4868
rect 17073 4924 17137 4928
rect 17073 4868 17077 4924
rect 17077 4868 17133 4924
rect 17133 4868 17137 4924
rect 17073 4864 17137 4868
rect 17153 4924 17217 4928
rect 17153 4868 17157 4924
rect 17157 4868 17213 4924
rect 17213 4868 17217 4924
rect 17153 4864 17217 4868
rect 17233 4924 17297 4928
rect 17233 4868 17237 4924
rect 17237 4868 17293 4924
rect 17293 4868 17297 4924
rect 17233 4864 17297 4868
rect 27687 4924 27751 4928
rect 27687 4868 27691 4924
rect 27691 4868 27747 4924
rect 27747 4868 27751 4924
rect 27687 4864 27751 4868
rect 27767 4924 27831 4928
rect 27767 4868 27771 4924
rect 27771 4868 27827 4924
rect 27827 4868 27831 4924
rect 27767 4864 27831 4868
rect 27847 4924 27911 4928
rect 27847 4868 27851 4924
rect 27851 4868 27907 4924
rect 27907 4868 27911 4924
rect 27847 4864 27911 4868
rect 27927 4924 27991 4928
rect 27927 4868 27931 4924
rect 27931 4868 27987 4924
rect 27987 4868 27991 4924
rect 27927 4864 27991 4868
rect 38381 4924 38445 4928
rect 38381 4868 38385 4924
rect 38385 4868 38441 4924
rect 38441 4868 38445 4924
rect 38381 4864 38445 4868
rect 38461 4924 38525 4928
rect 38461 4868 38465 4924
rect 38465 4868 38521 4924
rect 38521 4868 38525 4924
rect 38461 4864 38525 4868
rect 38541 4924 38605 4928
rect 38541 4868 38545 4924
rect 38545 4868 38601 4924
rect 38601 4868 38605 4924
rect 38541 4864 38605 4868
rect 38621 4924 38685 4928
rect 38621 4868 38625 4924
rect 38625 4868 38681 4924
rect 38681 4868 38685 4924
rect 38621 4864 38685 4868
rect 11646 4380 11710 4384
rect 11646 4324 11650 4380
rect 11650 4324 11706 4380
rect 11706 4324 11710 4380
rect 11646 4320 11710 4324
rect 11726 4380 11790 4384
rect 11726 4324 11730 4380
rect 11730 4324 11786 4380
rect 11786 4324 11790 4380
rect 11726 4320 11790 4324
rect 11806 4380 11870 4384
rect 11806 4324 11810 4380
rect 11810 4324 11866 4380
rect 11866 4324 11870 4380
rect 11806 4320 11870 4324
rect 11886 4380 11950 4384
rect 11886 4324 11890 4380
rect 11890 4324 11946 4380
rect 11946 4324 11950 4380
rect 11886 4320 11950 4324
rect 22340 4380 22404 4384
rect 22340 4324 22344 4380
rect 22344 4324 22400 4380
rect 22400 4324 22404 4380
rect 22340 4320 22404 4324
rect 22420 4380 22484 4384
rect 22420 4324 22424 4380
rect 22424 4324 22480 4380
rect 22480 4324 22484 4380
rect 22420 4320 22484 4324
rect 22500 4380 22564 4384
rect 22500 4324 22504 4380
rect 22504 4324 22560 4380
rect 22560 4324 22564 4380
rect 22500 4320 22564 4324
rect 22580 4380 22644 4384
rect 22580 4324 22584 4380
rect 22584 4324 22640 4380
rect 22640 4324 22644 4380
rect 22580 4320 22644 4324
rect 33034 4380 33098 4384
rect 33034 4324 33038 4380
rect 33038 4324 33094 4380
rect 33094 4324 33098 4380
rect 33034 4320 33098 4324
rect 33114 4380 33178 4384
rect 33114 4324 33118 4380
rect 33118 4324 33174 4380
rect 33174 4324 33178 4380
rect 33114 4320 33178 4324
rect 33194 4380 33258 4384
rect 33194 4324 33198 4380
rect 33198 4324 33254 4380
rect 33254 4324 33258 4380
rect 33194 4320 33258 4324
rect 33274 4380 33338 4384
rect 33274 4324 33278 4380
rect 33278 4324 33334 4380
rect 33334 4324 33338 4380
rect 33274 4320 33338 4324
rect 43728 4380 43792 4384
rect 43728 4324 43732 4380
rect 43732 4324 43788 4380
rect 43788 4324 43792 4380
rect 43728 4320 43792 4324
rect 43808 4380 43872 4384
rect 43808 4324 43812 4380
rect 43812 4324 43868 4380
rect 43868 4324 43872 4380
rect 43808 4320 43872 4324
rect 43888 4380 43952 4384
rect 43888 4324 43892 4380
rect 43892 4324 43948 4380
rect 43948 4324 43952 4380
rect 43888 4320 43952 4324
rect 43968 4380 44032 4384
rect 43968 4324 43972 4380
rect 43972 4324 44028 4380
rect 44028 4324 44032 4380
rect 43968 4320 44032 4324
rect 6299 3836 6363 3840
rect 6299 3780 6303 3836
rect 6303 3780 6359 3836
rect 6359 3780 6363 3836
rect 6299 3776 6363 3780
rect 6379 3836 6443 3840
rect 6379 3780 6383 3836
rect 6383 3780 6439 3836
rect 6439 3780 6443 3836
rect 6379 3776 6443 3780
rect 6459 3836 6523 3840
rect 6459 3780 6463 3836
rect 6463 3780 6519 3836
rect 6519 3780 6523 3836
rect 6459 3776 6523 3780
rect 6539 3836 6603 3840
rect 6539 3780 6543 3836
rect 6543 3780 6599 3836
rect 6599 3780 6603 3836
rect 6539 3776 6603 3780
rect 16993 3836 17057 3840
rect 16993 3780 16997 3836
rect 16997 3780 17053 3836
rect 17053 3780 17057 3836
rect 16993 3776 17057 3780
rect 17073 3836 17137 3840
rect 17073 3780 17077 3836
rect 17077 3780 17133 3836
rect 17133 3780 17137 3836
rect 17073 3776 17137 3780
rect 17153 3836 17217 3840
rect 17153 3780 17157 3836
rect 17157 3780 17213 3836
rect 17213 3780 17217 3836
rect 17153 3776 17217 3780
rect 17233 3836 17297 3840
rect 17233 3780 17237 3836
rect 17237 3780 17293 3836
rect 17293 3780 17297 3836
rect 17233 3776 17297 3780
rect 27687 3836 27751 3840
rect 27687 3780 27691 3836
rect 27691 3780 27747 3836
rect 27747 3780 27751 3836
rect 27687 3776 27751 3780
rect 27767 3836 27831 3840
rect 27767 3780 27771 3836
rect 27771 3780 27827 3836
rect 27827 3780 27831 3836
rect 27767 3776 27831 3780
rect 27847 3836 27911 3840
rect 27847 3780 27851 3836
rect 27851 3780 27907 3836
rect 27907 3780 27911 3836
rect 27847 3776 27911 3780
rect 27927 3836 27991 3840
rect 27927 3780 27931 3836
rect 27931 3780 27987 3836
rect 27987 3780 27991 3836
rect 27927 3776 27991 3780
rect 38381 3836 38445 3840
rect 38381 3780 38385 3836
rect 38385 3780 38441 3836
rect 38441 3780 38445 3836
rect 38381 3776 38445 3780
rect 38461 3836 38525 3840
rect 38461 3780 38465 3836
rect 38465 3780 38521 3836
rect 38521 3780 38525 3836
rect 38461 3776 38525 3780
rect 38541 3836 38605 3840
rect 38541 3780 38545 3836
rect 38545 3780 38601 3836
rect 38601 3780 38605 3836
rect 38541 3776 38605 3780
rect 38621 3836 38685 3840
rect 38621 3780 38625 3836
rect 38625 3780 38681 3836
rect 38681 3780 38685 3836
rect 38621 3776 38685 3780
rect 34468 3572 34532 3636
rect 11646 3292 11710 3296
rect 11646 3236 11650 3292
rect 11650 3236 11706 3292
rect 11706 3236 11710 3292
rect 11646 3232 11710 3236
rect 11726 3292 11790 3296
rect 11726 3236 11730 3292
rect 11730 3236 11786 3292
rect 11786 3236 11790 3292
rect 11726 3232 11790 3236
rect 11806 3292 11870 3296
rect 11806 3236 11810 3292
rect 11810 3236 11866 3292
rect 11866 3236 11870 3292
rect 11806 3232 11870 3236
rect 11886 3292 11950 3296
rect 11886 3236 11890 3292
rect 11890 3236 11946 3292
rect 11946 3236 11950 3292
rect 11886 3232 11950 3236
rect 22340 3292 22404 3296
rect 22340 3236 22344 3292
rect 22344 3236 22400 3292
rect 22400 3236 22404 3292
rect 22340 3232 22404 3236
rect 22420 3292 22484 3296
rect 22420 3236 22424 3292
rect 22424 3236 22480 3292
rect 22480 3236 22484 3292
rect 22420 3232 22484 3236
rect 22500 3292 22564 3296
rect 22500 3236 22504 3292
rect 22504 3236 22560 3292
rect 22560 3236 22564 3292
rect 22500 3232 22564 3236
rect 22580 3292 22644 3296
rect 22580 3236 22584 3292
rect 22584 3236 22640 3292
rect 22640 3236 22644 3292
rect 22580 3232 22644 3236
rect 33034 3292 33098 3296
rect 33034 3236 33038 3292
rect 33038 3236 33094 3292
rect 33094 3236 33098 3292
rect 33034 3232 33098 3236
rect 33114 3292 33178 3296
rect 33114 3236 33118 3292
rect 33118 3236 33174 3292
rect 33174 3236 33178 3292
rect 33114 3232 33178 3236
rect 33194 3292 33258 3296
rect 33194 3236 33198 3292
rect 33198 3236 33254 3292
rect 33254 3236 33258 3292
rect 33194 3232 33258 3236
rect 33274 3292 33338 3296
rect 33274 3236 33278 3292
rect 33278 3236 33334 3292
rect 33334 3236 33338 3292
rect 33274 3232 33338 3236
rect 43728 3292 43792 3296
rect 43728 3236 43732 3292
rect 43732 3236 43788 3292
rect 43788 3236 43792 3292
rect 43728 3232 43792 3236
rect 43808 3292 43872 3296
rect 43808 3236 43812 3292
rect 43812 3236 43868 3292
rect 43868 3236 43872 3292
rect 43808 3232 43872 3236
rect 43888 3292 43952 3296
rect 43888 3236 43892 3292
rect 43892 3236 43948 3292
rect 43948 3236 43952 3292
rect 43888 3232 43952 3236
rect 43968 3292 44032 3296
rect 43968 3236 43972 3292
rect 43972 3236 44028 3292
rect 44028 3236 44032 3292
rect 43968 3232 44032 3236
rect 21404 2756 21468 2820
rect 6299 2748 6363 2752
rect 6299 2692 6303 2748
rect 6303 2692 6359 2748
rect 6359 2692 6363 2748
rect 6299 2688 6363 2692
rect 6379 2748 6443 2752
rect 6379 2692 6383 2748
rect 6383 2692 6439 2748
rect 6439 2692 6443 2748
rect 6379 2688 6443 2692
rect 6459 2748 6523 2752
rect 6459 2692 6463 2748
rect 6463 2692 6519 2748
rect 6519 2692 6523 2748
rect 6459 2688 6523 2692
rect 6539 2748 6603 2752
rect 6539 2692 6543 2748
rect 6543 2692 6599 2748
rect 6599 2692 6603 2748
rect 6539 2688 6603 2692
rect 16993 2748 17057 2752
rect 16993 2692 16997 2748
rect 16997 2692 17053 2748
rect 17053 2692 17057 2748
rect 16993 2688 17057 2692
rect 17073 2748 17137 2752
rect 17073 2692 17077 2748
rect 17077 2692 17133 2748
rect 17133 2692 17137 2748
rect 17073 2688 17137 2692
rect 17153 2748 17217 2752
rect 17153 2692 17157 2748
rect 17157 2692 17213 2748
rect 17213 2692 17217 2748
rect 17153 2688 17217 2692
rect 17233 2748 17297 2752
rect 17233 2692 17237 2748
rect 17237 2692 17293 2748
rect 17293 2692 17297 2748
rect 17233 2688 17297 2692
rect 27687 2748 27751 2752
rect 27687 2692 27691 2748
rect 27691 2692 27747 2748
rect 27747 2692 27751 2748
rect 27687 2688 27751 2692
rect 27767 2748 27831 2752
rect 27767 2692 27771 2748
rect 27771 2692 27827 2748
rect 27827 2692 27831 2748
rect 27767 2688 27831 2692
rect 27847 2748 27911 2752
rect 27847 2692 27851 2748
rect 27851 2692 27907 2748
rect 27907 2692 27911 2748
rect 27847 2688 27911 2692
rect 27927 2748 27991 2752
rect 27927 2692 27931 2748
rect 27931 2692 27987 2748
rect 27987 2692 27991 2748
rect 27927 2688 27991 2692
rect 38381 2748 38445 2752
rect 38381 2692 38385 2748
rect 38385 2692 38441 2748
rect 38441 2692 38445 2748
rect 38381 2688 38445 2692
rect 38461 2748 38525 2752
rect 38461 2692 38465 2748
rect 38465 2692 38521 2748
rect 38521 2692 38525 2748
rect 38461 2688 38525 2692
rect 38541 2748 38605 2752
rect 38541 2692 38545 2748
rect 38545 2692 38601 2748
rect 38601 2692 38605 2748
rect 38541 2688 38605 2692
rect 38621 2748 38685 2752
rect 38621 2692 38625 2748
rect 38625 2692 38681 2748
rect 38681 2692 38685 2748
rect 38621 2688 38685 2692
rect 24900 2680 24964 2684
rect 24900 2624 24950 2680
rect 24950 2624 24964 2680
rect 24900 2620 24964 2624
rect 11646 2204 11710 2208
rect 11646 2148 11650 2204
rect 11650 2148 11706 2204
rect 11706 2148 11710 2204
rect 11646 2144 11710 2148
rect 11726 2204 11790 2208
rect 11726 2148 11730 2204
rect 11730 2148 11786 2204
rect 11786 2148 11790 2204
rect 11726 2144 11790 2148
rect 11806 2204 11870 2208
rect 11806 2148 11810 2204
rect 11810 2148 11866 2204
rect 11866 2148 11870 2204
rect 11806 2144 11870 2148
rect 11886 2204 11950 2208
rect 11886 2148 11890 2204
rect 11890 2148 11946 2204
rect 11946 2148 11950 2204
rect 11886 2144 11950 2148
rect 25084 2212 25148 2276
rect 22340 2204 22404 2208
rect 22340 2148 22344 2204
rect 22344 2148 22400 2204
rect 22400 2148 22404 2204
rect 22340 2144 22404 2148
rect 22420 2204 22484 2208
rect 22420 2148 22424 2204
rect 22424 2148 22480 2204
rect 22480 2148 22484 2204
rect 22420 2144 22484 2148
rect 22500 2204 22564 2208
rect 22500 2148 22504 2204
rect 22504 2148 22560 2204
rect 22560 2148 22564 2204
rect 22500 2144 22564 2148
rect 22580 2204 22644 2208
rect 22580 2148 22584 2204
rect 22584 2148 22640 2204
rect 22640 2148 22644 2204
rect 22580 2144 22644 2148
rect 33034 2204 33098 2208
rect 33034 2148 33038 2204
rect 33038 2148 33094 2204
rect 33094 2148 33098 2204
rect 33034 2144 33098 2148
rect 33114 2204 33178 2208
rect 33114 2148 33118 2204
rect 33118 2148 33174 2204
rect 33174 2148 33178 2204
rect 33114 2144 33178 2148
rect 33194 2204 33258 2208
rect 33194 2148 33198 2204
rect 33198 2148 33254 2204
rect 33254 2148 33258 2204
rect 33194 2144 33258 2148
rect 33274 2204 33338 2208
rect 33274 2148 33278 2204
rect 33278 2148 33334 2204
rect 33334 2148 33338 2204
rect 33274 2144 33338 2148
rect 43728 2204 43792 2208
rect 43728 2148 43732 2204
rect 43732 2148 43788 2204
rect 43788 2148 43792 2204
rect 43728 2144 43792 2148
rect 43808 2204 43872 2208
rect 43808 2148 43812 2204
rect 43812 2148 43868 2204
rect 43868 2148 43872 2204
rect 43808 2144 43872 2148
rect 43888 2204 43952 2208
rect 43888 2148 43892 2204
rect 43892 2148 43948 2204
rect 43948 2148 43952 2204
rect 43888 2144 43952 2148
rect 43968 2204 44032 2208
rect 43968 2148 43972 2204
rect 43972 2148 44028 2204
rect 44028 2148 44032 2204
rect 43968 2144 44032 2148
rect 6299 1660 6363 1664
rect 6299 1604 6303 1660
rect 6303 1604 6359 1660
rect 6359 1604 6363 1660
rect 6299 1600 6363 1604
rect 6379 1660 6443 1664
rect 6379 1604 6383 1660
rect 6383 1604 6439 1660
rect 6439 1604 6443 1660
rect 6379 1600 6443 1604
rect 6459 1660 6523 1664
rect 6459 1604 6463 1660
rect 6463 1604 6519 1660
rect 6519 1604 6523 1660
rect 6459 1600 6523 1604
rect 6539 1660 6603 1664
rect 6539 1604 6543 1660
rect 6543 1604 6599 1660
rect 6599 1604 6603 1660
rect 6539 1600 6603 1604
rect 16993 1660 17057 1664
rect 16993 1604 16997 1660
rect 16997 1604 17053 1660
rect 17053 1604 17057 1660
rect 16993 1600 17057 1604
rect 17073 1660 17137 1664
rect 17073 1604 17077 1660
rect 17077 1604 17133 1660
rect 17133 1604 17137 1660
rect 17073 1600 17137 1604
rect 17153 1660 17217 1664
rect 17153 1604 17157 1660
rect 17157 1604 17213 1660
rect 17213 1604 17217 1660
rect 17153 1600 17217 1604
rect 17233 1660 17297 1664
rect 17233 1604 17237 1660
rect 17237 1604 17293 1660
rect 17293 1604 17297 1660
rect 17233 1600 17297 1604
rect 27687 1660 27751 1664
rect 27687 1604 27691 1660
rect 27691 1604 27747 1660
rect 27747 1604 27751 1660
rect 27687 1600 27751 1604
rect 27767 1660 27831 1664
rect 27767 1604 27771 1660
rect 27771 1604 27827 1660
rect 27827 1604 27831 1660
rect 27767 1600 27831 1604
rect 27847 1660 27911 1664
rect 27847 1604 27851 1660
rect 27851 1604 27907 1660
rect 27907 1604 27911 1660
rect 27847 1600 27911 1604
rect 27927 1660 27991 1664
rect 27927 1604 27931 1660
rect 27931 1604 27987 1660
rect 27987 1604 27991 1660
rect 27927 1600 27991 1604
rect 38381 1660 38445 1664
rect 38381 1604 38385 1660
rect 38385 1604 38441 1660
rect 38441 1604 38445 1660
rect 38381 1600 38445 1604
rect 38461 1660 38525 1664
rect 38461 1604 38465 1660
rect 38465 1604 38521 1660
rect 38521 1604 38525 1660
rect 38461 1600 38525 1604
rect 38541 1660 38605 1664
rect 38541 1604 38545 1660
rect 38545 1604 38601 1660
rect 38601 1604 38605 1660
rect 38541 1600 38605 1604
rect 38621 1660 38685 1664
rect 38621 1604 38625 1660
rect 38625 1604 38681 1660
rect 38681 1604 38685 1660
rect 38621 1600 38685 1604
rect 21404 1260 21468 1324
rect 34468 1260 34532 1324
rect 11646 1116 11710 1120
rect 11646 1060 11650 1116
rect 11650 1060 11706 1116
rect 11706 1060 11710 1116
rect 11646 1056 11710 1060
rect 11726 1116 11790 1120
rect 11726 1060 11730 1116
rect 11730 1060 11786 1116
rect 11786 1060 11790 1116
rect 11726 1056 11790 1060
rect 11806 1116 11870 1120
rect 11806 1060 11810 1116
rect 11810 1060 11866 1116
rect 11866 1060 11870 1116
rect 11806 1056 11870 1060
rect 11886 1116 11950 1120
rect 11886 1060 11890 1116
rect 11890 1060 11946 1116
rect 11946 1060 11950 1116
rect 11886 1056 11950 1060
rect 22340 1116 22404 1120
rect 22340 1060 22344 1116
rect 22344 1060 22400 1116
rect 22400 1060 22404 1116
rect 22340 1056 22404 1060
rect 22420 1116 22484 1120
rect 22420 1060 22424 1116
rect 22424 1060 22480 1116
rect 22480 1060 22484 1116
rect 22420 1056 22484 1060
rect 22500 1116 22564 1120
rect 22500 1060 22504 1116
rect 22504 1060 22560 1116
rect 22560 1060 22564 1116
rect 22500 1056 22564 1060
rect 22580 1116 22644 1120
rect 22580 1060 22584 1116
rect 22584 1060 22640 1116
rect 22640 1060 22644 1116
rect 22580 1056 22644 1060
rect 33034 1116 33098 1120
rect 33034 1060 33038 1116
rect 33038 1060 33094 1116
rect 33094 1060 33098 1116
rect 33034 1056 33098 1060
rect 33114 1116 33178 1120
rect 33114 1060 33118 1116
rect 33118 1060 33174 1116
rect 33174 1060 33178 1116
rect 33114 1056 33178 1060
rect 33194 1116 33258 1120
rect 33194 1060 33198 1116
rect 33198 1060 33254 1116
rect 33254 1060 33258 1116
rect 33194 1056 33258 1060
rect 33274 1116 33338 1120
rect 33274 1060 33278 1116
rect 33278 1060 33334 1116
rect 33334 1060 33338 1116
rect 33274 1056 33338 1060
rect 43728 1116 43792 1120
rect 43728 1060 43732 1116
rect 43732 1060 43788 1116
rect 43788 1060 43792 1116
rect 43728 1056 43792 1060
rect 43808 1116 43872 1120
rect 43808 1060 43812 1116
rect 43812 1060 43868 1116
rect 43868 1060 43872 1116
rect 43808 1056 43872 1060
rect 43888 1116 43952 1120
rect 43888 1060 43892 1116
rect 43892 1060 43948 1116
rect 43948 1060 43952 1116
rect 43888 1056 43952 1060
rect 43968 1116 44032 1120
rect 43968 1060 43972 1116
rect 43972 1060 44028 1116
rect 44028 1060 44032 1116
rect 43968 1056 44032 1060
<< metal4 >>
rect 6291 8192 6611 8752
rect 6291 8128 6299 8192
rect 6363 8128 6379 8192
rect 6443 8128 6459 8192
rect 6523 8128 6539 8192
rect 6603 8128 6611 8192
rect 6291 7104 6611 8128
rect 6291 7040 6299 7104
rect 6363 7040 6379 7104
rect 6443 7040 6459 7104
rect 6523 7040 6539 7104
rect 6603 7040 6611 7104
rect 6291 6016 6611 7040
rect 6291 5952 6299 6016
rect 6363 5952 6379 6016
rect 6443 5952 6459 6016
rect 6523 5952 6539 6016
rect 6603 5952 6611 6016
rect 6291 4928 6611 5952
rect 6291 4864 6299 4928
rect 6363 4864 6379 4928
rect 6443 4864 6459 4928
rect 6523 4864 6539 4928
rect 6603 4864 6611 4928
rect 6291 3840 6611 4864
rect 6291 3776 6299 3840
rect 6363 3776 6379 3840
rect 6443 3776 6459 3840
rect 6523 3776 6539 3840
rect 6603 3776 6611 3840
rect 6291 2752 6611 3776
rect 6291 2688 6299 2752
rect 6363 2688 6379 2752
rect 6443 2688 6459 2752
rect 6523 2688 6539 2752
rect 6603 2688 6611 2752
rect 6291 1664 6611 2688
rect 6291 1600 6299 1664
rect 6363 1600 6379 1664
rect 6443 1600 6459 1664
rect 6523 1600 6539 1664
rect 6603 1600 6611 1664
rect 6291 1040 6611 1600
rect 11638 8736 11958 8752
rect 11638 8672 11646 8736
rect 11710 8672 11726 8736
rect 11790 8672 11806 8736
rect 11870 8672 11886 8736
rect 11950 8672 11958 8736
rect 11638 7648 11958 8672
rect 11638 7584 11646 7648
rect 11710 7584 11726 7648
rect 11790 7584 11806 7648
rect 11870 7584 11886 7648
rect 11950 7584 11958 7648
rect 11638 6560 11958 7584
rect 11638 6496 11646 6560
rect 11710 6496 11726 6560
rect 11790 6496 11806 6560
rect 11870 6496 11886 6560
rect 11950 6496 11958 6560
rect 11638 5472 11958 6496
rect 11638 5408 11646 5472
rect 11710 5408 11726 5472
rect 11790 5408 11806 5472
rect 11870 5408 11886 5472
rect 11950 5408 11958 5472
rect 11638 4384 11958 5408
rect 11638 4320 11646 4384
rect 11710 4320 11726 4384
rect 11790 4320 11806 4384
rect 11870 4320 11886 4384
rect 11950 4320 11958 4384
rect 11638 3296 11958 4320
rect 11638 3232 11646 3296
rect 11710 3232 11726 3296
rect 11790 3232 11806 3296
rect 11870 3232 11886 3296
rect 11950 3232 11958 3296
rect 11638 2208 11958 3232
rect 11638 2144 11646 2208
rect 11710 2144 11726 2208
rect 11790 2144 11806 2208
rect 11870 2144 11886 2208
rect 11950 2144 11958 2208
rect 11638 1120 11958 2144
rect 11638 1056 11646 1120
rect 11710 1056 11726 1120
rect 11790 1056 11806 1120
rect 11870 1056 11886 1120
rect 11950 1056 11958 1120
rect 11638 1040 11958 1056
rect 16985 8192 17305 8752
rect 16985 8128 16993 8192
rect 17057 8128 17073 8192
rect 17137 8128 17153 8192
rect 17217 8128 17233 8192
rect 17297 8128 17305 8192
rect 16985 7104 17305 8128
rect 16985 7040 16993 7104
rect 17057 7040 17073 7104
rect 17137 7040 17153 7104
rect 17217 7040 17233 7104
rect 17297 7040 17305 7104
rect 16985 6016 17305 7040
rect 16985 5952 16993 6016
rect 17057 5952 17073 6016
rect 17137 5952 17153 6016
rect 17217 5952 17233 6016
rect 17297 5952 17305 6016
rect 16985 4928 17305 5952
rect 16985 4864 16993 4928
rect 17057 4864 17073 4928
rect 17137 4864 17153 4928
rect 17217 4864 17233 4928
rect 17297 4864 17305 4928
rect 16985 3840 17305 4864
rect 16985 3776 16993 3840
rect 17057 3776 17073 3840
rect 17137 3776 17153 3840
rect 17217 3776 17233 3840
rect 17297 3776 17305 3840
rect 16985 2752 17305 3776
rect 22332 8736 22652 8752
rect 22332 8672 22340 8736
rect 22404 8672 22420 8736
rect 22484 8672 22500 8736
rect 22564 8672 22580 8736
rect 22644 8672 22652 8736
rect 22332 7648 22652 8672
rect 24899 8532 24965 8533
rect 24899 8468 24900 8532
rect 24964 8468 24965 8532
rect 24899 8467 24965 8468
rect 22332 7584 22340 7648
rect 22404 7584 22420 7648
rect 22484 7584 22500 7648
rect 22564 7584 22580 7648
rect 22644 7584 22652 7648
rect 22332 6560 22652 7584
rect 22332 6496 22340 6560
rect 22404 6496 22420 6560
rect 22484 6496 22500 6560
rect 22564 6496 22580 6560
rect 22644 6496 22652 6560
rect 22332 5472 22652 6496
rect 22332 5408 22340 5472
rect 22404 5408 22420 5472
rect 22484 5408 22500 5472
rect 22564 5408 22580 5472
rect 22644 5408 22652 5472
rect 22332 4384 22652 5408
rect 22332 4320 22340 4384
rect 22404 4320 22420 4384
rect 22484 4320 22500 4384
rect 22564 4320 22580 4384
rect 22644 4320 22652 4384
rect 22332 3296 22652 4320
rect 22332 3232 22340 3296
rect 22404 3232 22420 3296
rect 22484 3232 22500 3296
rect 22564 3232 22580 3296
rect 22644 3232 22652 3296
rect 21403 2820 21469 2821
rect 21403 2756 21404 2820
rect 21468 2756 21469 2820
rect 21403 2755 21469 2756
rect 16985 2688 16993 2752
rect 17057 2688 17073 2752
rect 17137 2688 17153 2752
rect 17217 2688 17233 2752
rect 17297 2688 17305 2752
rect 16985 1664 17305 2688
rect 16985 1600 16993 1664
rect 17057 1600 17073 1664
rect 17137 1600 17153 1664
rect 17217 1600 17233 1664
rect 17297 1600 17305 1664
rect 16985 1040 17305 1600
rect 21406 1325 21466 2755
rect 22332 2208 22652 3232
rect 24902 2685 24962 8467
rect 25083 8396 25149 8397
rect 25083 8332 25084 8396
rect 25148 8332 25149 8396
rect 25083 8331 25149 8332
rect 24899 2684 24965 2685
rect 24899 2620 24900 2684
rect 24964 2620 24965 2684
rect 24899 2619 24965 2620
rect 25086 2277 25146 8331
rect 27679 8192 27999 8752
rect 27679 8128 27687 8192
rect 27751 8128 27767 8192
rect 27831 8128 27847 8192
rect 27911 8128 27927 8192
rect 27991 8128 27999 8192
rect 27679 7104 27999 8128
rect 27679 7040 27687 7104
rect 27751 7040 27767 7104
rect 27831 7040 27847 7104
rect 27911 7040 27927 7104
rect 27991 7040 27999 7104
rect 27679 6016 27999 7040
rect 27679 5952 27687 6016
rect 27751 5952 27767 6016
rect 27831 5952 27847 6016
rect 27911 5952 27927 6016
rect 27991 5952 27999 6016
rect 27679 4928 27999 5952
rect 27679 4864 27687 4928
rect 27751 4864 27767 4928
rect 27831 4864 27847 4928
rect 27911 4864 27927 4928
rect 27991 4864 27999 4928
rect 27679 3840 27999 4864
rect 27679 3776 27687 3840
rect 27751 3776 27767 3840
rect 27831 3776 27847 3840
rect 27911 3776 27927 3840
rect 27991 3776 27999 3840
rect 27679 2752 27999 3776
rect 27679 2688 27687 2752
rect 27751 2688 27767 2752
rect 27831 2688 27847 2752
rect 27911 2688 27927 2752
rect 27991 2688 27999 2752
rect 25083 2276 25149 2277
rect 25083 2212 25084 2276
rect 25148 2212 25149 2276
rect 25083 2211 25149 2212
rect 22332 2144 22340 2208
rect 22404 2144 22420 2208
rect 22484 2144 22500 2208
rect 22564 2144 22580 2208
rect 22644 2144 22652 2208
rect 21403 1324 21469 1325
rect 21403 1260 21404 1324
rect 21468 1260 21469 1324
rect 21403 1259 21469 1260
rect 22332 1120 22652 2144
rect 22332 1056 22340 1120
rect 22404 1056 22420 1120
rect 22484 1056 22500 1120
rect 22564 1056 22580 1120
rect 22644 1056 22652 1120
rect 22332 1040 22652 1056
rect 27679 1664 27999 2688
rect 27679 1600 27687 1664
rect 27751 1600 27767 1664
rect 27831 1600 27847 1664
rect 27911 1600 27927 1664
rect 27991 1600 27999 1664
rect 27679 1040 27999 1600
rect 33026 8736 33346 8752
rect 33026 8672 33034 8736
rect 33098 8672 33114 8736
rect 33178 8672 33194 8736
rect 33258 8672 33274 8736
rect 33338 8672 33346 8736
rect 33026 7648 33346 8672
rect 33026 7584 33034 7648
rect 33098 7584 33114 7648
rect 33178 7584 33194 7648
rect 33258 7584 33274 7648
rect 33338 7584 33346 7648
rect 33026 6560 33346 7584
rect 33026 6496 33034 6560
rect 33098 6496 33114 6560
rect 33178 6496 33194 6560
rect 33258 6496 33274 6560
rect 33338 6496 33346 6560
rect 33026 5472 33346 6496
rect 33026 5408 33034 5472
rect 33098 5408 33114 5472
rect 33178 5408 33194 5472
rect 33258 5408 33274 5472
rect 33338 5408 33346 5472
rect 33026 4384 33346 5408
rect 33026 4320 33034 4384
rect 33098 4320 33114 4384
rect 33178 4320 33194 4384
rect 33258 4320 33274 4384
rect 33338 4320 33346 4384
rect 33026 3296 33346 4320
rect 38373 8192 38693 8752
rect 38373 8128 38381 8192
rect 38445 8128 38461 8192
rect 38525 8128 38541 8192
rect 38605 8128 38621 8192
rect 38685 8128 38693 8192
rect 38373 7104 38693 8128
rect 38373 7040 38381 7104
rect 38445 7040 38461 7104
rect 38525 7040 38541 7104
rect 38605 7040 38621 7104
rect 38685 7040 38693 7104
rect 38373 6016 38693 7040
rect 38373 5952 38381 6016
rect 38445 5952 38461 6016
rect 38525 5952 38541 6016
rect 38605 5952 38621 6016
rect 38685 5952 38693 6016
rect 38373 4928 38693 5952
rect 38373 4864 38381 4928
rect 38445 4864 38461 4928
rect 38525 4864 38541 4928
rect 38605 4864 38621 4928
rect 38685 4864 38693 4928
rect 38373 3840 38693 4864
rect 38373 3776 38381 3840
rect 38445 3776 38461 3840
rect 38525 3776 38541 3840
rect 38605 3776 38621 3840
rect 38685 3776 38693 3840
rect 34467 3636 34533 3637
rect 34467 3572 34468 3636
rect 34532 3572 34533 3636
rect 34467 3571 34533 3572
rect 33026 3232 33034 3296
rect 33098 3232 33114 3296
rect 33178 3232 33194 3296
rect 33258 3232 33274 3296
rect 33338 3232 33346 3296
rect 33026 2208 33346 3232
rect 33026 2144 33034 2208
rect 33098 2144 33114 2208
rect 33178 2144 33194 2208
rect 33258 2144 33274 2208
rect 33338 2144 33346 2208
rect 33026 1120 33346 2144
rect 34470 1325 34530 3571
rect 38373 2752 38693 3776
rect 38373 2688 38381 2752
rect 38445 2688 38461 2752
rect 38525 2688 38541 2752
rect 38605 2688 38621 2752
rect 38685 2688 38693 2752
rect 38373 1664 38693 2688
rect 38373 1600 38381 1664
rect 38445 1600 38461 1664
rect 38525 1600 38541 1664
rect 38605 1600 38621 1664
rect 38685 1600 38693 1664
rect 34467 1324 34533 1325
rect 34467 1260 34468 1324
rect 34532 1260 34533 1324
rect 34467 1259 34533 1260
rect 33026 1056 33034 1120
rect 33098 1056 33114 1120
rect 33178 1056 33194 1120
rect 33258 1056 33274 1120
rect 33338 1056 33346 1120
rect 33026 1040 33346 1056
rect 38373 1040 38693 1600
rect 43720 8736 44040 8752
rect 43720 8672 43728 8736
rect 43792 8672 43808 8736
rect 43872 8672 43888 8736
rect 43952 8672 43968 8736
rect 44032 8672 44040 8736
rect 43720 7648 44040 8672
rect 43720 7584 43728 7648
rect 43792 7584 43808 7648
rect 43872 7584 43888 7648
rect 43952 7584 43968 7648
rect 44032 7584 44040 7648
rect 43720 6560 44040 7584
rect 43720 6496 43728 6560
rect 43792 6496 43808 6560
rect 43872 6496 43888 6560
rect 43952 6496 43968 6560
rect 44032 6496 44040 6560
rect 43720 5472 44040 6496
rect 43720 5408 43728 5472
rect 43792 5408 43808 5472
rect 43872 5408 43888 5472
rect 43952 5408 43968 5472
rect 44032 5408 44040 5472
rect 43720 4384 44040 5408
rect 43720 4320 43728 4384
rect 43792 4320 43808 4384
rect 43872 4320 43888 4384
rect 43952 4320 43968 4384
rect 44032 4320 44040 4384
rect 43720 3296 44040 4320
rect 43720 3232 43728 3296
rect 43792 3232 43808 3296
rect 43872 3232 43888 3296
rect 43952 3232 43968 3296
rect 44032 3232 44040 3296
rect 43720 2208 44040 3232
rect 43720 2144 43728 2208
rect 43792 2144 43808 2208
rect 43872 2144 43888 2208
rect 43952 2144 43968 2208
rect 44032 2144 44040 2208
rect 43720 1120 44040 2144
rect 43720 1056 43728 1120
rect 43792 1056 43808 1120
rect 43872 1056 43888 1120
rect 43952 1056 43968 1120
rect 44032 1056 44040 1120
rect 43720 1040 44040 1056
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28796 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 4324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 35420 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 5060 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_218 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21160 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_231
timestamp 1688980957
transform 1 0 22356 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_275
timestamp 1688980957
transform 1 0 26404 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_299
timestamp 1688980957
transform 1 0 28612 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_303
timestamp 1688980957
transform 1 0 28980 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_371
timestamp 1688980957
transform 1 0 35236 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_390
timestamp 1688980957
transform 1 0 36984 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_442 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 41768 0 1 1088
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_461
timestamp 1688980957
transform 1 0 43516 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_62
timestamp 1688980957
transform 1 0 6808 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_74
timestamp 1688980957
transform 1 0 7912 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_86
timestamp 1688980957
transform 1 0 9016 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_98
timestamp 1688980957
transform 1 0 10120 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1688980957
transform 1 0 11224 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_140
timestamp 1688980957
transform 1 0 13984 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_145
timestamp 1688980957
transform 1 0 14444 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_204
timestamp 1688980957
transform 1 0 19872 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_233
timestamp 1688980957
transform 1 0 22540 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_262
timestamp 1688980957
transform 1 0 25208 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_275
timestamp 1688980957
transform 1 0 26404 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_299
timestamp 1688980957
transform 1 0 28612 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_310
timestamp 1688980957
transform 1 0 29624 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_321
timestamp 1688980957
transform 1 0 30636 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_371
timestamp 1688980957
transform 1 0 35236 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_386
timestamp 1688980957
transform 1 0 36616 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_399 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37812 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_412 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39008 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_420
timestamp 1688980957
transform 1 0 39744 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_425
timestamp 1688980957
transform 1 0 40204 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_431
timestamp 1688980957
transform 1 0 40756 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_435
timestamp 1688980957
transform 1 0 41124 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_461
timestamp 1688980957
transform 1 0 43516 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_144
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_156
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_162
timestamp 1688980957
transform 1 0 16008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_166
timestamp 1688980957
transform 1 0 16376 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_170
timestamp 1688980957
transform 1 0 16744 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_175
timestamp 1688980957
transform 1 0 17204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_224
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_235
timestamp 1688980957
transform 1 0 22724 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_240
timestamp 1688980957
transform 1 0 23184 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_256
timestamp 1688980957
transform 1 0 24656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_287
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_295
timestamp 1688980957
transform 1 0 28244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_306
timestamp 1688980957
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_332
timestamp 1688980957
transform 1 0 31648 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_336
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_344
timestamp 1688980957
transform 1 0 32752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_355
timestamp 1688980957
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_386
timestamp 1688980957
transform 1 0 36616 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_413
timestamp 1688980957
transform 1 0 39100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_429
timestamp 1688980957
transform 1 0 40572 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_450
timestamp 1688980957
transform 1 0 42504 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_202
timestamp 1688980957
transform 1 0 19688 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_214
timestamp 1688980957
transform 1 0 20792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_222
timestamp 1688980957
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_229
timestamp 1688980957
transform 1 0 22172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_241
timestamp 1688980957
transform 1 0 23276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_253
timestamp 1688980957
transform 1 0 24380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_265
timestamp 1688980957
transform 1 0 25484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_277
timestamp 1688980957
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_290
timestamp 1688980957
transform 1 0 27784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_302
timestamp 1688980957
transform 1 0 28888 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_310
timestamp 1688980957
transform 1 0 29624 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_322
timestamp 1688980957
transform 1 0 30728 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_334
timestamp 1688980957
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_461
timestamp 1688980957
transform 1 0 43516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_461
timestamp 1688980957
transform 1 0 43516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_461
timestamp 1688980957
transform 1 0 43516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_461
timestamp 1688980957
transform 1 0 43516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_461
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_457
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_461
timestamp 1688980957
transform 1 0 43516 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_21
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_37
timestamp 1688980957
transform 1 0 4508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_45
timestamp 1688980957
transform 1 0 5244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_76
timestamp 1688980957
transform 1 0 8096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_91
timestamp 1688980957
transform 1 0 9476 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_99
timestamp 1688980957
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_117
timestamp 1688980957
transform 1 0 11868 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_122
timestamp 1688980957
transform 1 0 12328 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_134
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_145
timestamp 1688980957
transform 1 0 14444 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_157
timestamp 1688980957
transform 1 0 15548 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_163
timestamp 1688980957
transform 1 0 16100 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_191
timestamp 1688980957
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_195
timestamp 1688980957
transform 1 0 19044 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_197
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_209
timestamp 1688980957
transform 1 0 20332 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_214
timestamp 1688980957
transform 1 0 20792 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1688980957
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_253
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_260
timestamp 1688980957
transform 1 0 25024 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_272
timestamp 1688980957
transform 1 0 26128 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_285
timestamp 1688980957
transform 1 0 27324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_297
timestamp 1688980957
transform 1 0 28428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_306
timestamp 1688980957
transform 1 0 29256 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_309
timestamp 1688980957
transform 1 0 29532 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_321
timestamp 1688980957
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_345
timestamp 1688980957
transform 1 0 32844 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_352
timestamp 1688980957
transform 1 0 33488 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_365
timestamp 1688980957
transform 1 0 34684 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_375
timestamp 1688980957
transform 1 0 35604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_387
timestamp 1688980957
transform 1 0 36708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_399
timestamp 1688980957
transform 1 0 37812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_411
timestamp 1688980957
transform 1 0 38916 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_419
timestamp 1688980957
transform 1 0 39652 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_427
timestamp 1688980957
transform 1 0 40388 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_439
timestamp 1688980957
transform 1 0 41492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_446
timestamp 1688980957
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_457
timestamp 1688980957
transform 1 0 43148 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36156 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38916 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 39192 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 39468 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 39836 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 40112 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 40388 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 40664 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 40940 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 41216 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 41492 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 36432 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 36708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 37260 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 37536 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 37812 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 38088 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 36340 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 38364 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 38640 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 5428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 5704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 9200 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1688980957
transform 1 0 9476 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1688980957
transform 1 0 9752 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 10028 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 6532 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 6624 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 6900 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 7176 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 10304 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 13156 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 13432 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 14904 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 10580 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 10856 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1688980957
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1688980957
transform 1 0 11776 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 12052 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1688980957
transform 1 0 12328 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1688980957
transform 1 0 12604 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 14352 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform 1 0 17480 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1688980957
transform 1 0 18032 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform 1 0 18584 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform 1 0 14628 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform 1 0 14904 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1688980957
transform 1 0 15456 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1688980957
transform 1 0 16008 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1688980957
transform 1 0 16928 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1688980957
transform 1 0 34316 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__00_
timestamp 1688980957
transform 1 0 22172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__01_
timestamp 1688980957
transform 1 0 22448 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__02_
timestamp 1688980957
transform 1 0 22724 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__03_
timestamp 1688980957
transform 1 0 23000 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__04_
timestamp 1688980957
transform 1 0 23276 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__05_
timestamp 1688980957
transform 1 0 23552 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__06_
timestamp 1688980957
transform 1 0 24104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__07_
timestamp 1688980957
transform 1 0 24380 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__08_
timestamp 1688980957
transform 1 0 19688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__09_
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__10_
timestamp 1688980957
transform 1 0 19228 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__11_
timestamp 1688980957
transform 1 0 20240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__12_
timestamp 1688980957
transform 1 0 20608 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__13_
timestamp 1688980957
transform 1 0 20884 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__14_
timestamp 1688980957
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__15_
timestamp 1688980957
transform 1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__16_
timestamp 1688980957
transform 1 0 24656 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__17_
timestamp 1688980957
transform 1 0 24932 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__18_
timestamp 1688980957
transform 1 0 27508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__19_
timestamp 1688980957
transform 1 0 28980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__20_
timestamp 1688980957
transform 1 0 28612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__21_
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__22_
timestamp 1688980957
transform 1 0 29808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__23_
timestamp 1688980957
transform 1 0 31740 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__24_
timestamp 1688980957
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__25_
timestamp 1688980957
transform 1 0 26588 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__26_
timestamp 1688980957
transform 1 0 27968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__27_
timestamp 1688980957
transform 1 0 29164 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__28_
timestamp 1688980957
transform 1 0 26680 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__29_
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__30_
timestamp 1688980957
transform 1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__31_
timestamp 1688980957
transform 1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__32_
timestamp 1688980957
transform 1 0 18952 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__33_
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__34_
timestamp 1688980957
transform 1 0 16284 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__35_
timestamp 1688980957
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__36_
timestamp 1688980957
transform 1 0 15732 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__37_
timestamp 1688980957
transform 1 0 15456 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__38_
timestamp 1688980957
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__39_
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__40_
timestamp 1688980957
transform 1 0 18676 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__41_
timestamp 1688980957
transform 1 0 18400 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__42_
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__43_
timestamp 1688980957
transform 1 0 17572 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__44_
timestamp 1688980957
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__45_
timestamp 1688980957
transform 1 0 17296 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__46_
timestamp 1688980957
transform 1 0 17020 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__47_
timestamp 1688980957
transform 1 0 16744 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__48_
timestamp 1688980957
transform 1 0 17848 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__49_
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__50_
timestamp 1688980957
transform 1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__51_
timestamp 1688980957
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output75 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24472 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 28704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1688980957
transform 1 0 31004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 32936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1688980957
transform 1 0 35236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 39836 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 41584 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1688980957
transform 1 0 43240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 5428 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1688980957
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1688980957
transform 1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1688980957
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1688980957
transform 1 0 18308 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1688980957
transform 1 0 20424 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1688980957
transform 1 0 22540 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1688980957
transform 1 0 19504 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 20056 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform 1 0 19504 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1688980957
transform 1 0 19872 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1688980957
transform 1 0 22908 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 23276 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1688980957
transform 1 0 23828 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 24748 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 25300 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 25852 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 26956 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 20608 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 21160 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1688980957
transform 1 0 20240 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1688980957
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 21988 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1688980957
transform 1 0 21344 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1688980957
transform 1 0 22540 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 25300 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 30084 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1688980957
transform 1 0 28336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 28704 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 30636 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1688980957
transform 1 0 30268 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform 1 0 31188 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 27508 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform 1 0 25852 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 28060 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform 1 0 26956 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1688980957
transform 1 0 26496 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 28060 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform 1 0 29532 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 27508 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1688980957
transform 1 0 29256 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 29716 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 34316 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 34684 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output133
timestamp 1688980957
transform 1 0 33212 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1688980957
transform 1 0 34868 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 33764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 35604 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 32108 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform 1 0 32660 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform 1 0 32108 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 30820 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 31372 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 33212 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 33764 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 32660 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1688980957
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 43884 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 43884 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 43884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 43884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 43884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 43884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 43884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 43884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 43884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 43884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 43884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform 1 0 29348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform 1 0 25300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 14168 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 16008 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform 1 0 18124 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 20792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 23828 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 26128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 29072 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 37536 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 37260 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 38088 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 38732 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 39928 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 40848 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 27600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 24748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 26404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 28704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 18584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 20516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 25024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 27232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 33488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 36340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 40664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 42228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 37168 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 34334 0 34390 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 37094 0 37150 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 37370 0 37426 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 37646 0 37702 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 37922 0 37978 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 38198 0 38254 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 38474 0 38530 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 38750 0 38806 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 39026 0 39082 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 39302 0 39358 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 39578 0 39634 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 34610 0 34666 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 34886 0 34942 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 35162 0 35218 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 35438 0 35494 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 35714 0 35770 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 35990 0 36046 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 36266 0 36322 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 36542 0 36598 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 36818 0 36874 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 3422 9840 3478 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 24582 9840 24638 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 26698 9840 26754 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 28814 9840 28870 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 30930 9840 30986 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 33046 9840 33102 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 35162 9840 35218 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 37278 9840 37334 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 39394 9840 39450 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 41510 9840 41566 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 43626 9840 43682 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 5538 9840 5594 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 7654 9840 7710 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 9770 9840 9826 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 11886 9840 11942 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 14002 9840 14058 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 16118 9840 16174 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 18234 9840 18290 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 20350 9840 20406 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 22466 9840 22522 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 5354 0 5410 160 0 FreeSans 224 90 0 0 N1END[0]
port 40 nsew signal input
flabel metal2 s 5630 0 5686 160 0 FreeSans 224 90 0 0 N1END[1]
port 41 nsew signal input
flabel metal2 s 5906 0 5962 160 0 FreeSans 224 90 0 0 N1END[2]
port 42 nsew signal input
flabel metal2 s 6182 0 6238 160 0 FreeSans 224 90 0 0 N1END[3]
port 43 nsew signal input
flabel metal2 s 8666 0 8722 160 0 FreeSans 224 90 0 0 N2END[0]
port 44 nsew signal input
flabel metal2 s 8942 0 8998 160 0 FreeSans 224 90 0 0 N2END[1]
port 45 nsew signal input
flabel metal2 s 9218 0 9274 160 0 FreeSans 224 90 0 0 N2END[2]
port 46 nsew signal input
flabel metal2 s 9494 0 9550 160 0 FreeSans 224 90 0 0 N2END[3]
port 47 nsew signal input
flabel metal2 s 9770 0 9826 160 0 FreeSans 224 90 0 0 N2END[4]
port 48 nsew signal input
flabel metal2 s 10046 0 10102 160 0 FreeSans 224 90 0 0 N2END[5]
port 49 nsew signal input
flabel metal2 s 10322 0 10378 160 0 FreeSans 224 90 0 0 N2END[6]
port 50 nsew signal input
flabel metal2 s 10598 0 10654 160 0 FreeSans 224 90 0 0 N2END[7]
port 51 nsew signal input
flabel metal2 s 6458 0 6514 160 0 FreeSans 224 90 0 0 N2MID[0]
port 52 nsew signal input
flabel metal2 s 6734 0 6790 160 0 FreeSans 224 90 0 0 N2MID[1]
port 53 nsew signal input
flabel metal2 s 7010 0 7066 160 0 FreeSans 224 90 0 0 N2MID[2]
port 54 nsew signal input
flabel metal2 s 7286 0 7342 160 0 FreeSans 224 90 0 0 N2MID[3]
port 55 nsew signal input
flabel metal2 s 7562 0 7618 160 0 FreeSans 224 90 0 0 N2MID[4]
port 56 nsew signal input
flabel metal2 s 7838 0 7894 160 0 FreeSans 224 90 0 0 N2MID[5]
port 57 nsew signal input
flabel metal2 s 8114 0 8170 160 0 FreeSans 224 90 0 0 N2MID[6]
port 58 nsew signal input
flabel metal2 s 8390 0 8446 160 0 FreeSans 224 90 0 0 N2MID[7]
port 59 nsew signal input
flabel metal2 s 10874 0 10930 160 0 FreeSans 224 90 0 0 N4END[0]
port 60 nsew signal input
flabel metal2 s 13634 0 13690 160 0 FreeSans 224 90 0 0 N4END[10]
port 61 nsew signal input
flabel metal2 s 13910 0 13966 160 0 FreeSans 224 90 0 0 N4END[11]
port 62 nsew signal input
flabel metal2 s 14186 0 14242 160 0 FreeSans 224 90 0 0 N4END[12]
port 63 nsew signal input
flabel metal2 s 14462 0 14518 160 0 FreeSans 224 90 0 0 N4END[13]
port 64 nsew signal input
flabel metal2 s 14738 0 14794 160 0 FreeSans 224 90 0 0 N4END[14]
port 65 nsew signal input
flabel metal2 s 15014 0 15070 160 0 FreeSans 224 90 0 0 N4END[15]
port 66 nsew signal input
flabel metal2 s 11150 0 11206 160 0 FreeSans 224 90 0 0 N4END[1]
port 67 nsew signal input
flabel metal2 s 11426 0 11482 160 0 FreeSans 224 90 0 0 N4END[2]
port 68 nsew signal input
flabel metal2 s 11702 0 11758 160 0 FreeSans 224 90 0 0 N4END[3]
port 69 nsew signal input
flabel metal2 s 11978 0 12034 160 0 FreeSans 224 90 0 0 N4END[4]
port 70 nsew signal input
flabel metal2 s 12254 0 12310 160 0 FreeSans 224 90 0 0 N4END[5]
port 71 nsew signal input
flabel metal2 s 12530 0 12586 160 0 FreeSans 224 90 0 0 N4END[6]
port 72 nsew signal input
flabel metal2 s 12806 0 12862 160 0 FreeSans 224 90 0 0 N4END[7]
port 73 nsew signal input
flabel metal2 s 13082 0 13138 160 0 FreeSans 224 90 0 0 N4END[8]
port 74 nsew signal input
flabel metal2 s 13358 0 13414 160 0 FreeSans 224 90 0 0 N4END[9]
port 75 nsew signal input
flabel metal2 s 15290 0 15346 160 0 FreeSans 224 90 0 0 NN4END[0]
port 76 nsew signal input
flabel metal2 s 18050 0 18106 160 0 FreeSans 224 90 0 0 NN4END[10]
port 77 nsew signal input
flabel metal2 s 18326 0 18382 160 0 FreeSans 224 90 0 0 NN4END[11]
port 78 nsew signal input
flabel metal2 s 18602 0 18658 160 0 FreeSans 224 90 0 0 NN4END[12]
port 79 nsew signal input
flabel metal2 s 18878 0 18934 160 0 FreeSans 224 90 0 0 NN4END[13]
port 80 nsew signal input
flabel metal2 s 19154 0 19210 160 0 FreeSans 224 90 0 0 NN4END[14]
port 81 nsew signal input
flabel metal2 s 19430 0 19486 160 0 FreeSans 224 90 0 0 NN4END[15]
port 82 nsew signal input
flabel metal2 s 15566 0 15622 160 0 FreeSans 224 90 0 0 NN4END[1]
port 83 nsew signal input
flabel metal2 s 15842 0 15898 160 0 FreeSans 224 90 0 0 NN4END[2]
port 84 nsew signal input
flabel metal2 s 16118 0 16174 160 0 FreeSans 224 90 0 0 NN4END[3]
port 85 nsew signal input
flabel metal2 s 16394 0 16450 160 0 FreeSans 224 90 0 0 NN4END[4]
port 86 nsew signal input
flabel metal2 s 16670 0 16726 160 0 FreeSans 224 90 0 0 NN4END[5]
port 87 nsew signal input
flabel metal2 s 16946 0 17002 160 0 FreeSans 224 90 0 0 NN4END[6]
port 88 nsew signal input
flabel metal2 s 17222 0 17278 160 0 FreeSans 224 90 0 0 NN4END[7]
port 89 nsew signal input
flabel metal2 s 17498 0 17554 160 0 FreeSans 224 90 0 0 NN4END[8]
port 90 nsew signal input
flabel metal2 s 17774 0 17830 160 0 FreeSans 224 90 0 0 NN4END[9]
port 91 nsew signal input
flabel metal2 s 19706 0 19762 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 92 nsew signal tristate
flabel metal2 s 19982 0 20038 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 93 nsew signal tristate
flabel metal2 s 20258 0 20314 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 94 nsew signal tristate
flabel metal2 s 20534 0 20590 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 95 nsew signal tristate
flabel metal2 s 23018 0 23074 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 96 nsew signal tristate
flabel metal2 s 23294 0 23350 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 97 nsew signal tristate
flabel metal2 s 23570 0 23626 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 98 nsew signal tristate
flabel metal2 s 23846 0 23902 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 99 nsew signal tristate
flabel metal2 s 24122 0 24178 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 100 nsew signal tristate
flabel metal2 s 24398 0 24454 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 101 nsew signal tristate
flabel metal2 s 24674 0 24730 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 102 nsew signal tristate
flabel metal2 s 24950 0 25006 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 103 nsew signal tristate
flabel metal2 s 20810 0 20866 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 104 nsew signal tristate
flabel metal2 s 21086 0 21142 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 105 nsew signal tristate
flabel metal2 s 21362 0 21418 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 106 nsew signal tristate
flabel metal2 s 21638 0 21694 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 107 nsew signal tristate
flabel metal2 s 21914 0 21970 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 108 nsew signal tristate
flabel metal2 s 22190 0 22246 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 109 nsew signal tristate
flabel metal2 s 22466 0 22522 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 110 nsew signal tristate
flabel metal2 s 22742 0 22798 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 111 nsew signal tristate
flabel metal2 s 25226 0 25282 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 112 nsew signal tristate
flabel metal2 s 27986 0 28042 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 113 nsew signal tristate
flabel metal2 s 28262 0 28318 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 114 nsew signal tristate
flabel metal2 s 28538 0 28594 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 115 nsew signal tristate
flabel metal2 s 28814 0 28870 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 116 nsew signal tristate
flabel metal2 s 29090 0 29146 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 117 nsew signal tristate
flabel metal2 s 29366 0 29422 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 118 nsew signal tristate
flabel metal2 s 25502 0 25558 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 119 nsew signal tristate
flabel metal2 s 25778 0 25834 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 120 nsew signal tristate
flabel metal2 s 26054 0 26110 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 121 nsew signal tristate
flabel metal2 s 26330 0 26386 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 122 nsew signal tristate
flabel metal2 s 26606 0 26662 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 123 nsew signal tristate
flabel metal2 s 26882 0 26938 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 124 nsew signal tristate
flabel metal2 s 27158 0 27214 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 125 nsew signal tristate
flabel metal2 s 27434 0 27490 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 126 nsew signal tristate
flabel metal2 s 27710 0 27766 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 127 nsew signal tristate
flabel metal2 s 29642 0 29698 160 0 FreeSans 224 90 0 0 SS4BEG[0]
port 128 nsew signal tristate
flabel metal2 s 32402 0 32458 160 0 FreeSans 224 90 0 0 SS4BEG[10]
port 129 nsew signal tristate
flabel metal2 s 32678 0 32734 160 0 FreeSans 224 90 0 0 SS4BEG[11]
port 130 nsew signal tristate
flabel metal2 s 32954 0 33010 160 0 FreeSans 224 90 0 0 SS4BEG[12]
port 131 nsew signal tristate
flabel metal2 s 33230 0 33286 160 0 FreeSans 224 90 0 0 SS4BEG[13]
port 132 nsew signal tristate
flabel metal2 s 33506 0 33562 160 0 FreeSans 224 90 0 0 SS4BEG[14]
port 133 nsew signal tristate
flabel metal2 s 33782 0 33838 160 0 FreeSans 224 90 0 0 SS4BEG[15]
port 134 nsew signal tristate
flabel metal2 s 29918 0 29974 160 0 FreeSans 224 90 0 0 SS4BEG[1]
port 135 nsew signal tristate
flabel metal2 s 30194 0 30250 160 0 FreeSans 224 90 0 0 SS4BEG[2]
port 136 nsew signal tristate
flabel metal2 s 30470 0 30526 160 0 FreeSans 224 90 0 0 SS4BEG[3]
port 137 nsew signal tristate
flabel metal2 s 30746 0 30802 160 0 FreeSans 224 90 0 0 SS4BEG[4]
port 138 nsew signal tristate
flabel metal2 s 31022 0 31078 160 0 FreeSans 224 90 0 0 SS4BEG[5]
port 139 nsew signal tristate
flabel metal2 s 31298 0 31354 160 0 FreeSans 224 90 0 0 SS4BEG[6]
port 140 nsew signal tristate
flabel metal2 s 31574 0 31630 160 0 FreeSans 224 90 0 0 SS4BEG[7]
port 141 nsew signal tristate
flabel metal2 s 31850 0 31906 160 0 FreeSans 224 90 0 0 SS4BEG[8]
port 142 nsew signal tristate
flabel metal2 s 32126 0 32182 160 0 FreeSans 224 90 0 0 SS4BEG[9]
port 143 nsew signal tristate
flabel metal2 s 34058 0 34114 160 0 FreeSans 224 90 0 0 UserCLK
port 144 nsew signal input
flabel metal2 s 1306 9840 1362 10000 0 FreeSans 224 90 0 0 UserCLKo
port 145 nsew signal tristate
flabel metal4 s 6291 1040 6611 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 16985 1040 17305 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 27679 1040 27999 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 38373 1040 38693 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 11638 1040 11958 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 22332 1040 22652 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 33026 1040 33346 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 43720 1040 44040 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
rlabel metal1 22494 8160 22494 8160 0 vccd1
rlabel via1 22572 8704 22572 8704 0 vssd1
rlabel metal2 34362 415 34362 415 0 FrameStrobe[0]
rlabel metal2 37175 68 37175 68 0 FrameStrobe[10]
rlabel metal2 37497 68 37497 68 0 FrameStrobe[11]
rlabel metal2 37773 68 37773 68 0 FrameStrobe[12]
rlabel metal2 37950 194 37950 194 0 FrameStrobe[13]
rlabel metal2 38325 68 38325 68 0 FrameStrobe[14]
rlabel metal2 38555 68 38555 68 0 FrameStrobe[15]
rlabel metal2 38877 68 38877 68 0 FrameStrobe[16]
rlabel metal2 39054 347 39054 347 0 FrameStrobe[17]
rlabel metal2 39330 738 39330 738 0 FrameStrobe[18]
rlabel metal2 39797 68 39797 68 0 FrameStrobe[19]
rlabel metal2 34737 68 34737 68 0 FrameStrobe[1]
rlabel metal2 34914 347 34914 347 0 FrameStrobe[2]
rlabel metal2 35289 68 35289 68 0 FrameStrobe[3]
rlabel metal2 35466 364 35466 364 0 FrameStrobe[4]
rlabel metal2 35795 68 35795 68 0 FrameStrobe[5]
rlabel metal2 36018 806 36018 806 0 FrameStrobe[6]
rlabel metal2 36347 68 36347 68 0 FrameStrobe[7]
rlabel metal2 36570 670 36570 670 0 FrameStrobe[8]
rlabel metal2 36846 160 36846 160 0 FrameStrobe[9]
rlabel metal1 3726 8602 3726 8602 0 FrameStrobe_O[0]
rlabel metal2 24610 9445 24610 9445 0 FrameStrobe_O[10]
rlabel metal1 26956 8602 26956 8602 0 FrameStrobe_O[11]
rlabel metal2 28842 9445 28842 9445 0 FrameStrobe_O[12]
rlabel metal1 31096 8602 31096 8602 0 FrameStrobe_O[13]
rlabel metal2 33074 9445 33074 9445 0 FrameStrobe_O[14]
rlabel metal1 35328 8602 35328 8602 0 FrameStrobe_O[15]
rlabel metal2 37306 9445 37306 9445 0 FrameStrobe_O[16]
rlabel metal2 39422 9224 39422 9224 0 FrameStrobe_O[17]
rlabel metal2 41538 9224 41538 9224 0 FrameStrobe_O[18]
rlabel metal1 43562 8602 43562 8602 0 FrameStrobe_O[19]
rlabel metal2 5566 9445 5566 9445 0 FrameStrobe_O[1]
rlabel metal1 7820 8602 7820 8602 0 FrameStrobe_O[2]
rlabel metal2 9798 9785 9798 9785 0 FrameStrobe_O[3]
rlabel metal1 12098 8602 12098 8602 0 FrameStrobe_O[4]
rlabel metal1 14168 8602 14168 8602 0 FrameStrobe_O[5]
rlabel metal1 16284 8602 16284 8602 0 FrameStrobe_O[6]
rlabel metal1 18400 8602 18400 8602 0 FrameStrobe_O[7]
rlabel metal1 20516 8602 20516 8602 0 FrameStrobe_O[8]
rlabel metal2 22770 9231 22770 9231 0 FrameStrobe_O[9]
rlabel metal1 27922 2414 27922 2414 0 FrameStrobe_O_i\[0\]
rlabel metal1 25300 2414 25300 2414 0 FrameStrobe_O_i\[10\]
rlabel metal1 28290 2890 28290 2890 0 FrameStrobe_O_i\[11\]
rlabel metal1 30360 2414 30360 2414 0 FrameStrobe_O_i\[12\]
rlabel metal1 31552 2410 31552 2410 0 FrameStrobe_O_i\[13\]
rlabel metal1 37582 2040 37582 2040 0 FrameStrobe_O_i\[14\]
rlabel metal1 36938 2074 36938 2074 0 FrameStrobe_O_i\[15\]
rlabel metal1 38042 2074 38042 2074 0 FrameStrobe_O_i\[16\]
rlabel metal1 39238 2074 39238 2074 0 FrameStrobe_O_i\[17\]
rlabel metal1 40434 2074 40434 2074 0 FrameStrobe_O_i\[18\]
rlabel metal1 42458 1938 42458 1938 0 FrameStrobe_O_i\[19\]
rlabel metal1 24794 2482 24794 2482 0 FrameStrobe_O_i\[1\]
rlabel metal1 26726 2822 26726 2822 0 FrameStrobe_O_i\[2\]
rlabel metal2 29118 2652 29118 2652 0 FrameStrobe_O_i\[3\]
rlabel metal1 24426 2380 24426 2380 0 FrameStrobe_O_i\[4\]
rlabel metal1 14260 2074 14260 2074 0 FrameStrobe_O_i\[5\]
rlabel metal1 16192 2074 16192 2074 0 FrameStrobe_O_i\[6\]
rlabel metal1 18492 2074 18492 2074 0 FrameStrobe_O_i\[7\]
rlabel metal1 20792 2414 20792 2414 0 FrameStrobe_O_i\[8\]
rlabel metal1 23736 2074 23736 2074 0 FrameStrobe_O_i\[9\]
rlabel metal2 5145 68 5145 68 0 N1END[0]
rlabel metal2 5658 415 5658 415 0 N1END[1]
rlabel metal2 5835 68 5835 68 0 N1END[2]
rlabel metal2 6111 68 6111 68 0 N1END[3]
rlabel metal2 8595 68 8595 68 0 N2END[0]
rlabel metal2 8970 670 8970 670 0 N2END[1]
rlabel metal2 9246 704 9246 704 0 N2END[2]
rlabel metal2 9522 670 9522 670 0 N2END[3]
rlabel metal2 9798 670 9798 670 0 N2END[4]
rlabel metal2 10074 398 10074 398 0 N2END[5]
rlabel metal2 10350 636 10350 636 0 N2END[6]
rlabel metal2 10626 398 10626 398 0 N2END[7]
rlabel metal2 6585 68 6585 68 0 N2MID[0]
rlabel metal2 6762 398 6762 398 0 N2MID[1]
rlabel metal1 6394 1292 6394 1292 0 N2MID[2]
rlabel metal2 6854 1377 6854 1377 0 N2MID[3]
rlabel metal2 7590 670 7590 670 0 N2MID[4]
rlabel metal2 7767 68 7767 68 0 N2MID[5]
rlabel metal2 8142 398 8142 398 0 N2MID[6]
rlabel metal2 8319 68 8319 68 0 N2MID[7]
rlabel metal2 10902 670 10902 670 0 N4END[0]
rlabel metal2 13715 68 13715 68 0 N4END[10]
rlabel metal2 13885 68 13885 68 0 N4END[11]
rlabel metal2 14115 68 14115 68 0 N4END[12]
rlabel metal2 14391 68 14391 68 0 N4END[13]
rlabel metal2 14766 670 14766 670 0 N4END[14]
rlabel metal2 15095 68 15095 68 0 N4END[15]
rlabel metal2 11178 347 11178 347 0 N4END[1]
rlabel metal2 11454 670 11454 670 0 N4END[2]
rlabel metal2 11730 398 11730 398 0 N4END[3]
rlabel metal2 12006 670 12006 670 0 N4END[4]
rlabel metal2 12229 68 12229 68 0 N4END[5]
rlabel metal2 12374 697 12374 697 0 N4END[6]
rlabel metal2 12735 68 12735 68 0 N4END[7]
rlabel metal2 13057 68 13057 68 0 N4END[8]
rlabel metal2 13287 68 13287 68 0 N4END[9]
rlabel metal2 15265 68 15265 68 0 NN4END[0]
rlabel metal2 18078 636 18078 636 0 NN4END[10]
rlabel metal2 18354 738 18354 738 0 NN4END[11]
rlabel metal2 18531 68 18531 68 0 NN4END[12]
rlabel metal2 18906 364 18906 364 0 NN4END[13]
rlabel metal2 19182 398 19182 398 0 NN4END[14]
rlabel metal2 19458 364 19458 364 0 NN4END[15]
rlabel metal2 15495 68 15495 68 0 NN4END[1]
rlabel metal2 15870 738 15870 738 0 NN4END[2]
rlabel metal2 16146 670 16146 670 0 NN4END[3]
rlabel metal2 16422 398 16422 398 0 NN4END[4]
rlabel metal2 16698 364 16698 364 0 NN4END[5]
rlabel metal2 16974 670 16974 670 0 NN4END[6]
rlabel metal2 17151 68 17151 68 0 NN4END[7]
rlabel metal2 17427 68 17427 68 0 NN4END[8]
rlabel metal2 17703 68 17703 68 0 NN4END[9]
rlabel metal2 19734 908 19734 908 0 S1BEG[0]
rlabel metal2 20010 908 20010 908 0 S1BEG[1]
rlabel metal2 20286 262 20286 262 0 S1BEG[2]
rlabel metal2 20463 68 20463 68 0 S1BEG[3]
rlabel metal2 23099 68 23099 68 0 S2BEG[0]
rlabel metal2 23322 806 23322 806 0 S2BEG[1]
rlabel metal2 23598 636 23598 636 0 S2BEG[2]
rlabel metal2 23874 687 23874 687 0 S2BEG[3]
rlabel metal2 24249 68 24249 68 0 S2BEG[4]
rlabel metal2 24426 228 24426 228 0 S2BEG[5]
rlabel metal2 24755 68 24755 68 0 S2BEG[6]
rlabel metal2 25077 68 25077 68 0 S2BEG[7]
rlabel metal2 20838 636 20838 636 0 S2BEGb[0]
rlabel metal2 21114 908 21114 908 0 S2BEGb[1]
rlabel metal2 21390 364 21390 364 0 S2BEGb[2]
rlabel metal2 21613 68 21613 68 0 S2BEGb[3]
rlabel metal2 21942 908 21942 908 0 S2BEGb[4]
rlabel metal2 22218 738 22218 738 0 S2BEGb[5]
rlabel metal2 22494 500 22494 500 0 S2BEGb[6]
rlabel metal2 22770 636 22770 636 0 S2BEGb[7]
rlabel metal2 25254 908 25254 908 0 S4BEG[0]
rlabel metal2 28067 68 28067 68 0 S4BEG[10]
rlabel metal2 28290 1180 28290 1180 0 S4BEG[11]
rlabel metal2 28566 942 28566 942 0 S4BEG[12]
rlabel metal2 28895 68 28895 68 0 S4BEG[13]
rlabel metal2 29217 68 29217 68 0 S4BEG[14]
rlabel metal2 29394 806 29394 806 0 S4BEG[15]
rlabel metal2 25530 347 25530 347 0 S4BEG[1]
rlabel metal2 25806 908 25806 908 0 S4BEG[2]
rlabel metal2 26082 500 26082 500 0 S4BEG[3]
rlabel metal2 26358 976 26358 976 0 S4BEG[4]
rlabel metal2 26687 68 26687 68 0 S4BEG[5]
rlabel metal2 26910 772 26910 772 0 S4BEG[6]
rlabel metal2 27186 347 27186 347 0 S4BEG[7]
rlabel metal2 27462 908 27462 908 0 S4BEG[8]
rlabel metal2 27738 806 27738 806 0 S4BEG[9]
rlabel metal2 29670 908 29670 908 0 SS4BEG[0]
rlabel metal2 32483 68 32483 68 0 SS4BEG[10]
rlabel metal2 32805 68 32805 68 0 SS4BEG[11]
rlabel metal2 32982 908 32982 908 0 SS4BEG[12]
rlabel metal2 33357 68 33357 68 0 SS4BEG[13]
rlabel metal2 33534 908 33534 908 0 SS4BEG[14]
rlabel metal2 33909 68 33909 68 0 SS4BEG[15]
rlabel metal1 32154 1462 32154 1462 0 SS4BEG[1]
rlabel metal1 31878 1292 31878 1292 0 SS4BEG[2]
rlabel metal1 31878 1802 31878 1802 0 SS4BEG[3]
rlabel metal2 30873 68 30873 68 0 SS4BEG[4]
rlabel metal2 31149 68 31149 68 0 SS4BEG[5]
rlabel metal2 31970 1632 31970 1632 0 SS4BEG[6]
rlabel metal2 31878 1360 31878 1360 0 SS4BEG[7]
rlabel metal2 31977 68 31977 68 0 SS4BEG[8]
rlabel metal2 32253 68 32253 68 0 SS4BEG[9]
rlabel metal2 34086 704 34086 704 0 UserCLK
rlabel metal2 1334 9173 1334 9173 0 UserCLKo
rlabel metal2 36202 1088 36202 1088 0 net1
rlabel metal1 40710 1530 40710 1530 0 net10
rlabel metal1 23874 1292 23874 1292 0 net100
rlabel metal1 24196 1326 24196 1326 0 net101
rlabel metal1 24794 1258 24794 1258 0 net102
rlabel metal1 25208 1258 25208 1258 0 net103
rlabel metal1 25392 1326 25392 1326 0 net104
rlabel metal1 26864 1326 26864 1326 0 net105
rlabel metal1 20562 1326 20562 1326 0 net106
rlabel metal1 20884 2006 20884 2006 0 net107
rlabel metal1 20286 1360 20286 1360 0 net108
rlabel metal1 21390 2448 21390 2448 0 net109
rlabel metal2 41538 1734 41538 1734 0 net11
rlabel metal1 21896 1938 21896 1938 0 net110
rlabel metal1 21436 1258 21436 1258 0 net111
rlabel metal1 21344 1326 21344 1326 0 net112
rlabel metal2 22034 1802 22034 1802 0 net113
rlabel metal1 25254 2006 25254 2006 0 net114
rlabel metal1 30084 1326 30084 1326 0 net115
rlabel metal1 28382 2380 28382 2380 0 net116
rlabel metal1 28750 2006 28750 2006 0 net117
rlabel metal1 30314 1258 30314 1258 0 net118
rlabel viali 30314 1940 30314 1940 0 net119
rlabel metal2 36662 1020 36662 1020 0 net12
rlabel metal1 31786 1224 31786 1224 0 net120
rlabel metal1 27591 1326 27591 1326 0 net121
rlabel metal1 25990 2040 25990 2040 0 net122
rlabel metal1 28014 1326 28014 1326 0 net123
rlabel metal1 27094 2040 27094 2040 0 net124
rlabel metal1 29210 1224 29210 1224 0 net125
rlabel metal1 27830 2006 27830 2006 0 net126
rlabel metal1 29578 1258 29578 1258 0 net127
rlabel metal1 28014 1938 28014 1938 0 net128
rlabel metal2 28980 2278 28980 2278 0 net129
rlabel metal2 36938 646 36938 646 0 net13
rlabel metal1 29624 1938 29624 1938 0 net130
rlabel metal1 34316 2006 34316 2006 0 net131
rlabel metal2 21850 748 21850 748 0 net132
rlabel metal1 15962 1972 15962 1972 0 net133
rlabel metal2 34914 3060 34914 3060 0 net134
rlabel metal1 32706 1904 32706 1904 0 net135
rlabel metal1 35420 1326 35420 1326 0 net136
rlabel metal2 19458 1088 19458 1088 0 net137
rlabel metal2 18906 1258 18906 1258 0 net138
rlabel metal1 31993 2006 31993 2006 0 net139
rlabel metal1 37306 1258 37306 1258 0 net14
rlabel metal1 19090 2312 19090 2312 0 net140
rlabel metal1 19826 1496 19826 1496 0 net141
rlabel metal3 26036 3128 26036 3128 0 net142
rlabel metal2 33948 4012 33948 4012 0 net143
rlabel metal1 17480 2074 17480 2074 0 net144
rlabel metal1 16928 2074 16928 2074 0 net145
rlabel metal1 9614 8568 9614 8568 0 net146
rlabel metal1 37766 1394 37766 1394 0 net15
rlabel metal2 37398 782 37398 782 0 net16
rlabel metal3 21597 1292 21597 1292 0 net17
rlabel metal2 18354 2023 18354 2023 0 net18
rlabel metal3 21620 340 21620 340 0 net19
rlabel metal2 34730 714 34730 714 0 net2
rlabel metal2 38870 1020 38870 1020 0 net20
rlabel metal1 5106 918 5106 918 0 net21
rlabel metal2 5382 2108 5382 2108 0 net22
rlabel metal2 5658 1088 5658 1088 0 net23
rlabel metal1 6118 476 6118 476 0 net24
rlabel metal1 8142 1190 8142 1190 0 net25
rlabel metal1 8602 646 8602 646 0 net26
rlabel metal1 8786 306 8786 306 0 net27
rlabel metal2 9154 646 9154 646 0 net28
rlabel metal1 20286 2448 20286 2448 0 net29
rlabel metal1 37559 3026 37559 3026 0 net3
rlabel metal1 19389 1938 19389 1938 0 net30
rlabel metal1 9982 884 9982 884 0 net31
rlabel metal2 10258 1190 10258 1190 0 net32
rlabel metal2 6762 3332 6762 3332 0 net33
rlabel metal2 6210 901 6210 901 0 net34
rlabel metal2 6578 765 6578 765 0 net35
rlabel metal2 6854 3094 6854 3094 0 net36
rlabel metal1 9890 816 9890 816 0 net37
rlabel via2 8326 1445 8326 1445 0 net38
rlabel metal1 7866 578 7866 578 0 net39
rlabel metal1 39468 1190 39468 1190 0 net4
rlabel metal1 8234 1530 8234 1530 0 net40
rlabel metal2 10994 969 10994 969 0 net41
rlabel metal2 17434 1751 17434 1751 0 net42
rlabel metal1 13432 1190 13432 1190 0 net43
rlabel metal2 13570 646 13570 646 0 net44
rlabel metal1 20470 2584 20470 2584 0 net45
rlabel metal2 25346 1360 25346 1360 0 net46
rlabel metal1 15778 1734 15778 1734 0 net47
rlabel metal2 10810 1751 10810 1751 0 net48
rlabel metal2 11270 1037 11270 1037 0 net49
rlabel metal2 39882 952 39882 952 0 net5
rlabel metal2 11362 2822 11362 2822 0 net50
rlabel metal1 11914 1190 11914 1190 0 net51
rlabel metal2 12006 3026 12006 3026 0 net52
rlabel metal2 12282 2244 12282 2244 0 net53
rlabel metal1 12558 1258 12558 1258 0 net54
rlabel metal2 12926 612 12926 612 0 net55
rlabel metal2 13294 748 13294 748 0 net56
rlabel metal1 14858 1462 14858 1462 0 net57
rlabel metal1 17434 1530 17434 1530 0 net58
rlabel metal2 17526 1513 17526 1513 0 net59
rlabel metal1 39974 1190 39974 1190 0 net6
rlabel metal1 18124 1530 18124 1530 0 net60
rlabel metal1 18078 1224 18078 1224 0 net61
rlabel metal1 19274 1292 19274 1292 0 net62
rlabel metal1 18906 1530 18906 1530 0 net63
rlabel metal2 14674 1972 14674 1972 0 net64
rlabel metal2 14950 1700 14950 1700 0 net65
rlabel metal1 15502 1530 15502 1530 0 net66
rlabel metal1 15686 1462 15686 1462 0 net67
rlabel metal1 16008 1190 16008 1190 0 net68
rlabel metal1 16238 1530 16238 1530 0 net69
rlabel metal1 40342 1190 40342 1190 0 net7
rlabel metal1 16468 1462 16468 1462 0 net70
rlabel metal1 16928 1190 16928 1190 0 net71
rlabel metal1 17066 1530 17066 1530 0 net72
rlabel metal2 34546 748 34546 748 0 net73
rlabel via2 4462 8347 4462 8347 0 net74
rlabel metal1 24840 8466 24840 8466 0 net75
rlabel metal1 27232 2618 27232 2618 0 net76
rlabel metal1 30130 2346 30130 2346 0 net77
rlabel metal1 31234 2618 31234 2618 0 net78
rlabel metal1 33304 8466 33304 8466 0 net79
rlabel metal2 40710 1530 40710 1530 0 net8
rlabel metal1 36133 8330 36133 8330 0 net80
rlabel metal1 37582 2618 37582 2618 0 net81
rlabel metal1 39744 2618 39744 2618 0 net82
rlabel metal1 41216 8466 41216 8466 0 net83
rlabel metal1 42780 2618 42780 2618 0 net84
rlabel via2 5566 8483 5566 8483 0 net85
rlabel metal1 7774 8432 7774 8432 0 net86
rlabel via1 9789 8466 9789 8466 0 net87
rlabel metal2 13938 8636 13938 8636 0 net88
rlabel metal2 14122 5542 14122 5542 0 net89
rlabel metal1 40526 1462 40526 1462 0 net9
rlabel metal1 16468 2618 16468 2618 0 net90
rlabel metal1 18630 2448 18630 2448 0 net91
rlabel metal2 20562 2689 20562 2689 0 net92
rlabel metal1 22770 8466 22770 8466 0 net93
rlabel metal1 19550 1972 19550 1972 0 net94
rlabel metal1 19136 1190 19136 1190 0 net95
rlabel metal2 19504 2788 19504 2788 0 net96
rlabel metal1 19872 1326 19872 1326 0 net97
rlabel metal1 22954 1360 22954 1360 0 net98
rlabel metal1 23322 1326 23322 1326 0 net99
<< properties >>
string FIXED_BBOX 0 0 45000 10000
<< end >>
